magic
tech gf180mcuD
magscale 1 10
timestamp 1699375940
<< metal1 >>
rect 6738 56590 6750 56642
rect 6802 56639 6814 56642
rect 7298 56639 7310 56642
rect 6802 56593 7310 56639
rect 6802 56590 6814 56593
rect 7298 56590 7310 56593
rect 7362 56590 7374 56642
rect 43698 56590 43710 56642
rect 43762 56639 43774 56642
rect 44370 56639 44382 56642
rect 43762 56593 44382 56639
rect 43762 56590 43774 56593
rect 44370 56590 44382 56593
rect 44434 56590 44446 56642
rect 56018 56590 56030 56642
rect 56082 56639 56094 56642
rect 57026 56639 57038 56642
rect 56082 56593 57038 56639
rect 56082 56590 56094 56593
rect 57026 56590 57038 56593
rect 57090 56590 57102 56642
rect 80658 56590 80670 56642
rect 80722 56639 80734 56642
rect 82226 56639 82238 56642
rect 80722 56593 82238 56639
rect 80722 56590 80734 56593
rect 82226 56590 82238 56593
rect 82290 56590 82302 56642
rect 92978 56590 92990 56642
rect 93042 56639 93054 56642
rect 93986 56639 93998 56642
rect 93042 56593 93998 56639
rect 93042 56590 93054 56593
rect 93986 56590 93998 56593
rect 94050 56590 94062 56642
rect 1344 56474 98560 56508
rect 1344 56422 8896 56474
rect 8948 56422 9020 56474
rect 9072 56422 9144 56474
rect 9196 56422 9268 56474
rect 9320 56422 17896 56474
rect 17948 56422 18020 56474
rect 18072 56422 18144 56474
rect 18196 56422 18268 56474
rect 18320 56422 26896 56474
rect 26948 56422 27020 56474
rect 27072 56422 27144 56474
rect 27196 56422 27268 56474
rect 27320 56422 35896 56474
rect 35948 56422 36020 56474
rect 36072 56422 36144 56474
rect 36196 56422 36268 56474
rect 36320 56422 44896 56474
rect 44948 56422 45020 56474
rect 45072 56422 45144 56474
rect 45196 56422 45268 56474
rect 45320 56422 53896 56474
rect 53948 56422 54020 56474
rect 54072 56422 54144 56474
rect 54196 56422 54268 56474
rect 54320 56422 62896 56474
rect 62948 56422 63020 56474
rect 63072 56422 63144 56474
rect 63196 56422 63268 56474
rect 63320 56422 71896 56474
rect 71948 56422 72020 56474
rect 72072 56422 72144 56474
rect 72196 56422 72268 56474
rect 72320 56422 80896 56474
rect 80948 56422 81020 56474
rect 81072 56422 81144 56474
rect 81196 56422 81268 56474
rect 81320 56422 89896 56474
rect 89948 56422 90020 56474
rect 90072 56422 90144 56474
rect 90196 56422 90268 56474
rect 90320 56422 98560 56474
rect 1344 56388 98560 56422
rect 32174 56306 32226 56318
rect 32174 56242 32226 56254
rect 57038 56306 57090 56318
rect 57038 56242 57090 56254
rect 93998 56306 94050 56318
rect 93998 56242 94050 56254
rect 97694 56306 97746 56318
rect 97694 56242 97746 56254
rect 2046 56194 2098 56206
rect 7298 56142 7310 56194
rect 7362 56142 7374 56194
rect 2046 56130 2098 56142
rect 1710 56082 1762 56094
rect 43934 56082 43986 56094
rect 8194 56030 8206 56082
rect 8258 56030 8270 56082
rect 20066 56030 20078 56082
rect 20130 56030 20142 56082
rect 32834 56030 32846 56082
rect 32898 56030 32910 56082
rect 1710 56018 1762 56030
rect 43934 56018 43986 56030
rect 56254 56082 56306 56094
rect 56254 56018 56306 56030
rect 68462 56082 68514 56094
rect 68462 56018 68514 56030
rect 81678 56082 81730 56094
rect 81678 56018 81730 56030
rect 93214 56082 93266 56094
rect 93214 56018 93266 56030
rect 96350 56082 96402 56094
rect 96350 56018 96402 56030
rect 96910 56082 96962 56094
rect 96910 56018 96962 56030
rect 98142 56082 98194 56094
rect 98142 56018 98194 56030
rect 2494 55970 2546 55982
rect 2494 55906 2546 55918
rect 8766 55970 8818 55982
rect 19170 55918 19182 55970
rect 19234 55918 19246 55970
rect 44370 55918 44382 55970
rect 44434 55918 44446 55970
rect 69010 55918 69022 55970
rect 69074 55918 69086 55970
rect 82226 55918 82238 55970
rect 82290 55918 82302 55970
rect 95890 55918 95902 55970
rect 95954 55918 95966 55970
rect 8766 55906 8818 55918
rect 1344 55690 98560 55724
rect 1344 55638 4396 55690
rect 4448 55638 4520 55690
rect 4572 55638 4644 55690
rect 4696 55638 4768 55690
rect 4820 55638 13396 55690
rect 13448 55638 13520 55690
rect 13572 55638 13644 55690
rect 13696 55638 13768 55690
rect 13820 55638 22396 55690
rect 22448 55638 22520 55690
rect 22572 55638 22644 55690
rect 22696 55638 22768 55690
rect 22820 55638 31396 55690
rect 31448 55638 31520 55690
rect 31572 55638 31644 55690
rect 31696 55638 31768 55690
rect 31820 55638 40396 55690
rect 40448 55638 40520 55690
rect 40572 55638 40644 55690
rect 40696 55638 40768 55690
rect 40820 55638 49396 55690
rect 49448 55638 49520 55690
rect 49572 55638 49644 55690
rect 49696 55638 49768 55690
rect 49820 55638 58396 55690
rect 58448 55638 58520 55690
rect 58572 55638 58644 55690
rect 58696 55638 58768 55690
rect 58820 55638 67396 55690
rect 67448 55638 67520 55690
rect 67572 55638 67644 55690
rect 67696 55638 67768 55690
rect 67820 55638 76396 55690
rect 76448 55638 76520 55690
rect 76572 55638 76644 55690
rect 76696 55638 76768 55690
rect 76820 55638 85396 55690
rect 85448 55638 85520 55690
rect 85572 55638 85644 55690
rect 85696 55638 85768 55690
rect 85820 55638 94396 55690
rect 94448 55638 94520 55690
rect 94572 55638 94644 55690
rect 94696 55638 94768 55690
rect 94820 55638 98560 55690
rect 1344 55604 98560 55638
rect 32050 55358 32062 55410
rect 32114 55358 32126 55410
rect 36418 55358 36430 55410
rect 36482 55358 36494 55410
rect 42578 55358 42590 55410
rect 42642 55358 42654 55410
rect 48066 55358 48078 55410
rect 48130 55358 48142 55410
rect 33182 55298 33234 55310
rect 37102 55298 37154 55310
rect 43710 55298 43762 55310
rect 29250 55246 29262 55298
rect 29314 55246 29326 55298
rect 33618 55246 33630 55298
rect 33682 55246 33694 55298
rect 39778 55246 39790 55298
rect 39842 55246 39854 55298
rect 33182 55234 33234 55246
rect 37102 55234 37154 55246
rect 43710 55234 43762 55246
rect 44270 55298 44322 55310
rect 45154 55246 45166 55298
rect 45218 55246 45230 55298
rect 55794 55246 55806 55298
rect 55858 55246 55870 55298
rect 66882 55246 66894 55298
rect 66946 55246 66958 55298
rect 97010 55246 97022 55298
rect 97074 55246 97086 55298
rect 44270 55234 44322 55246
rect 1710 55186 1762 55198
rect 1710 55122 1762 55134
rect 25454 55186 25506 55198
rect 25454 55122 25506 55134
rect 25790 55186 25842 55198
rect 25790 55122 25842 55134
rect 26126 55186 26178 55198
rect 26126 55122 26178 55134
rect 26462 55186 26514 55198
rect 32398 55186 32450 55198
rect 29922 55134 29934 55186
rect 29986 55134 29998 55186
rect 26462 55122 26514 55134
rect 32398 55122 32450 55134
rect 32734 55186 32786 55198
rect 42926 55186 42978 55198
rect 34290 55134 34302 55186
rect 34354 55134 34366 55186
rect 40450 55134 40462 55186
rect 40514 55134 40526 55186
rect 32734 55122 32786 55134
rect 42926 55122 42978 55134
rect 43262 55186 43314 55198
rect 56030 55186 56082 55198
rect 45938 55134 45950 55186
rect 46002 55134 46014 55186
rect 43262 55122 43314 55134
rect 56030 55122 56082 55134
rect 58494 55186 58546 55198
rect 58494 55122 58546 55134
rect 67118 55186 67170 55198
rect 67118 55122 67170 55134
rect 68350 55186 68402 55198
rect 98018 55134 98030 55186
rect 98082 55134 98094 55186
rect 68350 55122 68402 55134
rect 2046 55074 2098 55086
rect 2046 55010 2098 55022
rect 2494 55074 2546 55086
rect 2494 55010 2546 55022
rect 48638 55074 48690 55086
rect 48638 55010 48690 55022
rect 52222 55074 52274 55086
rect 52222 55010 52274 55022
rect 52670 55074 52722 55086
rect 52670 55010 52722 55022
rect 52782 55074 52834 55086
rect 52782 55010 52834 55022
rect 52894 55074 52946 55086
rect 52894 55010 52946 55022
rect 53118 55074 53170 55086
rect 53118 55010 53170 55022
rect 57262 55074 57314 55086
rect 57262 55010 57314 55022
rect 57486 55074 57538 55086
rect 57486 55010 57538 55022
rect 57598 55074 57650 55086
rect 57598 55010 57650 55022
rect 57710 55074 57762 55086
rect 57710 55010 57762 55022
rect 57934 55074 57986 55086
rect 57934 55010 57986 55022
rect 58382 55074 58434 55086
rect 58382 55010 58434 55022
rect 68686 55074 68738 55086
rect 68686 55010 68738 55022
rect 96574 55074 96626 55086
rect 96574 55010 96626 55022
rect 1344 54906 98560 54940
rect 1344 54854 8896 54906
rect 8948 54854 9020 54906
rect 9072 54854 9144 54906
rect 9196 54854 9268 54906
rect 9320 54854 17896 54906
rect 17948 54854 18020 54906
rect 18072 54854 18144 54906
rect 18196 54854 18268 54906
rect 18320 54854 26896 54906
rect 26948 54854 27020 54906
rect 27072 54854 27144 54906
rect 27196 54854 27268 54906
rect 27320 54854 35896 54906
rect 35948 54854 36020 54906
rect 36072 54854 36144 54906
rect 36196 54854 36268 54906
rect 36320 54854 44896 54906
rect 44948 54854 45020 54906
rect 45072 54854 45144 54906
rect 45196 54854 45268 54906
rect 45320 54854 53896 54906
rect 53948 54854 54020 54906
rect 54072 54854 54144 54906
rect 54196 54854 54268 54906
rect 54320 54854 62896 54906
rect 62948 54854 63020 54906
rect 63072 54854 63144 54906
rect 63196 54854 63268 54906
rect 63320 54854 71896 54906
rect 71948 54854 72020 54906
rect 72072 54854 72144 54906
rect 72196 54854 72268 54906
rect 72320 54854 80896 54906
rect 80948 54854 81020 54906
rect 81072 54854 81144 54906
rect 81196 54854 81268 54906
rect 81320 54854 89896 54906
rect 89948 54854 90020 54906
rect 90072 54854 90144 54906
rect 90196 54854 90268 54906
rect 90320 54854 98560 54906
rect 1344 54820 98560 54854
rect 40350 54738 40402 54750
rect 40350 54674 40402 54686
rect 41246 54738 41298 54750
rect 41246 54674 41298 54686
rect 41358 54738 41410 54750
rect 41358 54674 41410 54686
rect 48862 54738 48914 54750
rect 48862 54674 48914 54686
rect 49646 54738 49698 54750
rect 49646 54674 49698 54686
rect 82126 54738 82178 54750
rect 82126 54674 82178 54686
rect 44606 54626 44658 54638
rect 44606 54562 44658 54574
rect 47742 54626 47794 54638
rect 49758 54626 49810 54638
rect 47954 54574 47966 54626
rect 48018 54574 48030 54626
rect 51762 54574 51774 54626
rect 51826 54574 51838 54626
rect 56802 54574 56814 54626
rect 56866 54574 56878 54626
rect 57474 54574 57486 54626
rect 57538 54574 57550 54626
rect 60498 54574 60510 54626
rect 60562 54574 60574 54626
rect 47742 54562 47794 54574
rect 49758 54562 49810 54574
rect 40238 54514 40290 54526
rect 41470 54514 41522 54526
rect 45166 54514 45218 54526
rect 40898 54462 40910 54514
rect 40962 54462 40974 54514
rect 43250 54462 43262 54514
rect 43314 54462 43326 54514
rect 44818 54462 44830 54514
rect 44882 54462 44894 54514
rect 40238 54450 40290 54462
rect 41470 54450 41522 54462
rect 45166 54450 45218 54462
rect 47294 54514 47346 54526
rect 47294 54450 47346 54462
rect 48750 54514 48802 54526
rect 48750 54450 48802 54462
rect 48974 54514 49026 54526
rect 48974 54450 49026 54462
rect 49422 54514 49474 54526
rect 54350 54514 54402 54526
rect 50978 54462 50990 54514
rect 51042 54462 51054 54514
rect 49422 54450 49474 54462
rect 54350 54450 54402 54462
rect 55582 54514 55634 54526
rect 55582 54450 55634 54462
rect 56030 54514 56082 54526
rect 81790 54514 81842 54526
rect 56578 54462 56590 54514
rect 56642 54462 56654 54514
rect 61282 54462 61294 54514
rect 61346 54462 61358 54514
rect 56030 54450 56082 54462
rect 81790 54450 81842 54462
rect 35198 54402 35250 54414
rect 35198 54338 35250 54350
rect 36318 54402 36370 54414
rect 36318 54338 36370 54350
rect 36766 54402 36818 54414
rect 36766 54338 36818 54350
rect 39902 54402 39954 54414
rect 39902 54338 39954 54350
rect 41918 54402 41970 54414
rect 45502 54402 45554 54414
rect 44146 54350 44158 54402
rect 44210 54350 44222 54402
rect 41918 54338 41970 54350
rect 45502 54338 45554 54350
rect 45950 54402 46002 54414
rect 45950 54338 46002 54350
rect 48078 54402 48130 54414
rect 48078 54338 48130 54350
rect 50654 54402 50706 54414
rect 57822 54402 57874 54414
rect 61854 54402 61906 54414
rect 53890 54350 53902 54402
rect 53954 54350 53966 54402
rect 58370 54350 58382 54402
rect 58434 54350 58446 54402
rect 50654 54338 50706 54350
rect 57822 54338 57874 54350
rect 61854 54338 61906 54350
rect 65774 54402 65826 54414
rect 65774 54338 65826 54350
rect 81454 54402 81506 54414
rect 81454 54338 81506 54350
rect 44942 54290 44994 54302
rect 44942 54226 44994 54238
rect 47070 54290 47122 54302
rect 47070 54226 47122 54238
rect 54238 54290 54290 54302
rect 54238 54226 54290 54238
rect 1344 54122 98560 54156
rect 1344 54070 4396 54122
rect 4448 54070 4520 54122
rect 4572 54070 4644 54122
rect 4696 54070 4768 54122
rect 4820 54070 13396 54122
rect 13448 54070 13520 54122
rect 13572 54070 13644 54122
rect 13696 54070 13768 54122
rect 13820 54070 22396 54122
rect 22448 54070 22520 54122
rect 22572 54070 22644 54122
rect 22696 54070 22768 54122
rect 22820 54070 31396 54122
rect 31448 54070 31520 54122
rect 31572 54070 31644 54122
rect 31696 54070 31768 54122
rect 31820 54070 40396 54122
rect 40448 54070 40520 54122
rect 40572 54070 40644 54122
rect 40696 54070 40768 54122
rect 40820 54070 49396 54122
rect 49448 54070 49520 54122
rect 49572 54070 49644 54122
rect 49696 54070 49768 54122
rect 49820 54070 58396 54122
rect 58448 54070 58520 54122
rect 58572 54070 58644 54122
rect 58696 54070 58768 54122
rect 58820 54070 67396 54122
rect 67448 54070 67520 54122
rect 67572 54070 67644 54122
rect 67696 54070 67768 54122
rect 67820 54070 76396 54122
rect 76448 54070 76520 54122
rect 76572 54070 76644 54122
rect 76696 54070 76768 54122
rect 76820 54070 85396 54122
rect 85448 54070 85520 54122
rect 85572 54070 85644 54122
rect 85696 54070 85768 54122
rect 85820 54070 94396 54122
rect 94448 54070 94520 54122
rect 94572 54070 94644 54122
rect 94696 54070 94768 54122
rect 94820 54070 98560 54122
rect 1344 54036 98560 54070
rect 59278 53954 59330 53966
rect 59278 53890 59330 53902
rect 30046 53842 30098 53854
rect 30046 53778 30098 53790
rect 34526 53842 34578 53854
rect 34526 53778 34578 53790
rect 35310 53842 35362 53854
rect 35310 53778 35362 53790
rect 36318 53842 36370 53854
rect 59166 53842 59218 53854
rect 48738 53790 48750 53842
rect 48802 53790 48814 53842
rect 36318 53778 36370 53790
rect 59166 53778 59218 53790
rect 65326 53842 65378 53854
rect 65326 53778 65378 53790
rect 72830 53842 72882 53854
rect 72830 53778 72882 53790
rect 28478 53730 28530 53742
rect 35086 53730 35138 53742
rect 41694 53730 41746 53742
rect 29586 53678 29598 53730
rect 29650 53678 29662 53730
rect 35634 53678 35646 53730
rect 35698 53678 35710 53730
rect 37202 53678 37214 53730
rect 37266 53678 37278 53730
rect 38210 53678 38222 53730
rect 38274 53678 38286 53730
rect 41346 53678 41358 53730
rect 41410 53678 41422 53730
rect 28478 53666 28530 53678
rect 35086 53666 35138 53678
rect 41694 53666 41746 53678
rect 44942 53730 44994 53742
rect 56814 53730 56866 53742
rect 46050 53678 46062 53730
rect 46114 53678 46126 53730
rect 52770 53678 52782 53730
rect 52834 53678 52846 53730
rect 56578 53678 56590 53730
rect 56642 53678 56654 53730
rect 44942 53666 44994 53678
rect 56814 53666 56866 53678
rect 57486 53730 57538 53742
rect 57486 53666 57538 53678
rect 65214 53730 65266 53742
rect 66334 53730 66386 53742
rect 66782 53730 66834 53742
rect 65426 53678 65438 53730
rect 65490 53678 65502 53730
rect 65986 53678 65998 53730
rect 66050 53678 66062 53730
rect 66546 53678 66558 53730
rect 66610 53678 66622 53730
rect 65214 53666 65266 53678
rect 66334 53666 66386 53678
rect 66782 53666 66834 53678
rect 67118 53730 67170 53742
rect 69906 53678 69918 53730
rect 69970 53678 69982 53730
rect 96898 53678 96910 53730
rect 96962 53678 96974 53730
rect 67118 53666 67170 53678
rect 1710 53618 1762 53630
rect 1710 53554 1762 53566
rect 30830 53618 30882 53630
rect 30830 53554 30882 53566
rect 35870 53618 35922 53630
rect 40798 53618 40850 53630
rect 37314 53566 37326 53618
rect 37378 53566 37390 53618
rect 38882 53566 38894 53618
rect 38946 53566 38958 53618
rect 35870 53554 35922 53566
rect 40798 53554 40850 53566
rect 42254 53618 42306 53630
rect 64878 53618 64930 53630
rect 52882 53566 52894 53618
rect 52946 53566 52958 53618
rect 56466 53566 56478 53618
rect 56530 53566 56542 53618
rect 42254 53554 42306 53566
rect 64878 53554 64930 53566
rect 66670 53618 66722 53630
rect 66670 53554 66722 53566
rect 67230 53618 67282 53630
rect 70690 53566 70702 53618
rect 70754 53566 70766 53618
rect 98018 53566 98030 53618
rect 98082 53566 98094 53618
rect 67230 53554 67282 53566
rect 2046 53506 2098 53518
rect 2046 53442 2098 53454
rect 2494 53506 2546 53518
rect 2494 53442 2546 53454
rect 29262 53506 29314 53518
rect 29262 53442 29314 53454
rect 29934 53506 29986 53518
rect 29934 53442 29986 53454
rect 30158 53506 30210 53518
rect 30158 53442 30210 53454
rect 30718 53506 30770 53518
rect 30718 53442 30770 53454
rect 31278 53506 31330 53518
rect 31278 53442 31330 53454
rect 34414 53506 34466 53518
rect 34414 53442 34466 53454
rect 34638 53506 34690 53518
rect 34638 53442 34690 53454
rect 35422 53506 35474 53518
rect 35422 53442 35474 53454
rect 36206 53506 36258 53518
rect 43822 53506 43874 53518
rect 38322 53454 38334 53506
rect 38386 53454 38398 53506
rect 41234 53454 41246 53506
rect 41298 53454 41310 53506
rect 36206 53442 36258 53454
rect 43822 53442 43874 53454
rect 44270 53506 44322 53518
rect 44270 53442 44322 53454
rect 52110 53506 52162 53518
rect 57262 53506 57314 53518
rect 56354 53454 56366 53506
rect 56418 53454 56430 53506
rect 52110 53442 52162 53454
rect 57262 53442 57314 53454
rect 57374 53506 57426 53518
rect 57374 53442 57426 53454
rect 57934 53506 57986 53518
rect 57934 53442 57986 53454
rect 59054 53506 59106 53518
rect 59054 53442 59106 53454
rect 64542 53506 64594 53518
rect 64542 53442 64594 53454
rect 65662 53506 65714 53518
rect 65662 53442 65714 53454
rect 67678 53506 67730 53518
rect 67678 53442 67730 53454
rect 69582 53506 69634 53518
rect 69582 53442 69634 53454
rect 1344 53338 98560 53372
rect 1344 53286 8896 53338
rect 8948 53286 9020 53338
rect 9072 53286 9144 53338
rect 9196 53286 9268 53338
rect 9320 53286 17896 53338
rect 17948 53286 18020 53338
rect 18072 53286 18144 53338
rect 18196 53286 18268 53338
rect 18320 53286 26896 53338
rect 26948 53286 27020 53338
rect 27072 53286 27144 53338
rect 27196 53286 27268 53338
rect 27320 53286 35896 53338
rect 35948 53286 36020 53338
rect 36072 53286 36144 53338
rect 36196 53286 36268 53338
rect 36320 53286 44896 53338
rect 44948 53286 45020 53338
rect 45072 53286 45144 53338
rect 45196 53286 45268 53338
rect 45320 53286 53896 53338
rect 53948 53286 54020 53338
rect 54072 53286 54144 53338
rect 54196 53286 54268 53338
rect 54320 53286 62896 53338
rect 62948 53286 63020 53338
rect 63072 53286 63144 53338
rect 63196 53286 63268 53338
rect 63320 53286 71896 53338
rect 71948 53286 72020 53338
rect 72072 53286 72144 53338
rect 72196 53286 72268 53338
rect 72320 53286 80896 53338
rect 80948 53286 81020 53338
rect 81072 53286 81144 53338
rect 81196 53286 81268 53338
rect 81320 53286 89896 53338
rect 89948 53286 90020 53338
rect 90072 53286 90144 53338
rect 90196 53286 90268 53338
rect 90320 53286 98560 53338
rect 1344 53252 98560 53286
rect 29038 53170 29090 53182
rect 35534 53170 35586 53182
rect 33842 53118 33854 53170
rect 33906 53118 33918 53170
rect 29038 53106 29090 53118
rect 35534 53106 35586 53118
rect 35870 53170 35922 53182
rect 35870 53106 35922 53118
rect 36990 53170 37042 53182
rect 36990 53106 37042 53118
rect 39230 53170 39282 53182
rect 39230 53106 39282 53118
rect 39454 53170 39506 53182
rect 39454 53106 39506 53118
rect 48862 53170 48914 53182
rect 48862 53106 48914 53118
rect 48974 53170 49026 53182
rect 48974 53106 49026 53118
rect 51214 53170 51266 53182
rect 51214 53106 51266 53118
rect 51662 53170 51714 53182
rect 51662 53106 51714 53118
rect 60174 53170 60226 53182
rect 60174 53106 60226 53118
rect 2046 53058 2098 53070
rect 2046 52994 2098 53006
rect 27694 53058 27746 53070
rect 27694 52994 27746 53006
rect 29598 53058 29650 53070
rect 40910 53058 40962 53070
rect 50430 53058 50482 53070
rect 29810 53006 29822 53058
rect 29874 53006 29886 53058
rect 33730 53006 33742 53058
rect 33794 53006 33806 53058
rect 35186 53006 35198 53058
rect 35250 53006 35262 53058
rect 29598 52994 29650 53006
rect 35646 53002 35698 53014
rect 1710 52946 1762 52958
rect 1710 52882 1762 52894
rect 27918 52946 27970 52958
rect 27918 52882 27970 52894
rect 28142 52946 28194 52958
rect 28142 52882 28194 52894
rect 28590 52946 28642 52958
rect 28590 52882 28642 52894
rect 28814 52946 28866 52958
rect 28814 52882 28866 52894
rect 29150 52946 29202 52958
rect 31278 52946 31330 52958
rect 45490 53006 45502 53058
rect 45554 53006 45566 53058
rect 49746 53006 49758 53058
rect 49810 53006 49822 53058
rect 40910 52994 40962 53006
rect 50430 52994 50482 53006
rect 50766 53058 50818 53070
rect 50766 52994 50818 53006
rect 58046 53058 58098 53070
rect 58046 52994 58098 53006
rect 59502 53058 59554 53070
rect 65986 53006 65998 53058
rect 66050 53006 66062 53058
rect 59502 52994 59554 53006
rect 30370 52894 30382 52946
rect 30434 52894 30446 52946
rect 34290 52894 34302 52946
rect 34354 52894 34366 52946
rect 35298 52894 35310 52946
rect 35362 52894 35374 52946
rect 35646 52938 35698 52950
rect 36206 52946 36258 52958
rect 41358 52946 41410 52958
rect 49086 52946 49138 52958
rect 39666 52894 39678 52946
rect 39730 52894 39742 52946
rect 41122 52894 41134 52946
rect 41186 52894 41198 52946
rect 41570 52894 41582 52946
rect 41634 52894 41646 52946
rect 46610 52894 46622 52946
rect 46674 52894 46686 52946
rect 29150 52882 29202 52894
rect 31278 52882 31330 52894
rect 36206 52882 36258 52894
rect 41358 52882 41410 52894
rect 49086 52882 49138 52894
rect 49422 52946 49474 52958
rect 49422 52882 49474 52894
rect 50206 52946 50258 52958
rect 55582 52946 55634 52958
rect 68798 52946 68850 52958
rect 50978 52894 50990 52946
rect 51042 52894 51054 52946
rect 56914 52894 56926 52946
rect 56978 52894 56990 52946
rect 58930 52894 58942 52946
rect 58994 52894 59006 52946
rect 65202 52894 65214 52946
rect 65266 52894 65278 52946
rect 50206 52882 50258 52894
rect 55582 52882 55634 52894
rect 68798 52882 68850 52894
rect 2494 52834 2546 52846
rect 2494 52770 2546 52782
rect 28030 52834 28082 52846
rect 28030 52770 28082 52782
rect 29710 52834 29762 52846
rect 29710 52770 29762 52782
rect 30830 52834 30882 52846
rect 30830 52770 30882 52782
rect 36542 52834 36594 52846
rect 36542 52770 36594 52782
rect 38446 52834 38498 52846
rect 38446 52770 38498 52782
rect 38894 52834 38946 52846
rect 38894 52770 38946 52782
rect 39566 52834 39618 52846
rect 39566 52770 39618 52782
rect 40126 52834 40178 52846
rect 40126 52770 40178 52782
rect 41022 52834 41074 52846
rect 41022 52770 41074 52782
rect 48190 52834 48242 52846
rect 48190 52770 48242 52782
rect 50318 52834 50370 52846
rect 50318 52770 50370 52782
rect 50878 52834 50930 52846
rect 50878 52770 50930 52782
rect 52446 52834 52498 52846
rect 52446 52770 52498 52782
rect 55134 52834 55186 52846
rect 55134 52770 55186 52782
rect 56030 52834 56082 52846
rect 56030 52770 56082 52782
rect 68126 52834 68178 52846
rect 68126 52770 68178 52782
rect 28478 52722 28530 52734
rect 28478 52658 28530 52670
rect 30046 52722 30098 52734
rect 30046 52658 30098 52670
rect 49982 52722 50034 52734
rect 55010 52670 55022 52722
rect 55074 52719 55086 52722
rect 55570 52719 55582 52722
rect 55074 52673 55582 52719
rect 55074 52670 55086 52673
rect 55570 52670 55582 52673
rect 55634 52670 55646 52722
rect 49982 52658 50034 52670
rect 1344 52554 98560 52588
rect 1344 52502 4396 52554
rect 4448 52502 4520 52554
rect 4572 52502 4644 52554
rect 4696 52502 4768 52554
rect 4820 52502 13396 52554
rect 13448 52502 13520 52554
rect 13572 52502 13644 52554
rect 13696 52502 13768 52554
rect 13820 52502 22396 52554
rect 22448 52502 22520 52554
rect 22572 52502 22644 52554
rect 22696 52502 22768 52554
rect 22820 52502 31396 52554
rect 31448 52502 31520 52554
rect 31572 52502 31644 52554
rect 31696 52502 31768 52554
rect 31820 52502 40396 52554
rect 40448 52502 40520 52554
rect 40572 52502 40644 52554
rect 40696 52502 40768 52554
rect 40820 52502 49396 52554
rect 49448 52502 49520 52554
rect 49572 52502 49644 52554
rect 49696 52502 49768 52554
rect 49820 52502 58396 52554
rect 58448 52502 58520 52554
rect 58572 52502 58644 52554
rect 58696 52502 58768 52554
rect 58820 52502 67396 52554
rect 67448 52502 67520 52554
rect 67572 52502 67644 52554
rect 67696 52502 67768 52554
rect 67820 52502 76396 52554
rect 76448 52502 76520 52554
rect 76572 52502 76644 52554
rect 76696 52502 76768 52554
rect 76820 52502 85396 52554
rect 85448 52502 85520 52554
rect 85572 52502 85644 52554
rect 85696 52502 85768 52554
rect 85820 52502 94396 52554
rect 94448 52502 94520 52554
rect 94572 52502 94644 52554
rect 94696 52502 94768 52554
rect 94820 52502 98560 52554
rect 1344 52468 98560 52502
rect 27918 52386 27970 52398
rect 27918 52322 27970 52334
rect 28478 52386 28530 52398
rect 28478 52322 28530 52334
rect 33294 52386 33346 52398
rect 33294 52322 33346 52334
rect 41918 52386 41970 52398
rect 57822 52386 57874 52398
rect 48738 52334 48750 52386
rect 48802 52383 48814 52386
rect 49746 52383 49758 52386
rect 48802 52337 49758 52383
rect 48802 52334 48814 52337
rect 49746 52334 49758 52337
rect 49810 52334 49822 52386
rect 41918 52322 41970 52334
rect 57822 52322 57874 52334
rect 58494 52386 58546 52398
rect 58494 52322 58546 52334
rect 65998 52386 66050 52398
rect 65998 52322 66050 52334
rect 28366 52274 28418 52286
rect 22978 52222 22990 52274
rect 23042 52222 23054 52274
rect 25106 52222 25118 52274
rect 25170 52222 25182 52274
rect 28366 52210 28418 52222
rect 29262 52274 29314 52286
rect 31726 52274 31778 52286
rect 30034 52222 30046 52274
rect 30098 52222 30110 52274
rect 29262 52210 29314 52222
rect 31726 52210 31778 52222
rect 32174 52274 32226 52286
rect 32174 52210 32226 52222
rect 35758 52274 35810 52286
rect 35758 52210 35810 52222
rect 45614 52274 45666 52286
rect 45614 52210 45666 52222
rect 46734 52274 46786 52286
rect 48302 52274 48354 52286
rect 47170 52222 47182 52274
rect 47234 52222 47246 52274
rect 46734 52210 46786 52222
rect 48302 52210 48354 52222
rect 48750 52274 48802 52286
rect 48750 52210 48802 52222
rect 49198 52274 49250 52286
rect 50766 52274 50818 52286
rect 50194 52222 50206 52274
rect 50258 52222 50270 52274
rect 49198 52210 49250 52222
rect 50766 52210 50818 52222
rect 51214 52274 51266 52286
rect 51214 52210 51266 52222
rect 53342 52274 53394 52286
rect 53342 52210 53394 52222
rect 53790 52274 53842 52286
rect 58606 52274 58658 52286
rect 66110 52274 66162 52286
rect 55682 52222 55694 52274
rect 55746 52222 55758 52274
rect 60498 52222 60510 52274
rect 60562 52222 60574 52274
rect 62626 52222 62638 52274
rect 62690 52222 62702 52274
rect 53790 52210 53842 52222
rect 58606 52210 58658 52222
rect 66110 52210 66162 52222
rect 66558 52274 66610 52286
rect 66558 52210 66610 52222
rect 26350 52162 26402 52174
rect 25890 52110 25902 52162
rect 25954 52110 25966 52162
rect 26350 52098 26402 52110
rect 27582 52162 27634 52174
rect 27582 52098 27634 52110
rect 28142 52162 28194 52174
rect 28142 52098 28194 52110
rect 30158 52162 30210 52174
rect 33406 52162 33458 52174
rect 31266 52110 31278 52162
rect 31330 52110 31342 52162
rect 32946 52110 32958 52162
rect 33010 52110 33022 52162
rect 30158 52098 30210 52110
rect 33406 52098 33458 52110
rect 33742 52162 33794 52174
rect 33742 52098 33794 52110
rect 34190 52162 34242 52174
rect 34190 52098 34242 52110
rect 36206 52162 36258 52174
rect 45950 52162 46002 52174
rect 47742 52162 47794 52174
rect 43810 52110 43822 52162
rect 43874 52110 43886 52162
rect 46162 52110 46174 52162
rect 46226 52110 46238 52162
rect 36206 52098 36258 52110
rect 45950 52098 46002 52110
rect 47742 52098 47794 52110
rect 49646 52162 49698 52174
rect 56814 52162 56866 52174
rect 57598 52162 57650 52174
rect 63870 52162 63922 52174
rect 54338 52110 54350 52162
rect 54402 52110 54414 52162
rect 55346 52110 55358 52162
rect 55410 52110 55422 52162
rect 56578 52110 56590 52162
rect 56642 52110 56654 52162
rect 56914 52110 56926 52162
rect 56978 52110 56990 52162
rect 63410 52110 63422 52162
rect 63474 52110 63486 52162
rect 49646 52098 49698 52110
rect 56814 52098 56866 52110
rect 57598 52098 57650 52110
rect 63870 52098 63922 52110
rect 97694 52162 97746 52174
rect 97694 52098 97746 52110
rect 26910 52050 26962 52062
rect 26910 51986 26962 51998
rect 27806 52050 27858 52062
rect 49982 52050 50034 52062
rect 56366 52050 56418 52062
rect 29698 51998 29710 52050
rect 29762 51998 29774 52050
rect 31154 51998 31166 52050
rect 31218 51998 31230 52050
rect 54450 51998 54462 52050
rect 54514 51998 54526 52050
rect 56018 51998 56030 52050
rect 56082 51998 56094 52050
rect 27806 51986 27858 51998
rect 49982 51986 50034 51998
rect 56366 51986 56418 51998
rect 57934 52050 57986 52062
rect 57934 51986 57986 51998
rect 58158 52050 58210 52062
rect 58158 51986 58210 51998
rect 27022 51938 27074 51950
rect 27022 51874 27074 51886
rect 27134 51938 27186 51950
rect 27134 51874 27186 51886
rect 32958 51938 33010 51950
rect 32958 51874 33010 51886
rect 57150 51938 57202 51950
rect 57150 51874 57202 51886
rect 96910 51938 96962 51950
rect 96910 51874 96962 51886
rect 1344 51770 98560 51804
rect 1344 51718 8896 51770
rect 8948 51718 9020 51770
rect 9072 51718 9144 51770
rect 9196 51718 9268 51770
rect 9320 51718 17896 51770
rect 17948 51718 18020 51770
rect 18072 51718 18144 51770
rect 18196 51718 18268 51770
rect 18320 51718 26896 51770
rect 26948 51718 27020 51770
rect 27072 51718 27144 51770
rect 27196 51718 27268 51770
rect 27320 51718 35896 51770
rect 35948 51718 36020 51770
rect 36072 51718 36144 51770
rect 36196 51718 36268 51770
rect 36320 51718 44896 51770
rect 44948 51718 45020 51770
rect 45072 51718 45144 51770
rect 45196 51718 45268 51770
rect 45320 51718 53896 51770
rect 53948 51718 54020 51770
rect 54072 51718 54144 51770
rect 54196 51718 54268 51770
rect 54320 51718 62896 51770
rect 62948 51718 63020 51770
rect 63072 51718 63144 51770
rect 63196 51718 63268 51770
rect 63320 51718 71896 51770
rect 71948 51718 72020 51770
rect 72072 51718 72144 51770
rect 72196 51718 72268 51770
rect 72320 51718 80896 51770
rect 80948 51718 81020 51770
rect 81072 51718 81144 51770
rect 81196 51718 81268 51770
rect 81320 51718 89896 51770
rect 89948 51718 90020 51770
rect 90072 51718 90144 51770
rect 90196 51718 90268 51770
rect 90320 51718 98560 51770
rect 1344 51684 98560 51718
rect 28814 51602 28866 51614
rect 42702 51602 42754 51614
rect 37986 51550 37998 51602
rect 38050 51550 38062 51602
rect 28814 51538 28866 51550
rect 42702 51538 42754 51550
rect 43262 51602 43314 51614
rect 43262 51538 43314 51550
rect 43710 51602 43762 51614
rect 43710 51538 43762 51550
rect 44718 51602 44770 51614
rect 44718 51538 44770 51550
rect 47854 51602 47906 51614
rect 47854 51538 47906 51550
rect 50430 51602 50482 51614
rect 50430 51538 50482 51550
rect 55806 51602 55858 51614
rect 55806 51538 55858 51550
rect 57710 51602 57762 51614
rect 57710 51538 57762 51550
rect 62078 51602 62130 51614
rect 62078 51538 62130 51550
rect 90974 51602 91026 51614
rect 90974 51538 91026 51550
rect 2046 51490 2098 51502
rect 2046 51426 2098 51438
rect 11902 51490 11954 51502
rect 40910 51490 40962 51502
rect 38658 51438 38670 51490
rect 38722 51438 38734 51490
rect 11902 51426 11954 51438
rect 40910 51426 40962 51438
rect 41022 51490 41074 51502
rect 41022 51426 41074 51438
rect 41694 51490 41746 51502
rect 41694 51426 41746 51438
rect 47070 51490 47122 51502
rect 47070 51426 47122 51438
rect 70590 51490 70642 51502
rect 70590 51426 70642 51438
rect 71038 51490 71090 51502
rect 71038 51426 71090 51438
rect 71374 51490 71426 51502
rect 71374 51426 71426 51438
rect 77086 51490 77138 51502
rect 77086 51426 77138 51438
rect 1710 51378 1762 51390
rect 41246 51378 41298 51390
rect 38434 51326 38446 51378
rect 38498 51326 38510 51378
rect 39218 51326 39230 51378
rect 39282 51326 39294 51378
rect 39666 51326 39678 51378
rect 39730 51326 39742 51378
rect 1710 51314 1762 51326
rect 41246 51314 41298 51326
rect 41470 51378 41522 51390
rect 41470 51314 41522 51326
rect 42030 51378 42082 51390
rect 42030 51314 42082 51326
rect 42254 51378 42306 51390
rect 46174 51378 46226 51390
rect 44258 51326 44270 51378
rect 44322 51326 44334 51378
rect 42254 51314 42306 51326
rect 46174 51314 46226 51326
rect 46398 51378 46450 51390
rect 47406 51378 47458 51390
rect 62190 51378 62242 51390
rect 46722 51326 46734 51378
rect 46786 51326 46798 51378
rect 49970 51326 49982 51378
rect 50034 51326 50046 51378
rect 90738 51326 90750 51378
rect 90802 51326 90814 51378
rect 46398 51314 46450 51326
rect 47406 51314 47458 51326
rect 62190 51314 62242 51326
rect 2494 51266 2546 51278
rect 2494 51202 2546 51214
rect 39790 51266 39842 51278
rect 39790 51202 39842 51214
rect 40350 51266 40402 51278
rect 40350 51202 40402 51214
rect 42814 51266 42866 51278
rect 42814 51202 42866 51214
rect 55470 51266 55522 51278
rect 55470 51202 55522 51214
rect 55694 51266 55746 51278
rect 55694 51202 55746 51214
rect 57150 51266 57202 51278
rect 57150 51202 57202 51214
rect 61742 51266 61794 51278
rect 61742 51202 61794 51214
rect 76638 51266 76690 51278
rect 76638 51202 76690 51214
rect 41582 51154 41634 51166
rect 57138 51102 57150 51154
rect 57202 51151 57214 51154
rect 57474 51151 57486 51154
rect 57202 51105 57486 51151
rect 57202 51102 57214 51105
rect 57474 51102 57486 51105
rect 57538 51102 57550 51154
rect 41582 51090 41634 51102
rect 1344 50986 98560 51020
rect 1344 50934 4396 50986
rect 4448 50934 4520 50986
rect 4572 50934 4644 50986
rect 4696 50934 4768 50986
rect 4820 50934 13396 50986
rect 13448 50934 13520 50986
rect 13572 50934 13644 50986
rect 13696 50934 13768 50986
rect 13820 50934 22396 50986
rect 22448 50934 22520 50986
rect 22572 50934 22644 50986
rect 22696 50934 22768 50986
rect 22820 50934 31396 50986
rect 31448 50934 31520 50986
rect 31572 50934 31644 50986
rect 31696 50934 31768 50986
rect 31820 50934 40396 50986
rect 40448 50934 40520 50986
rect 40572 50934 40644 50986
rect 40696 50934 40768 50986
rect 40820 50934 49396 50986
rect 49448 50934 49520 50986
rect 49572 50934 49644 50986
rect 49696 50934 49768 50986
rect 49820 50934 58396 50986
rect 58448 50934 58520 50986
rect 58572 50934 58644 50986
rect 58696 50934 58768 50986
rect 58820 50934 67396 50986
rect 67448 50934 67520 50986
rect 67572 50934 67644 50986
rect 67696 50934 67768 50986
rect 67820 50934 76396 50986
rect 76448 50934 76520 50986
rect 76572 50934 76644 50986
rect 76696 50934 76768 50986
rect 76820 50934 85396 50986
rect 85448 50934 85520 50986
rect 85572 50934 85644 50986
rect 85696 50934 85768 50986
rect 85820 50934 94396 50986
rect 94448 50934 94520 50986
rect 94572 50934 94644 50986
rect 94696 50934 94768 50986
rect 94820 50934 98560 50986
rect 1344 50900 98560 50934
rect 27918 50818 27970 50830
rect 27918 50754 27970 50766
rect 29374 50818 29426 50830
rect 29374 50754 29426 50766
rect 32398 50818 32450 50830
rect 32398 50754 32450 50766
rect 44270 50818 44322 50830
rect 44270 50754 44322 50766
rect 49870 50818 49922 50830
rect 49870 50754 49922 50766
rect 38558 50706 38610 50718
rect 38558 50642 38610 50654
rect 39118 50706 39170 50718
rect 39118 50642 39170 50654
rect 39566 50706 39618 50718
rect 39566 50642 39618 50654
rect 55246 50706 55298 50718
rect 58606 50706 58658 50718
rect 57362 50654 57374 50706
rect 57426 50654 57438 50706
rect 55246 50642 55298 50654
rect 58606 50642 58658 50654
rect 74286 50706 74338 50718
rect 74286 50642 74338 50654
rect 16718 50594 16770 50606
rect 29934 50594 29986 50606
rect 17266 50542 17278 50594
rect 17330 50542 17342 50594
rect 16718 50530 16770 50542
rect 29934 50530 29986 50542
rect 39902 50594 39954 50606
rect 39902 50530 39954 50542
rect 40798 50594 40850 50606
rect 45502 50594 45554 50606
rect 41234 50542 41246 50594
rect 41298 50542 41310 50594
rect 40798 50530 40850 50542
rect 45502 50530 45554 50542
rect 46174 50594 46226 50606
rect 60398 50594 60450 50606
rect 70478 50594 70530 50606
rect 76974 50594 77026 50606
rect 46834 50542 46846 50594
rect 46898 50542 46910 50594
rect 58034 50542 58046 50594
rect 58098 50542 58110 50594
rect 60946 50542 60958 50594
rect 61010 50542 61022 50594
rect 70914 50542 70926 50594
rect 70978 50542 70990 50594
rect 76290 50542 76302 50594
rect 76354 50542 76366 50594
rect 77298 50542 77310 50594
rect 77362 50542 77374 50594
rect 46174 50530 46226 50542
rect 60398 50530 60450 50542
rect 70478 50530 70530 50542
rect 76974 50530 77026 50542
rect 1710 50482 1762 50494
rect 1710 50418 1762 50430
rect 2046 50482 2098 50494
rect 2046 50418 2098 50430
rect 2494 50482 2546 50494
rect 2494 50418 2546 50430
rect 16158 50482 16210 50494
rect 16158 50418 16210 50430
rect 19630 50482 19682 50494
rect 19630 50418 19682 50430
rect 20862 50482 20914 50494
rect 20862 50418 20914 50430
rect 28030 50482 28082 50494
rect 28030 50418 28082 50430
rect 29486 50482 29538 50494
rect 29486 50418 29538 50430
rect 32286 50482 32338 50494
rect 32286 50418 32338 50430
rect 32846 50482 32898 50494
rect 32846 50418 32898 50430
rect 40462 50482 40514 50494
rect 40462 50418 40514 50430
rect 46062 50482 46114 50494
rect 46062 50418 46114 50430
rect 49086 50482 49138 50494
rect 49086 50418 49138 50430
rect 63310 50482 63362 50494
rect 63310 50418 63362 50430
rect 64094 50482 64146 50494
rect 64094 50418 64146 50430
rect 64542 50482 64594 50494
rect 64542 50418 64594 50430
rect 73166 50482 73218 50494
rect 73166 50418 73218 50430
rect 73950 50482 74002 50494
rect 73950 50418 74002 50430
rect 76526 50482 76578 50494
rect 76526 50418 76578 50430
rect 79662 50482 79714 50494
rect 79662 50418 79714 50430
rect 80446 50482 80498 50494
rect 80446 50418 80498 50430
rect 96238 50482 96290 50494
rect 96238 50418 96290 50430
rect 96574 50482 96626 50494
rect 96574 50418 96626 50430
rect 5630 50370 5682 50382
rect 5630 50306 5682 50318
rect 16494 50370 16546 50382
rect 16494 50306 16546 50318
rect 20414 50370 20466 50382
rect 20414 50306 20466 50318
rect 28478 50370 28530 50382
rect 59950 50370 60002 50382
rect 43586 50318 43598 50370
rect 43650 50318 43662 50370
rect 28478 50306 28530 50318
rect 59950 50306 60002 50318
rect 65550 50370 65602 50382
rect 65550 50306 65602 50318
rect 86830 50370 86882 50382
rect 86830 50306 86882 50318
rect 1344 50202 98560 50236
rect 1344 50150 8896 50202
rect 8948 50150 9020 50202
rect 9072 50150 9144 50202
rect 9196 50150 9268 50202
rect 9320 50150 17896 50202
rect 17948 50150 18020 50202
rect 18072 50150 18144 50202
rect 18196 50150 18268 50202
rect 18320 50150 26896 50202
rect 26948 50150 27020 50202
rect 27072 50150 27144 50202
rect 27196 50150 27268 50202
rect 27320 50150 35896 50202
rect 35948 50150 36020 50202
rect 36072 50150 36144 50202
rect 36196 50150 36268 50202
rect 36320 50150 44896 50202
rect 44948 50150 45020 50202
rect 45072 50150 45144 50202
rect 45196 50150 45268 50202
rect 45320 50150 53896 50202
rect 53948 50150 54020 50202
rect 54072 50150 54144 50202
rect 54196 50150 54268 50202
rect 54320 50150 62896 50202
rect 62948 50150 63020 50202
rect 63072 50150 63144 50202
rect 63196 50150 63268 50202
rect 63320 50150 71896 50202
rect 71948 50150 72020 50202
rect 72072 50150 72144 50202
rect 72196 50150 72268 50202
rect 72320 50150 80896 50202
rect 80948 50150 81020 50202
rect 81072 50150 81144 50202
rect 81196 50150 81268 50202
rect 81320 50150 89896 50202
rect 89948 50150 90020 50202
rect 90072 50150 90144 50202
rect 90196 50150 90268 50202
rect 90320 50150 98560 50202
rect 1344 50116 98560 50150
rect 40350 50034 40402 50046
rect 8306 49982 8318 50034
rect 8370 49982 8382 50034
rect 40350 49970 40402 49982
rect 60958 50034 61010 50046
rect 69246 50034 69298 50046
rect 68114 49982 68126 50034
rect 68178 49982 68190 50034
rect 60958 49970 61010 49982
rect 69246 49970 69298 49982
rect 72382 50034 72434 50046
rect 72382 49970 72434 49982
rect 75742 50034 75794 50046
rect 75742 49970 75794 49982
rect 76862 50034 76914 50046
rect 76862 49970 76914 49982
rect 1934 49922 1986 49934
rect 1934 49858 1986 49870
rect 9550 49922 9602 49934
rect 9550 49858 9602 49870
rect 10110 49922 10162 49934
rect 10110 49858 10162 49870
rect 11342 49922 11394 49934
rect 11342 49858 11394 49870
rect 14478 49922 14530 49934
rect 64990 49922 65042 49934
rect 86270 49922 86322 49934
rect 26226 49870 26238 49922
rect 26290 49870 26302 49922
rect 29698 49870 29710 49922
rect 29762 49870 29774 49922
rect 37650 49870 37662 49922
rect 37714 49870 37726 49922
rect 51538 49870 51550 49922
rect 51602 49870 51614 49922
rect 62290 49870 62302 49922
rect 62354 49870 62366 49922
rect 62850 49870 62862 49922
rect 62914 49870 62926 49922
rect 72930 49870 72942 49922
rect 72994 49870 73006 49922
rect 73490 49870 73502 49922
rect 73554 49870 73566 49922
rect 77410 49870 77422 49922
rect 77474 49870 77486 49922
rect 77746 49870 77758 49922
rect 77810 49870 77822 49922
rect 14478 49858 14530 49870
rect 64990 49858 65042 49870
rect 86270 49858 86322 49870
rect 5518 49810 5570 49822
rect 42366 49810 42418 49822
rect 5842 49758 5854 49810
rect 5906 49758 5918 49810
rect 11666 49758 11678 49810
rect 11730 49758 11742 49810
rect 12114 49758 12126 49810
rect 12178 49758 12190 49810
rect 25554 49758 25566 49810
rect 25618 49758 25630 49810
rect 29026 49758 29038 49810
rect 29090 49758 29102 49810
rect 38434 49758 38446 49810
rect 38498 49758 38510 49810
rect 5518 49746 5570 49758
rect 42366 49746 42418 49758
rect 50430 49810 50482 49822
rect 61294 49810 61346 49822
rect 50754 49758 50766 49810
rect 50818 49758 50830 49810
rect 50430 49746 50482 49758
rect 61294 49746 61346 49758
rect 61742 49810 61794 49822
rect 65438 49810 65490 49822
rect 77198 49810 77250 49822
rect 64754 49758 64766 49810
rect 64818 49758 64830 49810
rect 65762 49758 65774 49810
rect 65826 49758 65838 49810
rect 86034 49758 86046 49810
rect 86098 49758 86110 49810
rect 96898 49758 96910 49810
rect 96962 49758 96974 49810
rect 61742 49746 61794 49758
rect 65438 49746 65490 49758
rect 77198 49746 77250 49758
rect 2494 49698 2546 49710
rect 32510 49698 32562 49710
rect 28466 49646 28478 49698
rect 28530 49646 28542 49698
rect 31938 49646 31950 49698
rect 32002 49646 32014 49698
rect 2494 49634 2546 49646
rect 32510 49634 32562 49646
rect 35534 49698 35586 49710
rect 35534 49634 35586 49646
rect 39006 49698 39058 49710
rect 60622 49698 60674 49710
rect 53778 49646 53790 49698
rect 53842 49646 53854 49698
rect 39006 49634 39058 49646
rect 60622 49634 60674 49646
rect 71262 49698 71314 49710
rect 71262 49634 71314 49646
rect 71710 49698 71762 49710
rect 71710 49634 71762 49646
rect 76190 49698 76242 49710
rect 76190 49634 76242 49646
rect 92430 49698 92482 49710
rect 98018 49646 98030 49698
rect 98082 49646 98094 49698
rect 92430 49634 92482 49646
rect 8990 49586 9042 49598
rect 8990 49522 9042 49534
rect 15262 49586 15314 49598
rect 15262 49522 15314 49534
rect 62078 49586 62130 49598
rect 62078 49522 62130 49534
rect 68910 49586 68962 49598
rect 68910 49522 68962 49534
rect 72718 49586 72770 49598
rect 72718 49522 72770 49534
rect 1344 49418 98560 49452
rect 1344 49366 4396 49418
rect 4448 49366 4520 49418
rect 4572 49366 4644 49418
rect 4696 49366 4768 49418
rect 4820 49366 13396 49418
rect 13448 49366 13520 49418
rect 13572 49366 13644 49418
rect 13696 49366 13768 49418
rect 13820 49366 22396 49418
rect 22448 49366 22520 49418
rect 22572 49366 22644 49418
rect 22696 49366 22768 49418
rect 22820 49366 31396 49418
rect 31448 49366 31520 49418
rect 31572 49366 31644 49418
rect 31696 49366 31768 49418
rect 31820 49366 40396 49418
rect 40448 49366 40520 49418
rect 40572 49366 40644 49418
rect 40696 49366 40768 49418
rect 40820 49366 49396 49418
rect 49448 49366 49520 49418
rect 49572 49366 49644 49418
rect 49696 49366 49768 49418
rect 49820 49366 58396 49418
rect 58448 49366 58520 49418
rect 58572 49366 58644 49418
rect 58696 49366 58768 49418
rect 58820 49366 67396 49418
rect 67448 49366 67520 49418
rect 67572 49366 67644 49418
rect 67696 49366 67768 49418
rect 67820 49366 76396 49418
rect 76448 49366 76520 49418
rect 76572 49366 76644 49418
rect 76696 49366 76768 49418
rect 76820 49366 85396 49418
rect 85448 49366 85520 49418
rect 85572 49366 85644 49418
rect 85696 49366 85768 49418
rect 85820 49366 94396 49418
rect 94448 49366 94520 49418
rect 94572 49366 94644 49418
rect 94696 49366 94768 49418
rect 94820 49366 98560 49418
rect 1344 49332 98560 49366
rect 64766 49250 64818 49262
rect 64766 49186 64818 49198
rect 86158 49250 86210 49262
rect 86158 49186 86210 49198
rect 29262 49138 29314 49150
rect 35086 49138 35138 49150
rect 32946 49086 32958 49138
rect 33010 49086 33022 49138
rect 29262 49074 29314 49086
rect 35086 49074 35138 49086
rect 35758 49138 35810 49150
rect 35758 49074 35810 49086
rect 61294 49138 61346 49150
rect 61294 49074 61346 49086
rect 63646 49138 63698 49150
rect 63646 49074 63698 49086
rect 77646 49138 77698 49150
rect 77646 49074 77698 49086
rect 79774 49138 79826 49150
rect 79774 49074 79826 49086
rect 90526 49138 90578 49150
rect 90526 49074 90578 49086
rect 8990 49026 9042 49038
rect 65102 49026 65154 49038
rect 9314 48974 9326 49026
rect 9378 48974 9390 49026
rect 32274 48974 32286 49026
rect 32338 48974 32350 49026
rect 8990 48962 9042 48974
rect 65102 48962 65154 48974
rect 72158 49026 72210 49038
rect 85822 49026 85874 49038
rect 85138 48974 85150 49026
rect 85202 48974 85214 49026
rect 72158 48962 72210 48974
rect 85822 48962 85874 48974
rect 86718 49026 86770 49038
rect 90190 49026 90242 49038
rect 87042 48974 87054 49026
rect 87106 48974 87118 49026
rect 86718 48962 86770 48974
rect 90190 48962 90242 48974
rect 92542 49026 92594 49038
rect 93090 48974 93102 49026
rect 93154 48974 93166 49026
rect 92542 48962 92594 48974
rect 1710 48914 1762 48926
rect 1710 48850 1762 48862
rect 2382 48914 2434 48926
rect 2382 48850 2434 48862
rect 3166 48914 3218 48926
rect 3166 48850 3218 48862
rect 64206 48914 64258 48926
rect 71822 48914 71874 48926
rect 92318 48914 92370 48926
rect 65314 48862 65326 48914
rect 65378 48862 65390 48914
rect 65874 48862 65886 48914
rect 65938 48862 65950 48914
rect 85026 48862 85038 48914
rect 85090 48862 85102 48914
rect 64206 48850 64258 48862
rect 71822 48850 71874 48862
rect 92318 48850 92370 48862
rect 95454 48914 95506 48926
rect 95454 48850 95506 48862
rect 2046 48802 2098 48814
rect 2046 48738 2098 48750
rect 2718 48802 2770 48814
rect 12462 48802 12514 48814
rect 11666 48750 11678 48802
rect 11730 48750 11742 48802
rect 2718 48738 2770 48750
rect 12462 48738 12514 48750
rect 14478 48802 14530 48814
rect 14478 48738 14530 48750
rect 20750 48802 20802 48814
rect 20750 48738 20802 48750
rect 55022 48802 55074 48814
rect 55022 48738 55074 48750
rect 56366 48802 56418 48814
rect 56366 48738 56418 48750
rect 73502 48802 73554 48814
rect 73502 48738 73554 48750
rect 73950 48802 74002 48814
rect 73950 48738 74002 48750
rect 80222 48802 80274 48814
rect 80222 48738 80274 48750
rect 84702 48802 84754 48814
rect 96238 48802 96290 48814
rect 89618 48750 89630 48802
rect 89682 48750 89694 48802
rect 84702 48738 84754 48750
rect 96238 48738 96290 48750
rect 1344 48634 98560 48668
rect 1344 48582 8896 48634
rect 8948 48582 9020 48634
rect 9072 48582 9144 48634
rect 9196 48582 9268 48634
rect 9320 48582 17896 48634
rect 17948 48582 18020 48634
rect 18072 48582 18144 48634
rect 18196 48582 18268 48634
rect 18320 48582 26896 48634
rect 26948 48582 27020 48634
rect 27072 48582 27144 48634
rect 27196 48582 27268 48634
rect 27320 48582 35896 48634
rect 35948 48582 36020 48634
rect 36072 48582 36144 48634
rect 36196 48582 36268 48634
rect 36320 48582 44896 48634
rect 44948 48582 45020 48634
rect 45072 48582 45144 48634
rect 45196 48582 45268 48634
rect 45320 48582 53896 48634
rect 53948 48582 54020 48634
rect 54072 48582 54144 48634
rect 54196 48582 54268 48634
rect 54320 48582 62896 48634
rect 62948 48582 63020 48634
rect 63072 48582 63144 48634
rect 63196 48582 63268 48634
rect 63320 48582 71896 48634
rect 71948 48582 72020 48634
rect 72072 48582 72144 48634
rect 72196 48582 72268 48634
rect 72320 48582 80896 48634
rect 80948 48582 81020 48634
rect 81072 48582 81144 48634
rect 81196 48582 81268 48634
rect 81320 48582 89896 48634
rect 89948 48582 90020 48634
rect 90072 48582 90144 48634
rect 90196 48582 90268 48634
rect 90320 48582 98560 48634
rect 1344 48548 98560 48582
rect 41022 48466 41074 48478
rect 53230 48466 53282 48478
rect 4722 48414 4734 48466
rect 4786 48414 4798 48466
rect 39890 48414 39902 48466
rect 39954 48414 39966 48466
rect 52322 48414 52334 48466
rect 52386 48414 52398 48466
rect 41022 48402 41074 48414
rect 53230 48402 53282 48414
rect 63870 48466 63922 48478
rect 63870 48402 63922 48414
rect 65326 48466 65378 48478
rect 96574 48466 96626 48478
rect 83122 48414 83134 48466
rect 83186 48414 83198 48466
rect 65326 48402 65378 48414
rect 96574 48402 96626 48414
rect 13582 48354 13634 48366
rect 13582 48290 13634 48302
rect 14254 48354 14306 48366
rect 19854 48354 19906 48366
rect 43486 48354 43538 48366
rect 14914 48302 14926 48354
rect 14978 48302 14990 48354
rect 20402 48302 20414 48354
rect 20466 48302 20478 48354
rect 14254 48290 14306 48302
rect 19854 48290 19906 48302
rect 43486 48290 43538 48302
rect 43934 48354 43986 48366
rect 43934 48290 43986 48302
rect 48974 48354 49026 48366
rect 48974 48290 49026 48302
rect 55694 48354 55746 48366
rect 64542 48354 64594 48366
rect 57362 48302 57374 48354
rect 57426 48302 57438 48354
rect 57810 48302 57822 48354
rect 57874 48302 57886 48354
rect 55694 48290 55746 48302
rect 64542 48290 64594 48302
rect 64878 48354 64930 48366
rect 64878 48290 64930 48302
rect 65102 48354 65154 48366
rect 65102 48290 65154 48302
rect 71038 48354 71090 48366
rect 71038 48290 71090 48302
rect 71374 48354 71426 48366
rect 73950 48354 74002 48366
rect 72930 48302 72942 48354
rect 72994 48302 73006 48354
rect 73490 48302 73502 48354
rect 73554 48302 73566 48354
rect 71374 48290 71426 48302
rect 73950 48290 74002 48302
rect 74174 48354 74226 48366
rect 74174 48290 74226 48302
rect 77198 48354 77250 48366
rect 77198 48290 77250 48302
rect 77646 48354 77698 48366
rect 83694 48354 83746 48366
rect 78306 48302 78318 48354
rect 78370 48302 78382 48354
rect 92530 48302 92542 48354
rect 92594 48302 92606 48354
rect 77646 48290 77698 48302
rect 83694 48290 83746 48302
rect 1822 48242 1874 48254
rect 15822 48242 15874 48254
rect 36766 48242 36818 48254
rect 44270 48242 44322 48254
rect 2146 48190 2158 48242
rect 2210 48190 2222 48242
rect 14018 48190 14030 48242
rect 14082 48190 14094 48242
rect 15026 48190 15038 48242
rect 15090 48190 15102 48242
rect 20290 48190 20302 48242
rect 20354 48190 20366 48242
rect 37314 48190 37326 48242
rect 37378 48190 37390 48242
rect 1822 48178 1874 48190
rect 15822 48178 15874 48190
rect 36766 48178 36818 48190
rect 44270 48178 44322 48190
rect 49198 48242 49250 48254
rect 56030 48242 56082 48254
rect 49858 48190 49870 48242
rect 49922 48190 49934 48242
rect 49198 48178 49250 48190
rect 56030 48178 56082 48190
rect 56702 48242 56754 48254
rect 71710 48242 71762 48254
rect 65538 48190 65550 48242
rect 65602 48190 65614 48242
rect 56702 48178 56754 48190
rect 71710 48178 71762 48190
rect 72382 48242 72434 48254
rect 72382 48178 72434 48190
rect 72718 48242 72770 48254
rect 72718 48178 72770 48190
rect 74398 48242 74450 48254
rect 76414 48242 76466 48254
rect 77422 48242 77474 48254
rect 78878 48242 78930 48254
rect 74610 48190 74622 48242
rect 74674 48190 74686 48242
rect 76962 48190 76974 48242
rect 77026 48190 77038 48242
rect 78082 48190 78094 48242
rect 78146 48190 78158 48242
rect 74398 48178 74450 48190
rect 76414 48178 76466 48190
rect 77422 48178 77474 48190
rect 78878 48178 78930 48190
rect 80222 48242 80274 48254
rect 91198 48242 91250 48254
rect 93102 48242 93154 48254
rect 80546 48190 80558 48242
rect 80610 48190 80622 48242
rect 92306 48190 92318 48242
rect 92370 48190 92382 48242
rect 80222 48178 80274 48190
rect 91198 48178 91250 48190
rect 93102 48178 93154 48190
rect 96238 48242 96290 48254
rect 96898 48190 96910 48242
rect 96962 48190 96974 48242
rect 96238 48178 96290 48190
rect 5630 48130 5682 48142
rect 5630 48066 5682 48078
rect 16494 48130 16546 48142
rect 16494 48066 16546 48078
rect 21086 48130 21138 48142
rect 21086 48066 21138 48078
rect 22094 48130 22146 48142
rect 22094 48066 22146 48078
rect 46398 48130 46450 48142
rect 46398 48066 46450 48078
rect 58382 48130 58434 48142
rect 58382 48066 58434 48078
rect 65214 48130 65266 48142
rect 65214 48066 65266 48078
rect 74286 48130 74338 48142
rect 74286 48066 74338 48078
rect 75966 48130 76018 48142
rect 75966 48066 76018 48078
rect 77310 48130 77362 48142
rect 77310 48066 77362 48078
rect 91646 48130 91698 48142
rect 98018 48078 98030 48130
rect 98082 48078 98094 48130
rect 91646 48066 91698 48078
rect 5294 48018 5346 48030
rect 5294 47954 5346 47966
rect 15486 48018 15538 48030
rect 15486 47954 15538 47966
rect 21422 48018 21474 48030
rect 21422 47954 21474 47966
rect 40462 48018 40514 48030
rect 40462 47954 40514 47966
rect 52894 48018 52946 48030
rect 52894 47954 52946 47966
rect 57038 48018 57090 48030
rect 57038 47954 57090 47966
rect 79214 48018 79266 48030
rect 79214 47954 79266 47966
rect 93438 48018 93490 48030
rect 93438 47954 93490 47966
rect 1344 47850 98560 47884
rect 1344 47798 4396 47850
rect 4448 47798 4520 47850
rect 4572 47798 4644 47850
rect 4696 47798 4768 47850
rect 4820 47798 13396 47850
rect 13448 47798 13520 47850
rect 13572 47798 13644 47850
rect 13696 47798 13768 47850
rect 13820 47798 22396 47850
rect 22448 47798 22520 47850
rect 22572 47798 22644 47850
rect 22696 47798 22768 47850
rect 22820 47798 31396 47850
rect 31448 47798 31520 47850
rect 31572 47798 31644 47850
rect 31696 47798 31768 47850
rect 31820 47798 40396 47850
rect 40448 47798 40520 47850
rect 40572 47798 40644 47850
rect 40696 47798 40768 47850
rect 40820 47798 49396 47850
rect 49448 47798 49520 47850
rect 49572 47798 49644 47850
rect 49696 47798 49768 47850
rect 49820 47798 58396 47850
rect 58448 47798 58520 47850
rect 58572 47798 58644 47850
rect 58696 47798 58768 47850
rect 58820 47798 67396 47850
rect 67448 47798 67520 47850
rect 67572 47798 67644 47850
rect 67696 47798 67768 47850
rect 67820 47798 76396 47850
rect 76448 47798 76520 47850
rect 76572 47798 76644 47850
rect 76696 47798 76768 47850
rect 76820 47798 85396 47850
rect 85448 47798 85520 47850
rect 85572 47798 85644 47850
rect 85696 47798 85768 47850
rect 85820 47798 94396 47850
rect 94448 47798 94520 47850
rect 94572 47798 94644 47850
rect 94696 47798 94768 47850
rect 94820 47798 98560 47850
rect 1344 47764 98560 47798
rect 44942 47682 44994 47694
rect 44942 47618 44994 47630
rect 74622 47682 74674 47694
rect 74622 47618 74674 47630
rect 35758 47570 35810 47582
rect 48750 47570 48802 47582
rect 38658 47518 38670 47570
rect 38722 47518 38734 47570
rect 35758 47506 35810 47518
rect 48750 47506 48802 47518
rect 54462 47570 54514 47582
rect 54462 47506 54514 47518
rect 74958 47570 75010 47582
rect 74958 47506 75010 47518
rect 77422 47570 77474 47582
rect 77422 47506 77474 47518
rect 10446 47458 10498 47470
rect 1810 47406 1822 47458
rect 1874 47406 1886 47458
rect 10446 47394 10498 47406
rect 14142 47458 14194 47470
rect 21198 47458 21250 47470
rect 33966 47458 34018 47470
rect 45278 47458 45330 47470
rect 49198 47458 49250 47470
rect 14690 47406 14702 47458
rect 14754 47406 14766 47458
rect 20514 47406 20526 47458
rect 20578 47406 20590 47458
rect 21746 47406 21758 47458
rect 21810 47406 21822 47458
rect 34626 47406 34638 47458
rect 34690 47406 34702 47458
rect 43250 47406 43262 47458
rect 43314 47406 43326 47458
rect 45938 47406 45950 47458
rect 46002 47406 46014 47458
rect 47394 47406 47406 47458
rect 47458 47406 47470 47458
rect 47730 47406 47742 47458
rect 47794 47406 47806 47458
rect 14142 47394 14194 47406
rect 21198 47394 21250 47406
rect 33966 47394 34018 47406
rect 45278 47394 45330 47406
rect 49198 47394 49250 47406
rect 54910 47458 54962 47470
rect 79214 47458 79266 47470
rect 55346 47406 55358 47458
rect 55410 47406 55422 47458
rect 71026 47406 71038 47458
rect 71090 47406 71102 47458
rect 71474 47406 71486 47458
rect 71538 47406 71550 47458
rect 92642 47406 92654 47458
rect 92706 47406 92718 47458
rect 54910 47394 54962 47406
rect 79214 47394 79266 47406
rect 2046 47346 2098 47358
rect 11342 47346 11394 47358
rect 9650 47294 9662 47346
rect 9714 47294 9726 47346
rect 10210 47294 10222 47346
rect 10274 47294 10286 47346
rect 2046 47282 2098 47294
rect 11342 47282 11394 47294
rect 20750 47346 20802 47358
rect 36430 47346 36482 47358
rect 34738 47294 34750 47346
rect 34802 47294 34814 47346
rect 20750 47282 20802 47294
rect 36430 47282 36482 47294
rect 37326 47346 37378 47358
rect 37326 47282 37378 47294
rect 37662 47346 37714 47358
rect 50542 47346 50594 47358
rect 46050 47294 46062 47346
rect 46114 47294 46126 47346
rect 46946 47294 46958 47346
rect 47010 47294 47022 47346
rect 37662 47282 37714 47294
rect 50542 47282 50594 47294
rect 50878 47346 50930 47358
rect 50878 47282 50930 47294
rect 57598 47346 57650 47358
rect 57598 47282 57650 47294
rect 79550 47346 79602 47358
rect 79550 47282 79602 47294
rect 86718 47346 86770 47358
rect 86718 47282 86770 47294
rect 87054 47346 87106 47358
rect 87054 47282 87106 47294
rect 92878 47346 92930 47358
rect 92878 47282 92930 47294
rect 2606 47234 2658 47246
rect 2606 47170 2658 47182
rect 9102 47234 9154 47246
rect 9102 47170 9154 47182
rect 10782 47234 10834 47246
rect 10782 47170 10834 47182
rect 11790 47234 11842 47246
rect 17838 47234 17890 47246
rect 17266 47182 17278 47234
rect 17330 47182 17342 47234
rect 11790 47170 11842 47182
rect 17838 47170 17890 47182
rect 18174 47234 18226 47246
rect 24894 47234 24946 47246
rect 24098 47182 24110 47234
rect 24162 47182 24174 47234
rect 18174 47170 18226 47182
rect 24894 47170 24946 47182
rect 31166 47234 31218 47246
rect 31166 47170 31218 47182
rect 33630 47234 33682 47246
rect 33630 47170 33682 47182
rect 35310 47234 35362 47246
rect 35310 47170 35362 47182
rect 43710 47234 43762 47246
rect 43710 47170 43762 47182
rect 44270 47234 44322 47246
rect 58382 47234 58434 47246
rect 47954 47182 47966 47234
rect 48018 47182 48030 47234
rect 48178 47182 48190 47234
rect 48242 47182 48254 47234
rect 44270 47170 44322 47182
rect 58382 47170 58434 47182
rect 60734 47234 60786 47246
rect 86382 47234 86434 47246
rect 74050 47182 74062 47234
rect 74114 47182 74126 47234
rect 60734 47170 60786 47182
rect 86382 47170 86434 47182
rect 1344 47066 98560 47100
rect 1344 47014 8896 47066
rect 8948 47014 9020 47066
rect 9072 47014 9144 47066
rect 9196 47014 9268 47066
rect 9320 47014 17896 47066
rect 17948 47014 18020 47066
rect 18072 47014 18144 47066
rect 18196 47014 18268 47066
rect 18320 47014 26896 47066
rect 26948 47014 27020 47066
rect 27072 47014 27144 47066
rect 27196 47014 27268 47066
rect 27320 47014 35896 47066
rect 35948 47014 36020 47066
rect 36072 47014 36144 47066
rect 36196 47014 36268 47066
rect 36320 47014 44896 47066
rect 44948 47014 45020 47066
rect 45072 47014 45144 47066
rect 45196 47014 45268 47066
rect 45320 47014 53896 47066
rect 53948 47014 54020 47066
rect 54072 47014 54144 47066
rect 54196 47014 54268 47066
rect 54320 47014 62896 47066
rect 62948 47014 63020 47066
rect 63072 47014 63144 47066
rect 63196 47014 63268 47066
rect 63320 47014 71896 47066
rect 71948 47014 72020 47066
rect 72072 47014 72144 47066
rect 72196 47014 72268 47066
rect 72320 47014 80896 47066
rect 80948 47014 81020 47066
rect 81072 47014 81144 47066
rect 81196 47014 81268 47066
rect 81320 47014 89896 47066
rect 89948 47014 90020 47066
rect 90072 47014 90144 47066
rect 90196 47014 90268 47066
rect 90320 47014 98560 47066
rect 1344 46980 98560 47014
rect 20974 46898 21026 46910
rect 31614 46898 31666 46910
rect 39118 46898 39170 46910
rect 5394 46846 5406 46898
rect 5458 46846 5470 46898
rect 28578 46846 28590 46898
rect 28642 46846 28654 46898
rect 38546 46846 38558 46898
rect 38610 46846 38622 46898
rect 20974 46834 21026 46846
rect 31614 46834 31666 46846
rect 39118 46834 39170 46846
rect 43038 46898 43090 46910
rect 43038 46834 43090 46846
rect 46958 46898 47010 46910
rect 46958 46834 47010 46846
rect 51438 46898 51490 46910
rect 51438 46834 51490 46846
rect 51886 46898 51938 46910
rect 51886 46834 51938 46846
rect 85038 46898 85090 46910
rect 85038 46834 85090 46846
rect 87278 46898 87330 46910
rect 87278 46834 87330 46846
rect 96574 46898 96626 46910
rect 96574 46834 96626 46846
rect 8654 46786 8706 46798
rect 8654 46722 8706 46734
rect 8990 46786 9042 46798
rect 8990 46722 9042 46734
rect 12350 46786 12402 46798
rect 32174 46786 32226 46798
rect 30370 46734 30382 46786
rect 30434 46734 30446 46786
rect 12350 46722 12402 46734
rect 32174 46722 32226 46734
rect 32510 46786 32562 46798
rect 46174 46786 46226 46798
rect 53566 46786 53618 46798
rect 61854 46786 61906 46798
rect 36754 46734 36766 46786
rect 36818 46734 36830 46786
rect 37874 46734 37886 46786
rect 37938 46734 37950 46786
rect 40002 46734 40014 46786
rect 40066 46734 40078 46786
rect 52434 46734 52446 46786
rect 52498 46734 52510 46786
rect 52994 46734 53006 46786
rect 53058 46734 53070 46786
rect 57250 46734 57262 46786
rect 57314 46734 57326 46786
rect 58370 46734 58382 46786
rect 58434 46734 58446 46786
rect 32510 46722 32562 46734
rect 46174 46722 46226 46734
rect 53566 46722 53618 46734
rect 61854 46722 61906 46734
rect 64990 46786 65042 46798
rect 67566 46786 67618 46798
rect 75294 46786 75346 46798
rect 78430 46786 78482 46798
rect 92206 46786 92258 46798
rect 65426 46734 65438 46786
rect 65490 46734 65502 46786
rect 73714 46734 73726 46786
rect 73778 46734 73790 46786
rect 76850 46734 76862 46786
rect 76914 46734 76926 46786
rect 86370 46734 86382 46786
rect 86434 46734 86446 46786
rect 86706 46734 86718 46786
rect 86770 46734 86782 46786
rect 64990 46722 65042 46734
rect 67566 46722 67618 46734
rect 75294 46722 75346 46734
rect 78430 46722 78482 46734
rect 92206 46722 92258 46734
rect 92542 46786 92594 46798
rect 92542 46722 92594 46734
rect 1822 46674 1874 46686
rect 1822 46610 1874 46622
rect 2494 46674 2546 46686
rect 25678 46674 25730 46686
rect 33294 46674 33346 46686
rect 43486 46674 43538 46686
rect 55246 46674 55298 46686
rect 62190 46674 62242 46686
rect 2818 46622 2830 46674
rect 2882 46622 2894 46674
rect 9538 46622 9550 46674
rect 9602 46622 9614 46674
rect 9986 46622 9998 46674
rect 10050 46622 10062 46674
rect 26114 46622 26126 46674
rect 26178 46622 26190 46674
rect 30594 46622 30606 46674
rect 30658 46622 30670 46674
rect 34738 46622 34750 46674
rect 34802 46622 34814 46674
rect 34962 46622 34974 46674
rect 35026 46622 35038 46674
rect 35634 46622 35646 46674
rect 35698 46622 35710 46674
rect 38210 46622 38222 46674
rect 38274 46622 38286 46674
rect 40226 46622 40238 46674
rect 40290 46622 40302 46674
rect 43922 46622 43934 46674
rect 43986 46622 43998 46674
rect 56578 46622 56590 46674
rect 56642 46622 56654 46674
rect 58482 46622 58494 46674
rect 58546 46622 58558 46674
rect 60050 46622 60062 46674
rect 60114 46622 60126 46674
rect 60386 46622 60398 46674
rect 60450 46622 60462 46674
rect 2494 46610 2546 46622
rect 25678 46610 25730 46622
rect 33294 46610 33346 46622
rect 43486 46610 43538 46622
rect 55246 46610 55298 46622
rect 62190 46610 62242 46622
rect 65214 46674 65266 46686
rect 91870 46674 91922 46686
rect 65762 46622 65774 46674
rect 65826 46622 65838 46674
rect 66434 46622 66446 46674
rect 66498 46622 66510 46674
rect 73938 46622 73950 46674
rect 74002 46622 74014 46674
rect 74498 46622 74510 46674
rect 74562 46622 74574 46674
rect 74946 46622 74958 46674
rect 75010 46622 75022 46674
rect 77074 46622 77086 46674
rect 77138 46622 77150 46674
rect 77634 46622 77646 46674
rect 77698 46622 77710 46674
rect 78082 46622 78094 46674
rect 78146 46622 78158 46674
rect 65214 46610 65266 46622
rect 91870 46610 91922 46622
rect 96238 46674 96290 46686
rect 96898 46622 96910 46674
rect 96962 46622 96974 46674
rect 96238 46610 96290 46622
rect 29150 46562 29202 46574
rect 29150 46498 29202 46510
rect 29822 46562 29874 46574
rect 29822 46498 29874 46510
rect 31166 46562 31218 46574
rect 31166 46498 31218 46510
rect 41022 46562 41074 46574
rect 41022 46498 41074 46510
rect 54238 46562 54290 46574
rect 54238 46498 54290 46510
rect 54686 46562 54738 46574
rect 54686 46498 54738 46510
rect 55582 46562 55634 46574
rect 55582 46498 55634 46510
rect 56030 46562 56082 46574
rect 56030 46498 56082 46510
rect 58270 46562 58322 46574
rect 58270 46498 58322 46510
rect 73390 46562 73442 46574
rect 73390 46498 73442 46510
rect 76638 46562 76690 46574
rect 76638 46498 76690 46510
rect 85486 46562 85538 46574
rect 98018 46510 98030 46562
rect 98082 46510 98094 46562
rect 85486 46498 85538 46510
rect 5966 46450 6018 46462
rect 5966 46386 6018 46398
rect 13134 46450 13186 46462
rect 13134 46386 13186 46398
rect 29486 46450 29538 46462
rect 29486 46386 29538 46398
rect 39454 46450 39506 46462
rect 39454 46386 39506 46398
rect 52222 46450 52274 46462
rect 66782 46450 66834 46462
rect 54226 46398 54238 46450
rect 54290 46447 54302 46450
rect 54674 46447 54686 46450
rect 54290 46401 54686 46447
rect 54290 46398 54302 46401
rect 54674 46398 54686 46401
rect 54738 46447 54750 46450
rect 55346 46447 55358 46450
rect 54738 46401 55358 46447
rect 54738 46398 54750 46401
rect 55346 46398 55358 46401
rect 55410 46398 55422 46450
rect 52222 46386 52274 46398
rect 66782 46386 66834 46398
rect 86942 46450 86994 46462
rect 86942 46386 86994 46398
rect 1344 46282 98560 46316
rect 1344 46230 4396 46282
rect 4448 46230 4520 46282
rect 4572 46230 4644 46282
rect 4696 46230 4768 46282
rect 4820 46230 13396 46282
rect 13448 46230 13520 46282
rect 13572 46230 13644 46282
rect 13696 46230 13768 46282
rect 13820 46230 22396 46282
rect 22448 46230 22520 46282
rect 22572 46230 22644 46282
rect 22696 46230 22768 46282
rect 22820 46230 31396 46282
rect 31448 46230 31520 46282
rect 31572 46230 31644 46282
rect 31696 46230 31768 46282
rect 31820 46230 40396 46282
rect 40448 46230 40520 46282
rect 40572 46230 40644 46282
rect 40696 46230 40768 46282
rect 40820 46230 49396 46282
rect 49448 46230 49520 46282
rect 49572 46230 49644 46282
rect 49696 46230 49768 46282
rect 49820 46230 58396 46282
rect 58448 46230 58520 46282
rect 58572 46230 58644 46282
rect 58696 46230 58768 46282
rect 58820 46230 67396 46282
rect 67448 46230 67520 46282
rect 67572 46230 67644 46282
rect 67696 46230 67768 46282
rect 67820 46230 76396 46282
rect 76448 46230 76520 46282
rect 76572 46230 76644 46282
rect 76696 46230 76768 46282
rect 76820 46230 85396 46282
rect 85448 46230 85520 46282
rect 85572 46230 85644 46282
rect 85696 46230 85768 46282
rect 85820 46230 94396 46282
rect 94448 46230 94520 46282
rect 94572 46230 94644 46282
rect 94696 46230 94768 46282
rect 94820 46230 98560 46282
rect 1344 46196 98560 46230
rect 34526 46114 34578 46126
rect 34526 46050 34578 46062
rect 73054 46114 73106 46126
rect 73054 46050 73106 46062
rect 89630 46114 89682 46126
rect 89630 46050 89682 46062
rect 14926 46002 14978 46014
rect 54126 46002 54178 46014
rect 50306 45950 50318 46002
rect 50370 45950 50382 46002
rect 14926 45938 14978 45950
rect 54126 45938 54178 45950
rect 77982 46002 78034 46014
rect 77982 45938 78034 45950
rect 79102 46002 79154 46014
rect 79102 45938 79154 45950
rect 89966 46002 90018 46014
rect 89966 45938 90018 45950
rect 27246 45890 27298 45902
rect 40686 45890 40738 45902
rect 60622 45890 60674 45902
rect 64878 45890 64930 45902
rect 30930 45838 30942 45890
rect 30994 45838 31006 45890
rect 31490 45838 31502 45890
rect 31554 45838 31566 45890
rect 47506 45838 47518 45890
rect 47570 45838 47582 45890
rect 49186 45838 49198 45890
rect 49250 45838 49262 45890
rect 55010 45838 55022 45890
rect 55074 45838 55086 45890
rect 57698 45838 57710 45890
rect 57762 45838 57774 45890
rect 58482 45838 58494 45890
rect 58546 45838 58558 45890
rect 59938 45838 59950 45890
rect 60002 45838 60014 45890
rect 61058 45838 61070 45890
rect 61122 45838 61134 45890
rect 27246 45826 27298 45838
rect 40686 45826 40738 45838
rect 60622 45826 60674 45838
rect 64878 45826 64930 45838
rect 68238 45890 68290 45902
rect 72718 45890 72770 45902
rect 68786 45838 68798 45890
rect 68850 45838 68862 45890
rect 68238 45826 68290 45838
rect 72718 45826 72770 45838
rect 72942 45890 72994 45902
rect 72942 45826 72994 45838
rect 77086 45890 77138 45902
rect 77086 45826 77138 45838
rect 77310 45890 77362 45902
rect 77310 45826 77362 45838
rect 77646 45890 77698 45902
rect 77646 45826 77698 45838
rect 79886 45890 79938 45902
rect 86158 45890 86210 45902
rect 91982 45890 92034 45902
rect 80434 45838 80446 45890
rect 80498 45838 80510 45890
rect 86482 45838 86494 45890
rect 86546 45838 86558 45890
rect 92530 45838 92542 45890
rect 92594 45838 92606 45890
rect 79886 45826 79938 45838
rect 86158 45826 86210 45838
rect 91982 45826 92034 45838
rect 1710 45778 1762 45790
rect 1710 45714 1762 45726
rect 25678 45778 25730 45790
rect 25678 45714 25730 45726
rect 26910 45778 26962 45790
rect 26910 45714 26962 45726
rect 29262 45778 29314 45790
rect 29262 45714 29314 45726
rect 30606 45778 30658 45790
rect 30606 45714 30658 45726
rect 33742 45778 33794 45790
rect 33742 45714 33794 45726
rect 38558 45778 38610 45790
rect 38558 45714 38610 45726
rect 40238 45778 40290 45790
rect 64542 45778 64594 45790
rect 48066 45726 48078 45778
rect 48130 45726 48142 45778
rect 49074 45726 49086 45778
rect 49138 45726 49150 45778
rect 55682 45726 55694 45778
rect 55746 45726 55758 45778
rect 56802 45726 56814 45778
rect 56866 45726 56878 45778
rect 40238 45714 40290 45726
rect 64542 45714 64594 45726
rect 79326 45778 79378 45790
rect 79326 45714 79378 45726
rect 82798 45778 82850 45790
rect 82798 45714 82850 45726
rect 2046 45666 2098 45678
rect 2046 45602 2098 45614
rect 2494 45666 2546 45678
rect 2494 45602 2546 45614
rect 3166 45666 3218 45678
rect 3166 45602 3218 45614
rect 21310 45666 21362 45678
rect 21310 45602 21362 45614
rect 39006 45666 39058 45678
rect 39006 45602 39058 45614
rect 39454 45666 39506 45678
rect 39454 45602 39506 45614
rect 39902 45666 39954 45678
rect 39902 45602 39954 45614
rect 54462 45666 54514 45678
rect 64094 45666 64146 45678
rect 56914 45614 56926 45666
rect 56978 45614 56990 45666
rect 63522 45614 63534 45666
rect 63586 45614 63598 45666
rect 54462 45602 54514 45614
rect 64094 45602 64146 45614
rect 64654 45666 64706 45678
rect 64654 45602 64706 45614
rect 65326 45666 65378 45678
rect 65326 45602 65378 45614
rect 67790 45666 67842 45678
rect 71934 45666 71986 45678
rect 71362 45614 71374 45666
rect 71426 45614 71438 45666
rect 67790 45602 67842 45614
rect 71934 45602 71986 45614
rect 73054 45666 73106 45678
rect 73054 45602 73106 45614
rect 77422 45666 77474 45678
rect 77422 45602 77474 45614
rect 79662 45666 79714 45678
rect 79662 45602 79714 45614
rect 83582 45666 83634 45678
rect 91310 45666 91362 45678
rect 95678 45666 95730 45678
rect 89058 45614 89070 45666
rect 89122 45614 89134 45666
rect 94994 45614 95006 45666
rect 95058 45614 95070 45666
rect 83582 45602 83634 45614
rect 91310 45602 91362 45614
rect 95678 45602 95730 45614
rect 1344 45498 98560 45532
rect 1344 45446 8896 45498
rect 8948 45446 9020 45498
rect 9072 45446 9144 45498
rect 9196 45446 9268 45498
rect 9320 45446 17896 45498
rect 17948 45446 18020 45498
rect 18072 45446 18144 45498
rect 18196 45446 18268 45498
rect 18320 45446 26896 45498
rect 26948 45446 27020 45498
rect 27072 45446 27144 45498
rect 27196 45446 27268 45498
rect 27320 45446 35896 45498
rect 35948 45446 36020 45498
rect 36072 45446 36144 45498
rect 36196 45446 36268 45498
rect 36320 45446 44896 45498
rect 44948 45446 45020 45498
rect 45072 45446 45144 45498
rect 45196 45446 45268 45498
rect 45320 45446 53896 45498
rect 53948 45446 54020 45498
rect 54072 45446 54144 45498
rect 54196 45446 54268 45498
rect 54320 45446 62896 45498
rect 62948 45446 63020 45498
rect 63072 45446 63144 45498
rect 63196 45446 63268 45498
rect 63320 45446 71896 45498
rect 71948 45446 72020 45498
rect 72072 45446 72144 45498
rect 72196 45446 72268 45498
rect 72320 45446 80896 45498
rect 80948 45446 81020 45498
rect 81072 45446 81144 45498
rect 81196 45446 81268 45498
rect 81320 45446 89896 45498
rect 89948 45446 90020 45498
rect 90072 45446 90144 45498
rect 90196 45446 90268 45498
rect 90320 45446 98560 45498
rect 1344 45412 98560 45446
rect 20302 45330 20354 45342
rect 5730 45278 5742 45330
rect 5794 45278 5806 45330
rect 20302 45266 20354 45278
rect 41022 45330 41074 45342
rect 41022 45266 41074 45278
rect 44494 45330 44546 45342
rect 44494 45266 44546 45278
rect 47294 45330 47346 45342
rect 47294 45266 47346 45278
rect 54462 45330 54514 45342
rect 54462 45266 54514 45278
rect 62414 45330 62466 45342
rect 62414 45266 62466 45278
rect 64542 45330 64594 45342
rect 64542 45266 64594 45278
rect 68574 45330 68626 45342
rect 68574 45266 68626 45278
rect 78654 45330 78706 45342
rect 78654 45266 78706 45278
rect 81006 45330 81058 45342
rect 81006 45266 81058 45278
rect 91198 45330 91250 45342
rect 91198 45266 91250 45278
rect 92878 45330 92930 45342
rect 92878 45266 92930 45278
rect 2046 45218 2098 45230
rect 2046 45154 2098 45166
rect 14254 45218 14306 45230
rect 14254 45154 14306 45166
rect 14590 45218 14642 45230
rect 19630 45218 19682 45230
rect 15474 45166 15486 45218
rect 15538 45166 15550 45218
rect 14590 45154 14642 45166
rect 19630 45154 19682 45166
rect 23438 45218 23490 45230
rect 23438 45154 23490 45166
rect 37438 45218 37490 45230
rect 43822 45218 43874 45230
rect 42018 45166 42030 45218
rect 42082 45166 42094 45218
rect 37438 45154 37490 45166
rect 43822 45154 43874 45166
rect 47518 45218 47570 45230
rect 47518 45154 47570 45166
rect 50206 45218 50258 45230
rect 50206 45154 50258 45166
rect 56926 45218 56978 45230
rect 56926 45154 56978 45166
rect 61294 45218 61346 45230
rect 76750 45218 76802 45230
rect 90638 45218 90690 45230
rect 63298 45166 63310 45218
rect 63362 45166 63374 45218
rect 71138 45166 71150 45218
rect 71202 45166 71214 45218
rect 77746 45166 77758 45218
rect 77810 45166 77822 45218
rect 91970 45166 91982 45218
rect 92034 45166 92046 45218
rect 61294 45154 61346 45166
rect 76750 45154 76802 45166
rect 90638 45154 90690 45166
rect 1710 45106 1762 45118
rect 1710 45042 1762 45054
rect 3054 45106 3106 45118
rect 14926 45106 14978 45118
rect 16494 45106 16546 45118
rect 20750 45106 20802 45118
rect 41358 45106 41410 45118
rect 47630 45106 47682 45118
rect 3378 45054 3390 45106
rect 3442 45054 3454 45106
rect 15362 45054 15374 45106
rect 15426 45054 15438 45106
rect 20066 45054 20078 45106
rect 20130 45054 20142 45106
rect 21074 45054 21086 45106
rect 21138 45054 21150 45106
rect 37986 45054 37998 45106
rect 38050 45054 38062 45106
rect 42130 45054 42142 45106
rect 42194 45054 42206 45106
rect 3054 45042 3106 45054
rect 14926 45042 14978 45054
rect 16494 45042 16546 45054
rect 20750 45042 20802 45054
rect 41358 45042 41410 45054
rect 47630 45042 47682 45054
rect 48078 45106 48130 45118
rect 48078 45042 48130 45054
rect 56590 45106 56642 45118
rect 56590 45042 56642 45054
rect 62750 45106 62802 45118
rect 68910 45106 68962 45118
rect 63522 45054 63534 45106
rect 63586 45054 63598 45106
rect 62750 45042 62802 45054
rect 68910 45042 68962 45054
rect 70142 45106 70194 45118
rect 70142 45042 70194 45054
rect 70478 45106 70530 45118
rect 78318 45106 78370 45118
rect 92542 45106 92594 45118
rect 71250 45054 71262 45106
rect 71314 45054 71326 45106
rect 77522 45054 77534 45106
rect 77586 45054 77598 45106
rect 91746 45054 91758 45106
rect 91810 45054 91822 45106
rect 70478 45042 70530 45054
rect 78318 45042 78370 45054
rect 92542 45042 92594 45054
rect 2494 44994 2546 45006
rect 2494 44930 2546 44942
rect 17614 44994 17666 45006
rect 42702 44994 42754 45006
rect 40002 44942 40014 44994
rect 40066 44942 40078 44994
rect 17614 44930 17666 44942
rect 42702 44930 42754 44942
rect 51662 44994 51714 45006
rect 51662 44930 51714 44942
rect 55918 44994 55970 45006
rect 55918 44930 55970 44942
rect 61742 44994 61794 45006
rect 61742 44930 61794 44942
rect 69470 44994 69522 45006
rect 69470 44930 69522 44942
rect 73614 44994 73666 45006
rect 73614 44930 73666 44942
rect 76302 44994 76354 45006
rect 76302 44930 76354 44942
rect 6526 44882 6578 44894
rect 6526 44818 6578 44830
rect 16158 44882 16210 44894
rect 16158 44818 16210 44830
rect 24222 44882 24274 44894
rect 24222 44818 24274 44830
rect 1344 44714 98560 44748
rect 1344 44662 4396 44714
rect 4448 44662 4520 44714
rect 4572 44662 4644 44714
rect 4696 44662 4768 44714
rect 4820 44662 13396 44714
rect 13448 44662 13520 44714
rect 13572 44662 13644 44714
rect 13696 44662 13768 44714
rect 13820 44662 22396 44714
rect 22448 44662 22520 44714
rect 22572 44662 22644 44714
rect 22696 44662 22768 44714
rect 22820 44662 31396 44714
rect 31448 44662 31520 44714
rect 31572 44662 31644 44714
rect 31696 44662 31768 44714
rect 31820 44662 40396 44714
rect 40448 44662 40520 44714
rect 40572 44662 40644 44714
rect 40696 44662 40768 44714
rect 40820 44662 49396 44714
rect 49448 44662 49520 44714
rect 49572 44662 49644 44714
rect 49696 44662 49768 44714
rect 49820 44662 58396 44714
rect 58448 44662 58520 44714
rect 58572 44662 58644 44714
rect 58696 44662 58768 44714
rect 58820 44662 67396 44714
rect 67448 44662 67520 44714
rect 67572 44662 67644 44714
rect 67696 44662 67768 44714
rect 67820 44662 76396 44714
rect 76448 44662 76520 44714
rect 76572 44662 76644 44714
rect 76696 44662 76768 44714
rect 76820 44662 85396 44714
rect 85448 44662 85520 44714
rect 85572 44662 85644 44714
rect 85696 44662 85768 44714
rect 85820 44662 94396 44714
rect 94448 44662 94520 44714
rect 94572 44662 94644 44714
rect 94696 44662 94768 44714
rect 94820 44662 98560 44714
rect 1344 44628 98560 44662
rect 41470 44546 41522 44558
rect 41470 44482 41522 44494
rect 45278 44546 45330 44558
rect 54910 44546 54962 44558
rect 46386 44494 46398 44546
rect 46450 44543 46462 44546
rect 46722 44543 46734 44546
rect 46450 44497 46734 44543
rect 46450 44494 46462 44497
rect 46722 44494 46734 44497
rect 46786 44494 46798 44546
rect 45278 44482 45330 44494
rect 54910 44482 54962 44494
rect 56366 44546 56418 44558
rect 56366 44482 56418 44494
rect 64430 44546 64482 44558
rect 64430 44482 64482 44494
rect 74062 44546 74114 44558
rect 74062 44482 74114 44494
rect 77982 44546 78034 44558
rect 77982 44482 78034 44494
rect 22542 44434 22594 44446
rect 22542 44370 22594 44382
rect 31054 44434 31106 44446
rect 31054 44370 31106 44382
rect 35982 44434 36034 44446
rect 35982 44370 36034 44382
rect 41806 44434 41858 44446
rect 54126 44434 54178 44446
rect 49074 44382 49086 44434
rect 49138 44382 49150 44434
rect 41806 44370 41858 44382
rect 54126 44370 54178 44382
rect 63086 44434 63138 44446
rect 63086 44370 63138 44382
rect 9438 44322 9490 44334
rect 8754 44270 8766 44322
rect 8818 44270 8830 44322
rect 9438 44258 9490 44270
rect 9774 44322 9826 44334
rect 11566 44322 11618 44334
rect 10210 44270 10222 44322
rect 10274 44270 10286 44322
rect 9774 44258 9826 44270
rect 11566 44258 11618 44270
rect 14254 44322 14306 44334
rect 22206 44322 22258 44334
rect 14802 44270 14814 44322
rect 14866 44270 14878 44322
rect 21746 44270 21758 44322
rect 21810 44270 21822 44322
rect 14254 44258 14306 44270
rect 22206 44258 22258 44270
rect 34190 44322 34242 44334
rect 37774 44322 37826 44334
rect 56702 44322 56754 44334
rect 34850 44270 34862 44322
rect 34914 44270 34926 44322
rect 38434 44270 38446 44322
rect 38498 44270 38510 44322
rect 45938 44270 45950 44322
rect 46002 44270 46014 44322
rect 48066 44270 48078 44322
rect 48130 44270 48142 44322
rect 51314 44270 51326 44322
rect 51378 44270 51390 44322
rect 55458 44270 55470 44322
rect 55522 44270 55534 44322
rect 34190 44258 34242 44270
rect 37774 44258 37826 44270
rect 56702 44258 56754 44270
rect 58494 44322 58546 44334
rect 58494 44258 58546 44270
rect 69694 44322 69746 44334
rect 69694 44258 69746 44270
rect 73614 44322 73666 44334
rect 73614 44258 73666 44270
rect 73838 44322 73890 44334
rect 74498 44270 74510 44322
rect 74562 44270 74574 44322
rect 75058 44270 75070 44322
rect 75122 44270 75134 44322
rect 77298 44270 77310 44322
rect 77362 44270 77374 44322
rect 96898 44270 96910 44322
rect 96962 44270 96974 44322
rect 73838 44258 73890 44270
rect 14030 44210 14082 44222
rect 44270 44210 44322 44222
rect 10322 44158 10334 44210
rect 10386 44158 10398 44210
rect 21410 44158 21422 44210
rect 21474 44158 21486 44210
rect 34962 44158 34974 44210
rect 35026 44158 35038 44210
rect 14030 44146 14082 44158
rect 44270 44146 44322 44158
rect 44942 44210 44994 44222
rect 47742 44210 47794 44222
rect 51998 44210 52050 44222
rect 46050 44158 46062 44210
rect 46114 44158 46126 44210
rect 48626 44158 48638 44210
rect 48690 44158 48702 44210
rect 49858 44158 49870 44210
rect 49922 44158 49934 44210
rect 44942 44146 44994 44158
rect 47742 44146 47794 44158
rect 51998 44146 52050 44158
rect 54574 44210 54626 44222
rect 78318 44210 78370 44222
rect 55682 44158 55694 44210
rect 55746 44158 55758 44210
rect 56914 44158 56926 44210
rect 56978 44158 56990 44210
rect 57474 44158 57486 44210
rect 57538 44158 57550 44210
rect 64642 44158 64654 44210
rect 64706 44158 64718 44210
rect 65202 44158 65214 44210
rect 65266 44158 65278 44210
rect 74050 44158 74062 44210
rect 74114 44158 74126 44210
rect 77410 44158 77422 44210
rect 77474 44158 77486 44210
rect 54574 44146 54626 44158
rect 78318 44146 78370 44158
rect 79774 44210 79826 44222
rect 79774 44146 79826 44158
rect 95566 44210 95618 44222
rect 95566 44146 95618 44158
rect 95902 44210 95954 44222
rect 95902 44146 95954 44158
rect 96238 44210 96290 44222
rect 96238 44146 96290 44158
rect 96574 44210 96626 44222
rect 98018 44158 98030 44210
rect 98082 44158 98094 44210
rect 96574 44146 96626 44158
rect 1822 44098 1874 44110
rect 1822 44034 1874 44046
rect 2606 44098 2658 44110
rect 2606 44034 2658 44046
rect 8318 44098 8370 44110
rect 8318 44034 8370 44046
rect 8990 44098 9042 44110
rect 8990 44034 9042 44046
rect 11118 44098 11170 44110
rect 17950 44098 18002 44110
rect 17378 44046 17390 44098
rect 17442 44046 17454 44098
rect 11118 44034 11170 44046
rect 17950 44034 18002 44046
rect 20750 44098 20802 44110
rect 20750 44034 20802 44046
rect 23102 44098 23154 44110
rect 23102 44034 23154 44046
rect 33854 44098 33906 44110
rect 33854 44034 33906 44046
rect 35534 44098 35586 44110
rect 43934 44098 43986 44110
rect 40898 44046 40910 44098
rect 40962 44046 40974 44098
rect 35534 44034 35586 44046
rect 43934 44034 43986 44046
rect 46734 44098 46786 44110
rect 46734 44034 46786 44046
rect 51662 44098 51714 44110
rect 51662 44034 51714 44046
rect 52894 44098 52946 44110
rect 52894 44034 52946 44046
rect 57934 44098 57986 44110
rect 57934 44034 57986 44046
rect 63534 44098 63586 44110
rect 63534 44034 63586 44046
rect 64094 44098 64146 44110
rect 64094 44034 64146 44046
rect 73054 44098 73106 44110
rect 73054 44034 73106 44046
rect 76638 44098 76690 44110
rect 76638 44034 76690 44046
rect 80110 44098 80162 44110
rect 80110 44034 80162 44046
rect 81118 44098 81170 44110
rect 81118 44034 81170 44046
rect 1344 43930 98560 43964
rect 1344 43878 8896 43930
rect 8948 43878 9020 43930
rect 9072 43878 9144 43930
rect 9196 43878 9268 43930
rect 9320 43878 17896 43930
rect 17948 43878 18020 43930
rect 18072 43878 18144 43930
rect 18196 43878 18268 43930
rect 18320 43878 26896 43930
rect 26948 43878 27020 43930
rect 27072 43878 27144 43930
rect 27196 43878 27268 43930
rect 27320 43878 35896 43930
rect 35948 43878 36020 43930
rect 36072 43878 36144 43930
rect 36196 43878 36268 43930
rect 36320 43878 44896 43930
rect 44948 43878 45020 43930
rect 45072 43878 45144 43930
rect 45196 43878 45268 43930
rect 45320 43878 53896 43930
rect 53948 43878 54020 43930
rect 54072 43878 54144 43930
rect 54196 43878 54268 43930
rect 54320 43878 62896 43930
rect 62948 43878 63020 43930
rect 63072 43878 63144 43930
rect 63196 43878 63268 43930
rect 63320 43878 71896 43930
rect 71948 43878 72020 43930
rect 72072 43878 72144 43930
rect 72196 43878 72268 43930
rect 72320 43878 80896 43930
rect 80948 43878 81020 43930
rect 81072 43878 81144 43930
rect 81196 43878 81268 43930
rect 81320 43878 89896 43930
rect 89948 43878 90020 43930
rect 90072 43878 90144 43930
rect 90196 43878 90268 43930
rect 90320 43878 98560 43930
rect 1344 43844 98560 43878
rect 55582 43762 55634 43774
rect 5394 43710 5406 43762
rect 5458 43710 5470 43762
rect 28578 43710 28590 43762
rect 28642 43710 28654 43762
rect 38658 43710 38670 43762
rect 38722 43710 38734 43762
rect 55582 43698 55634 43710
rect 60174 43762 60226 43774
rect 60174 43698 60226 43710
rect 71262 43762 71314 43774
rect 71262 43698 71314 43710
rect 75406 43762 75458 43774
rect 75406 43698 75458 43710
rect 77086 43762 77138 43774
rect 77086 43698 77138 43710
rect 2046 43650 2098 43662
rect 2046 43586 2098 43598
rect 6750 43650 6802 43662
rect 6750 43586 6802 43598
rect 7198 43650 7250 43662
rect 7198 43586 7250 43598
rect 12350 43650 12402 43662
rect 12350 43586 12402 43598
rect 13918 43650 13970 43662
rect 13918 43586 13970 43598
rect 25342 43650 25394 43662
rect 31726 43650 31778 43662
rect 30482 43598 30494 43650
rect 30546 43598 30558 43650
rect 25342 43586 25394 43598
rect 31726 43586 31778 43598
rect 33070 43650 33122 43662
rect 33070 43586 33122 43598
rect 33406 43650 33458 43662
rect 39678 43650 39730 43662
rect 37986 43598 37998 43650
rect 38050 43598 38062 43650
rect 33406 43586 33458 43598
rect 39678 43586 39730 43598
rect 43262 43650 43314 43662
rect 43262 43586 43314 43598
rect 46398 43650 46450 43662
rect 46398 43586 46450 43598
rect 47182 43650 47234 43662
rect 47182 43586 47234 43598
rect 52782 43650 52834 43662
rect 52782 43586 52834 43598
rect 53566 43650 53618 43662
rect 53566 43586 53618 43598
rect 53902 43650 53954 43662
rect 53902 43586 53954 43598
rect 56030 43650 56082 43662
rect 56030 43586 56082 43598
rect 59390 43650 59442 43662
rect 59390 43586 59442 43598
rect 62414 43650 62466 43662
rect 62414 43586 62466 43598
rect 63086 43650 63138 43662
rect 63086 43586 63138 43598
rect 63422 43650 63474 43662
rect 69918 43650 69970 43662
rect 65986 43598 65998 43650
rect 66050 43598 66062 43650
rect 63422 43586 63474 43598
rect 69918 43586 69970 43598
rect 70366 43650 70418 43662
rect 70366 43586 70418 43598
rect 71710 43650 71762 43662
rect 83694 43650 83746 43662
rect 73490 43598 73502 43650
rect 73554 43598 73566 43650
rect 76962 43598 76974 43650
rect 77026 43598 77038 43650
rect 71710 43586 71762 43598
rect 83694 43586 83746 43598
rect 84478 43650 84530 43662
rect 84478 43586 84530 43598
rect 86606 43650 86658 43662
rect 86606 43586 86658 43598
rect 91422 43650 91474 43662
rect 91422 43586 91474 43598
rect 94558 43650 94610 43662
rect 94558 43586 94610 43598
rect 2494 43538 2546 43550
rect 9438 43538 9490 43550
rect 25566 43538 25618 43550
rect 29262 43538 29314 43550
rect 1810 43486 1822 43538
rect 1874 43486 1886 43538
rect 2930 43486 2942 43538
rect 2994 43486 3006 43538
rect 10098 43486 10110 43538
rect 10162 43486 10174 43538
rect 26226 43486 26238 43538
rect 26290 43486 26302 43538
rect 2494 43474 2546 43486
rect 9438 43474 9490 43486
rect 25566 43474 25618 43486
rect 29262 43474 29314 43486
rect 29934 43538 29986 43550
rect 50094 43538 50146 43550
rect 56702 43538 56754 43550
rect 65438 43538 65490 43550
rect 30594 43486 30606 43538
rect 30658 43486 30670 43538
rect 34738 43486 34750 43538
rect 34802 43486 34814 43538
rect 35186 43486 35198 43538
rect 35250 43486 35262 43538
rect 35634 43486 35646 43538
rect 35698 43486 35710 43538
rect 35858 43486 35870 43538
rect 35922 43486 35934 43538
rect 38434 43486 38446 43538
rect 38498 43486 38510 43538
rect 43586 43486 43598 43538
rect 43650 43486 43662 43538
rect 44034 43486 44046 43538
rect 44098 43486 44110 43538
rect 50530 43486 50542 43538
rect 50594 43486 50606 43538
rect 57138 43486 57150 43538
rect 57202 43486 57214 43538
rect 29934 43474 29986 43486
rect 50094 43474 50146 43486
rect 56702 43474 56754 43486
rect 65438 43474 65490 43486
rect 65774 43538 65826 43550
rect 70702 43538 70754 43550
rect 66322 43486 66334 43538
rect 66386 43486 66398 43538
rect 66994 43486 67006 43538
rect 67058 43486 67070 43538
rect 65774 43474 65826 43486
rect 70702 43474 70754 43486
rect 72382 43538 72434 43550
rect 77198 43538 77250 43550
rect 73154 43486 73166 43538
rect 73218 43486 73230 43538
rect 75730 43486 75742 43538
rect 75794 43486 75806 43538
rect 76626 43486 76638 43538
rect 76690 43486 76702 43538
rect 72382 43474 72434 43486
rect 77198 43474 77250 43486
rect 80782 43538 80834 43550
rect 91646 43538 91698 43550
rect 81330 43486 81342 43538
rect 81394 43486 81406 43538
rect 92194 43486 92206 43538
rect 92258 43486 92270 43538
rect 80782 43474 80834 43486
rect 91646 43474 91698 43486
rect 31278 43426 31330 43438
rect 6290 43374 6302 43426
rect 6354 43374 6366 43426
rect 31278 43362 31330 43374
rect 32510 43426 32562 43438
rect 32510 43362 32562 43374
rect 39230 43426 39282 43438
rect 39230 43362 39282 43374
rect 64542 43426 64594 43438
rect 64542 43362 64594 43374
rect 64990 43426 65042 43438
rect 64990 43362 65042 43374
rect 72718 43426 72770 43438
rect 72718 43362 72770 43374
rect 74958 43426 75010 43438
rect 74958 43362 75010 43374
rect 80558 43426 80610 43438
rect 80558 43362 80610 43374
rect 90974 43426 91026 43438
rect 90974 43362 91026 43374
rect 5966 43314 6018 43326
rect 5966 43250 6018 43262
rect 13134 43314 13186 43326
rect 13134 43250 13186 43262
rect 29598 43314 29650 43326
rect 29598 43250 29650 43262
rect 66446 43314 66498 43326
rect 95342 43314 95394 43326
rect 74946 43262 74958 43314
rect 75010 43311 75022 43314
rect 75282 43311 75294 43314
rect 75010 43265 75294 43311
rect 75010 43262 75022 43265
rect 75282 43262 75294 43265
rect 75346 43262 75358 43314
rect 66446 43250 66498 43262
rect 95342 43250 95394 43262
rect 1344 43146 98560 43180
rect 1344 43094 4396 43146
rect 4448 43094 4520 43146
rect 4572 43094 4644 43146
rect 4696 43094 4768 43146
rect 4820 43094 13396 43146
rect 13448 43094 13520 43146
rect 13572 43094 13644 43146
rect 13696 43094 13768 43146
rect 13820 43094 22396 43146
rect 22448 43094 22520 43146
rect 22572 43094 22644 43146
rect 22696 43094 22768 43146
rect 22820 43094 31396 43146
rect 31448 43094 31520 43146
rect 31572 43094 31644 43146
rect 31696 43094 31768 43146
rect 31820 43094 40396 43146
rect 40448 43094 40520 43146
rect 40572 43094 40644 43146
rect 40696 43094 40768 43146
rect 40820 43094 49396 43146
rect 49448 43094 49520 43146
rect 49572 43094 49644 43146
rect 49696 43094 49768 43146
rect 49820 43094 58396 43146
rect 58448 43094 58520 43146
rect 58572 43094 58644 43146
rect 58696 43094 58768 43146
rect 58820 43094 67396 43146
rect 67448 43094 67520 43146
rect 67572 43094 67644 43146
rect 67696 43094 67768 43146
rect 67820 43094 76396 43146
rect 76448 43094 76520 43146
rect 76572 43094 76644 43146
rect 76696 43094 76768 43146
rect 76820 43094 85396 43146
rect 85448 43094 85520 43146
rect 85572 43094 85644 43146
rect 85696 43094 85768 43146
rect 85820 43094 94396 43146
rect 94448 43094 94520 43146
rect 94572 43094 94644 43146
rect 94696 43094 94768 43146
rect 94820 43094 98560 43146
rect 1344 43060 98560 43094
rect 35086 42978 35138 42990
rect 35086 42914 35138 42926
rect 65774 42978 65826 42990
rect 65774 42914 65826 42926
rect 73278 42978 73330 42990
rect 73278 42914 73330 42926
rect 92766 42978 92818 42990
rect 92766 42914 92818 42926
rect 29374 42866 29426 42878
rect 29374 42802 29426 42814
rect 31166 42866 31218 42878
rect 31166 42802 31218 42814
rect 61854 42866 61906 42878
rect 61854 42802 61906 42814
rect 14366 42754 14418 42766
rect 12674 42702 12686 42754
rect 12738 42702 12750 42754
rect 13794 42702 13806 42754
rect 13858 42702 13870 42754
rect 14366 42690 14418 42702
rect 18958 42754 19010 42766
rect 20190 42754 20242 42766
rect 19506 42702 19518 42754
rect 19570 42702 19582 42754
rect 18958 42690 19010 42702
rect 20190 42690 20242 42702
rect 27246 42754 27298 42766
rect 27246 42690 27298 42702
rect 31614 42754 31666 42766
rect 62302 42754 62354 42766
rect 69806 42754 69858 42766
rect 86606 42754 86658 42766
rect 90414 42754 90466 42766
rect 32050 42702 32062 42754
rect 32114 42702 32126 42754
rect 62738 42702 62750 42754
rect 62802 42702 62814 42754
rect 70242 42702 70254 42754
rect 70306 42702 70318 42754
rect 86930 42702 86942 42754
rect 86994 42702 87006 42754
rect 92306 42702 92318 42754
rect 92370 42702 92382 42754
rect 96898 42702 96910 42754
rect 96962 42702 96974 42754
rect 31614 42690 31666 42702
rect 62302 42690 62354 42702
rect 69806 42690 69858 42702
rect 86606 42690 86658 42702
rect 90414 42690 90466 42702
rect 1710 42642 1762 42654
rect 14702 42642 14754 42654
rect 26910 42642 26962 42654
rect 13570 42590 13582 42642
rect 13634 42590 13646 42642
rect 19394 42590 19406 42642
rect 19458 42590 19470 42642
rect 1710 42578 1762 42590
rect 14702 42578 14754 42590
rect 26910 42578 26962 42590
rect 34302 42642 34354 42654
rect 34302 42578 34354 42590
rect 77758 42642 77810 42654
rect 96238 42642 96290 42654
rect 91970 42590 91982 42642
rect 92034 42590 92046 42642
rect 77758 42578 77810 42590
rect 96238 42578 96290 42590
rect 96574 42642 96626 42654
rect 98018 42590 98030 42642
rect 98082 42590 98094 42642
rect 96574 42578 96626 42590
rect 2046 42530 2098 42542
rect 2046 42466 2098 42478
rect 2494 42530 2546 42542
rect 2494 42466 2546 42478
rect 2942 42530 2994 42542
rect 2942 42466 2994 42478
rect 12238 42530 12290 42542
rect 12238 42466 12290 42478
rect 12910 42530 12962 42542
rect 12910 42466 12962 42478
rect 15262 42530 15314 42542
rect 15262 42466 15314 42478
rect 20526 42530 20578 42542
rect 20526 42466 20578 42478
rect 21310 42530 21362 42542
rect 21310 42466 21362 42478
rect 21870 42530 21922 42542
rect 69358 42530 69410 42542
rect 75406 42530 75458 42542
rect 64978 42478 64990 42530
rect 65042 42478 65054 42530
rect 72482 42478 72494 42530
rect 72546 42478 72558 42530
rect 21870 42466 21922 42478
rect 69358 42466 69410 42478
rect 75406 42466 75458 42478
rect 78094 42530 78146 42542
rect 90078 42530 90130 42542
rect 89506 42478 89518 42530
rect 89570 42478 89582 42530
rect 78094 42466 78146 42478
rect 90078 42466 90130 42478
rect 90862 42530 90914 42542
rect 90862 42466 90914 42478
rect 91422 42530 91474 42542
rect 91422 42466 91474 42478
rect 93102 42530 93154 42542
rect 93102 42466 93154 42478
rect 1344 42362 98560 42396
rect 1344 42310 8896 42362
rect 8948 42310 9020 42362
rect 9072 42310 9144 42362
rect 9196 42310 9268 42362
rect 9320 42310 17896 42362
rect 17948 42310 18020 42362
rect 18072 42310 18144 42362
rect 18196 42310 18268 42362
rect 18320 42310 26896 42362
rect 26948 42310 27020 42362
rect 27072 42310 27144 42362
rect 27196 42310 27268 42362
rect 27320 42310 35896 42362
rect 35948 42310 36020 42362
rect 36072 42310 36144 42362
rect 36196 42310 36268 42362
rect 36320 42310 44896 42362
rect 44948 42310 45020 42362
rect 45072 42310 45144 42362
rect 45196 42310 45268 42362
rect 45320 42310 53896 42362
rect 53948 42310 54020 42362
rect 54072 42310 54144 42362
rect 54196 42310 54268 42362
rect 54320 42310 62896 42362
rect 62948 42310 63020 42362
rect 63072 42310 63144 42362
rect 63196 42310 63268 42362
rect 63320 42310 71896 42362
rect 71948 42310 72020 42362
rect 72072 42310 72144 42362
rect 72196 42310 72268 42362
rect 72320 42310 80896 42362
rect 80948 42310 81020 42362
rect 81072 42310 81144 42362
rect 81196 42310 81268 42362
rect 81320 42310 89896 42362
rect 89948 42310 90020 42362
rect 90072 42310 90144 42362
rect 90196 42310 90268 42362
rect 90320 42310 98560 42362
rect 1344 42276 98560 42310
rect 77534 42194 77586 42206
rect 5730 42142 5742 42194
rect 5794 42142 5806 42194
rect 16370 42142 16382 42194
rect 16434 42142 16446 42194
rect 77534 42130 77586 42142
rect 86830 42194 86882 42206
rect 86830 42130 86882 42142
rect 91982 42194 92034 42206
rect 91982 42130 92034 42142
rect 20414 42082 20466 42094
rect 20414 42018 20466 42030
rect 23550 42082 23602 42094
rect 23550 42018 23602 42030
rect 24446 42082 24498 42094
rect 24446 42018 24498 42030
rect 38558 42082 38610 42094
rect 38558 42018 38610 42030
rect 39230 42082 39282 42094
rect 39230 42018 39282 42030
rect 44046 42082 44098 42094
rect 44046 42018 44098 42030
rect 49646 42082 49698 42094
rect 58382 42082 58434 42094
rect 79102 42082 79154 42094
rect 57586 42030 57598 42082
rect 57650 42030 57662 42082
rect 78194 42030 78206 42082
rect 78258 42030 78270 42082
rect 78642 42030 78654 42082
rect 78706 42030 78718 42082
rect 88162 42030 88174 42082
rect 88226 42030 88238 42082
rect 49646 42018 49698 42030
rect 58382 42018 58434 42030
rect 79102 42018 79154 42030
rect 2830 41970 2882 41982
rect 13246 41970 13298 41982
rect 17502 41970 17554 41982
rect 3154 41918 3166 41970
rect 3218 41918 3230 41970
rect 13794 41918 13806 41970
rect 13858 41918 13870 41970
rect 2830 41906 2882 41918
rect 13246 41906 13298 41918
rect 17502 41906 17554 41918
rect 19742 41970 19794 41982
rect 20638 41970 20690 41982
rect 39566 41970 39618 41982
rect 20178 41918 20190 41970
rect 20242 41918 20254 41970
rect 21186 41918 21198 41970
rect 21250 41918 21262 41970
rect 19742 41906 19794 41918
rect 20638 41906 20690 41918
rect 39566 41906 39618 41918
rect 44494 41970 44546 41982
rect 44494 41906 44546 41918
rect 54238 41970 54290 41982
rect 54238 41906 54290 41918
rect 55582 41970 55634 41982
rect 67790 41970 67842 41982
rect 57474 41918 57486 41970
rect 57538 41918 57550 41970
rect 55582 41906 55634 41918
rect 67790 41906 67842 41918
rect 76862 41970 76914 41982
rect 76862 41906 76914 41918
rect 87166 41970 87218 41982
rect 88846 41970 88898 41982
rect 88386 41918 88398 41970
rect 88450 41918 88462 41970
rect 87166 41906 87218 41918
rect 88846 41906 88898 41918
rect 89182 41970 89234 41982
rect 89182 41906 89234 41918
rect 92318 41970 92370 41982
rect 92318 41906 92370 41918
rect 2158 41858 2210 41870
rect 2158 41794 2210 41806
rect 6638 41858 6690 41870
rect 6638 41794 6690 41806
rect 50318 41858 50370 41870
rect 50318 41794 50370 41806
rect 53342 41858 53394 41870
rect 53342 41794 53394 41806
rect 53790 41858 53842 41870
rect 53790 41794 53842 41806
rect 54686 41858 54738 41870
rect 54686 41794 54738 41806
rect 56030 41858 56082 41870
rect 56030 41794 56082 41806
rect 75966 41858 76018 41870
rect 75966 41794 76018 41806
rect 76414 41858 76466 41870
rect 76414 41794 76466 41806
rect 77870 41858 77922 41870
rect 77870 41794 77922 41806
rect 6302 41746 6354 41758
rect 6302 41682 6354 41694
rect 16942 41746 16994 41758
rect 16942 41682 16994 41694
rect 56702 41746 56754 41758
rect 56702 41682 56754 41694
rect 57038 41746 57090 41758
rect 57038 41682 57090 41694
rect 1344 41578 98560 41612
rect 1344 41526 4396 41578
rect 4448 41526 4520 41578
rect 4572 41526 4644 41578
rect 4696 41526 4768 41578
rect 4820 41526 13396 41578
rect 13448 41526 13520 41578
rect 13572 41526 13644 41578
rect 13696 41526 13768 41578
rect 13820 41526 22396 41578
rect 22448 41526 22520 41578
rect 22572 41526 22644 41578
rect 22696 41526 22768 41578
rect 22820 41526 31396 41578
rect 31448 41526 31520 41578
rect 31572 41526 31644 41578
rect 31696 41526 31768 41578
rect 31820 41526 40396 41578
rect 40448 41526 40520 41578
rect 40572 41526 40644 41578
rect 40696 41526 40768 41578
rect 40820 41526 49396 41578
rect 49448 41526 49520 41578
rect 49572 41526 49644 41578
rect 49696 41526 49768 41578
rect 49820 41526 58396 41578
rect 58448 41526 58520 41578
rect 58572 41526 58644 41578
rect 58696 41526 58768 41578
rect 58820 41526 67396 41578
rect 67448 41526 67520 41578
rect 67572 41526 67644 41578
rect 67696 41526 67768 41578
rect 67820 41526 76396 41578
rect 76448 41526 76520 41578
rect 76572 41526 76644 41578
rect 76696 41526 76768 41578
rect 76820 41526 85396 41578
rect 85448 41526 85520 41578
rect 85572 41526 85644 41578
rect 85696 41526 85768 41578
rect 85820 41526 94396 41578
rect 94448 41526 94520 41578
rect 94572 41526 94644 41578
rect 94696 41526 94768 41578
rect 94820 41526 98560 41578
rect 1344 41492 98560 41526
rect 53230 41410 53282 41422
rect 53230 41346 53282 41358
rect 81566 41410 81618 41422
rect 81566 41346 81618 41358
rect 33742 41298 33794 41310
rect 33742 41234 33794 41246
rect 42366 41298 42418 41310
rect 87614 41298 87666 41310
rect 76850 41246 76862 41298
rect 76914 41246 76926 41298
rect 42366 41234 42418 41246
rect 87614 41234 87666 41246
rect 34526 41186 34578 41198
rect 35870 41186 35922 41198
rect 35298 41134 35310 41186
rect 35362 41134 35374 41186
rect 34526 41122 34578 41134
rect 35870 41122 35922 41134
rect 38558 41186 38610 41198
rect 44718 41186 44770 41198
rect 63982 41186 64034 41198
rect 71038 41186 71090 41198
rect 75070 41186 75122 41198
rect 38994 41134 39006 41186
rect 39058 41134 39070 41186
rect 44034 41134 44046 41186
rect 44098 41134 44110 41186
rect 45266 41134 45278 41186
rect 45330 41134 45342 41186
rect 48850 41134 48862 41186
rect 48914 41134 48926 41186
rect 49522 41134 49534 41186
rect 49586 41134 49598 41186
rect 54562 41134 54574 41186
rect 54626 41134 54638 41186
rect 55682 41134 55694 41186
rect 55746 41134 55758 41186
rect 56130 41134 56142 41186
rect 56194 41134 56206 41186
rect 57026 41134 57038 41186
rect 57090 41134 57102 41186
rect 58930 41134 58942 41186
rect 58994 41134 59006 41186
rect 64642 41134 64654 41186
rect 64706 41134 64718 41186
rect 71586 41134 71598 41186
rect 71650 41134 71662 41186
rect 38558 41122 38610 41134
rect 44718 41122 44770 41134
rect 63982 41122 64034 41134
rect 71038 41122 71090 41134
rect 75070 41122 75122 41134
rect 76750 41186 76802 41198
rect 77970 41134 77982 41186
rect 78034 41134 78046 41186
rect 78418 41134 78430 41186
rect 78482 41134 78494 41186
rect 96898 41134 96910 41186
rect 96962 41134 96974 41186
rect 76750 41122 76802 41134
rect 1710 41074 1762 41086
rect 1710 41010 1762 41022
rect 2382 41074 2434 41086
rect 2382 41010 2434 41022
rect 8878 41074 8930 41086
rect 8878 41010 8930 41022
rect 19070 41074 19122 41086
rect 42030 41074 42082 41086
rect 35186 41022 35198 41074
rect 35250 41022 35262 41074
rect 19070 41010 19122 41022
rect 42030 41010 42082 41022
rect 44270 41074 44322 41086
rect 44270 41010 44322 41022
rect 47630 41074 47682 41086
rect 50990 41074 51042 41086
rect 63758 41074 63810 41086
rect 48738 41022 48750 41074
rect 48802 41022 48814 41074
rect 52658 41022 52670 41074
rect 52722 41022 52734 41074
rect 57810 41022 57822 41074
rect 57874 41022 57886 41074
rect 47630 41010 47682 41022
rect 50990 41010 51042 41022
rect 63758 41010 63810 41022
rect 70814 41074 70866 41086
rect 70814 41010 70866 41022
rect 74734 41074 74786 41086
rect 74734 41010 74786 41022
rect 76302 41074 76354 41086
rect 76302 41010 76354 41022
rect 76526 41074 76578 41086
rect 76526 41010 76578 41022
rect 76862 41074 76914 41086
rect 76862 41010 76914 41022
rect 96238 41074 96290 41086
rect 96238 41010 96290 41022
rect 96574 41074 96626 41086
rect 98018 41022 98030 41074
rect 98082 41022 98094 41074
rect 96574 41010 96626 41022
rect 2046 40962 2098 40974
rect 2046 40898 2098 40910
rect 2718 40962 2770 40974
rect 2718 40898 2770 40910
rect 3166 40962 3218 40974
rect 3166 40898 3218 40910
rect 5742 40962 5794 40974
rect 5742 40898 5794 40910
rect 9326 40962 9378 40974
rect 9326 40898 9378 40910
rect 25454 40962 25506 40974
rect 25454 40898 25506 40910
rect 31502 40962 31554 40974
rect 31502 40898 31554 40910
rect 33294 40962 33346 40974
rect 33294 40898 33346 40910
rect 34190 40962 34242 40974
rect 48414 40962 48466 40974
rect 50654 40962 50706 40974
rect 41458 40910 41470 40962
rect 41522 40910 41534 40962
rect 48962 40910 48974 40962
rect 49026 40910 49038 40962
rect 49970 40910 49982 40962
rect 50034 40910 50046 40962
rect 34190 40898 34242 40910
rect 48414 40898 48466 40910
rect 50654 40898 50706 40910
rect 52222 40962 52274 40974
rect 67678 40962 67730 40974
rect 59266 40910 59278 40962
rect 59330 40910 59342 40962
rect 66994 40910 67006 40962
rect 67058 40910 67070 40962
rect 52222 40898 52274 40910
rect 67678 40898 67730 40910
rect 68574 40962 68626 40974
rect 75630 40962 75682 40974
rect 74050 40910 74062 40962
rect 74114 40910 74126 40962
rect 68574 40898 68626 40910
rect 75630 40898 75682 40910
rect 77646 40962 77698 40974
rect 82574 40962 82626 40974
rect 80882 40910 80894 40962
rect 80946 40910 80958 40962
rect 77646 40898 77698 40910
rect 82574 40898 82626 40910
rect 84590 40962 84642 40974
rect 84590 40898 84642 40910
rect 1344 40794 98560 40828
rect 1344 40742 8896 40794
rect 8948 40742 9020 40794
rect 9072 40742 9144 40794
rect 9196 40742 9268 40794
rect 9320 40742 17896 40794
rect 17948 40742 18020 40794
rect 18072 40742 18144 40794
rect 18196 40742 18268 40794
rect 18320 40742 26896 40794
rect 26948 40742 27020 40794
rect 27072 40742 27144 40794
rect 27196 40742 27268 40794
rect 27320 40742 35896 40794
rect 35948 40742 36020 40794
rect 36072 40742 36144 40794
rect 36196 40742 36268 40794
rect 36320 40742 44896 40794
rect 44948 40742 45020 40794
rect 45072 40742 45144 40794
rect 45196 40742 45268 40794
rect 45320 40742 53896 40794
rect 53948 40742 54020 40794
rect 54072 40742 54144 40794
rect 54196 40742 54268 40794
rect 54320 40742 62896 40794
rect 62948 40742 63020 40794
rect 63072 40742 63144 40794
rect 63196 40742 63268 40794
rect 63320 40742 71896 40794
rect 71948 40742 72020 40794
rect 72072 40742 72144 40794
rect 72196 40742 72268 40794
rect 72320 40742 80896 40794
rect 80948 40742 81020 40794
rect 81072 40742 81144 40794
rect 81196 40742 81268 40794
rect 81320 40742 89896 40794
rect 89948 40742 90020 40794
rect 90072 40742 90144 40794
rect 90196 40742 90268 40794
rect 90320 40742 98560 40794
rect 1344 40708 98560 40742
rect 22654 40626 22706 40638
rect 4722 40574 4734 40626
rect 4786 40574 4798 40626
rect 8306 40574 8318 40626
rect 8370 40574 8382 40626
rect 12338 40574 12350 40626
rect 12402 40574 12414 40626
rect 21970 40574 21982 40626
rect 22034 40574 22046 40626
rect 22654 40562 22706 40574
rect 22990 40626 23042 40638
rect 31390 40626 31442 40638
rect 39902 40626 39954 40638
rect 28242 40574 28254 40626
rect 28306 40574 28318 40626
rect 38994 40574 39006 40626
rect 39058 40574 39070 40626
rect 22990 40562 23042 40574
rect 31390 40562 31442 40574
rect 39902 40562 39954 40574
rect 41022 40626 41074 40638
rect 41022 40562 41074 40574
rect 44830 40626 44882 40638
rect 44830 40562 44882 40574
rect 46510 40626 46562 40638
rect 46510 40562 46562 40574
rect 48862 40626 48914 40638
rect 53678 40626 53730 40638
rect 52546 40574 52558 40626
rect 52610 40574 52622 40626
rect 48862 40562 48914 40574
rect 53678 40562 53730 40574
rect 55358 40626 55410 40638
rect 55358 40562 55410 40574
rect 57822 40626 57874 40638
rect 61742 40626 61794 40638
rect 60946 40574 60958 40626
rect 61010 40574 61022 40626
rect 57822 40562 57874 40574
rect 61742 40562 61794 40574
rect 65214 40626 65266 40638
rect 65214 40562 65266 40574
rect 65998 40626 66050 40638
rect 65998 40562 66050 40574
rect 72270 40626 72322 40638
rect 72270 40562 72322 40574
rect 76302 40626 76354 40638
rect 85934 40626 85986 40638
rect 85362 40574 85374 40626
rect 85426 40574 85438 40626
rect 76302 40562 76354 40574
rect 85934 40562 85986 40574
rect 90750 40626 90802 40638
rect 90750 40562 90802 40574
rect 91422 40626 91474 40638
rect 96574 40626 96626 40638
rect 94770 40574 94782 40626
rect 94834 40574 94846 40626
rect 91422 40562 91474 40574
rect 96574 40562 96626 40574
rect 16830 40514 16882 40526
rect 30942 40514 30994 40526
rect 17602 40462 17614 40514
rect 17666 40462 17678 40514
rect 30370 40462 30382 40514
rect 30434 40462 30446 40514
rect 16830 40450 16882 40462
rect 30942 40450 30994 40462
rect 33070 40514 33122 40526
rect 33070 40450 33122 40462
rect 33406 40514 33458 40526
rect 33406 40450 33458 40462
rect 37998 40514 38050 40526
rect 42702 40514 42754 40526
rect 57038 40514 57090 40526
rect 41570 40462 41582 40514
rect 41634 40462 41646 40514
rect 42018 40462 42030 40514
rect 42082 40462 42094 40514
rect 45938 40462 45950 40514
rect 46002 40462 46014 40514
rect 54562 40462 54574 40514
rect 54626 40462 54638 40514
rect 37998 40450 38050 40462
rect 42702 40450 42754 40462
rect 57038 40450 57090 40462
rect 57374 40514 57426 40526
rect 86270 40514 86322 40526
rect 67106 40462 67118 40514
rect 67170 40462 67182 40514
rect 67442 40462 67454 40514
rect 67506 40462 67518 40514
rect 68114 40462 68126 40514
rect 68178 40462 68190 40514
rect 74162 40462 74174 40514
rect 74226 40462 74238 40514
rect 76514 40462 76526 40514
rect 76578 40462 76590 40514
rect 57374 40450 57426 40462
rect 86270 40450 86322 40462
rect 1822 40402 1874 40414
rect 5630 40402 5682 40414
rect 13582 40402 13634 40414
rect 18622 40402 18674 40414
rect 2146 40350 2158 40402
rect 2210 40350 2222 40402
rect 5954 40350 5966 40402
rect 6018 40350 6030 40402
rect 9538 40350 9550 40402
rect 9602 40350 9614 40402
rect 10098 40350 10110 40402
rect 10162 40350 10174 40402
rect 17490 40350 17502 40402
rect 17554 40350 17566 40402
rect 1822 40338 1874 40350
rect 5630 40338 5682 40350
rect 13582 40338 13634 40350
rect 18622 40338 18674 40350
rect 19182 40402 19234 40414
rect 25454 40402 25506 40414
rect 28926 40402 28978 40414
rect 19506 40350 19518 40402
rect 19570 40350 19582 40402
rect 25890 40350 25902 40402
rect 25954 40350 25966 40402
rect 19182 40338 19234 40350
rect 25454 40338 25506 40350
rect 28926 40338 28978 40350
rect 29598 40402 29650 40414
rect 39454 40402 39506 40414
rect 49422 40402 49474 40414
rect 53118 40402 53170 40414
rect 65550 40402 65602 40414
rect 30146 40350 30158 40402
rect 30210 40350 30222 40402
rect 34962 40350 34974 40402
rect 35026 40350 35038 40402
rect 35410 40350 35422 40402
rect 35474 40350 35486 40402
rect 35746 40350 35758 40402
rect 35810 40350 35822 40402
rect 36082 40350 36094 40402
rect 36146 40350 36158 40402
rect 38658 40350 38670 40402
rect 38722 40350 38734 40402
rect 45826 40350 45838 40402
rect 45890 40350 45902 40402
rect 50082 40350 50094 40402
rect 50146 40350 50158 40402
rect 54786 40350 54798 40402
rect 54850 40350 54862 40402
rect 58146 40350 58158 40402
rect 58210 40350 58222 40402
rect 58594 40350 58606 40402
rect 58658 40350 58670 40402
rect 29598 40338 29650 40350
rect 39454 40338 39506 40350
rect 49422 40338 49474 40350
rect 53118 40338 53170 40350
rect 65550 40338 65602 40350
rect 66558 40402 66610 40414
rect 71710 40402 71762 40414
rect 68226 40350 68238 40402
rect 68290 40350 68302 40402
rect 68898 40350 68910 40402
rect 68962 40350 68974 40402
rect 69346 40350 69358 40402
rect 69410 40350 69422 40402
rect 66558 40338 66610 40350
rect 71710 40338 71762 40350
rect 72606 40402 72658 40414
rect 72606 40338 72658 40350
rect 73166 40402 73218 40414
rect 82462 40402 82514 40414
rect 91870 40402 91922 40414
rect 95342 40402 95394 40414
rect 73938 40350 73950 40402
rect 74002 40350 74014 40402
rect 76626 40350 76638 40402
rect 76690 40350 76702 40402
rect 77410 40350 77422 40402
rect 77474 40350 77486 40402
rect 77746 40350 77758 40402
rect 77810 40350 77822 40402
rect 82786 40350 82798 40402
rect 82850 40350 82862 40402
rect 91186 40350 91198 40402
rect 91250 40350 91262 40402
rect 92194 40350 92206 40402
rect 92258 40350 92270 40402
rect 73166 40338 73218 40350
rect 82462 40338 82514 40350
rect 91870 40338 91922 40350
rect 95342 40338 95394 40350
rect 96238 40402 96290 40414
rect 96238 40338 96290 40350
rect 18286 40290 18338 40302
rect 18286 40226 18338 40238
rect 40350 40290 40402 40302
rect 40350 40226 40402 40238
rect 44382 40290 44434 40302
rect 44382 40226 44434 40238
rect 45166 40290 45218 40302
rect 45166 40226 45218 40238
rect 54014 40290 54066 40302
rect 54014 40226 54066 40238
rect 73502 40290 73554 40302
rect 73502 40226 73554 40238
rect 78094 40290 78146 40302
rect 78094 40226 78146 40238
rect 5294 40178 5346 40190
rect 5294 40114 5346 40126
rect 9102 40178 9154 40190
rect 9102 40114 9154 40126
rect 13134 40178 13186 40190
rect 13134 40114 13186 40126
rect 29262 40178 29314 40190
rect 29262 40114 29314 40126
rect 41358 40178 41410 40190
rect 41358 40114 41410 40126
rect 66894 40178 66946 40190
rect 66894 40114 66946 40126
rect 69694 40178 69746 40190
rect 69694 40114 69746 40126
rect 1344 40010 98560 40044
rect 1344 39958 4396 40010
rect 4448 39958 4520 40010
rect 4572 39958 4644 40010
rect 4696 39958 4768 40010
rect 4820 39958 13396 40010
rect 13448 39958 13520 40010
rect 13572 39958 13644 40010
rect 13696 39958 13768 40010
rect 13820 39958 22396 40010
rect 22448 39958 22520 40010
rect 22572 39958 22644 40010
rect 22696 39958 22768 40010
rect 22820 39958 31396 40010
rect 31448 39958 31520 40010
rect 31572 39958 31644 40010
rect 31696 39958 31768 40010
rect 31820 39958 40396 40010
rect 40448 39958 40520 40010
rect 40572 39958 40644 40010
rect 40696 39958 40768 40010
rect 40820 39958 49396 40010
rect 49448 39958 49520 40010
rect 49572 39958 49644 40010
rect 49696 39958 49768 40010
rect 49820 39958 58396 40010
rect 58448 39958 58520 40010
rect 58572 39958 58644 40010
rect 58696 39958 58768 40010
rect 58820 39958 67396 40010
rect 67448 39958 67520 40010
rect 67572 39958 67644 40010
rect 67696 39958 67768 40010
rect 67820 39958 76396 40010
rect 76448 39958 76520 40010
rect 76572 39958 76644 40010
rect 76696 39958 76768 40010
rect 76820 39958 85396 40010
rect 85448 39958 85520 40010
rect 85572 39958 85644 40010
rect 85696 39958 85768 40010
rect 85820 39958 94396 40010
rect 94448 39958 94520 40010
rect 94572 39958 94644 40010
rect 94696 39958 94768 40010
rect 94820 39958 98560 40010
rect 1344 39924 98560 39958
rect 12462 39842 12514 39854
rect 12462 39778 12514 39790
rect 34862 39842 34914 39854
rect 34862 39778 34914 39790
rect 9214 39730 9266 39742
rect 9214 39666 9266 39678
rect 29262 39730 29314 39742
rect 29262 39666 29314 39678
rect 30942 39730 30994 39742
rect 30942 39666 30994 39678
rect 37662 39730 37714 39742
rect 37662 39666 37714 39678
rect 48414 39730 48466 39742
rect 48414 39666 48466 39678
rect 53230 39730 53282 39742
rect 53230 39666 53282 39678
rect 53678 39730 53730 39742
rect 53678 39666 53730 39678
rect 67230 39730 67282 39742
rect 67230 39666 67282 39678
rect 67678 39730 67730 39742
rect 67678 39666 67730 39678
rect 69022 39730 69074 39742
rect 69022 39666 69074 39678
rect 82126 39730 82178 39742
rect 82126 39666 82178 39678
rect 82574 39730 82626 39742
rect 82574 39666 82626 39678
rect 90638 39730 90690 39742
rect 90638 39666 90690 39678
rect 31166 39618 31218 39630
rect 36542 39618 36594 39630
rect 1810 39566 1822 39618
rect 1874 39566 1886 39618
rect 11666 39566 11678 39618
rect 11730 39566 11742 39618
rect 18386 39566 18398 39618
rect 18450 39566 18462 39618
rect 26786 39566 26798 39618
rect 26850 39566 26862 39618
rect 31826 39566 31838 39618
rect 31890 39566 31902 39618
rect 31166 39554 31218 39566
rect 36542 39554 36594 39566
rect 37326 39618 37378 39630
rect 37326 39554 37378 39566
rect 68350 39618 68402 39630
rect 68350 39554 68402 39566
rect 68686 39618 68738 39630
rect 68686 39554 68738 39566
rect 82462 39618 82514 39630
rect 83918 39618 83970 39630
rect 83010 39566 83022 39618
rect 83074 39566 83086 39618
rect 82462 39554 82514 39566
rect 83918 39554 83970 39566
rect 84926 39618 84978 39630
rect 84926 39554 84978 39566
rect 85038 39618 85090 39630
rect 85598 39618 85650 39630
rect 85362 39566 85374 39618
rect 85426 39566 85438 39618
rect 85038 39554 85090 39566
rect 85598 39554 85650 39566
rect 86606 39618 86658 39630
rect 87154 39566 87166 39618
rect 87218 39566 87230 39618
rect 96898 39566 96910 39618
rect 96962 39566 96974 39618
rect 86606 39554 86658 39566
rect 2382 39506 2434 39518
rect 2382 39442 2434 39454
rect 5630 39506 5682 39518
rect 12798 39506 12850 39518
rect 11890 39454 11902 39506
rect 11954 39454 11966 39506
rect 5630 39442 5682 39454
rect 12798 39442 12850 39454
rect 13470 39506 13522 39518
rect 13470 39442 13522 39454
rect 19294 39506 19346 39518
rect 19294 39442 19346 39454
rect 26574 39506 26626 39518
rect 26574 39442 26626 39454
rect 36206 39506 36258 39518
rect 36206 39442 36258 39454
rect 36990 39506 37042 39518
rect 36990 39442 37042 39454
rect 37102 39506 37154 39518
rect 37102 39442 37154 39454
rect 68462 39506 68514 39518
rect 68462 39442 68514 39454
rect 84142 39506 84194 39518
rect 84142 39442 84194 39454
rect 84254 39506 84306 39518
rect 84254 39442 84306 39454
rect 84814 39506 84866 39518
rect 84814 39442 84866 39454
rect 85934 39506 85986 39518
rect 85934 39442 85986 39454
rect 86382 39506 86434 39518
rect 86382 39442 86434 39454
rect 92094 39506 92146 39518
rect 98018 39454 98030 39506
rect 98082 39454 98094 39506
rect 92094 39442 92146 39454
rect 2046 39394 2098 39406
rect 2046 39330 2098 39342
rect 11230 39394 11282 39406
rect 11230 39330 11282 39342
rect 13806 39394 13858 39406
rect 13806 39330 13858 39342
rect 14142 39394 14194 39406
rect 14142 39330 14194 39342
rect 18622 39394 18674 39406
rect 35870 39394 35922 39406
rect 34290 39342 34302 39394
rect 34354 39342 34366 39394
rect 18622 39330 18674 39342
rect 35870 39330 35922 39342
rect 36318 39394 36370 39406
rect 36318 39330 36370 39342
rect 66110 39394 66162 39406
rect 66110 39330 66162 39342
rect 72718 39394 72770 39406
rect 72718 39330 72770 39342
rect 82686 39394 82738 39406
rect 82686 39330 82738 39342
rect 83470 39394 83522 39406
rect 83470 39330 83522 39342
rect 85822 39394 85874 39406
rect 90302 39394 90354 39406
rect 89506 39342 89518 39394
rect 89570 39342 89582 39394
rect 85822 39330 85874 39342
rect 90302 39330 90354 39342
rect 1344 39226 98560 39260
rect 1344 39174 8896 39226
rect 8948 39174 9020 39226
rect 9072 39174 9144 39226
rect 9196 39174 9268 39226
rect 9320 39174 17896 39226
rect 17948 39174 18020 39226
rect 18072 39174 18144 39226
rect 18196 39174 18268 39226
rect 18320 39174 26896 39226
rect 26948 39174 27020 39226
rect 27072 39174 27144 39226
rect 27196 39174 27268 39226
rect 27320 39174 35896 39226
rect 35948 39174 36020 39226
rect 36072 39174 36144 39226
rect 36196 39174 36268 39226
rect 36320 39174 44896 39226
rect 44948 39174 45020 39226
rect 45072 39174 45144 39226
rect 45196 39174 45268 39226
rect 45320 39174 53896 39226
rect 53948 39174 54020 39226
rect 54072 39174 54144 39226
rect 54196 39174 54268 39226
rect 54320 39174 62896 39226
rect 62948 39174 63020 39226
rect 63072 39174 63144 39226
rect 63196 39174 63268 39226
rect 63320 39174 71896 39226
rect 71948 39174 72020 39226
rect 72072 39174 72144 39226
rect 72196 39174 72268 39226
rect 72320 39174 80896 39226
rect 80948 39174 81020 39226
rect 81072 39174 81144 39226
rect 81196 39174 81268 39226
rect 81320 39174 89896 39226
rect 89948 39174 90020 39226
rect 90072 39174 90144 39226
rect 90196 39174 90268 39226
rect 90320 39174 98560 39226
rect 1344 39140 98560 39174
rect 17502 39058 17554 39070
rect 16258 39006 16270 39058
rect 16322 39006 16334 39058
rect 17502 38994 17554 39006
rect 21086 39058 21138 39070
rect 21086 38994 21138 39006
rect 42142 39058 42194 39070
rect 42142 38994 42194 39006
rect 44494 39058 44546 39070
rect 44494 38994 44546 39006
rect 52894 39058 52946 39070
rect 52894 38994 52946 39006
rect 66670 39058 66722 39070
rect 66670 38994 66722 39006
rect 67118 39058 67170 39070
rect 67118 38994 67170 39006
rect 67902 39058 67954 39070
rect 67902 38994 67954 39006
rect 72494 39058 72546 39070
rect 72494 38994 72546 39006
rect 72942 39058 72994 39070
rect 72942 38994 72994 39006
rect 77310 39058 77362 39070
rect 77310 38994 77362 39006
rect 77870 39058 77922 39070
rect 77870 38994 77922 39006
rect 78542 39058 78594 39070
rect 78542 38994 78594 39006
rect 84366 39058 84418 39070
rect 84366 38994 84418 39006
rect 85262 39058 85314 39070
rect 85262 38994 85314 39006
rect 89742 39058 89794 39070
rect 89742 38994 89794 39006
rect 91982 39058 92034 39070
rect 91982 38994 92034 39006
rect 2382 38946 2434 38958
rect 2382 38882 2434 38894
rect 21646 38946 21698 38958
rect 21646 38882 21698 38894
rect 38558 38946 38610 38958
rect 38558 38882 38610 38894
rect 42590 38946 42642 38958
rect 42590 38882 42642 38894
rect 43822 38946 43874 38958
rect 43822 38882 43874 38894
rect 47742 38946 47794 38958
rect 47742 38882 47794 38894
rect 47966 38946 48018 38958
rect 47966 38882 48018 38894
rect 48078 38946 48130 38958
rect 53230 38946 53282 38958
rect 49298 38894 49310 38946
rect 49362 38894 49374 38946
rect 50530 38894 50542 38946
rect 50594 38894 50606 38946
rect 48078 38882 48130 38894
rect 53230 38882 53282 38894
rect 53902 38946 53954 38958
rect 53902 38882 53954 38894
rect 58382 38946 58434 38958
rect 76414 38946 76466 38958
rect 68002 38894 68014 38946
rect 68066 38894 68078 38946
rect 58382 38882 58434 38894
rect 76414 38882 76466 38894
rect 77534 38946 77586 38958
rect 77534 38882 77586 38894
rect 78990 38946 79042 38958
rect 78990 38882 79042 38894
rect 84702 38946 84754 38958
rect 84702 38882 84754 38894
rect 90190 38946 90242 38958
rect 90962 38894 90974 38946
rect 91026 38894 91038 38946
rect 91298 38894 91310 38946
rect 91362 38894 91374 38946
rect 90190 38882 90242 38894
rect 1822 38834 1874 38846
rect 1822 38770 1874 38782
rect 13358 38834 13410 38846
rect 48302 38834 48354 38846
rect 51886 38834 51938 38846
rect 13794 38782 13806 38834
rect 13858 38782 13870 38834
rect 48738 38782 48750 38834
rect 48802 38782 48814 38834
rect 13358 38770 13410 38782
rect 48302 38770 48354 38782
rect 51886 38770 51938 38782
rect 53566 38834 53618 38846
rect 53566 38770 53618 38782
rect 60174 38834 60226 38846
rect 60174 38770 60226 38782
rect 67790 38834 67842 38846
rect 77198 38834 77250 38846
rect 68338 38782 68350 38834
rect 68402 38782 68414 38834
rect 69010 38782 69022 38834
rect 69074 38782 69086 38834
rect 74834 38782 74846 38834
rect 74898 38782 74910 38834
rect 67790 38770 67842 38782
rect 77198 38770 77250 38782
rect 91646 38834 91698 38846
rect 91646 38770 91698 38782
rect 16830 38722 16882 38734
rect 16830 38658 16882 38670
rect 28814 38722 28866 38734
rect 28814 38658 28866 38670
rect 52446 38722 52498 38734
rect 52446 38658 52498 38670
rect 76862 38722 76914 38734
rect 76862 38658 76914 38670
rect 83694 38722 83746 38734
rect 83694 38658 83746 38670
rect 85710 38722 85762 38734
rect 85710 38658 85762 38670
rect 50094 38610 50146 38622
rect 50094 38546 50146 38558
rect 75294 38610 75346 38622
rect 83682 38558 83694 38610
rect 83746 38607 83758 38610
rect 84130 38607 84142 38610
rect 83746 38561 84142 38607
rect 83746 38558 83758 38561
rect 84130 38558 84142 38561
rect 84194 38558 84206 38610
rect 75294 38546 75346 38558
rect 1344 38442 98560 38476
rect 1344 38390 4396 38442
rect 4448 38390 4520 38442
rect 4572 38390 4644 38442
rect 4696 38390 4768 38442
rect 4820 38390 13396 38442
rect 13448 38390 13520 38442
rect 13572 38390 13644 38442
rect 13696 38390 13768 38442
rect 13820 38390 22396 38442
rect 22448 38390 22520 38442
rect 22572 38390 22644 38442
rect 22696 38390 22768 38442
rect 22820 38390 31396 38442
rect 31448 38390 31520 38442
rect 31572 38390 31644 38442
rect 31696 38390 31768 38442
rect 31820 38390 40396 38442
rect 40448 38390 40520 38442
rect 40572 38390 40644 38442
rect 40696 38390 40768 38442
rect 40820 38390 49396 38442
rect 49448 38390 49520 38442
rect 49572 38390 49644 38442
rect 49696 38390 49768 38442
rect 49820 38390 58396 38442
rect 58448 38390 58520 38442
rect 58572 38390 58644 38442
rect 58696 38390 58768 38442
rect 58820 38390 67396 38442
rect 67448 38390 67520 38442
rect 67572 38390 67644 38442
rect 67696 38390 67768 38442
rect 67820 38390 76396 38442
rect 76448 38390 76520 38442
rect 76572 38390 76644 38442
rect 76696 38390 76768 38442
rect 76820 38390 85396 38442
rect 85448 38390 85520 38442
rect 85572 38390 85644 38442
rect 85696 38390 85768 38442
rect 85820 38390 94396 38442
rect 94448 38390 94520 38442
rect 94572 38390 94644 38442
rect 94696 38390 94768 38442
rect 94820 38390 98560 38442
rect 1344 38356 98560 38390
rect 42030 38274 42082 38286
rect 42030 38210 42082 38222
rect 45278 38274 45330 38286
rect 60958 38274 61010 38286
rect 46386 38222 46398 38274
rect 46450 38271 46462 38274
rect 46722 38271 46734 38274
rect 46450 38225 46734 38271
rect 46450 38222 46462 38225
rect 46722 38222 46734 38225
rect 46786 38222 46798 38274
rect 45278 38210 45330 38222
rect 60958 38210 61010 38222
rect 76078 38274 76130 38286
rect 76078 38210 76130 38222
rect 33406 38162 33458 38174
rect 56702 38162 56754 38174
rect 75406 38162 75458 38174
rect 51538 38110 51550 38162
rect 51602 38110 51614 38162
rect 67666 38110 67678 38162
rect 67730 38110 67742 38162
rect 68786 38110 68798 38162
rect 68850 38110 68862 38162
rect 33406 38098 33458 38110
rect 56702 38098 56754 38110
rect 75406 38098 75458 38110
rect 87166 38162 87218 38174
rect 87166 38098 87218 38110
rect 21534 38050 21586 38062
rect 27694 38050 27746 38062
rect 34302 38050 34354 38062
rect 38558 38050 38610 38062
rect 52670 38050 52722 38062
rect 63310 38050 63362 38062
rect 68574 38050 68626 38062
rect 73166 38050 73218 38062
rect 20514 37998 20526 38050
rect 20578 37998 20590 38050
rect 21858 37998 21870 38050
rect 21922 37998 21934 38050
rect 28354 37998 28366 38050
rect 28418 37998 28430 38050
rect 35074 37998 35086 38050
rect 35138 37998 35150 38050
rect 38994 37998 39006 38050
rect 39058 37998 39070 38050
rect 42354 37998 42366 38050
rect 42418 37998 42430 38050
rect 45938 37998 45950 38050
rect 46002 37998 46014 38050
rect 48178 37998 48190 38050
rect 48242 37998 48254 38050
rect 49746 37998 49758 38050
rect 49810 37998 49822 38050
rect 53218 37998 53230 38050
rect 53282 37998 53294 38050
rect 63970 37998 63982 38050
rect 64034 37998 64046 38050
rect 72482 37998 72494 38050
rect 72546 37998 72558 38050
rect 21534 37986 21586 37998
rect 27694 37986 27746 37998
rect 34302 37986 34354 37998
rect 38558 37986 38610 37998
rect 52670 37986 52722 37998
rect 63310 37986 63362 37998
rect 68574 37986 68626 37998
rect 73166 37986 73218 37998
rect 73502 38050 73554 38062
rect 84926 38050 84978 38062
rect 73938 37998 73950 38050
rect 74002 37998 74014 38050
rect 76178 37998 76190 38050
rect 76242 37998 76254 38050
rect 76962 37998 76974 38050
rect 77026 37998 77038 38050
rect 77410 37998 77422 38050
rect 77474 37998 77486 38050
rect 78306 37998 78318 38050
rect 78370 37998 78382 38050
rect 78866 37998 78878 38050
rect 78930 37998 78942 38050
rect 79314 37998 79326 38050
rect 79378 37998 79390 38050
rect 73502 37986 73554 37998
rect 84926 37986 84978 37998
rect 85150 38050 85202 38062
rect 87490 37998 87502 38050
rect 87554 37998 87566 38050
rect 85150 37986 85202 37998
rect 1710 37938 1762 37950
rect 1710 37874 1762 37886
rect 20750 37938 20802 37950
rect 32958 37938 33010 37950
rect 36990 37938 37042 37950
rect 44270 37938 44322 37950
rect 28466 37886 28478 37938
rect 28530 37886 28542 37938
rect 34850 37886 34862 37938
rect 34914 37886 34926 37938
rect 43362 37886 43374 37938
rect 43426 37886 43438 37938
rect 20750 37874 20802 37886
rect 32958 37874 33010 37886
rect 36990 37874 37042 37886
rect 44270 37874 44322 37886
rect 44942 37938 44994 37950
rect 59278 37938 59330 37950
rect 46050 37886 46062 37938
rect 46114 37886 46126 37938
rect 48962 37886 48974 37938
rect 49026 37886 49038 37938
rect 49970 37886 49982 37938
rect 50034 37886 50046 37938
rect 44942 37874 44994 37886
rect 59278 37874 59330 37886
rect 60622 37938 60674 37950
rect 63086 37938 63138 37950
rect 61170 37886 61182 37938
rect 61234 37886 61246 37938
rect 61730 37886 61742 37938
rect 61794 37886 61806 37938
rect 60622 37874 60674 37886
rect 63086 37874 63138 37886
rect 68350 37938 68402 37950
rect 78542 37938 78594 37950
rect 74274 37886 74286 37938
rect 74338 37886 74350 37938
rect 76290 37886 76302 37938
rect 76354 37886 76366 37938
rect 68350 37874 68402 37886
rect 78542 37874 78594 37886
rect 81678 37938 81730 37950
rect 81678 37874 81730 37886
rect 85486 37938 85538 37950
rect 85486 37874 85538 37886
rect 96238 37938 96290 37950
rect 96238 37874 96290 37886
rect 96574 37938 96626 37950
rect 96574 37874 96626 37886
rect 2046 37826 2098 37838
rect 2046 37762 2098 37774
rect 2494 37826 2546 37838
rect 2494 37762 2546 37774
rect 5966 37826 6018 37838
rect 25006 37826 25058 37838
rect 24210 37774 24222 37826
rect 24274 37774 24286 37826
rect 5966 37762 6018 37774
rect 25006 37762 25058 37774
rect 26350 37826 26402 37838
rect 26350 37762 26402 37774
rect 27358 37826 27410 37838
rect 27358 37762 27410 37774
rect 29598 37826 29650 37838
rect 29598 37762 29650 37774
rect 30046 37826 30098 37838
rect 30046 37762 30098 37774
rect 33966 37826 34018 37838
rect 33966 37762 34018 37774
rect 35646 37826 35698 37838
rect 35646 37762 35698 37774
rect 37102 37826 37154 37838
rect 37102 37762 37154 37774
rect 37326 37826 37378 37838
rect 43934 37826 43986 37838
rect 41458 37774 41470 37826
rect 41522 37774 41534 37826
rect 37326 37762 37378 37774
rect 43934 37762 43986 37774
rect 46622 37826 46674 37838
rect 56366 37826 56418 37838
rect 55794 37774 55806 37826
rect 55858 37774 55870 37826
rect 46622 37762 46674 37774
rect 56366 37762 56418 37774
rect 58942 37826 58994 37838
rect 58942 37762 58994 37774
rect 59950 37826 60002 37838
rect 67006 37826 67058 37838
rect 66434 37774 66446 37826
rect 66498 37774 66510 37826
rect 59950 37762 60002 37774
rect 67006 37762 67058 37774
rect 67230 37826 67282 37838
rect 67230 37762 67282 37774
rect 68798 37826 68850 37838
rect 68798 37762 68850 37774
rect 68910 37826 68962 37838
rect 68910 37762 68962 37774
rect 71934 37826 71986 37838
rect 71934 37762 71986 37774
rect 72718 37826 72770 37838
rect 72718 37762 72770 37774
rect 74958 37826 75010 37838
rect 74958 37762 75010 37774
rect 82462 37826 82514 37838
rect 82462 37762 82514 37774
rect 83470 37826 83522 37838
rect 83470 37762 83522 37774
rect 84254 37826 84306 37838
rect 84254 37762 84306 37774
rect 84366 37826 84418 37838
rect 84366 37762 84418 37774
rect 84478 37826 84530 37838
rect 84478 37762 84530 37774
rect 85374 37826 85426 37838
rect 85374 37762 85426 37774
rect 85934 37826 85986 37838
rect 85934 37762 85986 37774
rect 88062 37826 88114 37838
rect 88062 37762 88114 37774
rect 1344 37658 98560 37692
rect 1344 37606 8896 37658
rect 8948 37606 9020 37658
rect 9072 37606 9144 37658
rect 9196 37606 9268 37658
rect 9320 37606 17896 37658
rect 17948 37606 18020 37658
rect 18072 37606 18144 37658
rect 18196 37606 18268 37658
rect 18320 37606 26896 37658
rect 26948 37606 27020 37658
rect 27072 37606 27144 37658
rect 27196 37606 27268 37658
rect 27320 37606 35896 37658
rect 35948 37606 36020 37658
rect 36072 37606 36144 37658
rect 36196 37606 36268 37658
rect 36320 37606 44896 37658
rect 44948 37606 45020 37658
rect 45072 37606 45144 37658
rect 45196 37606 45268 37658
rect 45320 37606 53896 37658
rect 53948 37606 54020 37658
rect 54072 37606 54144 37658
rect 54196 37606 54268 37658
rect 54320 37606 62896 37658
rect 62948 37606 63020 37658
rect 63072 37606 63144 37658
rect 63196 37606 63268 37658
rect 63320 37606 71896 37658
rect 71948 37606 72020 37658
rect 72072 37606 72144 37658
rect 72196 37606 72268 37658
rect 72320 37606 80896 37658
rect 80948 37606 81020 37658
rect 81072 37606 81144 37658
rect 81196 37606 81268 37658
rect 81320 37606 89896 37658
rect 89948 37606 90020 37658
rect 90072 37606 90144 37658
rect 90196 37606 90268 37658
rect 90320 37606 98560 37658
rect 1344 37572 98560 37606
rect 18398 37490 18450 37502
rect 18398 37426 18450 37438
rect 20190 37490 20242 37502
rect 20190 37426 20242 37438
rect 21646 37490 21698 37502
rect 39454 37490 39506 37502
rect 29138 37438 29150 37490
rect 29202 37438 29214 37490
rect 38546 37438 38558 37490
rect 38610 37438 38622 37490
rect 21646 37426 21698 37438
rect 39454 37426 39506 37438
rect 40462 37490 40514 37502
rect 40462 37426 40514 37438
rect 47182 37490 47234 37502
rect 53678 37490 53730 37502
rect 49858 37438 49870 37490
rect 49922 37438 49934 37490
rect 52098 37438 52110 37490
rect 52162 37438 52174 37490
rect 47182 37426 47234 37438
rect 53678 37426 53730 37438
rect 55358 37490 55410 37502
rect 55358 37426 55410 37438
rect 57934 37490 57986 37502
rect 61742 37490 61794 37502
rect 60946 37438 60958 37490
rect 61010 37438 61022 37490
rect 57934 37426 57986 37438
rect 61742 37426 61794 37438
rect 63870 37490 63922 37502
rect 63870 37426 63922 37438
rect 64430 37490 64482 37502
rect 64430 37426 64482 37438
rect 67790 37490 67842 37502
rect 67790 37426 67842 37438
rect 68238 37490 68290 37502
rect 75854 37490 75906 37502
rect 75282 37438 75294 37490
rect 75346 37438 75358 37490
rect 68238 37426 68290 37438
rect 75854 37426 75906 37438
rect 76862 37490 76914 37502
rect 76862 37426 76914 37438
rect 78654 37490 78706 37502
rect 88062 37490 88114 37502
rect 86818 37438 86830 37490
rect 86882 37438 86894 37490
rect 78654 37426 78706 37438
rect 88062 37426 88114 37438
rect 96462 37490 96514 37502
rect 96462 37426 96514 37438
rect 5070 37378 5122 37390
rect 5070 37314 5122 37326
rect 5854 37378 5906 37390
rect 5854 37314 5906 37326
rect 6078 37378 6130 37390
rect 6078 37314 6130 37326
rect 8318 37378 8370 37390
rect 8318 37314 8370 37326
rect 8654 37378 8706 37390
rect 8654 37314 8706 37326
rect 8990 37378 9042 37390
rect 8990 37314 9042 37326
rect 9662 37378 9714 37390
rect 15262 37378 15314 37390
rect 31726 37378 31778 37390
rect 10210 37326 10222 37378
rect 10274 37326 10286 37378
rect 10546 37326 10558 37378
rect 10610 37326 10622 37378
rect 20626 37326 20638 37378
rect 20690 37326 20702 37378
rect 9662 37314 9714 37326
rect 15262 37314 15314 37326
rect 31726 37314 31778 37326
rect 33070 37378 33122 37390
rect 33070 37314 33122 37326
rect 33406 37378 33458 37390
rect 43374 37378 43426 37390
rect 36866 37326 36878 37378
rect 36930 37326 36942 37378
rect 37986 37326 37998 37378
rect 38050 37326 38062 37378
rect 41906 37326 41918 37378
rect 41970 37326 41982 37378
rect 33406 37314 33458 37326
rect 43374 37314 43426 37326
rect 46398 37378 46450 37390
rect 46398 37314 46450 37326
rect 50654 37378 50706 37390
rect 90414 37378 90466 37390
rect 54226 37326 54238 37378
rect 54290 37326 54302 37378
rect 54562 37326 54574 37378
rect 54626 37326 54638 37378
rect 66322 37326 66334 37378
rect 66386 37326 66398 37378
rect 77634 37326 77646 37378
rect 77698 37326 77710 37378
rect 50654 37314 50706 37326
rect 90414 37314 90466 37326
rect 2382 37266 2434 37278
rect 15598 37266 15650 37278
rect 21310 37266 21362 37278
rect 2706 37214 2718 37266
rect 2770 37214 2782 37266
rect 6514 37214 6526 37266
rect 6578 37214 6590 37266
rect 20514 37214 20526 37266
rect 20578 37214 20590 37266
rect 2382 37202 2434 37214
rect 15598 37202 15650 37214
rect 21310 37202 21362 37214
rect 26238 37266 26290 37278
rect 29710 37266 29762 37278
rect 39790 37266 39842 37278
rect 26674 37214 26686 37266
rect 26738 37214 26750 37266
rect 29922 37214 29934 37266
rect 29986 37214 29998 37266
rect 34850 37214 34862 37266
rect 34914 37214 34926 37266
rect 35074 37214 35086 37266
rect 35138 37214 35150 37266
rect 35746 37214 35758 37266
rect 35810 37214 35822 37266
rect 38322 37214 38334 37266
rect 38386 37214 38398 37266
rect 26238 37202 26290 37214
rect 29710 37202 29762 37214
rect 39790 37202 39842 37214
rect 41022 37266 41074 37278
rect 41022 37202 41074 37214
rect 41358 37266 41410 37278
rect 50206 37266 50258 37278
rect 42018 37214 42030 37266
rect 42082 37214 42094 37266
rect 43586 37214 43598 37266
rect 43650 37214 43662 37266
rect 44034 37214 44046 37266
rect 44098 37214 44110 37266
rect 41358 37202 41410 37214
rect 50206 37202 50258 37214
rect 50430 37266 50482 37278
rect 64766 37266 64818 37278
rect 51538 37214 51550 37266
rect 51602 37214 51614 37266
rect 58146 37214 58158 37266
rect 58210 37214 58222 37266
rect 58706 37214 58718 37266
rect 58770 37214 58782 37266
rect 50430 37202 50482 37214
rect 64766 37202 64818 37214
rect 65214 37266 65266 37278
rect 65214 37202 65266 37214
rect 65550 37266 65602 37278
rect 72382 37266 72434 37278
rect 78318 37266 78370 37278
rect 96126 37266 96178 37278
rect 66098 37214 66110 37266
rect 66162 37214 66174 37266
rect 72706 37214 72718 37266
rect 72770 37214 72782 37266
rect 77522 37214 77534 37266
rect 77586 37214 77598 37266
rect 83906 37214 83918 37266
rect 83970 37214 83982 37266
rect 84354 37214 84366 37266
rect 84418 37214 84430 37266
rect 96898 37214 96910 37266
rect 96962 37214 96974 37266
rect 65550 37202 65602 37214
rect 72382 37202 72434 37214
rect 78318 37202 78370 37214
rect 96126 37202 96178 37214
rect 1822 37154 1874 37166
rect 1822 37090 1874 37102
rect 7086 37154 7138 37166
rect 7086 37090 7138 37102
rect 11342 37154 11394 37166
rect 11342 37090 11394 37102
rect 11902 37154 11954 37166
rect 11902 37090 11954 37102
rect 19630 37154 19682 37166
rect 19630 37090 19682 37102
rect 39118 37154 39170 37166
rect 39118 37090 39170 37102
rect 42702 37154 42754 37166
rect 42702 37090 42754 37102
rect 48974 37154 49026 37166
rect 48974 37090 49026 37102
rect 49422 37154 49474 37166
rect 49422 37090 49474 37102
rect 51214 37154 51266 37166
rect 51214 37090 51266 37102
rect 54014 37154 54066 37166
rect 54014 37090 54066 37102
rect 66894 37154 66946 37166
rect 66894 37090 66946 37102
rect 76190 37154 76242 37166
rect 98018 37102 98030 37154
rect 98082 37102 98094 37154
rect 76190 37090 76242 37102
rect 9998 37042 10050 37054
rect 9998 36978 10050 36990
rect 30942 37042 30994 37054
rect 30942 36978 30994 36990
rect 87502 37042 87554 37054
rect 87502 36978 87554 36990
rect 1344 36874 98560 36908
rect 1344 36822 4396 36874
rect 4448 36822 4520 36874
rect 4572 36822 4644 36874
rect 4696 36822 4768 36874
rect 4820 36822 13396 36874
rect 13448 36822 13520 36874
rect 13572 36822 13644 36874
rect 13696 36822 13768 36874
rect 13820 36822 22396 36874
rect 22448 36822 22520 36874
rect 22572 36822 22644 36874
rect 22696 36822 22768 36874
rect 22820 36822 31396 36874
rect 31448 36822 31520 36874
rect 31572 36822 31644 36874
rect 31696 36822 31768 36874
rect 31820 36822 40396 36874
rect 40448 36822 40520 36874
rect 40572 36822 40644 36874
rect 40696 36822 40768 36874
rect 40820 36822 49396 36874
rect 49448 36822 49520 36874
rect 49572 36822 49644 36874
rect 49696 36822 49768 36874
rect 49820 36822 58396 36874
rect 58448 36822 58520 36874
rect 58572 36822 58644 36874
rect 58696 36822 58768 36874
rect 58820 36822 67396 36874
rect 67448 36822 67520 36874
rect 67572 36822 67644 36874
rect 67696 36822 67768 36874
rect 67820 36822 76396 36874
rect 76448 36822 76520 36874
rect 76572 36822 76644 36874
rect 76696 36822 76768 36874
rect 76820 36822 85396 36874
rect 85448 36822 85520 36874
rect 85572 36822 85644 36874
rect 85696 36822 85768 36874
rect 85820 36822 94396 36874
rect 94448 36822 94520 36874
rect 94572 36822 94644 36874
rect 94696 36822 94768 36874
rect 94820 36822 98560 36874
rect 1344 36788 98560 36822
rect 18958 36706 19010 36718
rect 18958 36642 19010 36654
rect 35086 36706 35138 36718
rect 35086 36642 35138 36654
rect 53342 36706 53394 36718
rect 53342 36642 53394 36654
rect 3278 36594 3330 36606
rect 3278 36530 3330 36542
rect 7310 36594 7362 36606
rect 50878 36594 50930 36606
rect 46946 36542 46958 36594
rect 47010 36542 47022 36594
rect 7310 36530 7362 36542
rect 50878 36530 50930 36542
rect 51998 36594 52050 36606
rect 51998 36530 52050 36542
rect 56814 36594 56866 36606
rect 56814 36530 56866 36542
rect 64878 36594 64930 36606
rect 64878 36530 64930 36542
rect 67454 36594 67506 36606
rect 67454 36530 67506 36542
rect 68798 36594 68850 36606
rect 68798 36530 68850 36542
rect 77198 36594 77250 36606
rect 77198 36530 77250 36542
rect 1710 36482 1762 36494
rect 8654 36482 8706 36494
rect 12350 36482 12402 36494
rect 6738 36430 6750 36482
rect 6802 36430 6814 36482
rect 9202 36430 9214 36482
rect 9266 36430 9278 36482
rect 1710 36418 1762 36430
rect 8654 36418 8706 36430
rect 12350 36418 12402 36430
rect 14814 36482 14866 36494
rect 27470 36482 27522 36494
rect 15362 36430 15374 36482
rect 15426 36430 15438 36482
rect 19730 36430 19742 36482
rect 19794 36430 19806 36482
rect 14814 36418 14866 36430
rect 27470 36418 27522 36430
rect 31614 36482 31666 36494
rect 37326 36482 37378 36494
rect 51550 36482 51602 36494
rect 32050 36430 32062 36482
rect 32114 36430 32126 36482
rect 47730 36430 47742 36482
rect 47794 36430 47806 36482
rect 31614 36418 31666 36430
rect 37326 36418 37378 36430
rect 51550 36418 51602 36430
rect 52782 36482 52834 36494
rect 52782 36418 52834 36430
rect 53006 36482 53058 36494
rect 53006 36418 53058 36430
rect 53230 36482 53282 36494
rect 92206 36482 92258 36494
rect 69458 36430 69470 36482
rect 69522 36430 69534 36482
rect 53230 36418 53282 36430
rect 92206 36418 92258 36430
rect 92430 36482 92482 36494
rect 92430 36418 92482 36430
rect 14590 36370 14642 36382
rect 14590 36306 14642 36318
rect 17726 36370 17778 36382
rect 17726 36306 17778 36318
rect 18510 36370 18562 36382
rect 18510 36306 18562 36318
rect 27134 36370 27186 36382
rect 27134 36306 27186 36318
rect 36990 36370 37042 36382
rect 36990 36306 37042 36318
rect 37102 36370 37154 36382
rect 37102 36306 37154 36318
rect 37662 36370 37714 36382
rect 37662 36306 37714 36318
rect 46734 36370 46786 36382
rect 46734 36306 46786 36318
rect 53454 36370 53506 36382
rect 53454 36306 53506 36318
rect 67790 36370 67842 36382
rect 90526 36370 90578 36382
rect 69570 36318 69582 36370
rect 69634 36318 69646 36370
rect 67790 36306 67842 36318
rect 90526 36306 90578 36318
rect 96238 36370 96290 36382
rect 96238 36306 96290 36318
rect 96574 36370 96626 36382
rect 96574 36306 96626 36318
rect 2046 36258 2098 36270
rect 2046 36194 2098 36206
rect 2718 36258 2770 36270
rect 2718 36194 2770 36206
rect 6302 36258 6354 36270
rect 6302 36194 6354 36206
rect 8430 36258 8482 36270
rect 21310 36258 21362 36270
rect 11554 36206 11566 36258
rect 11618 36206 11630 36258
rect 8430 36194 8482 36206
rect 21310 36194 21362 36206
rect 29822 36258 29874 36270
rect 29822 36194 29874 36206
rect 31166 36258 31218 36270
rect 38894 36258 38946 36270
rect 34290 36206 34302 36258
rect 34354 36206 34366 36258
rect 31166 36194 31218 36206
rect 38894 36194 38946 36206
rect 45950 36258 46002 36270
rect 45950 36194 46002 36206
rect 46398 36258 46450 36270
rect 46398 36194 46450 36206
rect 48414 36258 48466 36270
rect 48414 36194 48466 36206
rect 48974 36258 49026 36270
rect 48974 36194 49026 36206
rect 53902 36258 53954 36270
rect 53902 36194 53954 36206
rect 68462 36258 68514 36270
rect 68462 36194 68514 36206
rect 78990 36258 79042 36270
rect 78990 36194 79042 36206
rect 90862 36258 90914 36270
rect 90862 36194 90914 36206
rect 91310 36258 91362 36270
rect 91858 36206 91870 36258
rect 91922 36206 91934 36258
rect 91310 36194 91362 36206
rect 1344 36090 98560 36124
rect 1344 36038 8896 36090
rect 8948 36038 9020 36090
rect 9072 36038 9144 36090
rect 9196 36038 9268 36090
rect 9320 36038 17896 36090
rect 17948 36038 18020 36090
rect 18072 36038 18144 36090
rect 18196 36038 18268 36090
rect 18320 36038 26896 36090
rect 26948 36038 27020 36090
rect 27072 36038 27144 36090
rect 27196 36038 27268 36090
rect 27320 36038 35896 36090
rect 35948 36038 36020 36090
rect 36072 36038 36144 36090
rect 36196 36038 36268 36090
rect 36320 36038 44896 36090
rect 44948 36038 45020 36090
rect 45072 36038 45144 36090
rect 45196 36038 45268 36090
rect 45320 36038 53896 36090
rect 53948 36038 54020 36090
rect 54072 36038 54144 36090
rect 54196 36038 54268 36090
rect 54320 36038 62896 36090
rect 62948 36038 63020 36090
rect 63072 36038 63144 36090
rect 63196 36038 63268 36090
rect 63320 36038 71896 36090
rect 71948 36038 72020 36090
rect 72072 36038 72144 36090
rect 72196 36038 72268 36090
rect 72320 36038 80896 36090
rect 80948 36038 81020 36090
rect 81072 36038 81144 36090
rect 81196 36038 81268 36090
rect 81320 36038 89896 36090
rect 89948 36038 90020 36090
rect 90072 36038 90144 36090
rect 90196 36038 90268 36090
rect 90320 36038 98560 36090
rect 1344 36004 98560 36038
rect 6638 35922 6690 35934
rect 5618 35870 5630 35922
rect 5682 35870 5694 35922
rect 6638 35858 6690 35870
rect 16494 35922 16546 35934
rect 16494 35858 16546 35870
rect 17502 35922 17554 35934
rect 17502 35858 17554 35870
rect 18622 35922 18674 35934
rect 18622 35858 18674 35870
rect 19742 35922 19794 35934
rect 19742 35858 19794 35870
rect 36766 35922 36818 35934
rect 36766 35858 36818 35870
rect 37326 35922 37378 35934
rect 37326 35858 37378 35870
rect 38670 35922 38722 35934
rect 38670 35858 38722 35870
rect 39118 35922 39170 35934
rect 39118 35858 39170 35870
rect 52446 35922 52498 35934
rect 57374 35922 57426 35934
rect 57138 35870 57150 35922
rect 57202 35870 57214 35922
rect 77982 35922 78034 35934
rect 52446 35858 52498 35870
rect 57374 35858 57426 35870
rect 68350 35866 68402 35878
rect 2046 35810 2098 35822
rect 22094 35810 22146 35822
rect 15474 35758 15486 35810
rect 15538 35758 15550 35810
rect 20290 35758 20302 35810
rect 20354 35758 20366 35810
rect 2046 35746 2098 35758
rect 22094 35746 22146 35758
rect 39566 35810 39618 35822
rect 39566 35746 39618 35758
rect 46510 35810 46562 35822
rect 53342 35810 53394 35822
rect 62974 35810 63026 35822
rect 47730 35758 47742 35810
rect 47794 35758 47806 35810
rect 49746 35758 49758 35810
rect 49810 35758 49822 35810
rect 53554 35758 53566 35810
rect 53618 35758 53630 35810
rect 77982 35858 78034 35870
rect 78206 35922 78258 35934
rect 78206 35858 78258 35870
rect 78430 35922 78482 35934
rect 78430 35858 78482 35870
rect 84254 35922 84306 35934
rect 84254 35858 84306 35870
rect 84590 35922 84642 35934
rect 93774 35922 93826 35934
rect 89842 35870 89854 35922
rect 89906 35870 89918 35922
rect 92978 35870 92990 35922
rect 93042 35870 93054 35922
rect 84590 35858 84642 35870
rect 93774 35858 93826 35870
rect 68350 35802 68402 35814
rect 68686 35810 68738 35822
rect 46510 35746 46562 35758
rect 53342 35746 53394 35758
rect 62974 35746 63026 35758
rect 68686 35746 68738 35758
rect 72382 35810 72434 35822
rect 72382 35746 72434 35758
rect 79102 35810 79154 35822
rect 79102 35746 79154 35758
rect 80222 35810 80274 35822
rect 80222 35746 80274 35758
rect 85486 35810 85538 35822
rect 85486 35746 85538 35758
rect 89294 35810 89346 35822
rect 89294 35746 89346 35758
rect 1710 35698 1762 35710
rect 1710 35634 1762 35646
rect 2718 35698 2770 35710
rect 6190 35698 6242 35710
rect 16158 35698 16210 35710
rect 21310 35698 21362 35710
rect 3042 35646 3054 35698
rect 3106 35646 3118 35698
rect 15362 35646 15374 35698
rect 15426 35646 15438 35698
rect 20178 35646 20190 35698
rect 20242 35646 20254 35698
rect 2718 35634 2770 35646
rect 6190 35634 6242 35646
rect 16158 35634 16210 35646
rect 21310 35634 21362 35646
rect 21758 35698 21810 35710
rect 21758 35634 21810 35646
rect 36654 35698 36706 35710
rect 36654 35634 36706 35646
rect 39006 35698 39058 35710
rect 39006 35634 39058 35646
rect 39342 35698 39394 35710
rect 53118 35698 53170 35710
rect 56030 35698 56082 35710
rect 47170 35646 47182 35698
rect 47234 35646 47246 35698
rect 48962 35646 48974 35698
rect 49026 35646 49038 35698
rect 53778 35646 53790 35698
rect 53842 35646 53854 35698
rect 39342 35634 39394 35646
rect 53118 35634 53170 35646
rect 56030 35634 56082 35646
rect 57150 35698 57202 35710
rect 57150 35634 57202 35646
rect 57598 35698 57650 35710
rect 57598 35634 57650 35646
rect 57822 35698 57874 35710
rect 57822 35634 57874 35646
rect 62638 35698 62690 35710
rect 78878 35698 78930 35710
rect 68114 35646 68126 35698
rect 68178 35646 68190 35698
rect 62638 35634 62690 35646
rect 78878 35634 78930 35646
rect 79998 35698 80050 35710
rect 79998 35634 80050 35646
rect 80334 35698 80386 35710
rect 80334 35634 80386 35646
rect 84702 35698 84754 35710
rect 84702 35634 84754 35646
rect 84814 35698 84866 35710
rect 84814 35634 84866 35646
rect 85262 35698 85314 35710
rect 85262 35634 85314 35646
rect 86046 35698 86098 35710
rect 86046 35634 86098 35646
rect 90302 35698 90354 35710
rect 96910 35698 96962 35710
rect 90738 35646 90750 35698
rect 90802 35646 90814 35698
rect 90302 35634 90354 35646
rect 96910 35634 96962 35646
rect 14926 35586 14978 35598
rect 14926 35522 14978 35534
rect 36206 35586 36258 35598
rect 36206 35522 36258 35534
rect 45054 35586 45106 35598
rect 45502 35586 45554 35598
rect 45378 35534 45390 35586
rect 45442 35534 45454 35586
rect 45054 35522 45106 35534
rect 20974 35474 21026 35486
rect 20974 35410 21026 35422
rect 36766 35474 36818 35486
rect 45393 35471 45439 35534
rect 45502 35522 45554 35534
rect 45950 35586 46002 35598
rect 45950 35522 46002 35534
rect 56702 35586 56754 35598
rect 56702 35522 56754 35534
rect 78318 35586 78370 35598
rect 78318 35522 78370 35534
rect 80782 35586 80834 35598
rect 80782 35522 80834 35534
rect 89070 35586 89122 35598
rect 89070 35522 89122 35534
rect 46286 35474 46338 35486
rect 45938 35471 45950 35474
rect 45393 35425 45950 35471
rect 45938 35422 45950 35425
rect 46002 35422 46014 35474
rect 36766 35410 36818 35422
rect 46286 35410 46338 35422
rect 46622 35474 46674 35486
rect 46622 35410 46674 35422
rect 54126 35474 54178 35486
rect 54126 35410 54178 35422
rect 89518 35474 89570 35486
rect 89518 35410 89570 35422
rect 97694 35474 97746 35486
rect 97694 35410 97746 35422
rect 1344 35306 98560 35340
rect 1344 35254 4396 35306
rect 4448 35254 4520 35306
rect 4572 35254 4644 35306
rect 4696 35254 4768 35306
rect 4820 35254 13396 35306
rect 13448 35254 13520 35306
rect 13572 35254 13644 35306
rect 13696 35254 13768 35306
rect 13820 35254 22396 35306
rect 22448 35254 22520 35306
rect 22572 35254 22644 35306
rect 22696 35254 22768 35306
rect 22820 35254 31396 35306
rect 31448 35254 31520 35306
rect 31572 35254 31644 35306
rect 31696 35254 31768 35306
rect 31820 35254 40396 35306
rect 40448 35254 40520 35306
rect 40572 35254 40644 35306
rect 40696 35254 40768 35306
rect 40820 35254 49396 35306
rect 49448 35254 49520 35306
rect 49572 35254 49644 35306
rect 49696 35254 49768 35306
rect 49820 35254 58396 35306
rect 58448 35254 58520 35306
rect 58572 35254 58644 35306
rect 58696 35254 58768 35306
rect 58820 35254 67396 35306
rect 67448 35254 67520 35306
rect 67572 35254 67644 35306
rect 67696 35254 67768 35306
rect 67820 35254 76396 35306
rect 76448 35254 76520 35306
rect 76572 35254 76644 35306
rect 76696 35254 76768 35306
rect 76820 35254 85396 35306
rect 85448 35254 85520 35306
rect 85572 35254 85644 35306
rect 85696 35254 85768 35306
rect 85820 35254 94396 35306
rect 94448 35254 94520 35306
rect 94572 35254 94644 35306
rect 94696 35254 94768 35306
rect 94820 35254 98560 35306
rect 1344 35220 98560 35254
rect 44046 35138 44098 35150
rect 44046 35074 44098 35086
rect 52782 35138 52834 35150
rect 52782 35074 52834 35086
rect 71934 35138 71986 35150
rect 71934 35074 71986 35086
rect 81566 35138 81618 35150
rect 81566 35074 81618 35086
rect 20750 35026 20802 35038
rect 20750 34962 20802 34974
rect 35310 35026 35362 35038
rect 35310 34962 35362 34974
rect 39006 35026 39058 35038
rect 39006 34962 39058 34974
rect 51662 35026 51714 35038
rect 51662 34962 51714 34974
rect 52110 35026 52162 35038
rect 52110 34962 52162 34974
rect 89966 35026 90018 35038
rect 89966 34962 90018 34974
rect 5518 34914 5570 34926
rect 21198 34914 21250 34926
rect 35870 34914 35922 34926
rect 6066 34862 6078 34914
rect 6130 34862 6142 34914
rect 21858 34862 21870 34914
rect 21922 34862 21934 34914
rect 5518 34850 5570 34862
rect 21198 34850 21250 34862
rect 35870 34850 35922 34862
rect 38670 34914 38722 34926
rect 38670 34850 38722 34862
rect 39118 34914 39170 34926
rect 52558 34914 52610 34926
rect 45490 34862 45502 34914
rect 45554 34862 45566 34914
rect 46050 34862 46062 34914
rect 46114 34862 46126 34914
rect 47282 34862 47294 34914
rect 47346 34862 47358 34914
rect 51090 34862 51102 34914
rect 51154 34862 51166 34914
rect 39118 34850 39170 34862
rect 52558 34850 52610 34862
rect 55246 34914 55298 34926
rect 58942 34914 58994 34926
rect 55794 34862 55806 34914
rect 55858 34862 55870 34914
rect 55246 34850 55298 34862
rect 58942 34850 58994 34862
rect 61630 34914 61682 34926
rect 68462 34914 68514 34926
rect 78094 34914 78146 34926
rect 61954 34862 61966 34914
rect 62018 34862 62030 34914
rect 68898 34862 68910 34914
rect 68962 34862 68974 34914
rect 72146 34862 72158 34914
rect 72210 34862 72222 34914
rect 72706 34862 72718 34914
rect 72770 34862 72782 34914
rect 78418 34862 78430 34914
rect 78482 34862 78494 34914
rect 84578 34862 84590 34914
rect 84642 34862 84654 34914
rect 85026 34862 85038 34914
rect 85090 34862 85102 34914
rect 61630 34850 61682 34862
rect 68462 34850 68514 34862
rect 78094 34850 78146 34862
rect 1710 34802 1762 34814
rect 1710 34738 1762 34750
rect 5070 34802 5122 34814
rect 5070 34738 5122 34750
rect 24894 34802 24946 34814
rect 24894 34738 24946 34750
rect 35758 34802 35810 34814
rect 44942 34802 44994 34814
rect 36978 34750 36990 34802
rect 37042 34750 37054 34802
rect 40786 34750 40798 34802
rect 40850 34750 40862 34802
rect 43026 34750 43038 34802
rect 43090 34750 43102 34802
rect 35758 34738 35810 34750
rect 44942 34738 44994 34750
rect 46846 34802 46898 34814
rect 46846 34738 46898 34750
rect 48414 34802 48466 34814
rect 48414 34738 48466 34750
rect 49870 34802 49922 34814
rect 49870 34738 49922 34750
rect 53118 34802 53170 34814
rect 53118 34738 53170 34750
rect 55022 34802 55074 34814
rect 77646 34802 77698 34814
rect 65426 34750 65438 34802
rect 65490 34750 65502 34802
rect 55022 34738 55074 34750
rect 77646 34738 77698 34750
rect 80782 34802 80834 34814
rect 80782 34738 80834 34750
rect 88174 34802 88226 34814
rect 88174 34738 88226 34750
rect 96238 34802 96290 34814
rect 96238 34738 96290 34750
rect 96574 34802 96626 34814
rect 96574 34738 96626 34750
rect 2046 34690 2098 34702
rect 2046 34626 2098 34638
rect 2382 34690 2434 34702
rect 2382 34626 2434 34638
rect 2942 34690 2994 34702
rect 9214 34690 9266 34702
rect 8642 34638 8654 34690
rect 8706 34638 8718 34690
rect 2942 34626 2994 34638
rect 9214 34626 9266 34638
rect 11342 34690 11394 34702
rect 26238 34690 26290 34702
rect 24210 34638 24222 34690
rect 24274 34638 24286 34690
rect 11342 34626 11394 34638
rect 26238 34626 26290 34638
rect 27470 34690 27522 34702
rect 27470 34626 27522 34638
rect 35534 34690 35586 34702
rect 35534 34626 35586 34638
rect 36430 34690 36482 34702
rect 36430 34626 36482 34638
rect 41246 34690 41298 34702
rect 41246 34626 41298 34638
rect 46958 34690 47010 34702
rect 46958 34626 47010 34638
rect 50318 34690 50370 34702
rect 50318 34626 50370 34638
rect 52894 34690 52946 34702
rect 52894 34626 52946 34638
rect 54686 34690 54738 34702
rect 67902 34690 67954 34702
rect 75742 34690 75794 34702
rect 58146 34638 58158 34690
rect 58210 34638 58222 34690
rect 71138 34638 71150 34690
rect 71202 34638 71214 34690
rect 75170 34638 75182 34690
rect 75234 34638 75246 34690
rect 54686 34626 54738 34638
rect 67902 34626 67954 34638
rect 75742 34626 75794 34638
rect 76414 34690 76466 34702
rect 76414 34626 76466 34638
rect 84366 34690 84418 34702
rect 87378 34638 87390 34690
rect 87442 34638 87454 34690
rect 84366 34626 84418 34638
rect 1344 34522 98560 34556
rect 1344 34470 8896 34522
rect 8948 34470 9020 34522
rect 9072 34470 9144 34522
rect 9196 34470 9268 34522
rect 9320 34470 17896 34522
rect 17948 34470 18020 34522
rect 18072 34470 18144 34522
rect 18196 34470 18268 34522
rect 18320 34470 26896 34522
rect 26948 34470 27020 34522
rect 27072 34470 27144 34522
rect 27196 34470 27268 34522
rect 27320 34470 35896 34522
rect 35948 34470 36020 34522
rect 36072 34470 36144 34522
rect 36196 34470 36268 34522
rect 36320 34470 44896 34522
rect 44948 34470 45020 34522
rect 45072 34470 45144 34522
rect 45196 34470 45268 34522
rect 45320 34470 53896 34522
rect 53948 34470 54020 34522
rect 54072 34470 54144 34522
rect 54196 34470 54268 34522
rect 54320 34470 62896 34522
rect 62948 34470 63020 34522
rect 63072 34470 63144 34522
rect 63196 34470 63268 34522
rect 63320 34470 71896 34522
rect 71948 34470 72020 34522
rect 72072 34470 72144 34522
rect 72196 34470 72268 34522
rect 72320 34470 80896 34522
rect 80948 34470 81020 34522
rect 81072 34470 81144 34522
rect 81196 34470 81268 34522
rect 81320 34470 89896 34522
rect 89948 34470 90020 34522
rect 90072 34470 90144 34522
rect 90196 34470 90268 34522
rect 90320 34470 98560 34522
rect 1344 34436 98560 34470
rect 37102 34354 37154 34366
rect 4722 34302 4734 34354
rect 4786 34302 4798 34354
rect 30146 34302 30158 34354
rect 30210 34302 30222 34354
rect 37102 34290 37154 34302
rect 38670 34354 38722 34366
rect 38670 34290 38722 34302
rect 39566 34354 39618 34366
rect 39566 34290 39618 34302
rect 41022 34354 41074 34366
rect 41022 34290 41074 34302
rect 41470 34354 41522 34366
rect 41470 34290 41522 34302
rect 46286 34354 46338 34366
rect 50430 34354 50482 34366
rect 47954 34302 47966 34354
rect 48018 34302 48030 34354
rect 46286 34290 46338 34302
rect 50430 34290 50482 34302
rect 50990 34354 51042 34366
rect 55694 34354 55746 34366
rect 51538 34302 51550 34354
rect 51602 34302 51614 34354
rect 50990 34290 51042 34302
rect 55694 34290 55746 34302
rect 61630 34354 61682 34366
rect 61630 34290 61682 34302
rect 62190 34354 62242 34366
rect 62190 34290 62242 34302
rect 64654 34354 64706 34366
rect 64654 34290 64706 34302
rect 72494 34354 72546 34366
rect 72494 34290 72546 34302
rect 72830 34354 72882 34366
rect 72830 34290 72882 34302
rect 74510 34354 74562 34366
rect 74510 34290 74562 34302
rect 85374 34354 85426 34366
rect 85374 34290 85426 34302
rect 85822 34354 85874 34366
rect 85822 34290 85874 34302
rect 14030 34242 14082 34254
rect 14030 34178 14082 34190
rect 20862 34242 20914 34254
rect 20862 34178 20914 34190
rect 30942 34242 30994 34254
rect 30942 34178 30994 34190
rect 32510 34242 32562 34254
rect 32510 34178 32562 34190
rect 35870 34242 35922 34254
rect 35870 34178 35922 34190
rect 40238 34242 40290 34254
rect 40238 34178 40290 34190
rect 47518 34242 47570 34254
rect 55358 34242 55410 34254
rect 63758 34242 63810 34254
rect 52658 34190 52670 34242
rect 52722 34190 52734 34242
rect 57362 34190 57374 34242
rect 57426 34190 57438 34242
rect 57698 34190 57710 34242
rect 57762 34190 57774 34242
rect 63074 34190 63086 34242
rect 63138 34190 63150 34242
rect 47518 34178 47570 34190
rect 55358 34178 55410 34190
rect 63758 34178 63810 34190
rect 76190 34242 76242 34254
rect 76190 34178 76242 34190
rect 76526 34242 76578 34254
rect 76526 34178 76578 34190
rect 85934 34242 85986 34254
rect 85934 34178 85986 34190
rect 1822 34130 1874 34142
rect 11342 34130 11394 34142
rect 27358 34130 27410 34142
rect 32958 34130 33010 34142
rect 39790 34130 39842 34142
rect 2258 34078 2270 34130
rect 2322 34078 2334 34130
rect 11778 34078 11790 34130
rect 11842 34078 11854 34130
rect 27794 34078 27806 34130
rect 27858 34078 27870 34130
rect 33506 34078 33518 34130
rect 33570 34078 33582 34130
rect 38994 34078 39006 34130
rect 39058 34078 39070 34130
rect 39330 34078 39342 34130
rect 39394 34078 39406 34130
rect 1822 34066 1874 34078
rect 11342 34066 11394 34078
rect 27358 34066 27410 34078
rect 32958 34066 33010 34078
rect 39790 34066 39842 34078
rect 40126 34130 40178 34142
rect 47294 34130 47346 34142
rect 46834 34078 46846 34130
rect 46898 34078 46910 34130
rect 40126 34066 40178 34078
rect 47294 34066 47346 34078
rect 47406 34130 47458 34142
rect 49758 34130 49810 34142
rect 49298 34078 49310 34130
rect 49362 34078 49374 34130
rect 47406 34066 47458 34078
rect 49758 34066 49810 34078
rect 50094 34130 50146 34142
rect 56030 34130 56082 34142
rect 52322 34078 52334 34130
rect 52386 34078 52398 34130
rect 50094 34066 50146 34078
rect 56030 34066 56082 34078
rect 56814 34130 56866 34142
rect 64318 34130 64370 34142
rect 62962 34078 62974 34130
rect 63026 34078 63038 34130
rect 56814 34066 56866 34078
rect 64318 34066 64370 34078
rect 64654 34130 64706 34142
rect 64654 34066 64706 34078
rect 64878 34130 64930 34142
rect 64878 34066 64930 34078
rect 65438 34130 65490 34142
rect 65438 34066 65490 34078
rect 72718 34130 72770 34142
rect 72718 34066 72770 34078
rect 72942 34130 72994 34142
rect 72942 34066 72994 34078
rect 73390 34130 73442 34142
rect 73390 34066 73442 34078
rect 74286 34130 74338 34142
rect 74286 34066 74338 34078
rect 74622 34130 74674 34142
rect 74622 34066 74674 34078
rect 96574 34130 96626 34142
rect 97010 34078 97022 34130
rect 97074 34078 97086 34130
rect 96574 34066 96626 34078
rect 5294 34018 5346 34030
rect 5294 33954 5346 33966
rect 5630 34018 5682 34030
rect 5630 33954 5682 33966
rect 27022 34018 27074 34030
rect 27022 33954 27074 33966
rect 31390 34018 31442 34030
rect 31390 33954 31442 33966
rect 32174 34018 32226 34030
rect 32174 33954 32226 33966
rect 38222 34018 38274 34030
rect 44606 34018 44658 34030
rect 39442 33966 39454 34018
rect 39506 33966 39518 34018
rect 38222 33954 38274 33966
rect 44606 33954 44658 33966
rect 45278 34018 45330 34030
rect 61070 34018 61122 34030
rect 48850 33966 48862 34018
rect 48914 33966 48926 34018
rect 45278 33954 45330 33966
rect 61070 33954 61122 33966
rect 73726 34018 73778 34030
rect 73726 33954 73778 33966
rect 75070 34018 75122 34030
rect 75070 33954 75122 33966
rect 14814 33906 14866 33918
rect 14814 33842 14866 33854
rect 57150 33906 57202 33918
rect 57150 33842 57202 33854
rect 62526 33906 62578 33918
rect 62526 33842 62578 33854
rect 85822 33906 85874 33918
rect 85822 33842 85874 33854
rect 97694 33906 97746 33918
rect 97694 33842 97746 33854
rect 1344 33738 98560 33772
rect 1344 33686 4396 33738
rect 4448 33686 4520 33738
rect 4572 33686 4644 33738
rect 4696 33686 4768 33738
rect 4820 33686 13396 33738
rect 13448 33686 13520 33738
rect 13572 33686 13644 33738
rect 13696 33686 13768 33738
rect 13820 33686 22396 33738
rect 22448 33686 22520 33738
rect 22572 33686 22644 33738
rect 22696 33686 22768 33738
rect 22820 33686 31396 33738
rect 31448 33686 31520 33738
rect 31572 33686 31644 33738
rect 31696 33686 31768 33738
rect 31820 33686 40396 33738
rect 40448 33686 40520 33738
rect 40572 33686 40644 33738
rect 40696 33686 40768 33738
rect 40820 33686 49396 33738
rect 49448 33686 49520 33738
rect 49572 33686 49644 33738
rect 49696 33686 49768 33738
rect 49820 33686 58396 33738
rect 58448 33686 58520 33738
rect 58572 33686 58644 33738
rect 58696 33686 58768 33738
rect 58820 33686 67396 33738
rect 67448 33686 67520 33738
rect 67572 33686 67644 33738
rect 67696 33686 67768 33738
rect 67820 33686 76396 33738
rect 76448 33686 76520 33738
rect 76572 33686 76644 33738
rect 76696 33686 76768 33738
rect 76820 33686 85396 33738
rect 85448 33686 85520 33738
rect 85572 33686 85644 33738
rect 85696 33686 85768 33738
rect 85820 33686 94396 33738
rect 94448 33686 94520 33738
rect 94572 33686 94644 33738
rect 94696 33686 94768 33738
rect 94820 33686 98560 33738
rect 1344 33652 98560 33686
rect 45502 33570 45554 33582
rect 45502 33506 45554 33518
rect 14590 33458 14642 33470
rect 14590 33394 14642 33406
rect 19070 33458 19122 33470
rect 19070 33394 19122 33406
rect 45950 33458 46002 33470
rect 45950 33394 46002 33406
rect 53230 33458 53282 33470
rect 53230 33394 53282 33406
rect 60846 33458 60898 33470
rect 60846 33394 60898 33406
rect 67006 33458 67058 33470
rect 67006 33394 67058 33406
rect 15822 33346 15874 33358
rect 15026 33294 15038 33346
rect 15090 33294 15102 33346
rect 15822 33282 15874 33294
rect 16718 33346 16770 33358
rect 20302 33346 20354 33358
rect 19618 33294 19630 33346
rect 19682 33294 19694 33346
rect 16718 33282 16770 33294
rect 20302 33282 20354 33294
rect 20638 33346 20690 33358
rect 38894 33346 38946 33358
rect 45054 33346 45106 33358
rect 21522 33294 21534 33346
rect 21586 33294 21598 33346
rect 39330 33294 39342 33346
rect 39394 33294 39406 33346
rect 44258 33294 44270 33346
rect 44322 33294 44334 33346
rect 20638 33282 20690 33294
rect 38894 33282 38946 33294
rect 45054 33282 45106 33294
rect 45166 33346 45218 33358
rect 45166 33282 45218 33294
rect 45390 33346 45442 33358
rect 48862 33346 48914 33358
rect 48514 33294 48526 33346
rect 48578 33294 48590 33346
rect 45390 33282 45442 33294
rect 48862 33282 48914 33294
rect 61854 33346 61906 33358
rect 61854 33282 61906 33294
rect 63198 33346 63250 33358
rect 63522 33294 63534 33346
rect 63586 33294 63598 33346
rect 63198 33282 63250 33294
rect 1710 33234 1762 33246
rect 1710 33170 1762 33182
rect 2494 33234 2546 33246
rect 43934 33234 43986 33246
rect 15138 33182 15150 33234
rect 15202 33182 15214 33234
rect 19506 33182 19518 33234
rect 19570 33182 19582 33234
rect 2494 33170 2546 33182
rect 43934 33170 43986 33182
rect 47406 33234 47458 33246
rect 47406 33170 47458 33182
rect 49422 33234 49474 33246
rect 62066 33182 62078 33234
rect 62130 33182 62142 33234
rect 62514 33182 62526 33234
rect 62578 33182 62590 33234
rect 49422 33170 49474 33182
rect 2046 33122 2098 33134
rect 2046 33058 2098 33070
rect 8878 33122 8930 33134
rect 8878 33058 8930 33070
rect 16158 33122 16210 33134
rect 16158 33058 16210 33070
rect 21310 33122 21362 33134
rect 21310 33058 21362 33070
rect 32510 33122 32562 33134
rect 32510 33058 32562 33070
rect 38558 33122 38610 33134
rect 42366 33122 42418 33134
rect 41794 33070 41806 33122
rect 41858 33070 41870 33122
rect 38558 33058 38610 33070
rect 42366 33058 42418 33070
rect 44046 33122 44098 33134
rect 44046 33058 44098 33070
rect 46398 33122 46450 33134
rect 56366 33122 56418 33134
rect 50418 33070 50430 33122
rect 50482 33070 50494 33122
rect 46398 33058 46450 33070
rect 56366 33058 56418 33070
rect 61518 33122 61570 33134
rect 66670 33122 66722 33134
rect 66098 33070 66110 33122
rect 66162 33070 66174 33122
rect 61518 33058 61570 33070
rect 66670 33058 66722 33070
rect 1344 32954 98560 32988
rect 1344 32902 8896 32954
rect 8948 32902 9020 32954
rect 9072 32902 9144 32954
rect 9196 32902 9268 32954
rect 9320 32902 17896 32954
rect 17948 32902 18020 32954
rect 18072 32902 18144 32954
rect 18196 32902 18268 32954
rect 18320 32902 26896 32954
rect 26948 32902 27020 32954
rect 27072 32902 27144 32954
rect 27196 32902 27268 32954
rect 27320 32902 35896 32954
rect 35948 32902 36020 32954
rect 36072 32902 36144 32954
rect 36196 32902 36268 32954
rect 36320 32902 44896 32954
rect 44948 32902 45020 32954
rect 45072 32902 45144 32954
rect 45196 32902 45268 32954
rect 45320 32902 53896 32954
rect 53948 32902 54020 32954
rect 54072 32902 54144 32954
rect 54196 32902 54268 32954
rect 54320 32902 62896 32954
rect 62948 32902 63020 32954
rect 63072 32902 63144 32954
rect 63196 32902 63268 32954
rect 63320 32902 71896 32954
rect 71948 32902 72020 32954
rect 72072 32902 72144 32954
rect 72196 32902 72268 32954
rect 72320 32902 80896 32954
rect 80948 32902 81020 32954
rect 81072 32902 81144 32954
rect 81196 32902 81268 32954
rect 81320 32902 89896 32954
rect 89948 32902 90020 32954
rect 90072 32902 90144 32954
rect 90196 32902 90268 32954
rect 90320 32902 98560 32954
rect 1344 32868 98560 32902
rect 13134 32786 13186 32798
rect 38894 32786 38946 32798
rect 29026 32734 29038 32786
rect 29090 32734 29102 32786
rect 13134 32722 13186 32734
rect 38894 32722 38946 32734
rect 41022 32786 41074 32798
rect 41022 32722 41074 32734
rect 41470 32786 41522 32798
rect 41470 32722 41522 32734
rect 46174 32786 46226 32798
rect 46174 32722 46226 32734
rect 47854 32786 47906 32798
rect 47854 32722 47906 32734
rect 48302 32786 48354 32798
rect 53118 32786 53170 32798
rect 52546 32734 52558 32786
rect 52610 32734 52622 32786
rect 48302 32722 48354 32734
rect 53118 32722 53170 32734
rect 55246 32786 55298 32798
rect 55246 32722 55298 32734
rect 55694 32786 55746 32798
rect 55694 32722 55746 32734
rect 59838 32786 59890 32798
rect 59838 32722 59890 32734
rect 60734 32786 60786 32798
rect 60734 32722 60786 32734
rect 61182 32786 61234 32798
rect 61182 32722 61234 32734
rect 63758 32786 63810 32798
rect 63758 32722 63810 32734
rect 2046 32674 2098 32686
rect 2046 32610 2098 32622
rect 8542 32674 8594 32686
rect 8542 32610 8594 32622
rect 12350 32674 12402 32686
rect 12350 32610 12402 32622
rect 14814 32674 14866 32686
rect 14814 32610 14866 32622
rect 15150 32674 15202 32686
rect 15150 32610 15202 32622
rect 15486 32674 15538 32686
rect 15486 32610 15538 32622
rect 20302 32674 20354 32686
rect 20302 32610 20354 32622
rect 23438 32674 23490 32686
rect 23438 32610 23490 32622
rect 29710 32674 29762 32686
rect 29710 32610 29762 32622
rect 35982 32674 36034 32686
rect 35982 32610 36034 32622
rect 39230 32674 39282 32686
rect 46398 32674 46450 32686
rect 44034 32622 44046 32674
rect 44098 32622 44110 32674
rect 39230 32610 39282 32622
rect 46398 32610 46450 32622
rect 49198 32674 49250 32686
rect 56030 32674 56082 32686
rect 54562 32622 54574 32674
rect 54626 32622 54638 32674
rect 57250 32622 57262 32674
rect 57314 32622 57326 32674
rect 57810 32622 57822 32674
rect 57874 32622 57886 32674
rect 61394 32622 61406 32674
rect 61458 32622 61470 32674
rect 63298 32622 63310 32674
rect 63362 32622 63374 32674
rect 49198 32610 49250 32622
rect 56030 32610 56082 32622
rect 1710 32562 1762 32574
rect 1710 32498 1762 32510
rect 9102 32562 9154 32574
rect 20526 32562 20578 32574
rect 26126 32562 26178 32574
rect 35870 32562 35922 32574
rect 9538 32510 9550 32562
rect 9602 32510 9614 32562
rect 9986 32510 9998 32562
rect 10050 32510 10062 32562
rect 21186 32510 21198 32562
rect 21250 32510 21262 32562
rect 26450 32510 26462 32562
rect 26514 32510 26526 32562
rect 9102 32498 9154 32510
rect 20526 32498 20578 32510
rect 26126 32498 26178 32510
rect 35870 32498 35922 32510
rect 36206 32562 36258 32574
rect 36206 32498 36258 32510
rect 39342 32562 39394 32574
rect 39342 32498 39394 32510
rect 39678 32562 39730 32574
rect 45726 32562 45778 32574
rect 39890 32510 39902 32562
rect 39954 32510 39966 32562
rect 40226 32510 40238 32562
rect 40290 32510 40302 32562
rect 43810 32510 43822 32562
rect 43874 32510 43886 32562
rect 39678 32498 39730 32510
rect 45726 32498 45778 32510
rect 46510 32562 46562 32574
rect 46510 32498 46562 32510
rect 49422 32562 49474 32574
rect 53790 32562 53842 32574
rect 57038 32562 57090 32574
rect 62974 32562 63026 32574
rect 50082 32510 50094 32562
rect 50146 32510 50158 32562
rect 54450 32510 54462 32562
rect 54514 32510 54526 32562
rect 61730 32510 61742 32562
rect 61794 32510 61806 32562
rect 62514 32510 62526 32562
rect 62578 32510 62590 32562
rect 49422 32498 49474 32510
rect 53790 32498 53842 32510
rect 57038 32498 57090 32510
rect 62974 32498 63026 32510
rect 2494 32450 2546 32462
rect 2494 32386 2546 32398
rect 25790 32450 25842 32462
rect 25790 32386 25842 32398
rect 30158 32450 30210 32462
rect 30158 32386 30210 32398
rect 38446 32450 38498 32462
rect 60286 32450 60338 32462
rect 64878 32450 64930 32462
rect 44594 32398 44606 32450
rect 44658 32398 44670 32450
rect 63074 32398 63086 32450
rect 63138 32398 63150 32450
rect 38446 32386 38498 32398
rect 60286 32386 60338 32398
rect 64878 32386 64930 32398
rect 24222 32338 24274 32350
rect 24222 32274 24274 32286
rect 53454 32338 53506 32350
rect 53454 32274 53506 32286
rect 56702 32338 56754 32350
rect 56702 32274 56754 32286
rect 1344 32170 98560 32204
rect 1344 32118 4396 32170
rect 4448 32118 4520 32170
rect 4572 32118 4644 32170
rect 4696 32118 4768 32170
rect 4820 32118 13396 32170
rect 13448 32118 13520 32170
rect 13572 32118 13644 32170
rect 13696 32118 13768 32170
rect 13820 32118 22396 32170
rect 22448 32118 22520 32170
rect 22572 32118 22644 32170
rect 22696 32118 22768 32170
rect 22820 32118 31396 32170
rect 31448 32118 31520 32170
rect 31572 32118 31644 32170
rect 31696 32118 31768 32170
rect 31820 32118 40396 32170
rect 40448 32118 40520 32170
rect 40572 32118 40644 32170
rect 40696 32118 40768 32170
rect 40820 32118 49396 32170
rect 49448 32118 49520 32170
rect 49572 32118 49644 32170
rect 49696 32118 49768 32170
rect 49820 32118 58396 32170
rect 58448 32118 58520 32170
rect 58572 32118 58644 32170
rect 58696 32118 58768 32170
rect 58820 32118 67396 32170
rect 67448 32118 67520 32170
rect 67572 32118 67644 32170
rect 67696 32118 67768 32170
rect 67820 32118 76396 32170
rect 76448 32118 76520 32170
rect 76572 32118 76644 32170
rect 76696 32118 76768 32170
rect 76820 32118 85396 32170
rect 85448 32118 85520 32170
rect 85572 32118 85644 32170
rect 85696 32118 85768 32170
rect 85820 32118 94396 32170
rect 94448 32118 94520 32170
rect 94572 32118 94644 32170
rect 94696 32118 94768 32170
rect 94820 32118 98560 32170
rect 1344 32084 98560 32118
rect 42366 32002 42418 32014
rect 64094 32002 64146 32014
rect 43362 31950 43374 32002
rect 43426 31950 43438 32002
rect 42366 31938 42418 31950
rect 64094 31938 64146 31950
rect 9214 31890 9266 31902
rect 9214 31826 9266 31838
rect 38894 31890 38946 31902
rect 38894 31826 38946 31838
rect 42926 31890 42978 31902
rect 53118 31890 53170 31902
rect 45826 31838 45838 31890
rect 45890 31838 45902 31890
rect 42926 31826 42978 31838
rect 53118 31826 53170 31838
rect 64430 31890 64482 31902
rect 64430 31826 64482 31838
rect 68574 31890 68626 31902
rect 68574 31826 68626 31838
rect 5518 31778 5570 31790
rect 14590 31778 14642 31790
rect 27134 31778 27186 31790
rect 6066 31726 6078 31778
rect 6130 31726 6142 31778
rect 14914 31726 14926 31778
rect 14978 31726 14990 31778
rect 5518 31714 5570 31726
rect 14590 31714 14642 31726
rect 27134 31714 27186 31726
rect 36206 31778 36258 31790
rect 43598 31778 43650 31790
rect 39218 31726 39230 31778
rect 39282 31726 39294 31778
rect 41458 31726 41470 31778
rect 41522 31726 41534 31778
rect 36206 31714 36258 31726
rect 43598 31714 43650 31726
rect 44046 31778 44098 31790
rect 51214 31778 51266 31790
rect 44818 31726 44830 31778
rect 44882 31726 44894 31778
rect 46498 31726 46510 31778
rect 46562 31726 46574 31778
rect 44046 31714 44098 31726
rect 51214 31714 51266 31726
rect 56142 31778 56194 31790
rect 56142 31714 56194 31726
rect 60398 31778 60450 31790
rect 65774 31778 65826 31790
rect 61058 31726 61070 31778
rect 61122 31726 61134 31778
rect 60398 31714 60450 31726
rect 65774 31714 65826 31726
rect 69246 31778 69298 31790
rect 69794 31726 69806 31778
rect 69858 31726 69870 31778
rect 96898 31726 96910 31778
rect 96962 31726 96974 31778
rect 69246 31714 69298 31726
rect 1710 31666 1762 31678
rect 1710 31602 1762 31614
rect 5070 31666 5122 31678
rect 5070 31602 5122 31614
rect 18062 31666 18114 31678
rect 18062 31602 18114 31614
rect 35870 31666 35922 31678
rect 35870 31602 35922 31614
rect 36318 31666 36370 31678
rect 36318 31602 36370 31614
rect 36542 31666 36594 31678
rect 50878 31666 50930 31678
rect 40674 31614 40686 31666
rect 40738 31614 40750 31666
rect 41570 31614 41582 31666
rect 41634 31614 41646 31666
rect 45378 31614 45390 31666
rect 45442 31614 45454 31666
rect 36542 31602 36594 31614
rect 50878 31602 50930 31614
rect 59950 31666 60002 31678
rect 59950 31602 60002 31614
rect 65102 31666 65154 31678
rect 65102 31602 65154 31614
rect 69022 31666 69074 31678
rect 69022 31602 69074 31614
rect 72942 31666 72994 31678
rect 72942 31602 72994 31614
rect 74062 31666 74114 31678
rect 98018 31614 98030 31666
rect 98082 31614 98094 31666
rect 74062 31602 74114 31614
rect 2046 31554 2098 31566
rect 2046 31490 2098 31502
rect 2382 31554 2434 31566
rect 2382 31490 2434 31502
rect 2942 31554 2994 31566
rect 18398 31554 18450 31566
rect 8642 31502 8654 31554
rect 8706 31502 8718 31554
rect 17490 31502 17502 31554
rect 17554 31502 17566 31554
rect 2942 31490 2994 31502
rect 18398 31490 18450 31502
rect 26798 31554 26850 31566
rect 26798 31490 26850 31502
rect 27470 31554 27522 31566
rect 27470 31490 27522 31502
rect 30046 31554 30098 31566
rect 30046 31490 30098 31502
rect 32734 31554 32786 31566
rect 32734 31490 32786 31502
rect 38446 31554 38498 31566
rect 38446 31490 38498 31502
rect 55806 31554 55858 31566
rect 55806 31490 55858 31502
rect 56478 31554 56530 31566
rect 65214 31554 65266 31566
rect 63522 31502 63534 31554
rect 63586 31502 63598 31554
rect 56478 31490 56530 31502
rect 65214 31490 65266 31502
rect 65326 31554 65378 31566
rect 65326 31490 65378 31502
rect 65998 31554 66050 31566
rect 65998 31490 66050 31502
rect 66558 31554 66610 31566
rect 74398 31554 74450 31566
rect 72146 31502 72158 31554
rect 72210 31502 72222 31554
rect 66558 31490 66610 31502
rect 74398 31490 74450 31502
rect 96686 31554 96738 31566
rect 96686 31490 96738 31502
rect 1344 31386 98560 31420
rect 1344 31334 8896 31386
rect 8948 31334 9020 31386
rect 9072 31334 9144 31386
rect 9196 31334 9268 31386
rect 9320 31334 17896 31386
rect 17948 31334 18020 31386
rect 18072 31334 18144 31386
rect 18196 31334 18268 31386
rect 18320 31334 26896 31386
rect 26948 31334 27020 31386
rect 27072 31334 27144 31386
rect 27196 31334 27268 31386
rect 27320 31334 35896 31386
rect 35948 31334 36020 31386
rect 36072 31334 36144 31386
rect 36196 31334 36268 31386
rect 36320 31334 44896 31386
rect 44948 31334 45020 31386
rect 45072 31334 45144 31386
rect 45196 31334 45268 31386
rect 45320 31334 53896 31386
rect 53948 31334 54020 31386
rect 54072 31334 54144 31386
rect 54196 31334 54268 31386
rect 54320 31334 62896 31386
rect 62948 31334 63020 31386
rect 63072 31334 63144 31386
rect 63196 31334 63268 31386
rect 63320 31334 71896 31386
rect 71948 31334 72020 31386
rect 72072 31334 72144 31386
rect 72196 31334 72268 31386
rect 72320 31334 80896 31386
rect 80948 31334 81020 31386
rect 81072 31334 81144 31386
rect 81196 31334 81268 31386
rect 81320 31334 89896 31386
rect 89948 31334 90020 31386
rect 90072 31334 90144 31386
rect 90196 31334 90268 31386
rect 90320 31334 98560 31386
rect 1344 31300 98560 31334
rect 19966 31218 20018 31230
rect 30606 31218 30658 31230
rect 4722 31166 4734 31218
rect 4786 31166 4798 31218
rect 29362 31166 29374 31218
rect 29426 31166 29438 31218
rect 19966 31154 20018 31166
rect 30606 31154 30658 31166
rect 38894 31218 38946 31230
rect 38894 31154 38946 31166
rect 39790 31218 39842 31230
rect 39790 31154 39842 31166
rect 42702 31218 42754 31230
rect 42702 31154 42754 31166
rect 61182 31218 61234 31230
rect 68910 31218 68962 31230
rect 67890 31166 67902 31218
rect 67954 31166 67966 31218
rect 61182 31154 61234 31166
rect 68910 31154 68962 31166
rect 69806 31218 69858 31230
rect 69806 31154 69858 31166
rect 69918 31218 69970 31230
rect 69918 31154 69970 31166
rect 70702 31218 70754 31230
rect 70702 31154 70754 31166
rect 72382 31218 72434 31230
rect 72382 31154 72434 31166
rect 72942 31218 72994 31230
rect 72942 31154 72994 31166
rect 20862 31106 20914 31118
rect 20862 31042 20914 31054
rect 23998 31106 24050 31118
rect 35870 31106 35922 31118
rect 46846 31106 46898 31118
rect 31042 31054 31054 31106
rect 31106 31054 31118 31106
rect 43810 31054 43822 31106
rect 43874 31054 43886 31106
rect 45042 31054 45054 31106
rect 45106 31054 45118 31106
rect 23998 31042 24050 31054
rect 35870 31042 35922 31054
rect 46846 31042 46898 31054
rect 69470 31106 69522 31118
rect 69470 31042 69522 31054
rect 69694 31106 69746 31118
rect 69694 31042 69746 31054
rect 1822 30994 1874 31006
rect 20414 30994 20466 31006
rect 2146 30942 2158 30994
rect 2210 30942 2222 30994
rect 1822 30930 1874 30942
rect 20414 30930 20466 30942
rect 21086 30994 21138 31006
rect 26462 30994 26514 31006
rect 32958 30994 33010 31006
rect 39678 30994 39730 31006
rect 21634 30942 21646 30994
rect 21698 30942 21710 30994
rect 26786 30942 26798 30994
rect 26850 30942 26862 30994
rect 30930 30942 30942 30994
rect 30994 30942 31006 30994
rect 33506 30942 33518 30994
rect 33570 30942 33582 30994
rect 21086 30930 21138 30942
rect 26462 30930 26514 30942
rect 32958 30930 33010 30942
rect 39678 30930 39730 30942
rect 40014 30994 40066 31006
rect 46398 30994 46450 31006
rect 61518 30994 61570 31006
rect 44034 30942 44046 30994
rect 44098 30942 44110 30994
rect 47170 30942 47182 30994
rect 47234 30942 47246 30994
rect 40014 30930 40066 30942
rect 46398 30930 46450 30942
rect 61518 30930 61570 30942
rect 65102 30994 65154 31006
rect 70366 30994 70418 31006
rect 65426 30942 65438 30994
rect 65490 30942 65502 30994
rect 65102 30930 65154 30942
rect 70366 30930 70418 30942
rect 72494 30994 72546 31006
rect 72494 30930 72546 30942
rect 14702 30882 14754 30894
rect 14702 30818 14754 30830
rect 31726 30882 31778 30894
rect 31726 30818 31778 30830
rect 39454 30882 39506 30894
rect 46958 30882 47010 30894
rect 44482 30830 44494 30882
rect 44546 30830 44558 30882
rect 39454 30818 39506 30830
rect 46958 30818 47010 30830
rect 5294 30770 5346 30782
rect 5294 30706 5346 30718
rect 24782 30770 24834 30782
rect 24782 30706 24834 30718
rect 29934 30770 29986 30782
rect 29934 30706 29986 30718
rect 32062 30770 32114 30782
rect 32062 30706 32114 30718
rect 36654 30770 36706 30782
rect 68574 30770 68626 30782
rect 39218 30718 39230 30770
rect 39282 30767 39294 30770
rect 39442 30767 39454 30770
rect 39282 30721 39454 30767
rect 39282 30718 39294 30721
rect 39442 30718 39454 30721
rect 39506 30718 39518 30770
rect 36654 30706 36706 30718
rect 68574 30706 68626 30718
rect 72382 30770 72434 30782
rect 72382 30706 72434 30718
rect 1344 30602 98560 30636
rect 1344 30550 4396 30602
rect 4448 30550 4520 30602
rect 4572 30550 4644 30602
rect 4696 30550 4768 30602
rect 4820 30550 13396 30602
rect 13448 30550 13520 30602
rect 13572 30550 13644 30602
rect 13696 30550 13768 30602
rect 13820 30550 22396 30602
rect 22448 30550 22520 30602
rect 22572 30550 22644 30602
rect 22696 30550 22768 30602
rect 22820 30550 31396 30602
rect 31448 30550 31520 30602
rect 31572 30550 31644 30602
rect 31696 30550 31768 30602
rect 31820 30550 40396 30602
rect 40448 30550 40520 30602
rect 40572 30550 40644 30602
rect 40696 30550 40768 30602
rect 40820 30550 49396 30602
rect 49448 30550 49520 30602
rect 49572 30550 49644 30602
rect 49696 30550 49768 30602
rect 49820 30550 58396 30602
rect 58448 30550 58520 30602
rect 58572 30550 58644 30602
rect 58696 30550 58768 30602
rect 58820 30550 67396 30602
rect 67448 30550 67520 30602
rect 67572 30550 67644 30602
rect 67696 30550 67768 30602
rect 67820 30550 76396 30602
rect 76448 30550 76520 30602
rect 76572 30550 76644 30602
rect 76696 30550 76768 30602
rect 76820 30550 85396 30602
rect 85448 30550 85520 30602
rect 85572 30550 85644 30602
rect 85696 30550 85768 30602
rect 85820 30550 94396 30602
rect 94448 30550 94520 30602
rect 94572 30550 94644 30602
rect 94696 30550 94768 30602
rect 94820 30550 98560 30602
rect 1344 30516 98560 30550
rect 27918 30434 27970 30446
rect 27918 30370 27970 30382
rect 28254 30434 28306 30446
rect 28254 30370 28306 30382
rect 15934 30322 15986 30334
rect 43026 30270 43038 30322
rect 43090 30270 43102 30322
rect 85138 30270 85150 30322
rect 85202 30270 85214 30322
rect 15934 30258 15986 30270
rect 8878 30210 8930 30222
rect 26238 30210 26290 30222
rect 30270 30210 30322 30222
rect 32734 30210 32786 30222
rect 9426 30158 9438 30210
rect 9490 30158 9502 30210
rect 15138 30158 15150 30210
rect 15202 30158 15214 30210
rect 27234 30158 27246 30210
rect 27298 30158 27310 30210
rect 31826 30158 31838 30210
rect 31890 30158 31902 30210
rect 8878 30146 8930 30158
rect 26238 30146 26290 30158
rect 30270 30146 30322 30158
rect 32734 30146 32786 30158
rect 42142 30210 42194 30222
rect 42142 30146 42194 30158
rect 44158 30210 44210 30222
rect 49758 30210 49810 30222
rect 66446 30210 66498 30222
rect 45042 30158 45054 30210
rect 45106 30158 45118 30210
rect 47058 30158 47070 30210
rect 47122 30158 47134 30210
rect 52658 30158 52670 30210
rect 52722 30158 52734 30210
rect 44158 30146 44210 30158
rect 49758 30146 49810 30158
rect 66446 30146 66498 30158
rect 72494 30210 72546 30222
rect 72494 30146 72546 30158
rect 83470 30210 83522 30222
rect 84466 30158 84478 30210
rect 84530 30158 84542 30210
rect 96898 30158 96910 30210
rect 96962 30158 96974 30210
rect 83470 30146 83522 30158
rect 1710 30098 1762 30110
rect 1710 30034 1762 30046
rect 8654 30098 8706 30110
rect 8654 30034 8706 30046
rect 14702 30098 14754 30110
rect 16270 30098 16322 30110
rect 32062 30098 32114 30110
rect 15362 30046 15374 30098
rect 15426 30046 15438 30098
rect 27122 30046 27134 30098
rect 27186 30046 27198 30098
rect 14702 30034 14754 30046
rect 16270 30034 16322 30046
rect 32062 30034 32114 30046
rect 36990 30098 37042 30110
rect 36990 30034 37042 30046
rect 37102 30098 37154 30110
rect 37102 30034 37154 30046
rect 41582 30098 41634 30110
rect 41582 30034 41634 30046
rect 43598 30098 43650 30110
rect 43598 30034 43650 30046
rect 45614 30098 45666 30110
rect 45614 30034 45666 30046
rect 47630 30098 47682 30110
rect 47630 30034 47682 30046
rect 49198 30098 49250 30110
rect 49198 30034 49250 30046
rect 66670 30098 66722 30110
rect 66670 30034 66722 30046
rect 66782 30098 66834 30110
rect 66782 30034 66834 30046
rect 67230 30098 67282 30110
rect 67230 30034 67282 30046
rect 72830 30098 72882 30110
rect 72830 30034 72882 30046
rect 96686 30098 96738 30110
rect 98018 30046 98030 30098
rect 98082 30046 98094 30098
rect 96686 30034 96738 30046
rect 2046 29986 2098 29998
rect 2046 29922 2098 29934
rect 2494 29986 2546 29998
rect 12574 29986 12626 29998
rect 12002 29934 12014 29986
rect 12066 29934 12078 29986
rect 2494 29922 2546 29934
rect 12574 29922 12626 29934
rect 13918 29986 13970 29998
rect 13918 29922 13970 29934
rect 14366 29986 14418 29998
rect 14366 29922 14418 29934
rect 16830 29986 16882 29998
rect 16830 29922 16882 29934
rect 26686 29986 26738 29998
rect 26686 29922 26738 29934
rect 33182 29986 33234 29998
rect 33182 29922 33234 29934
rect 37326 29986 37378 29998
rect 49310 29986 49362 29998
rect 46722 29934 46734 29986
rect 46786 29934 46798 29986
rect 37326 29922 37378 29934
rect 49310 29922 49362 29934
rect 50206 29986 50258 29998
rect 50206 29922 50258 29934
rect 52110 29986 52162 29998
rect 59042 29934 59054 29986
rect 59106 29934 59118 29986
rect 52110 29922 52162 29934
rect 1344 29818 98560 29852
rect 1344 29766 8896 29818
rect 8948 29766 9020 29818
rect 9072 29766 9144 29818
rect 9196 29766 9268 29818
rect 9320 29766 17896 29818
rect 17948 29766 18020 29818
rect 18072 29766 18144 29818
rect 18196 29766 18268 29818
rect 18320 29766 26896 29818
rect 26948 29766 27020 29818
rect 27072 29766 27144 29818
rect 27196 29766 27268 29818
rect 27320 29766 35896 29818
rect 35948 29766 36020 29818
rect 36072 29766 36144 29818
rect 36196 29766 36268 29818
rect 36320 29766 44896 29818
rect 44948 29766 45020 29818
rect 45072 29766 45144 29818
rect 45196 29766 45268 29818
rect 45320 29766 53896 29818
rect 53948 29766 54020 29818
rect 54072 29766 54144 29818
rect 54196 29766 54268 29818
rect 54320 29766 62896 29818
rect 62948 29766 63020 29818
rect 63072 29766 63144 29818
rect 63196 29766 63268 29818
rect 63320 29766 71896 29818
rect 71948 29766 72020 29818
rect 72072 29766 72144 29818
rect 72196 29766 72268 29818
rect 72320 29766 80896 29818
rect 80948 29766 81020 29818
rect 81072 29766 81144 29818
rect 81196 29766 81268 29818
rect 81320 29766 89896 29818
rect 89948 29766 90020 29818
rect 90072 29766 90144 29818
rect 90196 29766 90268 29818
rect 90320 29766 98560 29818
rect 1344 29732 98560 29766
rect 22430 29650 22482 29662
rect 5058 29598 5070 29650
rect 5122 29598 5134 29650
rect 21522 29598 21534 29650
rect 21586 29598 21598 29650
rect 22430 29586 22482 29598
rect 39342 29650 39394 29662
rect 39342 29586 39394 29598
rect 39790 29650 39842 29662
rect 39790 29586 39842 29598
rect 44046 29650 44098 29662
rect 46174 29650 46226 29662
rect 44482 29598 44494 29650
rect 44546 29598 44558 29650
rect 44046 29586 44098 29598
rect 46174 29586 46226 29598
rect 46286 29650 46338 29662
rect 68798 29650 68850 29662
rect 53106 29598 53118 29650
rect 53170 29598 53182 29650
rect 46286 29586 46338 29598
rect 68798 29586 68850 29598
rect 69694 29650 69746 29662
rect 69694 29586 69746 29598
rect 1934 29538 1986 29550
rect 1934 29474 1986 29486
rect 16158 29538 16210 29550
rect 16158 29474 16210 29486
rect 18174 29538 18226 29550
rect 18174 29474 18226 29486
rect 38782 29538 38834 29550
rect 44158 29538 44210 29550
rect 43138 29486 43150 29538
rect 43202 29486 43214 29538
rect 38782 29474 38834 29486
rect 44158 29474 44210 29486
rect 54238 29538 54290 29550
rect 54238 29474 54290 29486
rect 56030 29538 56082 29550
rect 56030 29474 56082 29486
rect 56926 29538 56978 29550
rect 56926 29474 56978 29486
rect 57598 29538 57650 29550
rect 57598 29474 57650 29486
rect 2158 29426 2210 29438
rect 13470 29426 13522 29438
rect 17726 29426 17778 29438
rect 2706 29374 2718 29426
rect 2770 29374 2782 29426
rect 13906 29374 13918 29426
rect 13970 29374 13982 29426
rect 2158 29362 2210 29374
rect 13470 29362 13522 29374
rect 17726 29362 17778 29374
rect 18398 29426 18450 29438
rect 42478 29426 42530 29438
rect 45502 29426 45554 29438
rect 46062 29426 46114 29438
rect 18946 29374 18958 29426
rect 19010 29374 19022 29426
rect 43250 29374 43262 29426
rect 43314 29374 43326 29426
rect 44706 29374 44718 29426
rect 44770 29374 44782 29426
rect 45826 29374 45838 29426
rect 45890 29374 45902 29426
rect 18398 29362 18450 29374
rect 42478 29362 42530 29374
rect 45502 29362 45554 29374
rect 46062 29362 46114 29374
rect 46398 29426 46450 29438
rect 46398 29362 46450 29374
rect 46958 29426 47010 29438
rect 46958 29362 47010 29374
rect 50206 29426 50258 29438
rect 56814 29426 56866 29438
rect 50530 29374 50542 29426
rect 50594 29374 50606 29426
rect 50206 29362 50258 29374
rect 56814 29362 56866 29374
rect 57150 29426 57202 29438
rect 57150 29362 57202 29374
rect 68574 29426 68626 29438
rect 68574 29362 68626 29374
rect 69246 29426 69298 29438
rect 69246 29362 69298 29374
rect 75854 29426 75906 29438
rect 75854 29362 75906 29374
rect 13022 29314 13074 29326
rect 13022 29250 13074 29262
rect 68350 29314 68402 29326
rect 68350 29250 68402 29262
rect 68686 29314 68738 29326
rect 68686 29250 68738 29262
rect 5854 29202 5906 29214
rect 5854 29138 5906 29150
rect 16942 29202 16994 29214
rect 16942 29138 16994 29150
rect 22094 29202 22146 29214
rect 22094 29138 22146 29150
rect 42142 29202 42194 29214
rect 42142 29138 42194 29150
rect 44046 29202 44098 29214
rect 44046 29138 44098 29150
rect 53678 29202 53730 29214
rect 53678 29138 53730 29150
rect 1344 29034 98560 29068
rect 1344 28982 4396 29034
rect 4448 28982 4520 29034
rect 4572 28982 4644 29034
rect 4696 28982 4768 29034
rect 4820 28982 13396 29034
rect 13448 28982 13520 29034
rect 13572 28982 13644 29034
rect 13696 28982 13768 29034
rect 13820 28982 22396 29034
rect 22448 28982 22520 29034
rect 22572 28982 22644 29034
rect 22696 28982 22768 29034
rect 22820 28982 31396 29034
rect 31448 28982 31520 29034
rect 31572 28982 31644 29034
rect 31696 28982 31768 29034
rect 31820 28982 40396 29034
rect 40448 28982 40520 29034
rect 40572 28982 40644 29034
rect 40696 28982 40768 29034
rect 40820 28982 49396 29034
rect 49448 28982 49520 29034
rect 49572 28982 49644 29034
rect 49696 28982 49768 29034
rect 49820 28982 58396 29034
rect 58448 28982 58520 29034
rect 58572 28982 58644 29034
rect 58696 28982 58768 29034
rect 58820 28982 67396 29034
rect 67448 28982 67520 29034
rect 67572 28982 67644 29034
rect 67696 28982 67768 29034
rect 67820 28982 76396 29034
rect 76448 28982 76520 29034
rect 76572 28982 76644 29034
rect 76696 28982 76768 29034
rect 76820 28982 85396 29034
rect 85448 28982 85520 29034
rect 85572 28982 85644 29034
rect 85696 28982 85768 29034
rect 85820 28982 94396 29034
rect 94448 28982 94520 29034
rect 94572 28982 94644 29034
rect 94696 28982 94768 29034
rect 94820 28982 98560 29034
rect 1344 28948 98560 28982
rect 45054 28866 45106 28878
rect 45054 28802 45106 28814
rect 54910 28866 54962 28878
rect 54910 28802 54962 28814
rect 58942 28866 58994 28878
rect 58942 28802 58994 28814
rect 61182 28866 61234 28878
rect 61182 28802 61234 28814
rect 61742 28866 61794 28878
rect 61742 28802 61794 28814
rect 75406 28866 75458 28878
rect 75406 28802 75458 28814
rect 2494 28754 2546 28766
rect 2494 28690 2546 28702
rect 24222 28754 24274 28766
rect 24222 28690 24274 28702
rect 25902 28754 25954 28766
rect 60734 28754 60786 28766
rect 46498 28702 46510 28754
rect 46562 28702 46574 28754
rect 25902 28690 25954 28702
rect 60734 28690 60786 28702
rect 67342 28754 67394 28766
rect 76738 28702 76750 28754
rect 76802 28702 76814 28754
rect 67342 28690 67394 28702
rect 1710 28642 1762 28654
rect 1710 28578 1762 28590
rect 13806 28642 13858 28654
rect 26238 28642 26290 28654
rect 25442 28590 25454 28642
rect 25506 28590 25518 28642
rect 13806 28578 13858 28590
rect 26238 28578 26290 28590
rect 26798 28642 26850 28654
rect 26798 28578 26850 28590
rect 29262 28642 29314 28654
rect 29262 28578 29314 28590
rect 41694 28642 41746 28654
rect 41694 28578 41746 28590
rect 44382 28642 44434 28654
rect 47406 28642 47458 28654
rect 45826 28590 45838 28642
rect 45890 28590 45902 28642
rect 46834 28590 46846 28642
rect 46898 28590 46910 28642
rect 44382 28578 44434 28590
rect 47406 28578 47458 28590
rect 47742 28642 47794 28654
rect 62302 28642 62354 28654
rect 55346 28590 55358 28642
rect 55410 28590 55422 28642
rect 55794 28590 55806 28642
rect 55858 28590 55870 28642
rect 47742 28578 47794 28590
rect 62302 28578 62354 28590
rect 63198 28642 63250 28654
rect 63198 28578 63250 28590
rect 63646 28642 63698 28654
rect 63646 28578 63698 28590
rect 64430 28642 64482 28654
rect 64430 28578 64482 28590
rect 68238 28642 68290 28654
rect 71934 28642 71986 28654
rect 68786 28590 68798 28642
rect 68850 28590 68862 28642
rect 68238 28578 68290 28590
rect 71934 28578 71986 28590
rect 72382 28642 72434 28654
rect 96574 28642 96626 28654
rect 97694 28642 97746 28654
rect 77410 28590 77422 28642
rect 77474 28590 77486 28642
rect 97010 28590 97022 28642
rect 97074 28590 97086 28642
rect 72382 28578 72434 28590
rect 96574 28578 96626 28590
rect 97694 28578 97746 28590
rect 2046 28530 2098 28542
rect 30270 28530 30322 28542
rect 25218 28478 25230 28530
rect 25282 28478 25294 28530
rect 2046 28466 2098 28478
rect 30270 28466 30322 28478
rect 30606 28530 30658 28542
rect 30606 28466 30658 28478
rect 55022 28530 55074 28542
rect 55022 28466 55074 28478
rect 61070 28530 61122 28542
rect 61070 28466 61122 28478
rect 61182 28530 61234 28542
rect 61742 28530 61794 28542
rect 61182 28466 61234 28478
rect 61630 28474 61682 28486
rect 7422 28418 7474 28430
rect 7422 28354 7474 28366
rect 24670 28418 24722 28430
rect 24670 28354 24722 28366
rect 30942 28418 30994 28430
rect 30942 28354 30994 28366
rect 35422 28418 35474 28430
rect 35422 28354 35474 28366
rect 41358 28418 41410 28430
rect 41358 28354 41410 28366
rect 48078 28418 48130 28430
rect 48078 28354 48130 28366
rect 48526 28418 48578 28430
rect 48526 28354 48578 28366
rect 54574 28418 54626 28430
rect 54574 28354 54626 28366
rect 54910 28418 54962 28430
rect 61742 28466 61794 28478
rect 62974 28530 63026 28542
rect 62974 28466 63026 28478
rect 67790 28530 67842 28542
rect 67790 28466 67842 28478
rect 71150 28530 71202 28542
rect 71150 28466 71202 28478
rect 72718 28530 72770 28542
rect 72718 28466 72770 28478
rect 74174 28530 74226 28542
rect 74386 28478 74398 28530
rect 74450 28478 74462 28530
rect 74174 28466 74226 28478
rect 58146 28366 58158 28418
rect 58210 28366 58222 28418
rect 61630 28410 61682 28422
rect 63086 28418 63138 28430
rect 54910 28354 54962 28366
rect 63086 28354 63138 28366
rect 63870 28418 63922 28430
rect 63870 28354 63922 28366
rect 77758 28418 77810 28430
rect 77758 28354 77810 28366
rect 1344 28250 98560 28284
rect 1344 28198 8896 28250
rect 8948 28198 9020 28250
rect 9072 28198 9144 28250
rect 9196 28198 9268 28250
rect 9320 28198 17896 28250
rect 17948 28198 18020 28250
rect 18072 28198 18144 28250
rect 18196 28198 18268 28250
rect 18320 28198 26896 28250
rect 26948 28198 27020 28250
rect 27072 28198 27144 28250
rect 27196 28198 27268 28250
rect 27320 28198 35896 28250
rect 35948 28198 36020 28250
rect 36072 28198 36144 28250
rect 36196 28198 36268 28250
rect 36320 28198 44896 28250
rect 44948 28198 45020 28250
rect 45072 28198 45144 28250
rect 45196 28198 45268 28250
rect 45320 28198 53896 28250
rect 53948 28198 54020 28250
rect 54072 28198 54144 28250
rect 54196 28198 54268 28250
rect 54320 28198 62896 28250
rect 62948 28198 63020 28250
rect 63072 28198 63144 28250
rect 63196 28198 63268 28250
rect 63320 28198 71896 28250
rect 71948 28198 72020 28250
rect 72072 28198 72144 28250
rect 72196 28198 72268 28250
rect 72320 28198 80896 28250
rect 80948 28198 81020 28250
rect 81072 28198 81144 28250
rect 81196 28198 81268 28250
rect 81320 28198 89896 28250
rect 89948 28198 90020 28250
rect 90072 28198 90144 28250
rect 90196 28198 90268 28250
rect 90320 28198 98560 28250
rect 1344 28164 98560 28198
rect 14478 28082 14530 28094
rect 33182 28082 33234 28094
rect 5058 28030 5070 28082
rect 5122 28030 5134 28082
rect 28242 28030 28254 28082
rect 28306 28030 28318 28082
rect 32050 28030 32062 28082
rect 32114 28030 32126 28082
rect 14478 28018 14530 28030
rect 33182 28018 33234 28030
rect 39902 28082 39954 28094
rect 44494 28082 44546 28094
rect 52894 28082 52946 28094
rect 43922 28030 43934 28082
rect 43986 28030 43998 28082
rect 51762 28030 51774 28082
rect 51826 28030 51838 28082
rect 39902 28018 39954 28030
rect 44494 28018 44546 28030
rect 52894 28018 52946 28030
rect 55022 28082 55074 28094
rect 66222 28082 66274 28094
rect 59602 28030 59614 28082
rect 59666 28030 59678 28082
rect 55022 28018 55074 28030
rect 66222 28018 66274 28030
rect 70478 28082 70530 28094
rect 70478 28018 70530 28030
rect 70702 28082 70754 28094
rect 70702 28018 70754 28030
rect 75742 28082 75794 28094
rect 75742 28018 75794 28030
rect 1934 27970 1986 27982
rect 14142 27970 14194 27982
rect 12450 27918 12462 27970
rect 12514 27918 12526 27970
rect 1934 27906 1986 27918
rect 14142 27906 14194 27918
rect 24670 27970 24722 27982
rect 24670 27906 24722 27918
rect 34862 27970 34914 27982
rect 34862 27906 34914 27918
rect 37998 27970 38050 27982
rect 37998 27906 38050 27918
rect 40350 27970 40402 27982
rect 40350 27906 40402 27918
rect 60174 27970 60226 27982
rect 60174 27906 60226 27918
rect 65662 27970 65714 27982
rect 65662 27906 65714 27918
rect 70814 27970 70866 27982
rect 70814 27906 70866 27918
rect 71262 27970 71314 27982
rect 71262 27906 71314 27918
rect 78878 27970 78930 27982
rect 78878 27906 78930 27918
rect 2158 27858 2210 27870
rect 13022 27858 13074 27870
rect 2706 27806 2718 27858
rect 2770 27806 2782 27858
rect 6066 27806 6078 27858
rect 6130 27806 6142 27858
rect 12226 27806 12238 27858
rect 12290 27806 12302 27858
rect 2158 27794 2210 27806
rect 13022 27794 13074 27806
rect 13358 27858 13410 27870
rect 13358 27794 13410 27806
rect 13806 27858 13858 27870
rect 25118 27858 25170 27870
rect 29150 27858 29202 27870
rect 35310 27858 35362 27870
rect 40798 27858 40850 27870
rect 48638 27858 48690 27870
rect 52446 27858 52498 27870
rect 24434 27806 24446 27858
rect 24498 27806 24510 27858
rect 25666 27806 25678 27858
rect 25730 27806 25742 27858
rect 29586 27806 29598 27858
rect 29650 27806 29662 27858
rect 35634 27806 35646 27858
rect 35698 27806 35710 27858
rect 41346 27806 41358 27858
rect 41410 27806 41422 27858
rect 46386 27806 46398 27858
rect 46450 27806 46462 27858
rect 49186 27806 49198 27858
rect 49250 27806 49262 27858
rect 13806 27794 13858 27806
rect 25118 27794 25170 27806
rect 29150 27794 29202 27806
rect 35310 27794 35362 27806
rect 40798 27794 40850 27806
rect 48638 27794 48690 27806
rect 52446 27794 52498 27806
rect 56478 27858 56530 27870
rect 65774 27858 65826 27870
rect 76190 27858 76242 27870
rect 57138 27806 57150 27858
rect 57202 27806 57214 27858
rect 73602 27806 73614 27858
rect 73666 27806 73678 27858
rect 76514 27806 76526 27858
rect 76578 27806 76590 27858
rect 56478 27794 56530 27806
rect 65774 27794 65826 27806
rect 76190 27794 76242 27806
rect 11790 27746 11842 27758
rect 46846 27746 46898 27758
rect 6738 27694 6750 27746
rect 6802 27694 6814 27746
rect 45714 27694 45726 27746
rect 45778 27694 45790 27746
rect 11790 27682 11842 27694
rect 46846 27682 46898 27694
rect 56030 27746 56082 27758
rect 56030 27682 56082 27694
rect 73166 27746 73218 27758
rect 74610 27694 74622 27746
rect 74674 27694 74686 27746
rect 73166 27682 73218 27694
rect 5854 27634 5906 27646
rect 5854 27570 5906 27582
rect 28814 27634 28866 27646
rect 28814 27570 28866 27582
rect 32622 27634 32674 27646
rect 32622 27570 32674 27582
rect 38782 27634 38834 27646
rect 38782 27570 38834 27582
rect 65662 27634 65714 27646
rect 65662 27570 65714 27582
rect 79662 27634 79714 27646
rect 79662 27570 79714 27582
rect 1344 27466 98560 27500
rect 1344 27414 4396 27466
rect 4448 27414 4520 27466
rect 4572 27414 4644 27466
rect 4696 27414 4768 27466
rect 4820 27414 13396 27466
rect 13448 27414 13520 27466
rect 13572 27414 13644 27466
rect 13696 27414 13768 27466
rect 13820 27414 22396 27466
rect 22448 27414 22520 27466
rect 22572 27414 22644 27466
rect 22696 27414 22768 27466
rect 22820 27414 31396 27466
rect 31448 27414 31520 27466
rect 31572 27414 31644 27466
rect 31696 27414 31768 27466
rect 31820 27414 40396 27466
rect 40448 27414 40520 27466
rect 40572 27414 40644 27466
rect 40696 27414 40768 27466
rect 40820 27414 49396 27466
rect 49448 27414 49520 27466
rect 49572 27414 49644 27466
rect 49696 27414 49768 27466
rect 49820 27414 58396 27466
rect 58448 27414 58520 27466
rect 58572 27414 58644 27466
rect 58696 27414 58768 27466
rect 58820 27414 67396 27466
rect 67448 27414 67520 27466
rect 67572 27414 67644 27466
rect 67696 27414 67768 27466
rect 67820 27414 76396 27466
rect 76448 27414 76520 27466
rect 76572 27414 76644 27466
rect 76696 27414 76768 27466
rect 76820 27414 85396 27466
rect 85448 27414 85520 27466
rect 85572 27414 85644 27466
rect 85696 27414 85768 27466
rect 85820 27414 94396 27466
rect 94448 27414 94520 27466
rect 94572 27414 94644 27466
rect 94696 27414 94768 27466
rect 94820 27414 98560 27466
rect 1344 27380 98560 27414
rect 17390 27298 17442 27310
rect 17390 27234 17442 27246
rect 31502 27298 31554 27310
rect 31502 27234 31554 27246
rect 37326 27298 37378 27310
rect 37326 27234 37378 27246
rect 56926 27298 56978 27310
rect 56926 27234 56978 27246
rect 57262 27298 57314 27310
rect 57262 27234 57314 27246
rect 57934 27298 57986 27310
rect 57934 27234 57986 27246
rect 66222 27298 66274 27310
rect 66222 27234 66274 27246
rect 17726 27186 17778 27198
rect 17726 27122 17778 27134
rect 20750 27186 20802 27198
rect 20750 27122 20802 27134
rect 29486 27186 29538 27198
rect 29486 27122 29538 27134
rect 29934 27186 29986 27198
rect 29934 27122 29986 27134
rect 32062 27186 32114 27198
rect 32062 27122 32114 27134
rect 37550 27186 37602 27198
rect 37550 27122 37602 27134
rect 38110 27186 38162 27198
rect 38110 27122 38162 27134
rect 53678 27186 53730 27198
rect 53678 27122 53730 27134
rect 59950 27186 60002 27198
rect 59950 27122 60002 27134
rect 73838 27186 73890 27198
rect 73838 27122 73890 27134
rect 76414 27186 76466 27198
rect 76414 27122 76466 27134
rect 96574 27186 96626 27198
rect 96574 27122 96626 27134
rect 1710 27074 1762 27086
rect 7310 27074 7362 27086
rect 13918 27074 13970 27086
rect 21758 27074 21810 27086
rect 31166 27074 31218 27086
rect 60846 27074 60898 27086
rect 2594 27022 2606 27074
rect 2658 27022 2670 27074
rect 7634 27022 7646 27074
rect 7698 27022 7710 27074
rect 14242 27022 14254 27074
rect 14306 27022 14318 27074
rect 30370 27022 30382 27074
rect 30434 27022 30446 27074
rect 35410 27022 35422 27074
rect 35474 27022 35486 27074
rect 57810 27022 57822 27074
rect 57874 27022 57886 27074
rect 1710 27010 1762 27022
rect 7310 27010 7362 27022
rect 13918 27010 13970 27022
rect 21758 27010 21810 27022
rect 31166 27010 31218 27022
rect 60846 27010 60898 27022
rect 61070 27074 61122 27086
rect 61070 27010 61122 27022
rect 61630 27074 61682 27086
rect 61630 27010 61682 27022
rect 62750 27074 62802 27086
rect 67230 27074 67282 27086
rect 76302 27074 76354 27086
rect 63074 27022 63086 27074
rect 63138 27022 63150 27074
rect 74274 27022 74286 27074
rect 74338 27022 74350 27074
rect 62750 27010 62802 27022
rect 67230 27010 67282 27022
rect 76302 27010 76354 27022
rect 76974 27074 77026 27086
rect 76974 27010 77026 27022
rect 77310 27074 77362 27086
rect 77310 27010 77362 27022
rect 96910 27074 96962 27086
rect 96910 27010 96962 27022
rect 2046 26962 2098 26974
rect 2046 26898 2098 26910
rect 3166 26962 3218 26974
rect 3166 26898 3218 26910
rect 5742 26962 5794 26974
rect 5742 26898 5794 26910
rect 9998 26962 10050 26974
rect 9998 26898 10050 26910
rect 16606 26962 16658 26974
rect 35646 26962 35698 26974
rect 60510 26962 60562 26974
rect 21970 26910 21982 26962
rect 22034 26910 22046 26962
rect 22306 26910 22318 26962
rect 22370 26910 22382 26962
rect 30482 26910 30494 26962
rect 30546 26910 30558 26962
rect 57922 26910 57934 26962
rect 57986 26910 57998 26962
rect 16606 26898 16658 26910
rect 35646 26898 35698 26910
rect 60510 26898 60562 26910
rect 60622 26962 60674 26974
rect 60622 26898 60674 26910
rect 61182 26962 61234 26974
rect 61182 26898 61234 26910
rect 61742 26962 61794 26974
rect 61742 26898 61794 26910
rect 61966 26962 62018 26974
rect 61966 26898 62018 26910
rect 62302 26962 62354 26974
rect 62302 26898 62354 26910
rect 65438 26962 65490 26974
rect 65438 26898 65490 26910
rect 67566 26962 67618 26974
rect 77534 26962 77586 26974
rect 75282 26910 75294 26962
rect 75346 26910 75358 26962
rect 67566 26898 67618 26910
rect 77534 26898 77586 26910
rect 77646 26962 77698 26974
rect 77646 26898 77698 26910
rect 78094 26962 78146 26974
rect 78094 26898 78146 26910
rect 97694 26962 97746 26974
rect 97694 26898 97746 26910
rect 2382 26850 2434 26862
rect 2382 26786 2434 26798
rect 10782 26850 10834 26862
rect 10782 26786 10834 26798
rect 19742 26850 19794 26862
rect 19742 26786 19794 26798
rect 21422 26850 21474 26862
rect 21422 26786 21474 26798
rect 23102 26850 23154 26862
rect 54238 26850 54290 26862
rect 36978 26798 36990 26850
rect 37042 26798 37054 26850
rect 23102 26786 23154 26798
rect 54238 26786 54290 26798
rect 57038 26850 57090 26862
rect 57038 26786 57090 26798
rect 61406 26850 61458 26862
rect 61406 26786 61458 26798
rect 76526 26850 76578 26862
rect 76526 26786 76578 26798
rect 1344 26682 98560 26716
rect 1344 26630 8896 26682
rect 8948 26630 9020 26682
rect 9072 26630 9144 26682
rect 9196 26630 9268 26682
rect 9320 26630 17896 26682
rect 17948 26630 18020 26682
rect 18072 26630 18144 26682
rect 18196 26630 18268 26682
rect 18320 26630 26896 26682
rect 26948 26630 27020 26682
rect 27072 26630 27144 26682
rect 27196 26630 27268 26682
rect 27320 26630 35896 26682
rect 35948 26630 36020 26682
rect 36072 26630 36144 26682
rect 36196 26630 36268 26682
rect 36320 26630 44896 26682
rect 44948 26630 45020 26682
rect 45072 26630 45144 26682
rect 45196 26630 45268 26682
rect 45320 26630 53896 26682
rect 53948 26630 54020 26682
rect 54072 26630 54144 26682
rect 54196 26630 54268 26682
rect 54320 26630 62896 26682
rect 62948 26630 63020 26682
rect 63072 26630 63144 26682
rect 63196 26630 63268 26682
rect 63320 26630 71896 26682
rect 71948 26630 72020 26682
rect 72072 26630 72144 26682
rect 72196 26630 72268 26682
rect 72320 26630 80896 26682
rect 80948 26630 81020 26682
rect 81072 26630 81144 26682
rect 81196 26630 81268 26682
rect 81320 26630 89896 26682
rect 89948 26630 90020 26682
rect 90072 26630 90144 26682
rect 90196 26630 90268 26682
rect 90320 26630 98560 26682
rect 1344 26596 98560 26630
rect 2494 26514 2546 26526
rect 2494 26450 2546 26462
rect 11454 26514 11506 26526
rect 11454 26450 11506 26462
rect 12014 26514 12066 26526
rect 12014 26450 12066 26462
rect 19182 26514 19234 26526
rect 23102 26514 23154 26526
rect 53566 26514 53618 26526
rect 22306 26462 22318 26514
rect 22370 26462 22382 26514
rect 52994 26462 53006 26514
rect 53058 26462 53070 26514
rect 19182 26450 19234 26462
rect 23102 26450 23154 26462
rect 53566 26450 53618 26462
rect 57598 26514 57650 26526
rect 57598 26450 57650 26462
rect 59614 26514 59666 26526
rect 59614 26450 59666 26462
rect 60062 26514 60114 26526
rect 60062 26450 60114 26462
rect 60846 26514 60898 26526
rect 60846 26450 60898 26462
rect 67118 26514 67170 26526
rect 67118 26450 67170 26462
rect 72494 26514 72546 26526
rect 72494 26450 72546 26462
rect 74734 26514 74786 26526
rect 74734 26450 74786 26462
rect 1934 26402 1986 26414
rect 1934 26338 1986 26350
rect 5294 26402 5346 26414
rect 5294 26338 5346 26350
rect 26686 26402 26738 26414
rect 26686 26338 26738 26350
rect 49646 26402 49698 26414
rect 58494 26402 58546 26414
rect 53778 26350 53790 26402
rect 53842 26350 53854 26402
rect 49646 26338 49698 26350
rect 58494 26338 58546 26350
rect 59950 26402 60002 26414
rect 59950 26338 60002 26350
rect 66670 26402 66722 26414
rect 66670 26338 66722 26350
rect 67342 26402 67394 26414
rect 67342 26338 67394 26350
rect 68126 26402 68178 26414
rect 68126 26338 68178 26350
rect 72718 26402 72770 26414
rect 72718 26338 72770 26350
rect 73502 26402 73554 26414
rect 73502 26338 73554 26350
rect 77086 26402 77138 26414
rect 77086 26338 77138 26350
rect 84254 26402 84306 26414
rect 84254 26338 84306 26350
rect 19630 26290 19682 26302
rect 49870 26290 49922 26302
rect 57038 26290 57090 26302
rect 20066 26238 20078 26290
rect 20130 26238 20142 26290
rect 26450 26238 26462 26290
rect 26514 26238 26526 26290
rect 50418 26238 50430 26290
rect 50482 26238 50494 26290
rect 19630 26226 19682 26238
rect 49870 26226 49922 26238
rect 57038 26226 57090 26238
rect 57934 26290 57986 26302
rect 57934 26226 57986 26238
rect 62302 26290 62354 26302
rect 62302 26226 62354 26238
rect 67790 26290 67842 26302
rect 67790 26226 67842 26238
rect 73166 26290 73218 26302
rect 75058 26238 75070 26290
rect 75122 26238 75134 26290
rect 84018 26238 84030 26290
rect 84082 26238 84094 26290
rect 73166 26226 73218 26238
rect 54798 26178 54850 26190
rect 10882 26126 10894 26178
rect 10946 26126 10958 26178
rect 54798 26114 54850 26126
rect 67230 26178 67282 26190
rect 67230 26114 67282 26126
rect 72606 26178 72658 26190
rect 77982 26178 78034 26190
rect 75730 26126 75742 26178
rect 75794 26126 75806 26178
rect 72606 26114 72658 26126
rect 77982 26114 78034 26126
rect 60062 26066 60114 26078
rect 60062 26002 60114 26014
rect 1344 25898 98560 25932
rect 1344 25846 4396 25898
rect 4448 25846 4520 25898
rect 4572 25846 4644 25898
rect 4696 25846 4768 25898
rect 4820 25846 13396 25898
rect 13448 25846 13520 25898
rect 13572 25846 13644 25898
rect 13696 25846 13768 25898
rect 13820 25846 22396 25898
rect 22448 25846 22520 25898
rect 22572 25846 22644 25898
rect 22696 25846 22768 25898
rect 22820 25846 31396 25898
rect 31448 25846 31520 25898
rect 31572 25846 31644 25898
rect 31696 25846 31768 25898
rect 31820 25846 40396 25898
rect 40448 25846 40520 25898
rect 40572 25846 40644 25898
rect 40696 25846 40768 25898
rect 40820 25846 49396 25898
rect 49448 25846 49520 25898
rect 49572 25846 49644 25898
rect 49696 25846 49768 25898
rect 49820 25846 58396 25898
rect 58448 25846 58520 25898
rect 58572 25846 58644 25898
rect 58696 25846 58768 25898
rect 58820 25846 67396 25898
rect 67448 25846 67520 25898
rect 67572 25846 67644 25898
rect 67696 25846 67768 25898
rect 67820 25846 76396 25898
rect 76448 25846 76520 25898
rect 76572 25846 76644 25898
rect 76696 25846 76768 25898
rect 76820 25846 85396 25898
rect 85448 25846 85520 25898
rect 85572 25846 85644 25898
rect 85696 25846 85768 25898
rect 85820 25846 94396 25898
rect 94448 25846 94520 25898
rect 94572 25846 94644 25898
rect 94696 25846 94768 25898
rect 94820 25846 98560 25898
rect 1344 25812 98560 25846
rect 27246 25730 27298 25742
rect 48414 25730 48466 25742
rect 35410 25678 35422 25730
rect 35474 25678 35486 25730
rect 27246 25666 27298 25678
rect 48414 25666 48466 25678
rect 57710 25730 57762 25742
rect 76066 25678 76078 25730
rect 76130 25727 76142 25730
rect 76738 25727 76750 25730
rect 76130 25681 76750 25727
rect 76130 25678 76142 25681
rect 76738 25678 76750 25681
rect 76802 25727 76814 25730
rect 77074 25727 77086 25730
rect 76802 25681 77086 25727
rect 76802 25678 76814 25681
rect 77074 25678 77086 25681
rect 77138 25678 77150 25730
rect 57710 25666 57762 25678
rect 25230 25618 25282 25630
rect 25230 25554 25282 25566
rect 25678 25618 25730 25630
rect 25678 25554 25730 25566
rect 53454 25618 53506 25630
rect 53454 25554 53506 25566
rect 58046 25618 58098 25630
rect 58046 25554 58098 25566
rect 65774 25618 65826 25630
rect 65774 25554 65826 25566
rect 69358 25618 69410 25630
rect 69358 25554 69410 25566
rect 76750 25618 76802 25630
rect 76750 25554 76802 25566
rect 5518 25506 5570 25518
rect 9214 25506 9266 25518
rect 6066 25454 6078 25506
rect 6130 25454 6142 25506
rect 5518 25442 5570 25454
rect 9214 25442 9266 25454
rect 11342 25506 11394 25518
rect 11342 25442 11394 25454
rect 20638 25506 20690 25518
rect 26910 25506 26962 25518
rect 26226 25454 26238 25506
rect 26290 25454 26302 25506
rect 20638 25442 20690 25454
rect 26910 25442 26962 25454
rect 34862 25506 34914 25518
rect 34862 25442 34914 25454
rect 35086 25506 35138 25518
rect 43150 25506 43202 25518
rect 44718 25506 44770 25518
rect 54238 25506 54290 25518
rect 62302 25506 62354 25518
rect 38882 25454 38894 25506
rect 38946 25454 38958 25506
rect 43362 25454 43374 25506
rect 43426 25454 43438 25506
rect 45266 25454 45278 25506
rect 45330 25454 45342 25506
rect 54562 25454 54574 25506
rect 54626 25454 54638 25506
rect 35086 25442 35138 25454
rect 43150 25442 43202 25454
rect 44718 25442 44770 25454
rect 54238 25442 54290 25454
rect 62302 25442 62354 25454
rect 62974 25506 63026 25518
rect 62974 25442 63026 25454
rect 64990 25506 65042 25518
rect 64990 25442 65042 25454
rect 65326 25506 65378 25518
rect 65326 25442 65378 25454
rect 68574 25506 68626 25518
rect 68574 25442 68626 25454
rect 68910 25506 68962 25518
rect 68910 25442 68962 25454
rect 72046 25506 72098 25518
rect 76302 25506 76354 25518
rect 72594 25454 72606 25506
rect 72658 25454 72670 25506
rect 72046 25442 72098 25454
rect 76302 25442 76354 25454
rect 77310 25506 77362 25518
rect 77310 25442 77362 25454
rect 77422 25506 77474 25518
rect 77422 25442 77474 25454
rect 77534 25506 77586 25518
rect 78430 25506 78482 25518
rect 77858 25454 77870 25506
rect 77922 25454 77934 25506
rect 78754 25454 78766 25506
rect 78818 25454 78830 25506
rect 77534 25442 77586 25454
rect 78430 25442 78482 25454
rect 1710 25394 1762 25406
rect 1710 25330 1762 25342
rect 2046 25394 2098 25406
rect 2046 25330 2098 25342
rect 2494 25394 2546 25406
rect 2494 25330 2546 25342
rect 8430 25394 8482 25406
rect 12350 25394 12402 25406
rect 10546 25342 10558 25394
rect 10610 25342 10622 25394
rect 11106 25342 11118 25394
rect 11170 25342 11182 25394
rect 8430 25330 8482 25342
rect 12350 25330 12402 25342
rect 20302 25394 20354 25406
rect 33070 25394 33122 25406
rect 26114 25342 26126 25394
rect 26178 25342 26190 25394
rect 20302 25330 20354 25342
rect 33070 25330 33122 25342
rect 43038 25394 43090 25406
rect 43038 25330 43090 25342
rect 43822 25394 43874 25406
rect 43822 25330 43874 25342
rect 44270 25394 44322 25406
rect 44270 25330 44322 25342
rect 71822 25394 71874 25406
rect 71822 25330 71874 25342
rect 81118 25394 81170 25406
rect 81118 25330 81170 25342
rect 9550 25282 9602 25294
rect 9550 25218 9602 25230
rect 11678 25282 11730 25294
rect 11678 25218 11730 25230
rect 12686 25282 12738 25294
rect 12686 25218 12738 25230
rect 27694 25282 27746 25294
rect 27694 25218 27746 25230
rect 28254 25282 28306 25294
rect 28254 25218 28306 25230
rect 33406 25282 33458 25294
rect 33406 25218 33458 25230
rect 34078 25282 34130 25294
rect 34078 25218 34130 25230
rect 34526 25282 34578 25294
rect 34526 25218 34578 25230
rect 39118 25282 39170 25294
rect 39118 25218 39170 25230
rect 39454 25282 39506 25294
rect 39454 25218 39506 25230
rect 42702 25282 42754 25294
rect 61854 25282 61906 25294
rect 47618 25230 47630 25282
rect 47682 25230 47694 25282
rect 57138 25230 57150 25282
rect 57202 25230 57214 25282
rect 42702 25218 42754 25230
rect 61854 25218 61906 25230
rect 62414 25282 62466 25294
rect 62414 25218 62466 25230
rect 62526 25282 62578 25294
rect 62526 25218 62578 25230
rect 63310 25282 63362 25294
rect 63310 25218 63362 25230
rect 65214 25282 65266 25294
rect 65214 25218 65266 25230
rect 68798 25282 68850 25294
rect 75742 25282 75794 25294
rect 75058 25230 75070 25282
rect 75122 25230 75134 25282
rect 68798 25218 68850 25230
rect 75742 25218 75794 25230
rect 81902 25282 81954 25294
rect 81902 25218 81954 25230
rect 1344 25114 98560 25148
rect 1344 25062 8896 25114
rect 8948 25062 9020 25114
rect 9072 25062 9144 25114
rect 9196 25062 9268 25114
rect 9320 25062 17896 25114
rect 17948 25062 18020 25114
rect 18072 25062 18144 25114
rect 18196 25062 18268 25114
rect 18320 25062 26896 25114
rect 26948 25062 27020 25114
rect 27072 25062 27144 25114
rect 27196 25062 27268 25114
rect 27320 25062 35896 25114
rect 35948 25062 36020 25114
rect 36072 25062 36144 25114
rect 36196 25062 36268 25114
rect 36320 25062 44896 25114
rect 44948 25062 45020 25114
rect 45072 25062 45144 25114
rect 45196 25062 45268 25114
rect 45320 25062 53896 25114
rect 53948 25062 54020 25114
rect 54072 25062 54144 25114
rect 54196 25062 54268 25114
rect 54320 25062 62896 25114
rect 62948 25062 63020 25114
rect 63072 25062 63144 25114
rect 63196 25062 63268 25114
rect 63320 25062 71896 25114
rect 71948 25062 72020 25114
rect 72072 25062 72144 25114
rect 72196 25062 72268 25114
rect 72320 25062 80896 25114
rect 80948 25062 81020 25114
rect 81072 25062 81144 25114
rect 81196 25062 81268 25114
rect 81320 25062 89896 25114
rect 89948 25062 90020 25114
rect 90072 25062 90144 25114
rect 90196 25062 90268 25114
rect 90320 25062 98560 25114
rect 1344 25028 98560 25062
rect 5294 24946 5346 24958
rect 11902 24946 11954 24958
rect 30158 24946 30210 24958
rect 4722 24894 4734 24946
rect 4786 24894 4798 24946
rect 10322 24894 10334 24946
rect 10386 24894 10398 24946
rect 29362 24894 29374 24946
rect 29426 24894 29438 24946
rect 5294 24882 5346 24894
rect 11902 24882 11954 24894
rect 30158 24882 30210 24894
rect 32062 24946 32114 24958
rect 32062 24882 32114 24894
rect 39566 24946 39618 24958
rect 39566 24882 39618 24894
rect 43038 24946 43090 24958
rect 43038 24882 43090 24894
rect 43374 24946 43426 24958
rect 43374 24882 43426 24894
rect 44270 24946 44322 24958
rect 44270 24882 44322 24894
rect 60174 24946 60226 24958
rect 60174 24882 60226 24894
rect 60622 24946 60674 24958
rect 60622 24882 60674 24894
rect 66334 24946 66386 24958
rect 66334 24882 66386 24894
rect 70254 24946 70306 24958
rect 70254 24882 70306 24894
rect 74174 24946 74226 24958
rect 74174 24882 74226 24894
rect 75070 24946 75122 24958
rect 75070 24882 75122 24894
rect 76974 24946 77026 24958
rect 76974 24882 77026 24894
rect 77758 24946 77810 24958
rect 77758 24882 77810 24894
rect 77870 24946 77922 24958
rect 77870 24882 77922 24894
rect 78094 24946 78146 24958
rect 78094 24882 78146 24894
rect 78542 24946 78594 24958
rect 78542 24882 78594 24894
rect 12462 24834 12514 24846
rect 10882 24782 10894 24834
rect 10946 24782 10958 24834
rect 12462 24770 12514 24782
rect 15598 24834 15650 24846
rect 15598 24770 15650 24782
rect 16606 24834 16658 24846
rect 16606 24770 16658 24782
rect 30494 24834 30546 24846
rect 30494 24770 30546 24782
rect 32510 24834 32562 24846
rect 32510 24770 32562 24782
rect 35870 24834 35922 24846
rect 35870 24770 35922 24782
rect 37550 24834 37602 24846
rect 60510 24834 60562 24846
rect 38546 24782 38558 24834
rect 38610 24782 38622 24834
rect 37550 24770 37602 24782
rect 60510 24770 60562 24782
rect 69470 24834 69522 24846
rect 69470 24770 69522 24782
rect 74398 24834 74450 24846
rect 74398 24770 74450 24782
rect 74510 24834 74562 24846
rect 74510 24770 74562 24782
rect 83134 24834 83186 24846
rect 83134 24770 83186 24782
rect 83470 24834 83522 24846
rect 83470 24770 83522 24782
rect 1822 24722 1874 24734
rect 5630 24722 5682 24734
rect 12686 24722 12738 24734
rect 26462 24722 26514 24734
rect 32958 24722 33010 24734
rect 36654 24722 36706 24734
rect 43486 24722 43538 24734
rect 78206 24722 78258 24734
rect 2258 24670 2270 24722
rect 2322 24670 2334 24722
rect 9762 24670 9774 24722
rect 9826 24670 9838 24722
rect 11666 24670 11678 24722
rect 11730 24670 11742 24722
rect 13234 24670 13246 24722
rect 13298 24670 13310 24722
rect 27010 24670 27022 24722
rect 27074 24670 27086 24722
rect 33618 24670 33630 24722
rect 33682 24670 33694 24722
rect 38434 24670 38446 24722
rect 38498 24670 38510 24722
rect 66658 24670 66670 24722
rect 66722 24670 66734 24722
rect 67218 24670 67230 24722
rect 67282 24670 67294 24722
rect 96898 24670 96910 24722
rect 96962 24670 96974 24722
rect 1822 24658 1874 24670
rect 5630 24658 5682 24670
rect 12686 24658 12738 24670
rect 26462 24658 26514 24670
rect 32958 24658 33010 24670
rect 36654 24658 36706 24670
rect 43486 24658 43538 24670
rect 78206 24658 78258 24670
rect 38110 24610 38162 24622
rect 38110 24546 38162 24558
rect 40238 24610 40290 24622
rect 98018 24558 98030 24610
rect 98082 24558 98094 24610
rect 40238 24546 40290 24558
rect 16382 24498 16434 24510
rect 16382 24434 16434 24446
rect 39230 24498 39282 24510
rect 39230 24434 39282 24446
rect 60622 24498 60674 24510
rect 60622 24434 60674 24446
rect 1344 24330 98560 24364
rect 1344 24278 4396 24330
rect 4448 24278 4520 24330
rect 4572 24278 4644 24330
rect 4696 24278 4768 24330
rect 4820 24278 13396 24330
rect 13448 24278 13520 24330
rect 13572 24278 13644 24330
rect 13696 24278 13768 24330
rect 13820 24278 22396 24330
rect 22448 24278 22520 24330
rect 22572 24278 22644 24330
rect 22696 24278 22768 24330
rect 22820 24278 31396 24330
rect 31448 24278 31520 24330
rect 31572 24278 31644 24330
rect 31696 24278 31768 24330
rect 31820 24278 40396 24330
rect 40448 24278 40520 24330
rect 40572 24278 40644 24330
rect 40696 24278 40768 24330
rect 40820 24278 49396 24330
rect 49448 24278 49520 24330
rect 49572 24278 49644 24330
rect 49696 24278 49768 24330
rect 49820 24278 58396 24330
rect 58448 24278 58520 24330
rect 58572 24278 58644 24330
rect 58696 24278 58768 24330
rect 58820 24278 67396 24330
rect 67448 24278 67520 24330
rect 67572 24278 67644 24330
rect 67696 24278 67768 24330
rect 67820 24278 76396 24330
rect 76448 24278 76520 24330
rect 76572 24278 76644 24330
rect 76696 24278 76768 24330
rect 76820 24278 85396 24330
rect 85448 24278 85520 24330
rect 85572 24278 85644 24330
rect 85696 24278 85768 24330
rect 85820 24278 94396 24330
rect 94448 24278 94520 24330
rect 94572 24278 94644 24330
rect 94696 24278 94768 24330
rect 94820 24278 98560 24330
rect 1344 24244 98560 24278
rect 33854 24162 33906 24174
rect 33854 24098 33906 24110
rect 34190 24162 34242 24174
rect 34190 24098 34242 24110
rect 3614 24050 3666 24062
rect 19630 24050 19682 24062
rect 11218 23998 11230 24050
rect 11282 23998 11294 24050
rect 3614 23986 3666 23998
rect 19630 23986 19682 23998
rect 20302 24050 20354 24062
rect 20302 23986 20354 23998
rect 34750 24050 34802 24062
rect 34750 23986 34802 23998
rect 59390 24050 59442 24062
rect 59390 23986 59442 23998
rect 1710 23938 1762 23950
rect 15822 23938 15874 23950
rect 22206 23938 22258 23950
rect 10882 23886 10894 23938
rect 10946 23886 10958 23938
rect 16146 23886 16158 23938
rect 16210 23886 16222 23938
rect 21522 23886 21534 23938
rect 21586 23886 21598 23938
rect 1710 23874 1762 23886
rect 15822 23874 15874 23886
rect 22206 23874 22258 23886
rect 38894 23938 38946 23950
rect 60510 23938 60562 23950
rect 39218 23886 39230 23938
rect 39282 23886 39294 23938
rect 38894 23874 38946 23886
rect 60510 23874 60562 23886
rect 61742 23938 61794 23950
rect 71150 23938 71202 23950
rect 62178 23886 62190 23938
rect 62242 23886 62254 23938
rect 61742 23874 61794 23886
rect 71150 23874 71202 23886
rect 76302 23938 76354 23950
rect 76302 23874 76354 23886
rect 2382 23826 2434 23838
rect 32622 23826 32674 23838
rect 59726 23826 59778 23838
rect 10434 23774 10446 23826
rect 10498 23774 10510 23826
rect 21410 23774 21422 23826
rect 21474 23774 21486 23826
rect 33058 23774 33070 23826
rect 33122 23774 33134 23826
rect 33506 23774 33518 23826
rect 33570 23774 33582 23826
rect 2382 23762 2434 23774
rect 32622 23762 32674 23774
rect 59726 23762 59778 23774
rect 59838 23826 59890 23838
rect 59838 23762 59890 23774
rect 61070 23826 61122 23838
rect 61070 23762 61122 23774
rect 61182 23826 61234 23838
rect 61182 23762 61234 23774
rect 2046 23714 2098 23726
rect 2046 23650 2098 23662
rect 2718 23714 2770 23726
rect 2718 23650 2770 23662
rect 3166 23714 3218 23726
rect 3166 23650 3218 23662
rect 12462 23714 12514 23726
rect 19294 23714 19346 23726
rect 18722 23662 18734 23714
rect 18786 23662 18798 23714
rect 12462 23650 12514 23662
rect 19294 23650 19346 23662
rect 20638 23714 20690 23726
rect 20638 23650 20690 23662
rect 22542 23714 22594 23726
rect 22542 23650 22594 23662
rect 23102 23714 23154 23726
rect 23102 23650 23154 23662
rect 26910 23714 26962 23726
rect 26910 23650 26962 23662
rect 32174 23714 32226 23726
rect 32174 23650 32226 23662
rect 38446 23714 38498 23726
rect 42366 23714 42418 23726
rect 41570 23662 41582 23714
rect 41634 23662 41646 23714
rect 38446 23650 38498 23662
rect 42366 23650 42418 23662
rect 60062 23714 60114 23726
rect 60062 23650 60114 23662
rect 60622 23714 60674 23726
rect 60622 23650 60674 23662
rect 60846 23714 60898 23726
rect 60846 23650 60898 23662
rect 61406 23714 61458 23726
rect 65214 23714 65266 23726
rect 64642 23662 64654 23714
rect 64706 23662 64718 23714
rect 61406 23650 61458 23662
rect 65214 23650 65266 23662
rect 65550 23714 65602 23726
rect 65550 23650 65602 23662
rect 71486 23714 71538 23726
rect 71486 23650 71538 23662
rect 76638 23714 76690 23726
rect 76638 23650 76690 23662
rect 1344 23546 98560 23580
rect 1344 23494 8896 23546
rect 8948 23494 9020 23546
rect 9072 23494 9144 23546
rect 9196 23494 9268 23546
rect 9320 23494 17896 23546
rect 17948 23494 18020 23546
rect 18072 23494 18144 23546
rect 18196 23494 18268 23546
rect 18320 23494 26896 23546
rect 26948 23494 27020 23546
rect 27072 23494 27144 23546
rect 27196 23494 27268 23546
rect 27320 23494 35896 23546
rect 35948 23494 36020 23546
rect 36072 23494 36144 23546
rect 36196 23494 36268 23546
rect 36320 23494 44896 23546
rect 44948 23494 45020 23546
rect 45072 23494 45144 23546
rect 45196 23494 45268 23546
rect 45320 23494 53896 23546
rect 53948 23494 54020 23546
rect 54072 23494 54144 23546
rect 54196 23494 54268 23546
rect 54320 23494 62896 23546
rect 62948 23494 63020 23546
rect 63072 23494 63144 23546
rect 63196 23494 63268 23546
rect 63320 23494 71896 23546
rect 71948 23494 72020 23546
rect 72072 23494 72144 23546
rect 72196 23494 72268 23546
rect 72320 23494 80896 23546
rect 80948 23494 81020 23546
rect 81072 23494 81144 23546
rect 81196 23494 81268 23546
rect 81320 23494 89896 23546
rect 89948 23494 90020 23546
rect 90072 23494 90144 23546
rect 90196 23494 90268 23546
rect 90320 23494 98560 23546
rect 1344 23460 98560 23494
rect 6078 23378 6130 23390
rect 26350 23378 26402 23390
rect 30606 23378 30658 23390
rect 4722 23326 4734 23378
rect 4786 23326 4798 23378
rect 10098 23326 10110 23378
rect 10162 23326 10174 23378
rect 29474 23326 29486 23378
rect 29538 23326 29550 23378
rect 6078 23314 6130 23326
rect 26350 23314 26402 23326
rect 30606 23314 30658 23326
rect 60286 23378 60338 23390
rect 60286 23314 60338 23326
rect 60846 23378 60898 23390
rect 60846 23314 60898 23326
rect 62302 23378 62354 23390
rect 62302 23314 62354 23326
rect 62526 23378 62578 23390
rect 62526 23314 62578 23326
rect 63310 23378 63362 23390
rect 63310 23314 63362 23326
rect 65998 23378 66050 23390
rect 73502 23378 73554 23390
rect 69794 23326 69806 23378
rect 69858 23326 69870 23378
rect 65998 23314 66050 23326
rect 73502 23314 73554 23326
rect 77422 23378 77474 23390
rect 77422 23314 77474 23326
rect 77982 23378 78034 23390
rect 77982 23314 78034 23326
rect 81006 23378 81058 23390
rect 81006 23314 81058 23326
rect 82238 23378 82290 23390
rect 82238 23314 82290 23326
rect 96574 23378 96626 23390
rect 96574 23314 96626 23326
rect 5294 23266 5346 23278
rect 5294 23202 5346 23214
rect 5630 23266 5682 23278
rect 20302 23266 20354 23278
rect 10210 23214 10222 23266
rect 10274 23214 10286 23266
rect 5630 23202 5682 23214
rect 20302 23202 20354 23214
rect 23438 23266 23490 23278
rect 23438 23202 23490 23214
rect 46062 23266 46114 23278
rect 46062 23202 46114 23214
rect 66334 23266 66386 23278
rect 66334 23202 66386 23214
rect 66670 23266 66722 23278
rect 66670 23202 66722 23214
rect 72942 23266 72994 23278
rect 72942 23202 72994 23214
rect 73726 23266 73778 23278
rect 73726 23202 73778 23214
rect 74510 23266 74562 23278
rect 74510 23202 74562 23214
rect 77758 23266 77810 23278
rect 77758 23202 77810 23214
rect 78654 23266 78706 23278
rect 78654 23202 78706 23214
rect 85710 23266 85762 23278
rect 85710 23202 85762 23214
rect 1822 23154 1874 23166
rect 24222 23154 24274 23166
rect 2258 23102 2270 23154
rect 2322 23102 2334 23154
rect 10882 23102 10894 23154
rect 10946 23102 10958 23154
rect 20626 23102 20638 23154
rect 20690 23102 20702 23154
rect 21186 23102 21198 23154
rect 21250 23102 21262 23154
rect 1822 23090 1874 23102
rect 24222 23090 24274 23102
rect 26574 23154 26626 23166
rect 45166 23154 45218 23166
rect 27122 23102 27134 23154
rect 27186 23102 27198 23154
rect 26574 23090 26626 23102
rect 45166 23090 45218 23102
rect 45950 23154 46002 23166
rect 45950 23090 46002 23102
rect 46286 23154 46338 23166
rect 46286 23090 46338 23102
rect 62974 23154 63026 23166
rect 62974 23090 63026 23102
rect 67118 23154 67170 23166
rect 74174 23154 74226 23166
rect 67554 23102 67566 23154
rect 67618 23102 67630 23154
rect 67118 23090 67170 23102
rect 74174 23090 74226 23102
rect 78430 23154 78482 23166
rect 78430 23090 78482 23102
rect 82014 23154 82066 23166
rect 82014 23090 82066 23102
rect 82126 23154 82178 23166
rect 82126 23090 82178 23102
rect 82686 23154 82738 23166
rect 82686 23090 82738 23102
rect 83022 23154 83074 23166
rect 83346 23102 83358 23154
rect 83410 23102 83422 23154
rect 96898 23102 96910 23154
rect 96962 23102 96974 23154
rect 83022 23090 83074 23102
rect 45614 23042 45666 23054
rect 45614 22978 45666 22990
rect 62414 23042 62466 23054
rect 62414 22978 62466 22990
rect 73614 23042 73666 23054
rect 73614 22978 73666 22990
rect 77870 23042 77922 23054
rect 77870 22978 77922 22990
rect 81454 23042 81506 23054
rect 98018 22990 98030 23042
rect 98082 22990 98094 23042
rect 81454 22978 81506 22990
rect 30270 22930 30322 22942
rect 30270 22866 30322 22878
rect 70590 22930 70642 22942
rect 70590 22866 70642 22878
rect 86494 22930 86546 22942
rect 86494 22866 86546 22878
rect 1344 22762 98560 22796
rect 1344 22710 4396 22762
rect 4448 22710 4520 22762
rect 4572 22710 4644 22762
rect 4696 22710 4768 22762
rect 4820 22710 13396 22762
rect 13448 22710 13520 22762
rect 13572 22710 13644 22762
rect 13696 22710 13768 22762
rect 13820 22710 22396 22762
rect 22448 22710 22520 22762
rect 22572 22710 22644 22762
rect 22696 22710 22768 22762
rect 22820 22710 31396 22762
rect 31448 22710 31520 22762
rect 31572 22710 31644 22762
rect 31696 22710 31768 22762
rect 31820 22710 40396 22762
rect 40448 22710 40520 22762
rect 40572 22710 40644 22762
rect 40696 22710 40768 22762
rect 40820 22710 49396 22762
rect 49448 22710 49520 22762
rect 49572 22710 49644 22762
rect 49696 22710 49768 22762
rect 49820 22710 58396 22762
rect 58448 22710 58520 22762
rect 58572 22710 58644 22762
rect 58696 22710 58768 22762
rect 58820 22710 67396 22762
rect 67448 22710 67520 22762
rect 67572 22710 67644 22762
rect 67696 22710 67768 22762
rect 67820 22710 76396 22762
rect 76448 22710 76520 22762
rect 76572 22710 76644 22762
rect 76696 22710 76768 22762
rect 76820 22710 85396 22762
rect 85448 22710 85520 22762
rect 85572 22710 85644 22762
rect 85696 22710 85768 22762
rect 85820 22710 94396 22762
rect 94448 22710 94520 22762
rect 94572 22710 94644 22762
rect 94696 22710 94768 22762
rect 94820 22710 98560 22762
rect 1344 22676 98560 22710
rect 9214 22594 9266 22606
rect 9214 22530 9266 22542
rect 65662 22594 65714 22606
rect 65662 22530 65714 22542
rect 9550 22482 9602 22494
rect 9550 22418 9602 22430
rect 38110 22482 38162 22494
rect 38110 22418 38162 22430
rect 68462 22482 68514 22494
rect 68462 22418 68514 22430
rect 69918 22482 69970 22494
rect 69918 22418 69970 22430
rect 76302 22482 76354 22494
rect 76302 22418 76354 22430
rect 77758 22482 77810 22494
rect 77758 22418 77810 22430
rect 21646 22370 21698 22382
rect 39342 22370 39394 22382
rect 5618 22318 5630 22370
rect 5682 22318 5694 22370
rect 6066 22318 6078 22370
rect 6130 22318 6142 22370
rect 10882 22318 10894 22370
rect 10946 22318 10958 22370
rect 33618 22318 33630 22370
rect 33682 22318 33694 22370
rect 38546 22318 38558 22370
rect 38610 22318 38622 22370
rect 21646 22306 21698 22318
rect 39342 22306 39394 22318
rect 64318 22370 64370 22382
rect 68350 22370 68402 22382
rect 64642 22318 64654 22370
rect 64706 22318 64718 22370
rect 64318 22306 64370 22318
rect 68350 22306 68402 22318
rect 68574 22370 68626 22382
rect 69134 22370 69186 22382
rect 78206 22370 78258 22382
rect 82574 22370 82626 22382
rect 68898 22318 68910 22370
rect 68962 22318 68974 22370
rect 72146 22318 72158 22370
rect 72210 22318 72222 22370
rect 72706 22318 72718 22370
rect 72770 22318 72782 22370
rect 78530 22318 78542 22370
rect 78594 22318 78606 22370
rect 68574 22306 68626 22318
rect 69134 22306 69186 22318
rect 78206 22306 78258 22318
rect 82574 22306 82626 22318
rect 84926 22370 84978 22382
rect 84926 22306 84978 22318
rect 1710 22258 1762 22270
rect 1710 22194 1762 22206
rect 2382 22258 2434 22270
rect 2382 22194 2434 22206
rect 8430 22258 8482 22270
rect 21310 22258 21362 22270
rect 67118 22258 67170 22270
rect 10770 22206 10782 22258
rect 10834 22206 10846 22258
rect 27794 22206 27806 22258
rect 27858 22206 27870 22258
rect 28578 22206 28590 22258
rect 28642 22206 28654 22258
rect 38658 22206 38670 22258
rect 38722 22206 38734 22258
rect 8430 22194 8482 22206
rect 21310 22194 21362 22206
rect 67118 22194 67170 22206
rect 69358 22258 69410 22270
rect 69358 22194 69410 22206
rect 69470 22258 69522 22270
rect 69470 22194 69522 22206
rect 83134 22258 83186 22270
rect 83134 22194 83186 22206
rect 84590 22258 84642 22270
rect 84590 22194 84642 22206
rect 84814 22258 84866 22270
rect 84814 22194 84866 22206
rect 2046 22146 2098 22158
rect 2046 22082 2098 22094
rect 2942 22146 2994 22158
rect 14590 22146 14642 22158
rect 11666 22094 11678 22146
rect 11730 22094 11742 22146
rect 2942 22082 2994 22094
rect 14590 22082 14642 22094
rect 14926 22146 14978 22158
rect 14926 22082 14978 22094
rect 29150 22146 29202 22158
rect 29150 22082 29202 22094
rect 29710 22146 29762 22158
rect 29710 22082 29762 22094
rect 33854 22146 33906 22158
rect 33854 22082 33906 22094
rect 34190 22146 34242 22158
rect 34190 22082 34242 22094
rect 39678 22146 39730 22158
rect 39678 22082 39730 22094
rect 40126 22146 40178 22158
rect 40126 22082 40178 22094
rect 61854 22146 61906 22158
rect 61854 22082 61906 22094
rect 70366 22146 70418 22158
rect 75742 22146 75794 22158
rect 81678 22146 81730 22158
rect 75058 22094 75070 22146
rect 75122 22094 75134 22146
rect 80882 22094 80894 22146
rect 80946 22094 80958 22146
rect 70366 22082 70418 22094
rect 75742 22082 75794 22094
rect 81678 22082 81730 22094
rect 84366 22146 84418 22158
rect 84366 22082 84418 22094
rect 1344 21978 98560 22012
rect 1344 21926 8896 21978
rect 8948 21926 9020 21978
rect 9072 21926 9144 21978
rect 9196 21926 9268 21978
rect 9320 21926 17896 21978
rect 17948 21926 18020 21978
rect 18072 21926 18144 21978
rect 18196 21926 18268 21978
rect 18320 21926 26896 21978
rect 26948 21926 27020 21978
rect 27072 21926 27144 21978
rect 27196 21926 27268 21978
rect 27320 21926 35896 21978
rect 35948 21926 36020 21978
rect 36072 21926 36144 21978
rect 36196 21926 36268 21978
rect 36320 21926 44896 21978
rect 44948 21926 45020 21978
rect 45072 21926 45144 21978
rect 45196 21926 45268 21978
rect 45320 21926 53896 21978
rect 53948 21926 54020 21978
rect 54072 21926 54144 21978
rect 54196 21926 54268 21978
rect 54320 21926 62896 21978
rect 62948 21926 63020 21978
rect 63072 21926 63144 21978
rect 63196 21926 63268 21978
rect 63320 21926 71896 21978
rect 71948 21926 72020 21978
rect 72072 21926 72144 21978
rect 72196 21926 72268 21978
rect 72320 21926 80896 21978
rect 80948 21926 81020 21978
rect 81072 21926 81144 21978
rect 81196 21926 81268 21978
rect 81320 21926 89896 21978
rect 89948 21926 90020 21978
rect 90072 21926 90144 21978
rect 90196 21926 90268 21978
rect 90320 21926 98560 21978
rect 1344 21892 98560 21926
rect 8990 21810 9042 21822
rect 43374 21810 43426 21822
rect 13010 21758 13022 21810
rect 13074 21758 13086 21810
rect 31938 21758 31950 21810
rect 32002 21758 32014 21810
rect 8990 21746 9042 21758
rect 43374 21746 43426 21758
rect 43822 21810 43874 21822
rect 43822 21746 43874 21758
rect 64318 21810 64370 21822
rect 64318 21746 64370 21758
rect 74958 21810 75010 21822
rect 74958 21746 75010 21758
rect 80222 21810 80274 21822
rect 80222 21746 80274 21758
rect 96574 21810 96626 21822
rect 96574 21746 96626 21758
rect 2046 21698 2098 21710
rect 2046 21634 2098 21646
rect 9886 21698 9938 21710
rect 9886 21634 9938 21646
rect 13806 21698 13858 21710
rect 13806 21634 13858 21646
rect 14590 21698 14642 21710
rect 25230 21698 25282 21710
rect 15138 21646 15150 21698
rect 15202 21646 15214 21698
rect 15586 21646 15598 21698
rect 15650 21646 15662 21698
rect 14590 21634 14642 21646
rect 25230 21634 25282 21646
rect 36206 21698 36258 21710
rect 36206 21634 36258 21646
rect 39342 21698 39394 21710
rect 39342 21634 39394 21646
rect 64542 21698 64594 21710
rect 64542 21634 64594 21646
rect 64654 21698 64706 21710
rect 64654 21634 64706 21646
rect 65102 21698 65154 21710
rect 65102 21634 65154 21646
rect 75182 21698 75234 21710
rect 75182 21634 75234 21646
rect 80446 21698 80498 21710
rect 80446 21634 80498 21646
rect 87054 21698 87106 21710
rect 87054 21634 87106 21646
rect 87390 21698 87442 21710
rect 87390 21634 87442 21646
rect 1710 21586 1762 21598
rect 10110 21586 10162 21598
rect 16158 21586 16210 21598
rect 29038 21586 29090 21598
rect 43710 21586 43762 21598
rect 6402 21534 6414 21586
rect 6466 21534 6478 21586
rect 10658 21534 10670 21586
rect 10722 21534 10734 21586
rect 14354 21534 14366 21586
rect 14418 21534 14430 21586
rect 17826 21534 17838 21586
rect 17890 21534 17902 21586
rect 27346 21534 27358 21586
rect 27410 21534 27422 21586
rect 29362 21534 29374 21586
rect 29426 21534 29438 21586
rect 33394 21534 33406 21586
rect 33458 21534 33470 21586
rect 33842 21534 33854 21586
rect 33906 21534 33918 21586
rect 39106 21534 39118 21586
rect 39170 21534 39182 21586
rect 1710 21522 1762 21534
rect 10110 21522 10162 21534
rect 16158 21522 16210 21534
rect 29038 21522 29090 21534
rect 43710 21522 43762 21534
rect 75294 21586 75346 21598
rect 75294 21522 75346 21534
rect 80558 21586 80610 21598
rect 80558 21522 80610 21534
rect 81006 21586 81058 21598
rect 96898 21534 96910 21586
rect 96962 21534 96974 21586
rect 81006 21522 81058 21534
rect 2494 21474 2546 21486
rect 2494 21410 2546 21422
rect 6862 21474 6914 21486
rect 6862 21410 6914 21422
rect 16830 21474 16882 21486
rect 16830 21410 16882 21422
rect 17502 21474 17554 21486
rect 26574 21474 26626 21486
rect 18722 21422 18734 21474
rect 18786 21422 18798 21474
rect 17502 21410 17554 21422
rect 26574 21410 26626 21422
rect 27022 21474 27074 21486
rect 27022 21410 27074 21422
rect 28366 21474 28418 21486
rect 28366 21410 28418 21422
rect 75742 21474 75794 21486
rect 98018 21422 98030 21474
rect 98082 21422 98094 21474
rect 75742 21410 75794 21422
rect 5854 21362 5906 21374
rect 5854 21298 5906 21310
rect 15822 21362 15874 21374
rect 15822 21298 15874 21310
rect 32510 21362 32562 21374
rect 32510 21298 32562 21310
rect 36990 21362 37042 21374
rect 36990 21298 37042 21310
rect 43822 21362 43874 21374
rect 43822 21298 43874 21310
rect 1344 21194 98560 21228
rect 1344 21142 4396 21194
rect 4448 21142 4520 21194
rect 4572 21142 4644 21194
rect 4696 21142 4768 21194
rect 4820 21142 13396 21194
rect 13448 21142 13520 21194
rect 13572 21142 13644 21194
rect 13696 21142 13768 21194
rect 13820 21142 22396 21194
rect 22448 21142 22520 21194
rect 22572 21142 22644 21194
rect 22696 21142 22768 21194
rect 22820 21142 31396 21194
rect 31448 21142 31520 21194
rect 31572 21142 31644 21194
rect 31696 21142 31768 21194
rect 31820 21142 40396 21194
rect 40448 21142 40520 21194
rect 40572 21142 40644 21194
rect 40696 21142 40768 21194
rect 40820 21142 49396 21194
rect 49448 21142 49520 21194
rect 49572 21142 49644 21194
rect 49696 21142 49768 21194
rect 49820 21142 58396 21194
rect 58448 21142 58520 21194
rect 58572 21142 58644 21194
rect 58696 21142 58768 21194
rect 58820 21142 67396 21194
rect 67448 21142 67520 21194
rect 67572 21142 67644 21194
rect 67696 21142 67768 21194
rect 67820 21142 76396 21194
rect 76448 21142 76520 21194
rect 76572 21142 76644 21194
rect 76696 21142 76768 21194
rect 76820 21142 85396 21194
rect 85448 21142 85520 21194
rect 85572 21142 85644 21194
rect 85696 21142 85768 21194
rect 85820 21142 94396 21194
rect 94448 21142 94520 21194
rect 94572 21142 94644 21194
rect 94696 21142 94768 21194
rect 94820 21142 98560 21194
rect 1344 21108 98560 21142
rect 9886 21026 9938 21038
rect 9886 20962 9938 20974
rect 30158 21026 30210 21038
rect 30158 20962 30210 20974
rect 34750 21026 34802 21038
rect 34750 20962 34802 20974
rect 42926 21026 42978 21038
rect 42926 20962 42978 20974
rect 65214 21026 65266 21038
rect 65214 20962 65266 20974
rect 74846 21026 74898 21038
rect 74846 20962 74898 20974
rect 4286 20914 4338 20926
rect 4286 20850 4338 20862
rect 18398 20914 18450 20926
rect 18398 20850 18450 20862
rect 18734 20914 18786 20926
rect 18734 20850 18786 20862
rect 32622 20914 32674 20926
rect 32622 20850 32674 20862
rect 33070 20914 33122 20926
rect 33070 20850 33122 20862
rect 39006 20914 39058 20926
rect 39006 20850 39058 20862
rect 43486 20914 43538 20926
rect 43486 20850 43538 20862
rect 55470 20914 55522 20926
rect 55470 20850 55522 20862
rect 56702 20914 56754 20926
rect 56702 20850 56754 20862
rect 65550 20914 65602 20926
rect 65550 20850 65602 20862
rect 73726 20914 73778 20926
rect 73726 20850 73778 20862
rect 80670 20914 80722 20926
rect 80670 20850 80722 20862
rect 84366 20914 84418 20926
rect 84366 20850 84418 20862
rect 6190 20802 6242 20814
rect 14926 20802 14978 20814
rect 22990 20802 23042 20814
rect 4610 20750 4622 20802
rect 4674 20750 4686 20802
rect 6738 20750 6750 20802
rect 6802 20750 6814 20802
rect 15250 20750 15262 20802
rect 15314 20750 15326 20802
rect 6190 20738 6242 20750
rect 14926 20738 14978 20750
rect 22990 20738 23042 20750
rect 24222 20802 24274 20814
rect 24222 20738 24274 20750
rect 25118 20802 25170 20814
rect 28590 20802 28642 20814
rect 34414 20802 34466 20814
rect 25554 20750 25566 20802
rect 25618 20750 25630 20802
rect 29138 20750 29150 20802
rect 29202 20750 29214 20802
rect 33730 20750 33742 20802
rect 33794 20750 33806 20802
rect 25118 20738 25170 20750
rect 28590 20738 28642 20750
rect 34414 20738 34466 20750
rect 39230 20802 39282 20814
rect 43822 20802 43874 20814
rect 39778 20750 39790 20802
rect 39842 20750 39854 20802
rect 39230 20738 39282 20750
rect 43822 20738 43874 20750
rect 56030 20802 56082 20814
rect 56030 20738 56082 20750
rect 56366 20802 56418 20814
rect 56366 20738 56418 20750
rect 61742 20802 61794 20814
rect 72046 20802 72098 20814
rect 62178 20750 62190 20802
rect 62242 20750 62254 20802
rect 61742 20738 61794 20750
rect 72046 20738 72098 20750
rect 72718 20802 72770 20814
rect 84926 20802 84978 20814
rect 74162 20750 74174 20802
rect 74226 20750 74238 20802
rect 72718 20738 72770 20750
rect 84926 20738 84978 20750
rect 85598 20802 85650 20814
rect 85598 20738 85650 20750
rect 5070 20690 5122 20702
rect 5070 20626 5122 20638
rect 5966 20690 6018 20702
rect 5966 20626 6018 20638
rect 9102 20690 9154 20702
rect 27806 20690 27858 20702
rect 42142 20690 42194 20702
rect 23426 20638 23438 20690
rect 23490 20638 23502 20690
rect 23986 20638 23998 20690
rect 24050 20638 24062 20690
rect 33618 20638 33630 20690
rect 33682 20638 33694 20690
rect 9102 20626 9154 20638
rect 27806 20626 27858 20638
rect 42142 20626 42194 20638
rect 43934 20690 43986 20702
rect 43934 20626 43986 20638
rect 56142 20690 56194 20702
rect 56142 20626 56194 20638
rect 1934 20578 1986 20590
rect 19070 20578 19122 20590
rect 17826 20526 17838 20578
rect 17890 20526 17902 20578
rect 1934 20514 1986 20526
rect 19070 20514 19122 20526
rect 24558 20578 24610 20590
rect 24558 20514 24610 20526
rect 44158 20578 44210 20590
rect 72158 20578 72210 20590
rect 64642 20526 64654 20578
rect 64706 20526 64718 20578
rect 44158 20514 44210 20526
rect 72158 20514 72210 20526
rect 72270 20578 72322 20590
rect 72270 20514 72322 20526
rect 73054 20578 73106 20590
rect 73054 20514 73106 20526
rect 76302 20578 76354 20590
rect 76302 20514 76354 20526
rect 85038 20578 85090 20590
rect 85038 20514 85090 20526
rect 85150 20578 85202 20590
rect 85150 20514 85202 20526
rect 1344 20410 98560 20444
rect 1344 20358 8896 20410
rect 8948 20358 9020 20410
rect 9072 20358 9144 20410
rect 9196 20358 9268 20410
rect 9320 20358 17896 20410
rect 17948 20358 18020 20410
rect 18072 20358 18144 20410
rect 18196 20358 18268 20410
rect 18320 20358 26896 20410
rect 26948 20358 27020 20410
rect 27072 20358 27144 20410
rect 27196 20358 27268 20410
rect 27320 20358 35896 20410
rect 35948 20358 36020 20410
rect 36072 20358 36144 20410
rect 36196 20358 36268 20410
rect 36320 20358 44896 20410
rect 44948 20358 45020 20410
rect 45072 20358 45144 20410
rect 45196 20358 45268 20410
rect 45320 20358 53896 20410
rect 53948 20358 54020 20410
rect 54072 20358 54144 20410
rect 54196 20358 54268 20410
rect 54320 20358 62896 20410
rect 62948 20358 63020 20410
rect 63072 20358 63144 20410
rect 63196 20358 63268 20410
rect 63320 20358 71896 20410
rect 71948 20358 72020 20410
rect 72072 20358 72144 20410
rect 72196 20358 72268 20410
rect 72320 20358 80896 20410
rect 80948 20358 81020 20410
rect 81072 20358 81144 20410
rect 81196 20358 81268 20410
rect 81320 20358 89896 20410
rect 89948 20358 90020 20410
rect 90072 20358 90144 20410
rect 90196 20358 90268 20410
rect 90320 20358 98560 20410
rect 1344 20324 98560 20358
rect 18174 20242 18226 20254
rect 25566 20242 25618 20254
rect 21746 20190 21758 20242
rect 21810 20190 21822 20242
rect 18174 20178 18226 20190
rect 25566 20178 25618 20190
rect 28926 20242 28978 20254
rect 28926 20178 28978 20190
rect 73166 20242 73218 20254
rect 73166 20178 73218 20190
rect 75518 20242 75570 20254
rect 75518 20178 75570 20190
rect 76302 20242 76354 20254
rect 76302 20178 76354 20190
rect 81230 20242 81282 20254
rect 81230 20178 81282 20190
rect 81902 20242 81954 20254
rect 81902 20178 81954 20190
rect 86046 20242 86098 20254
rect 86046 20178 86098 20190
rect 4510 20130 4562 20142
rect 4510 20066 4562 20078
rect 5294 20130 5346 20142
rect 5294 20066 5346 20078
rect 22430 20130 22482 20142
rect 22430 20066 22482 20078
rect 28478 20130 28530 20142
rect 28478 20066 28530 20078
rect 29374 20130 29426 20142
rect 29374 20066 29426 20078
rect 39902 20130 39954 20142
rect 39902 20066 39954 20078
rect 40126 20130 40178 20142
rect 40126 20066 40178 20078
rect 40238 20130 40290 20142
rect 40238 20066 40290 20078
rect 65886 20130 65938 20142
rect 65886 20066 65938 20078
rect 66222 20130 66274 20142
rect 66222 20066 66274 20078
rect 71038 20130 71090 20142
rect 71038 20066 71090 20078
rect 73390 20130 73442 20142
rect 73390 20066 73442 20078
rect 73502 20130 73554 20142
rect 75966 20130 76018 20142
rect 75058 20078 75070 20130
rect 75122 20078 75134 20130
rect 73502 20066 73554 20078
rect 75966 20066 76018 20078
rect 78094 20130 78146 20142
rect 78094 20066 78146 20078
rect 78206 20130 78258 20142
rect 78206 20066 78258 20078
rect 78766 20130 78818 20142
rect 78766 20066 78818 20078
rect 82910 20130 82962 20142
rect 82910 20066 82962 20078
rect 83246 20130 83298 20142
rect 83246 20066 83298 20078
rect 83358 20130 83410 20142
rect 83358 20066 83410 20078
rect 85598 20130 85650 20142
rect 85598 20066 85650 20078
rect 85822 20130 85874 20142
rect 85822 20066 85874 20078
rect 1822 20018 1874 20030
rect 18958 20018 19010 20030
rect 40462 20018 40514 20030
rect 2146 19966 2158 20018
rect 2210 19966 2222 20018
rect 5730 19966 5742 20018
rect 5794 19966 5806 20018
rect 19282 19966 19294 20018
rect 19346 19966 19358 20018
rect 25330 19966 25342 20018
rect 25394 19966 25406 20018
rect 1822 19954 1874 19966
rect 18958 19954 19010 19966
rect 40462 19954 40514 19966
rect 76526 20018 76578 20030
rect 76526 19954 76578 19966
rect 76974 20018 77026 20030
rect 76974 19954 77026 19966
rect 81006 20018 81058 20030
rect 81006 19954 81058 19966
rect 81678 20018 81730 20030
rect 81678 19954 81730 19966
rect 83022 20018 83074 20030
rect 83022 19954 83074 19966
rect 85486 20018 85538 20030
rect 85486 19954 85538 19966
rect 6078 19906 6130 19918
rect 6078 19842 6130 19854
rect 7310 19906 7362 19918
rect 7310 19842 7362 19854
rect 18510 19906 18562 19918
rect 18510 19842 18562 19854
rect 73054 19906 73106 19918
rect 73054 19842 73106 19854
rect 76414 19906 76466 19918
rect 76414 19842 76466 19854
rect 77422 19906 77474 19918
rect 77422 19842 77474 19854
rect 80446 19906 80498 19918
rect 80446 19842 80498 19854
rect 81118 19906 81170 19918
rect 81118 19842 81170 19854
rect 84702 19906 84754 19918
rect 84702 19842 84754 19854
rect 85262 19906 85314 19918
rect 85262 19842 85314 19854
rect 74510 19794 74562 19806
rect 74510 19730 74562 19742
rect 78094 19794 78146 19806
rect 78094 19730 78146 19742
rect 1344 19626 98560 19660
rect 1344 19574 4396 19626
rect 4448 19574 4520 19626
rect 4572 19574 4644 19626
rect 4696 19574 4768 19626
rect 4820 19574 13396 19626
rect 13448 19574 13520 19626
rect 13572 19574 13644 19626
rect 13696 19574 13768 19626
rect 13820 19574 22396 19626
rect 22448 19574 22520 19626
rect 22572 19574 22644 19626
rect 22696 19574 22768 19626
rect 22820 19574 31396 19626
rect 31448 19574 31520 19626
rect 31572 19574 31644 19626
rect 31696 19574 31768 19626
rect 31820 19574 40396 19626
rect 40448 19574 40520 19626
rect 40572 19574 40644 19626
rect 40696 19574 40768 19626
rect 40820 19574 49396 19626
rect 49448 19574 49520 19626
rect 49572 19574 49644 19626
rect 49696 19574 49768 19626
rect 49820 19574 58396 19626
rect 58448 19574 58520 19626
rect 58572 19574 58644 19626
rect 58696 19574 58768 19626
rect 58820 19574 67396 19626
rect 67448 19574 67520 19626
rect 67572 19574 67644 19626
rect 67696 19574 67768 19626
rect 67820 19574 76396 19626
rect 76448 19574 76520 19626
rect 76572 19574 76644 19626
rect 76696 19574 76768 19626
rect 76820 19574 85396 19626
rect 85448 19574 85520 19626
rect 85572 19574 85644 19626
rect 85696 19574 85768 19626
rect 85820 19574 94396 19626
rect 94448 19574 94520 19626
rect 94572 19574 94644 19626
rect 94696 19574 94768 19626
rect 94820 19574 98560 19626
rect 1344 19540 98560 19574
rect 74398 19458 74450 19470
rect 74398 19394 74450 19406
rect 79774 19458 79826 19470
rect 79774 19394 79826 19406
rect 89070 19458 89122 19470
rect 89070 19394 89122 19406
rect 3166 19346 3218 19358
rect 3166 19282 3218 19294
rect 6078 19346 6130 19358
rect 6078 19282 6130 19294
rect 6526 19346 6578 19358
rect 6526 19282 6578 19294
rect 74734 19346 74786 19358
rect 74734 19282 74786 19294
rect 75630 19346 75682 19358
rect 75630 19282 75682 19294
rect 1710 19234 1762 19246
rect 44270 19234 44322 19246
rect 40002 19182 40014 19234
rect 40066 19182 40078 19234
rect 1710 19170 1762 19182
rect 44270 19170 44322 19182
rect 70926 19234 70978 19246
rect 76078 19234 76130 19246
rect 80110 19234 80162 19246
rect 85598 19234 85650 19246
rect 71362 19182 71374 19234
rect 71426 19182 71438 19234
rect 76626 19182 76638 19234
rect 76690 19182 76702 19234
rect 80546 19182 80558 19234
rect 80610 19182 80622 19234
rect 86034 19182 86046 19234
rect 86098 19182 86110 19234
rect 96898 19182 96910 19234
rect 96962 19182 96974 19234
rect 70926 19170 70978 19182
rect 76078 19170 76130 19182
rect 80110 19170 80162 19182
rect 85598 19170 85650 19182
rect 2382 19122 2434 19134
rect 2382 19058 2434 19070
rect 2718 19122 2770 19134
rect 96686 19122 96738 19134
rect 42018 19070 42030 19122
rect 42082 19070 42094 19122
rect 98018 19070 98030 19122
rect 98082 19070 98094 19122
rect 2718 19058 2770 19070
rect 96686 19058 96738 19070
rect 2046 19010 2098 19022
rect 83582 19010 83634 19022
rect 73826 18958 73838 19010
rect 73890 18958 73902 19010
rect 79202 18958 79214 19010
rect 79266 18958 79278 19010
rect 82786 18958 82798 19010
rect 82850 18958 82862 19010
rect 2046 18946 2098 18958
rect 83582 18946 83634 18958
rect 85150 19010 85202 19022
rect 88274 18958 88286 19010
rect 88338 18958 88350 19010
rect 85150 18946 85202 18958
rect 1344 18842 98560 18876
rect 1344 18790 8896 18842
rect 8948 18790 9020 18842
rect 9072 18790 9144 18842
rect 9196 18790 9268 18842
rect 9320 18790 17896 18842
rect 17948 18790 18020 18842
rect 18072 18790 18144 18842
rect 18196 18790 18268 18842
rect 18320 18790 26896 18842
rect 26948 18790 27020 18842
rect 27072 18790 27144 18842
rect 27196 18790 27268 18842
rect 27320 18790 35896 18842
rect 35948 18790 36020 18842
rect 36072 18790 36144 18842
rect 36196 18790 36268 18842
rect 36320 18790 44896 18842
rect 44948 18790 45020 18842
rect 45072 18790 45144 18842
rect 45196 18790 45268 18842
rect 45320 18790 53896 18842
rect 53948 18790 54020 18842
rect 54072 18790 54144 18842
rect 54196 18790 54268 18842
rect 54320 18790 62896 18842
rect 62948 18790 63020 18842
rect 63072 18790 63144 18842
rect 63196 18790 63268 18842
rect 63320 18790 71896 18842
rect 71948 18790 72020 18842
rect 72072 18790 72144 18842
rect 72196 18790 72268 18842
rect 72320 18790 80896 18842
rect 80948 18790 81020 18842
rect 81072 18790 81144 18842
rect 81196 18790 81268 18842
rect 81320 18790 89896 18842
rect 89948 18790 90020 18842
rect 90072 18790 90144 18842
rect 90196 18790 90268 18842
rect 90320 18790 98560 18842
rect 1344 18756 98560 18790
rect 79662 18674 79714 18686
rect 79662 18610 79714 18622
rect 75182 18562 75234 18574
rect 75182 18498 75234 18510
rect 75518 18562 75570 18574
rect 75518 18498 75570 18510
rect 80222 18562 80274 18574
rect 80222 18498 80274 18510
rect 80558 18562 80610 18574
rect 80558 18498 80610 18510
rect 89966 18562 90018 18574
rect 89966 18498 90018 18510
rect 90302 18562 90354 18574
rect 90302 18498 90354 18510
rect 2158 18450 2210 18462
rect 2158 18386 2210 18398
rect 1344 18058 98560 18092
rect 1344 18006 4396 18058
rect 4448 18006 4520 18058
rect 4572 18006 4644 18058
rect 4696 18006 4768 18058
rect 4820 18006 13396 18058
rect 13448 18006 13520 18058
rect 13572 18006 13644 18058
rect 13696 18006 13768 18058
rect 13820 18006 22396 18058
rect 22448 18006 22520 18058
rect 22572 18006 22644 18058
rect 22696 18006 22768 18058
rect 22820 18006 31396 18058
rect 31448 18006 31520 18058
rect 31572 18006 31644 18058
rect 31696 18006 31768 18058
rect 31820 18006 40396 18058
rect 40448 18006 40520 18058
rect 40572 18006 40644 18058
rect 40696 18006 40768 18058
rect 40820 18006 49396 18058
rect 49448 18006 49520 18058
rect 49572 18006 49644 18058
rect 49696 18006 49768 18058
rect 49820 18006 58396 18058
rect 58448 18006 58520 18058
rect 58572 18006 58644 18058
rect 58696 18006 58768 18058
rect 58820 18006 67396 18058
rect 67448 18006 67520 18058
rect 67572 18006 67644 18058
rect 67696 18006 67768 18058
rect 67820 18006 76396 18058
rect 76448 18006 76520 18058
rect 76572 18006 76644 18058
rect 76696 18006 76768 18058
rect 76820 18006 85396 18058
rect 85448 18006 85520 18058
rect 85572 18006 85644 18058
rect 85696 18006 85768 18058
rect 85820 18006 94396 18058
rect 94448 18006 94520 18058
rect 94572 18006 94644 18058
rect 94696 18006 94768 18058
rect 94820 18006 98560 18058
rect 1344 17972 98560 18006
rect 85710 17666 85762 17678
rect 96898 17614 96910 17666
rect 96962 17614 96974 17666
rect 85710 17602 85762 17614
rect 1710 17554 1762 17566
rect 1710 17490 1762 17502
rect 2046 17554 2098 17566
rect 2046 17490 2098 17502
rect 2494 17554 2546 17566
rect 98018 17502 98030 17554
rect 98082 17502 98094 17554
rect 2494 17490 2546 17502
rect 86046 17442 86098 17454
rect 86046 17378 86098 17390
rect 96686 17442 96738 17454
rect 96686 17378 96738 17390
rect 1344 17274 98560 17308
rect 1344 17222 8896 17274
rect 8948 17222 9020 17274
rect 9072 17222 9144 17274
rect 9196 17222 9268 17274
rect 9320 17222 17896 17274
rect 17948 17222 18020 17274
rect 18072 17222 18144 17274
rect 18196 17222 18268 17274
rect 18320 17222 26896 17274
rect 26948 17222 27020 17274
rect 27072 17222 27144 17274
rect 27196 17222 27268 17274
rect 27320 17222 35896 17274
rect 35948 17222 36020 17274
rect 36072 17222 36144 17274
rect 36196 17222 36268 17274
rect 36320 17222 44896 17274
rect 44948 17222 45020 17274
rect 45072 17222 45144 17274
rect 45196 17222 45268 17274
rect 45320 17222 53896 17274
rect 53948 17222 54020 17274
rect 54072 17222 54144 17274
rect 54196 17222 54268 17274
rect 54320 17222 62896 17274
rect 62948 17222 63020 17274
rect 63072 17222 63144 17274
rect 63196 17222 63268 17274
rect 63320 17222 71896 17274
rect 71948 17222 72020 17274
rect 72072 17222 72144 17274
rect 72196 17222 72268 17274
rect 72320 17222 80896 17274
rect 80948 17222 81020 17274
rect 81072 17222 81144 17274
rect 81196 17222 81268 17274
rect 81320 17222 89896 17274
rect 89948 17222 90020 17274
rect 90072 17222 90144 17274
rect 90196 17222 90268 17274
rect 90320 17222 98560 17274
rect 1344 17188 98560 17222
rect 2046 17106 2098 17118
rect 2046 17042 2098 17054
rect 1710 16882 1762 16894
rect 1710 16818 1762 16830
rect 2494 16882 2546 16894
rect 2494 16818 2546 16830
rect 1344 16490 98560 16524
rect 1344 16438 4396 16490
rect 4448 16438 4520 16490
rect 4572 16438 4644 16490
rect 4696 16438 4768 16490
rect 4820 16438 13396 16490
rect 13448 16438 13520 16490
rect 13572 16438 13644 16490
rect 13696 16438 13768 16490
rect 13820 16438 22396 16490
rect 22448 16438 22520 16490
rect 22572 16438 22644 16490
rect 22696 16438 22768 16490
rect 22820 16438 31396 16490
rect 31448 16438 31520 16490
rect 31572 16438 31644 16490
rect 31696 16438 31768 16490
rect 31820 16438 40396 16490
rect 40448 16438 40520 16490
rect 40572 16438 40644 16490
rect 40696 16438 40768 16490
rect 40820 16438 49396 16490
rect 49448 16438 49520 16490
rect 49572 16438 49644 16490
rect 49696 16438 49768 16490
rect 49820 16438 58396 16490
rect 58448 16438 58520 16490
rect 58572 16438 58644 16490
rect 58696 16438 58768 16490
rect 58820 16438 67396 16490
rect 67448 16438 67520 16490
rect 67572 16438 67644 16490
rect 67696 16438 67768 16490
rect 67820 16438 76396 16490
rect 76448 16438 76520 16490
rect 76572 16438 76644 16490
rect 76696 16438 76768 16490
rect 76820 16438 85396 16490
rect 85448 16438 85520 16490
rect 85572 16438 85644 16490
rect 85696 16438 85768 16490
rect 85820 16438 94396 16490
rect 94448 16438 94520 16490
rect 94572 16438 94644 16490
rect 94696 16438 94768 16490
rect 94820 16438 98560 16490
rect 1344 16404 98560 16438
rect 96686 16098 96738 16110
rect 96898 16046 96910 16098
rect 96962 16046 96974 16098
rect 96686 16034 96738 16046
rect 98018 15934 98030 15986
rect 98082 15934 98094 15986
rect 1344 15706 98560 15740
rect 1344 15654 8896 15706
rect 8948 15654 9020 15706
rect 9072 15654 9144 15706
rect 9196 15654 9268 15706
rect 9320 15654 17896 15706
rect 17948 15654 18020 15706
rect 18072 15654 18144 15706
rect 18196 15654 18268 15706
rect 18320 15654 26896 15706
rect 26948 15654 27020 15706
rect 27072 15654 27144 15706
rect 27196 15654 27268 15706
rect 27320 15654 35896 15706
rect 35948 15654 36020 15706
rect 36072 15654 36144 15706
rect 36196 15654 36268 15706
rect 36320 15654 44896 15706
rect 44948 15654 45020 15706
rect 45072 15654 45144 15706
rect 45196 15654 45268 15706
rect 45320 15654 53896 15706
rect 53948 15654 54020 15706
rect 54072 15654 54144 15706
rect 54196 15654 54268 15706
rect 54320 15654 62896 15706
rect 62948 15654 63020 15706
rect 63072 15654 63144 15706
rect 63196 15654 63268 15706
rect 63320 15654 71896 15706
rect 71948 15654 72020 15706
rect 72072 15654 72144 15706
rect 72196 15654 72268 15706
rect 72320 15654 80896 15706
rect 80948 15654 81020 15706
rect 81072 15654 81144 15706
rect 81196 15654 81268 15706
rect 81320 15654 89896 15706
rect 89948 15654 90020 15706
rect 90072 15654 90144 15706
rect 90196 15654 90268 15706
rect 90320 15654 98560 15706
rect 1344 15620 98560 15654
rect 42242 15374 42254 15426
rect 42306 15374 42318 15426
rect 44594 15374 44606 15426
rect 44658 15374 44670 15426
rect 41682 15262 41694 15314
rect 41746 15262 41758 15314
rect 43026 15262 43038 15314
rect 43090 15262 43102 15314
rect 44818 15262 44830 15314
rect 44882 15262 44894 15314
rect 41134 15202 41186 15214
rect 41134 15138 41186 15150
rect 43934 15202 43986 15214
rect 43934 15138 43986 15150
rect 79662 15202 79714 15214
rect 79662 15138 79714 15150
rect 80334 15202 80386 15214
rect 80334 15138 80386 15150
rect 82798 15202 82850 15214
rect 82798 15138 82850 15150
rect 1344 14922 98560 14956
rect 1344 14870 4396 14922
rect 4448 14870 4520 14922
rect 4572 14870 4644 14922
rect 4696 14870 4768 14922
rect 4820 14870 13396 14922
rect 13448 14870 13520 14922
rect 13572 14870 13644 14922
rect 13696 14870 13768 14922
rect 13820 14870 22396 14922
rect 22448 14870 22520 14922
rect 22572 14870 22644 14922
rect 22696 14870 22768 14922
rect 22820 14870 31396 14922
rect 31448 14870 31520 14922
rect 31572 14870 31644 14922
rect 31696 14870 31768 14922
rect 31820 14870 40396 14922
rect 40448 14870 40520 14922
rect 40572 14870 40644 14922
rect 40696 14870 40768 14922
rect 40820 14870 49396 14922
rect 49448 14870 49520 14922
rect 49572 14870 49644 14922
rect 49696 14870 49768 14922
rect 49820 14870 58396 14922
rect 58448 14870 58520 14922
rect 58572 14870 58644 14922
rect 58696 14870 58768 14922
rect 58820 14870 67396 14922
rect 67448 14870 67520 14922
rect 67572 14870 67644 14922
rect 67696 14870 67768 14922
rect 67820 14870 76396 14922
rect 76448 14870 76520 14922
rect 76572 14870 76644 14922
rect 76696 14870 76768 14922
rect 76820 14870 85396 14922
rect 85448 14870 85520 14922
rect 85572 14870 85644 14922
rect 85696 14870 85768 14922
rect 85820 14870 94396 14922
rect 94448 14870 94520 14922
rect 94572 14870 94644 14922
rect 94696 14870 94768 14922
rect 94820 14870 98560 14922
rect 1344 14836 98560 14870
rect 46622 14642 46674 14654
rect 46622 14578 46674 14590
rect 44942 14530 44994 14542
rect 82798 14530 82850 14542
rect 21410 14478 21422 14530
rect 21474 14478 21486 14530
rect 45378 14478 45390 14530
rect 45442 14478 45454 14530
rect 46722 14478 46734 14530
rect 46786 14478 46798 14530
rect 47058 14478 47070 14530
rect 47122 14478 47134 14530
rect 70018 14478 70030 14530
rect 70082 14478 70094 14530
rect 71698 14478 71710 14530
rect 71762 14478 71774 14530
rect 74162 14478 74174 14530
rect 74226 14478 74238 14530
rect 78418 14478 78430 14530
rect 78482 14478 78494 14530
rect 80546 14478 80558 14530
rect 80610 14478 80622 14530
rect 81890 14478 81902 14530
rect 81954 14478 81966 14530
rect 96898 14478 96910 14530
rect 96962 14478 96974 14530
rect 44942 14466 44994 14478
rect 82798 14466 82850 14478
rect 83134 14418 83186 14430
rect 70578 14366 70590 14418
rect 70642 14366 70654 14418
rect 74162 14366 74174 14418
rect 74226 14366 74238 14418
rect 78306 14366 78318 14418
rect 78370 14366 78382 14418
rect 81666 14366 81678 14418
rect 81730 14366 81742 14418
rect 98018 14366 98030 14418
rect 98082 14366 98094 14418
rect 83134 14354 83186 14366
rect 20750 14306 20802 14318
rect 44270 14306 44322 14318
rect 74622 14306 74674 14318
rect 27682 14254 27694 14306
rect 27746 14254 27758 14306
rect 73938 14254 73950 14306
rect 74002 14254 74014 14306
rect 20750 14242 20802 14254
rect 44270 14242 44322 14254
rect 74622 14242 74674 14254
rect 75070 14306 75122 14318
rect 82226 14254 82238 14306
rect 82290 14254 82302 14306
rect 75070 14242 75122 14254
rect 1344 14138 98560 14172
rect 1344 14086 8896 14138
rect 8948 14086 9020 14138
rect 9072 14086 9144 14138
rect 9196 14086 9268 14138
rect 9320 14086 17896 14138
rect 17948 14086 18020 14138
rect 18072 14086 18144 14138
rect 18196 14086 18268 14138
rect 18320 14086 26896 14138
rect 26948 14086 27020 14138
rect 27072 14086 27144 14138
rect 27196 14086 27268 14138
rect 27320 14086 35896 14138
rect 35948 14086 36020 14138
rect 36072 14086 36144 14138
rect 36196 14086 36268 14138
rect 36320 14086 44896 14138
rect 44948 14086 45020 14138
rect 45072 14086 45144 14138
rect 45196 14086 45268 14138
rect 45320 14086 53896 14138
rect 53948 14086 54020 14138
rect 54072 14086 54144 14138
rect 54196 14086 54268 14138
rect 54320 14086 62896 14138
rect 62948 14086 63020 14138
rect 63072 14086 63144 14138
rect 63196 14086 63268 14138
rect 63320 14086 71896 14138
rect 71948 14086 72020 14138
rect 72072 14086 72144 14138
rect 72196 14086 72268 14138
rect 72320 14086 80896 14138
rect 80948 14086 81020 14138
rect 81072 14086 81144 14138
rect 81196 14086 81268 14138
rect 81320 14086 89896 14138
rect 89948 14086 90020 14138
rect 90072 14086 90144 14138
rect 90196 14086 90268 14138
rect 90320 14086 98560 14138
rect 1344 14052 98560 14086
rect 2046 13970 2098 13982
rect 2046 13906 2098 13918
rect 55582 13970 55634 13982
rect 55582 13906 55634 13918
rect 55134 13858 55186 13870
rect 72270 13858 72322 13870
rect 59042 13806 59054 13858
rect 59106 13806 59118 13858
rect 61842 13806 61854 13858
rect 61906 13806 61918 13858
rect 55134 13794 55186 13806
rect 72270 13794 72322 13806
rect 72606 13858 72658 13870
rect 80210 13806 80222 13858
rect 80274 13806 80286 13858
rect 72606 13794 72658 13806
rect 1710 13746 1762 13758
rect 74062 13746 74114 13758
rect 82798 13746 82850 13758
rect 34850 13694 34862 13746
rect 34914 13694 34926 13746
rect 43138 13694 43150 13746
rect 43202 13694 43214 13746
rect 51650 13694 51662 13746
rect 51714 13694 51726 13746
rect 52098 13694 52110 13746
rect 52162 13694 52174 13746
rect 52994 13694 53006 13746
rect 53058 13694 53070 13746
rect 53442 13694 53454 13746
rect 53506 13694 53518 13746
rect 54562 13694 54574 13746
rect 54626 13694 54638 13746
rect 58818 13694 58830 13746
rect 58882 13694 58894 13746
rect 60498 13694 60510 13746
rect 60562 13694 60574 13746
rect 61954 13694 61966 13746
rect 62018 13694 62030 13746
rect 75506 13694 75518 13746
rect 75570 13694 75582 13746
rect 76962 13694 76974 13746
rect 77026 13694 77038 13746
rect 77298 13694 77310 13746
rect 77362 13694 77374 13746
rect 77970 13694 77982 13746
rect 78034 13694 78046 13746
rect 80098 13694 80110 13746
rect 80162 13694 80174 13746
rect 81778 13694 81790 13746
rect 81842 13694 81854 13746
rect 83570 13694 83582 13746
rect 83634 13694 83646 13746
rect 1710 13682 1762 13694
rect 74062 13682 74114 13694
rect 82798 13682 82850 13694
rect 2494 13634 2546 13646
rect 51214 13634 51266 13646
rect 37202 13582 37214 13634
rect 37266 13582 37278 13634
rect 44258 13582 44270 13634
rect 44322 13582 44334 13634
rect 2494 13570 2546 13582
rect 51214 13570 51266 13582
rect 52334 13634 52386 13646
rect 52334 13570 52386 13582
rect 61070 13634 61122 13646
rect 79326 13634 79378 13646
rect 75394 13582 75406 13634
rect 75458 13582 75470 13634
rect 78866 13582 78878 13634
rect 78930 13582 78942 13634
rect 61070 13570 61122 13582
rect 79326 13570 79378 13582
rect 82686 13634 82738 13646
rect 82686 13570 82738 13582
rect 1344 13354 98560 13388
rect 1344 13302 4396 13354
rect 4448 13302 4520 13354
rect 4572 13302 4644 13354
rect 4696 13302 4768 13354
rect 4820 13302 13396 13354
rect 13448 13302 13520 13354
rect 13572 13302 13644 13354
rect 13696 13302 13768 13354
rect 13820 13302 22396 13354
rect 22448 13302 22520 13354
rect 22572 13302 22644 13354
rect 22696 13302 22768 13354
rect 22820 13302 31396 13354
rect 31448 13302 31520 13354
rect 31572 13302 31644 13354
rect 31696 13302 31768 13354
rect 31820 13302 40396 13354
rect 40448 13302 40520 13354
rect 40572 13302 40644 13354
rect 40696 13302 40768 13354
rect 40820 13302 49396 13354
rect 49448 13302 49520 13354
rect 49572 13302 49644 13354
rect 49696 13302 49768 13354
rect 49820 13302 58396 13354
rect 58448 13302 58520 13354
rect 58572 13302 58644 13354
rect 58696 13302 58768 13354
rect 58820 13302 67396 13354
rect 67448 13302 67520 13354
rect 67572 13302 67644 13354
rect 67696 13302 67768 13354
rect 67820 13302 76396 13354
rect 76448 13302 76520 13354
rect 76572 13302 76644 13354
rect 76696 13302 76768 13354
rect 76820 13302 85396 13354
rect 85448 13302 85520 13354
rect 85572 13302 85644 13354
rect 85696 13302 85768 13354
rect 85820 13302 94396 13354
rect 94448 13302 94520 13354
rect 94572 13302 94644 13354
rect 94696 13302 94768 13354
rect 94820 13302 98560 13354
rect 1344 13268 98560 13302
rect 45390 13074 45442 13086
rect 80434 13022 80446 13074
rect 80498 13022 80510 13074
rect 45390 13010 45442 13022
rect 37202 12910 37214 12962
rect 37266 12910 37278 12962
rect 46946 12910 46958 12962
rect 47010 12910 47022 12962
rect 48066 12910 48078 12962
rect 48130 12910 48142 12962
rect 50082 12910 50094 12962
rect 50146 12910 50158 12962
rect 66098 12910 66110 12962
rect 66162 12910 66174 12962
rect 73826 12910 73838 12962
rect 73890 12910 73902 12962
rect 82226 12910 82238 12962
rect 82290 12910 82302 12962
rect 41458 12798 41470 12850
rect 41522 12798 41534 12850
rect 47170 12798 47182 12850
rect 47234 12798 47246 12850
rect 49522 12798 49534 12850
rect 49586 12798 49598 12850
rect 61058 12798 61070 12850
rect 61122 12798 61134 12850
rect 69682 12798 69694 12850
rect 69746 12798 69758 12850
rect 47854 12738 47906 12750
rect 47854 12674 47906 12686
rect 50878 12738 50930 12750
rect 50878 12674 50930 12686
rect 51326 12738 51378 12750
rect 51326 12674 51378 12686
rect 66558 12738 66610 12750
rect 66558 12674 66610 12686
rect 74286 12738 74338 12750
rect 74286 12674 74338 12686
rect 1344 12570 98560 12604
rect 1344 12518 8896 12570
rect 8948 12518 9020 12570
rect 9072 12518 9144 12570
rect 9196 12518 9268 12570
rect 9320 12518 17896 12570
rect 17948 12518 18020 12570
rect 18072 12518 18144 12570
rect 18196 12518 18268 12570
rect 18320 12518 26896 12570
rect 26948 12518 27020 12570
rect 27072 12518 27144 12570
rect 27196 12518 27268 12570
rect 27320 12518 35896 12570
rect 35948 12518 36020 12570
rect 36072 12518 36144 12570
rect 36196 12518 36268 12570
rect 36320 12518 44896 12570
rect 44948 12518 45020 12570
rect 45072 12518 45144 12570
rect 45196 12518 45268 12570
rect 45320 12518 53896 12570
rect 53948 12518 54020 12570
rect 54072 12518 54144 12570
rect 54196 12518 54268 12570
rect 54320 12518 62896 12570
rect 62948 12518 63020 12570
rect 63072 12518 63144 12570
rect 63196 12518 63268 12570
rect 63320 12518 71896 12570
rect 71948 12518 72020 12570
rect 72072 12518 72144 12570
rect 72196 12518 72268 12570
rect 72320 12518 80896 12570
rect 80948 12518 81020 12570
rect 81072 12518 81144 12570
rect 81196 12518 81268 12570
rect 81320 12518 89896 12570
rect 89948 12518 90020 12570
rect 90072 12518 90144 12570
rect 90196 12518 90268 12570
rect 90320 12518 98560 12570
rect 1344 12484 98560 12518
rect 96574 12290 96626 12302
rect 2034 12238 2046 12290
rect 2098 12238 2110 12290
rect 48850 12238 48862 12290
rect 48914 12238 48926 12290
rect 52770 12238 52782 12290
rect 52834 12238 52846 12290
rect 60386 12238 60398 12290
rect 60450 12238 60462 12290
rect 68450 12238 68462 12290
rect 68514 12238 68526 12290
rect 71698 12238 71710 12290
rect 71762 12238 71774 12290
rect 96574 12226 96626 12238
rect 1710 12178 1762 12190
rect 40002 12126 40014 12178
rect 40066 12126 40078 12178
rect 42690 12126 42702 12178
rect 42754 12126 42766 12178
rect 48738 12126 48750 12178
rect 48802 12126 48814 12178
rect 51090 12126 51102 12178
rect 51154 12126 51166 12178
rect 52434 12126 52446 12178
rect 52498 12126 52510 12178
rect 63746 12126 63758 12178
rect 63810 12126 63822 12178
rect 67890 12126 67902 12178
rect 67954 12126 67966 12178
rect 69682 12126 69694 12178
rect 69746 12126 69758 12178
rect 71474 12126 71486 12178
rect 71538 12126 71550 12178
rect 76066 12126 76078 12178
rect 76130 12126 76142 12178
rect 80098 12126 80110 12178
rect 80162 12126 80174 12178
rect 81330 12126 81342 12178
rect 81394 12126 81406 12178
rect 82562 12126 82574 12178
rect 82626 12126 82638 12178
rect 83458 12126 83470 12178
rect 83522 12126 83534 12178
rect 96898 12126 96910 12178
rect 96962 12126 96974 12178
rect 1710 12114 1762 12126
rect 2494 12066 2546 12078
rect 48190 12066 48242 12078
rect 36866 12014 36878 12066
rect 36930 12014 36942 12066
rect 44370 12014 44382 12066
rect 44434 12014 44446 12066
rect 2494 12002 2546 12014
rect 48190 12002 48242 12014
rect 51326 12066 51378 12078
rect 51326 12002 51378 12014
rect 70142 12066 70194 12078
rect 78878 12066 78930 12078
rect 72482 12014 72494 12066
rect 72546 12014 72558 12066
rect 70142 12002 70194 12014
rect 78878 12002 78930 12014
rect 79326 12066 79378 12078
rect 83794 12014 83806 12066
rect 83858 12014 83870 12066
rect 98018 12014 98030 12066
rect 98082 12014 98094 12066
rect 79326 12002 79378 12014
rect 83906 11902 83918 11954
rect 83970 11902 83982 11954
rect 1344 11786 98560 11820
rect 1344 11734 4396 11786
rect 4448 11734 4520 11786
rect 4572 11734 4644 11786
rect 4696 11734 4768 11786
rect 4820 11734 13396 11786
rect 13448 11734 13520 11786
rect 13572 11734 13644 11786
rect 13696 11734 13768 11786
rect 13820 11734 22396 11786
rect 22448 11734 22520 11786
rect 22572 11734 22644 11786
rect 22696 11734 22768 11786
rect 22820 11734 31396 11786
rect 31448 11734 31520 11786
rect 31572 11734 31644 11786
rect 31696 11734 31768 11786
rect 31820 11734 40396 11786
rect 40448 11734 40520 11786
rect 40572 11734 40644 11786
rect 40696 11734 40768 11786
rect 40820 11734 49396 11786
rect 49448 11734 49520 11786
rect 49572 11734 49644 11786
rect 49696 11734 49768 11786
rect 49820 11734 58396 11786
rect 58448 11734 58520 11786
rect 58572 11734 58644 11786
rect 58696 11734 58768 11786
rect 58820 11734 67396 11786
rect 67448 11734 67520 11786
rect 67572 11734 67644 11786
rect 67696 11734 67768 11786
rect 67820 11734 76396 11786
rect 76448 11734 76520 11786
rect 76572 11734 76644 11786
rect 76696 11734 76768 11786
rect 76820 11734 85396 11786
rect 85448 11734 85520 11786
rect 85572 11734 85644 11786
rect 85696 11734 85768 11786
rect 85820 11734 94396 11786
rect 94448 11734 94520 11786
rect 94572 11734 94644 11786
rect 94696 11734 94768 11786
rect 94820 11734 98560 11786
rect 1344 11700 98560 11734
rect 67566 11618 67618 11630
rect 67566 11554 67618 11566
rect 62190 11506 62242 11518
rect 71138 11454 71150 11506
rect 71202 11454 71214 11506
rect 62190 11442 62242 11454
rect 31154 11342 31166 11394
rect 31218 11342 31230 11394
rect 38994 11342 39006 11394
rect 39058 11342 39070 11394
rect 46386 11342 46398 11394
rect 46450 11342 46462 11394
rect 56130 11342 56142 11394
rect 56194 11342 56206 11394
rect 58146 11342 58158 11394
rect 58210 11342 58222 11394
rect 59378 11342 59390 11394
rect 59442 11342 59454 11394
rect 63634 11342 63646 11394
rect 63698 11342 63710 11394
rect 73602 11342 73614 11394
rect 73666 11342 73678 11394
rect 81890 11342 81902 11394
rect 81954 11342 81966 11394
rect 1710 11282 1762 11294
rect 33954 11230 33966 11282
rect 34018 11230 34030 11282
rect 41010 11230 41022 11282
rect 41074 11230 41086 11282
rect 47058 11230 47070 11282
rect 47122 11230 47134 11282
rect 56690 11230 56702 11282
rect 56754 11230 56766 11282
rect 58034 11230 58046 11282
rect 58098 11230 58110 11282
rect 59154 11230 59166 11282
rect 59218 11230 59230 11282
rect 1710 11218 1762 11230
rect 2046 11170 2098 11182
rect 2046 11106 2098 11118
rect 2494 11170 2546 11182
rect 2494 11106 2546 11118
rect 60622 11170 60674 11182
rect 60622 11106 60674 11118
rect 61070 11170 61122 11182
rect 78194 11118 78206 11170
rect 78258 11118 78270 11170
rect 61070 11106 61122 11118
rect 1344 11002 98560 11036
rect 1344 10950 8896 11002
rect 8948 10950 9020 11002
rect 9072 10950 9144 11002
rect 9196 10950 9268 11002
rect 9320 10950 17896 11002
rect 17948 10950 18020 11002
rect 18072 10950 18144 11002
rect 18196 10950 18268 11002
rect 18320 10950 26896 11002
rect 26948 10950 27020 11002
rect 27072 10950 27144 11002
rect 27196 10950 27268 11002
rect 27320 10950 35896 11002
rect 35948 10950 36020 11002
rect 36072 10950 36144 11002
rect 36196 10950 36268 11002
rect 36320 10950 44896 11002
rect 44948 10950 45020 11002
rect 45072 10950 45144 11002
rect 45196 10950 45268 11002
rect 45320 10950 53896 11002
rect 53948 10950 54020 11002
rect 54072 10950 54144 11002
rect 54196 10950 54268 11002
rect 54320 10950 62896 11002
rect 62948 10950 63020 11002
rect 63072 10950 63144 11002
rect 63196 10950 63268 11002
rect 63320 10950 71896 11002
rect 71948 10950 72020 11002
rect 72072 10950 72144 11002
rect 72196 10950 72268 11002
rect 72320 10950 80896 11002
rect 80948 10950 81020 11002
rect 81072 10950 81144 11002
rect 81196 10950 81268 11002
rect 81320 10950 89896 11002
rect 89948 10950 90020 11002
rect 90072 10950 90144 11002
rect 90196 10950 90268 11002
rect 90320 10950 98560 11002
rect 1344 10916 98560 10950
rect 65538 10782 65550 10834
rect 65602 10782 65614 10834
rect 77870 10722 77922 10734
rect 76066 10670 76078 10722
rect 76130 10670 76142 10722
rect 77870 10658 77922 10670
rect 78206 10722 78258 10734
rect 78206 10658 78258 10670
rect 96686 10722 96738 10734
rect 96686 10658 96738 10670
rect 35298 10558 35310 10610
rect 35362 10558 35374 10610
rect 47170 10558 47182 10610
rect 47234 10558 47246 10610
rect 53218 10558 53230 10610
rect 53282 10558 53294 10610
rect 59938 10558 59950 10610
rect 60002 10558 60014 10610
rect 69682 10558 69694 10610
rect 69746 10558 69758 10610
rect 72594 10558 72606 10610
rect 72658 10558 72670 10610
rect 81554 10558 81566 10610
rect 81618 10558 81630 10610
rect 96898 10558 96910 10610
rect 96962 10558 96974 10610
rect 38098 10446 38110 10498
rect 38162 10446 38174 10498
rect 43698 10446 43710 10498
rect 43762 10446 43774 10498
rect 50418 10446 50430 10498
rect 50482 10446 50494 10498
rect 63522 10446 63534 10498
rect 63586 10446 63598 10498
rect 85138 10446 85150 10498
rect 85202 10446 85214 10498
rect 98018 10446 98030 10498
rect 98082 10446 98094 10498
rect 1344 10218 98560 10252
rect 1344 10166 4396 10218
rect 4448 10166 4520 10218
rect 4572 10166 4644 10218
rect 4696 10166 4768 10218
rect 4820 10166 13396 10218
rect 13448 10166 13520 10218
rect 13572 10166 13644 10218
rect 13696 10166 13768 10218
rect 13820 10166 22396 10218
rect 22448 10166 22520 10218
rect 22572 10166 22644 10218
rect 22696 10166 22768 10218
rect 22820 10166 31396 10218
rect 31448 10166 31520 10218
rect 31572 10166 31644 10218
rect 31696 10166 31768 10218
rect 31820 10166 40396 10218
rect 40448 10166 40520 10218
rect 40572 10166 40644 10218
rect 40696 10166 40768 10218
rect 40820 10166 49396 10218
rect 49448 10166 49520 10218
rect 49572 10166 49644 10218
rect 49696 10166 49768 10218
rect 49820 10166 58396 10218
rect 58448 10166 58520 10218
rect 58572 10166 58644 10218
rect 58696 10166 58768 10218
rect 58820 10166 67396 10218
rect 67448 10166 67520 10218
rect 67572 10166 67644 10218
rect 67696 10166 67768 10218
rect 67820 10166 76396 10218
rect 76448 10166 76520 10218
rect 76572 10166 76644 10218
rect 76696 10166 76768 10218
rect 76820 10166 85396 10218
rect 85448 10166 85520 10218
rect 85572 10166 85644 10218
rect 85696 10166 85768 10218
rect 85820 10166 94396 10218
rect 94448 10166 94520 10218
rect 94572 10166 94644 10218
rect 94696 10166 94768 10218
rect 94820 10166 98560 10218
rect 1344 10132 98560 10166
rect 45054 9938 45106 9950
rect 45054 9874 45106 9886
rect 46062 9938 46114 9950
rect 54674 9886 54686 9938
rect 54738 9886 54750 9938
rect 46062 9874 46114 9886
rect 35410 9774 35422 9826
rect 35474 9774 35486 9826
rect 38994 9774 39006 9826
rect 39058 9774 39070 9826
rect 47058 9774 47070 9826
rect 47122 9774 47134 9826
rect 52770 9774 52782 9826
rect 52834 9774 52846 9826
rect 64306 9774 64318 9826
rect 64370 9774 64382 9826
rect 75058 9774 75070 9826
rect 75122 9774 75134 9826
rect 81442 9774 81454 9826
rect 81506 9774 81518 9826
rect 88946 9774 88958 9826
rect 89010 9774 89022 9826
rect 1710 9714 1762 9726
rect 1710 9650 1762 9662
rect 2494 9714 2546 9726
rect 31938 9662 31950 9714
rect 32002 9662 32014 9714
rect 41010 9662 41022 9714
rect 41074 9662 41086 9714
rect 48962 9662 48974 9714
rect 49026 9662 49038 9714
rect 62402 9662 62414 9714
rect 62466 9662 62478 9714
rect 70690 9662 70702 9714
rect 70754 9662 70766 9714
rect 77298 9662 77310 9714
rect 77362 9662 77374 9714
rect 84354 9662 84366 9714
rect 84418 9662 84430 9714
rect 2494 9650 2546 9662
rect 45166 9602 45218 9614
rect 2034 9550 2046 9602
rect 2098 9550 2110 9602
rect 45166 9538 45218 9550
rect 45950 9602 46002 9614
rect 45950 9538 46002 9550
rect 1344 9434 98560 9468
rect 1344 9382 8896 9434
rect 8948 9382 9020 9434
rect 9072 9382 9144 9434
rect 9196 9382 9268 9434
rect 9320 9382 17896 9434
rect 17948 9382 18020 9434
rect 18072 9382 18144 9434
rect 18196 9382 18268 9434
rect 18320 9382 26896 9434
rect 26948 9382 27020 9434
rect 27072 9382 27144 9434
rect 27196 9382 27268 9434
rect 27320 9382 35896 9434
rect 35948 9382 36020 9434
rect 36072 9382 36144 9434
rect 36196 9382 36268 9434
rect 36320 9382 44896 9434
rect 44948 9382 45020 9434
rect 45072 9382 45144 9434
rect 45196 9382 45268 9434
rect 45320 9382 53896 9434
rect 53948 9382 54020 9434
rect 54072 9382 54144 9434
rect 54196 9382 54268 9434
rect 54320 9382 62896 9434
rect 62948 9382 63020 9434
rect 63072 9382 63144 9434
rect 63196 9382 63268 9434
rect 63320 9382 71896 9434
rect 71948 9382 72020 9434
rect 72072 9382 72144 9434
rect 72196 9382 72268 9434
rect 72320 9382 80896 9434
rect 80948 9382 81020 9434
rect 81072 9382 81144 9434
rect 81196 9382 81268 9434
rect 81320 9382 89896 9434
rect 89948 9382 90020 9434
rect 90072 9382 90144 9434
rect 90196 9382 90268 9434
rect 90320 9382 98560 9434
rect 1344 9348 98560 9382
rect 96686 9266 96738 9278
rect 96686 9202 96738 9214
rect 96910 9266 96962 9278
rect 96910 9202 96962 9214
rect 48862 9154 48914 9166
rect 48862 9090 48914 9102
rect 49198 9154 49250 9166
rect 80658 9102 80670 9154
rect 80722 9102 80734 9154
rect 49198 9090 49250 9102
rect 50206 9042 50258 9054
rect 31826 8990 31838 9042
rect 31890 8990 31902 9042
rect 35522 8990 35534 9042
rect 35586 8990 35598 9042
rect 43138 8990 43150 9042
rect 43202 8990 43214 9042
rect 50530 8990 50542 9042
rect 50594 8990 50606 9042
rect 63074 8990 63086 9042
rect 63138 8990 63150 9042
rect 68898 8990 68910 9042
rect 68962 8990 68974 9042
rect 76066 8990 76078 9042
rect 76130 8990 76142 9042
rect 84018 8990 84030 9042
rect 84082 8990 84094 9042
rect 50206 8978 50258 8990
rect 34526 8930 34578 8942
rect 42702 8930 42754 8942
rect 49758 8930 49810 8942
rect 30146 8878 30158 8930
rect 30210 8878 30222 8930
rect 37202 8878 37214 8930
rect 37266 8878 37278 8930
rect 45938 8878 45950 8930
rect 46002 8878 46014 8930
rect 54562 8878 54574 8930
rect 54626 8878 54638 8930
rect 59826 8878 59838 8930
rect 59890 8878 59902 8930
rect 65538 8878 65550 8930
rect 65602 8878 65614 8930
rect 72482 8878 72494 8930
rect 72546 8878 72558 8930
rect 34526 8866 34578 8878
rect 42702 8866 42754 8878
rect 49758 8866 49810 8878
rect 48750 8818 48802 8830
rect 48750 8754 48802 8766
rect 50094 8818 50146 8830
rect 50094 8754 50146 8766
rect 97694 8818 97746 8830
rect 97694 8754 97746 8766
rect 1344 8650 98560 8684
rect 1344 8598 4396 8650
rect 4448 8598 4520 8650
rect 4572 8598 4644 8650
rect 4696 8598 4768 8650
rect 4820 8598 13396 8650
rect 13448 8598 13520 8650
rect 13572 8598 13644 8650
rect 13696 8598 13768 8650
rect 13820 8598 22396 8650
rect 22448 8598 22520 8650
rect 22572 8598 22644 8650
rect 22696 8598 22768 8650
rect 22820 8598 31396 8650
rect 31448 8598 31520 8650
rect 31572 8598 31644 8650
rect 31696 8598 31768 8650
rect 31820 8598 40396 8650
rect 40448 8598 40520 8650
rect 40572 8598 40644 8650
rect 40696 8598 40768 8650
rect 40820 8598 49396 8650
rect 49448 8598 49520 8650
rect 49572 8598 49644 8650
rect 49696 8598 49768 8650
rect 49820 8598 58396 8650
rect 58448 8598 58520 8650
rect 58572 8598 58644 8650
rect 58696 8598 58768 8650
rect 58820 8598 67396 8650
rect 67448 8598 67520 8650
rect 67572 8598 67644 8650
rect 67696 8598 67768 8650
rect 67820 8598 76396 8650
rect 76448 8598 76520 8650
rect 76572 8598 76644 8650
rect 76696 8598 76768 8650
rect 76820 8598 85396 8650
rect 85448 8598 85520 8650
rect 85572 8598 85644 8650
rect 85696 8598 85768 8650
rect 85820 8598 94396 8650
rect 94448 8598 94520 8650
rect 94572 8598 94644 8650
rect 94696 8598 94768 8650
rect 94820 8598 98560 8650
rect 1344 8564 98560 8598
rect 58830 8370 58882 8382
rect 45714 8318 45726 8370
rect 45778 8318 45790 8370
rect 81442 8318 81454 8370
rect 81506 8367 81518 8370
rect 81778 8367 81790 8370
rect 81506 8321 81790 8367
rect 81506 8318 81518 8321
rect 81778 8318 81790 8321
rect 81842 8318 81854 8370
rect 58830 8306 58882 8318
rect 45838 8258 45890 8270
rect 58942 8258 58994 8270
rect 36418 8206 36430 8258
rect 36482 8206 36494 8258
rect 40002 8206 40014 8258
rect 40066 8206 40078 8258
rect 45378 8206 45390 8258
rect 45442 8206 45454 8258
rect 46274 8206 46286 8258
rect 46338 8206 46350 8258
rect 51874 8206 51886 8258
rect 51938 8206 51950 8258
rect 52658 8206 52670 8258
rect 52722 8206 52734 8258
rect 45838 8194 45890 8206
rect 58942 8194 58994 8206
rect 59166 8258 59218 8270
rect 61954 8206 61966 8258
rect 62018 8206 62030 8258
rect 69010 8206 69022 8258
rect 69074 8206 69086 8258
rect 81442 8206 81454 8258
rect 81506 8206 81518 8258
rect 88050 8206 88062 8258
rect 88114 8206 88126 8258
rect 59166 8194 59218 8206
rect 44830 8146 44882 8158
rect 34290 8094 34302 8146
rect 34354 8094 34366 8146
rect 44034 8094 44046 8146
rect 44098 8094 44110 8146
rect 48626 8094 48638 8146
rect 48690 8094 48702 8146
rect 54674 8094 54686 8146
rect 54738 8094 54750 8146
rect 63858 8094 63870 8146
rect 63922 8094 63934 8146
rect 71362 8094 71374 8146
rect 71426 8094 71438 8146
rect 76402 8094 76414 8146
rect 76466 8094 76478 8146
rect 86146 8094 86158 8146
rect 86210 8094 86222 8146
rect 44830 8082 44882 8094
rect 58830 8034 58882 8046
rect 58830 7970 58882 7982
rect 66222 8034 66274 8046
rect 66222 7970 66274 7982
rect 81902 8034 81954 8046
rect 81902 7970 81954 7982
rect 1344 7866 98560 7900
rect 1344 7814 8896 7866
rect 8948 7814 9020 7866
rect 9072 7814 9144 7866
rect 9196 7814 9268 7866
rect 9320 7814 17896 7866
rect 17948 7814 18020 7866
rect 18072 7814 18144 7866
rect 18196 7814 18268 7866
rect 18320 7814 26896 7866
rect 26948 7814 27020 7866
rect 27072 7814 27144 7866
rect 27196 7814 27268 7866
rect 27320 7814 35896 7866
rect 35948 7814 36020 7866
rect 36072 7814 36144 7866
rect 36196 7814 36268 7866
rect 36320 7814 44896 7866
rect 44948 7814 45020 7866
rect 45072 7814 45144 7866
rect 45196 7814 45268 7866
rect 45320 7814 53896 7866
rect 53948 7814 54020 7866
rect 54072 7814 54144 7866
rect 54196 7814 54268 7866
rect 54320 7814 62896 7866
rect 62948 7814 63020 7866
rect 63072 7814 63144 7866
rect 63196 7814 63268 7866
rect 63320 7814 71896 7866
rect 71948 7814 72020 7866
rect 72072 7814 72144 7866
rect 72196 7814 72268 7866
rect 72320 7814 80896 7866
rect 80948 7814 81020 7866
rect 81072 7814 81144 7866
rect 81196 7814 81268 7866
rect 81320 7814 89896 7866
rect 89948 7814 90020 7866
rect 90072 7814 90144 7866
rect 90196 7814 90268 7866
rect 90320 7814 98560 7866
rect 1344 7780 98560 7814
rect 42478 7698 42530 7710
rect 42478 7634 42530 7646
rect 48974 7698 49026 7710
rect 48974 7634 49026 7646
rect 49870 7698 49922 7710
rect 49870 7634 49922 7646
rect 33518 7586 33570 7598
rect 30034 7534 30046 7586
rect 30098 7534 30110 7586
rect 33518 7522 33570 7534
rect 34302 7586 34354 7598
rect 34302 7522 34354 7534
rect 34638 7586 34690 7598
rect 34638 7522 34690 7534
rect 41246 7586 41298 7598
rect 62190 7586 62242 7598
rect 59266 7534 59278 7586
rect 59330 7534 59342 7586
rect 66434 7534 66446 7586
rect 66498 7534 66510 7586
rect 90850 7534 90862 7586
rect 90914 7534 90926 7586
rect 41246 7522 41298 7534
rect 62190 7522 62242 7534
rect 42142 7474 42194 7486
rect 32498 7422 32510 7474
rect 32562 7422 32574 7474
rect 40114 7422 40126 7474
rect 40178 7422 40190 7474
rect 42142 7410 42194 7422
rect 42478 7474 42530 7486
rect 71038 7474 71090 7486
rect 42914 7422 42926 7474
rect 42978 7422 42990 7474
rect 50306 7422 50318 7474
rect 50370 7422 50382 7474
rect 51986 7422 51998 7474
rect 52050 7422 52062 7474
rect 56578 7422 56590 7474
rect 56642 7422 56654 7474
rect 64642 7422 64654 7474
rect 64706 7422 64718 7474
rect 42478 7410 42530 7422
rect 71038 7410 71090 7422
rect 71374 7474 71426 7486
rect 77186 7422 77198 7474
rect 77250 7422 77262 7474
rect 78306 7422 78318 7474
rect 78370 7422 78382 7474
rect 84018 7422 84030 7474
rect 84082 7422 84094 7474
rect 87938 7422 87950 7474
rect 88002 7422 88014 7474
rect 71374 7410 71426 7422
rect 1822 7362 1874 7374
rect 70366 7362 70418 7374
rect 38322 7310 38334 7362
rect 38386 7310 38398 7362
rect 45378 7310 45390 7362
rect 45442 7310 45454 7362
rect 53778 7310 53790 7362
rect 53842 7310 53854 7362
rect 74050 7310 74062 7362
rect 74114 7310 74126 7362
rect 77970 7310 77982 7362
rect 78034 7310 78046 7362
rect 81554 7310 81566 7362
rect 81618 7310 81630 7362
rect 1822 7298 1874 7310
rect 70366 7298 70418 7310
rect 34190 7250 34242 7262
rect 34190 7186 34242 7198
rect 34750 7250 34802 7262
rect 34750 7186 34802 7198
rect 41694 7250 41746 7262
rect 41694 7186 41746 7198
rect 42366 7250 42418 7262
rect 42366 7186 42418 7198
rect 71150 7250 71202 7262
rect 71150 7186 71202 7198
rect 71486 7250 71538 7262
rect 71486 7186 71538 7198
rect 1344 7082 98560 7116
rect 1344 7030 4396 7082
rect 4448 7030 4520 7082
rect 4572 7030 4644 7082
rect 4696 7030 4768 7082
rect 4820 7030 13396 7082
rect 13448 7030 13520 7082
rect 13572 7030 13644 7082
rect 13696 7030 13768 7082
rect 13820 7030 22396 7082
rect 22448 7030 22520 7082
rect 22572 7030 22644 7082
rect 22696 7030 22768 7082
rect 22820 7030 31396 7082
rect 31448 7030 31520 7082
rect 31572 7030 31644 7082
rect 31696 7030 31768 7082
rect 31820 7030 40396 7082
rect 40448 7030 40520 7082
rect 40572 7030 40644 7082
rect 40696 7030 40768 7082
rect 40820 7030 49396 7082
rect 49448 7030 49520 7082
rect 49572 7030 49644 7082
rect 49696 7030 49768 7082
rect 49820 7030 58396 7082
rect 58448 7030 58520 7082
rect 58572 7030 58644 7082
rect 58696 7030 58768 7082
rect 58820 7030 67396 7082
rect 67448 7030 67520 7082
rect 67572 7030 67644 7082
rect 67696 7030 67768 7082
rect 67820 7030 76396 7082
rect 76448 7030 76520 7082
rect 76572 7030 76644 7082
rect 76696 7030 76768 7082
rect 76820 7030 85396 7082
rect 85448 7030 85520 7082
rect 85572 7030 85644 7082
rect 85696 7030 85768 7082
rect 85820 7030 94396 7082
rect 94448 7030 94520 7082
rect 94572 7030 94644 7082
rect 94696 7030 94768 7082
rect 94820 7030 98560 7082
rect 1344 6996 98560 7030
rect 37102 6914 37154 6926
rect 37102 6850 37154 6862
rect 37326 6914 37378 6926
rect 37326 6850 37378 6862
rect 37438 6914 37490 6926
rect 59726 6914 59778 6926
rect 59266 6862 59278 6914
rect 59330 6911 59342 6914
rect 59490 6911 59502 6914
rect 59330 6865 59502 6911
rect 59330 6862 59342 6865
rect 59490 6862 59502 6865
rect 59554 6862 59566 6914
rect 37438 6850 37490 6862
rect 59726 6850 59778 6862
rect 46274 6750 46286 6802
rect 46338 6750 46350 6802
rect 51874 6750 51886 6802
rect 51938 6750 51950 6802
rect 64306 6750 64318 6802
rect 64370 6750 64382 6802
rect 87938 6750 87950 6802
rect 88002 6750 88014 6802
rect 2270 6690 2322 6702
rect 25902 6690 25954 6702
rect 45614 6690 45666 6702
rect 59838 6690 59890 6702
rect 73950 6690 74002 6702
rect 25106 6638 25118 6690
rect 25170 6638 25182 6690
rect 26786 6638 26798 6690
rect 26850 6638 26862 6690
rect 28354 6638 28366 6690
rect 28418 6638 28430 6690
rect 35634 6638 35646 6690
rect 35698 6638 35710 6690
rect 44258 6638 44270 6690
rect 44322 6638 44334 6690
rect 46050 6638 46062 6690
rect 46114 6638 46126 6690
rect 47842 6638 47854 6690
rect 47906 6638 47918 6690
rect 54338 6638 54350 6690
rect 54402 6638 54414 6690
rect 60498 6638 60510 6690
rect 60562 6638 60574 6690
rect 72706 6638 72718 6690
rect 72770 6638 72782 6690
rect 2270 6626 2322 6638
rect 25902 6626 25954 6638
rect 45614 6626 45666 6638
rect 59838 6626 59890 6638
rect 73950 6626 74002 6638
rect 74062 6690 74114 6702
rect 96686 6690 96738 6702
rect 76178 6638 76190 6690
rect 76242 6638 76254 6690
rect 84018 6638 84030 6690
rect 84082 6638 84094 6690
rect 96898 6638 96910 6690
rect 96962 6638 96974 6690
rect 74062 6626 74114 6638
rect 96686 6626 96738 6638
rect 36990 6578 37042 6590
rect 81790 6578 81842 6590
rect 27906 6526 27918 6578
rect 27970 6526 27982 6578
rect 34402 6526 34414 6578
rect 34466 6526 34478 6578
rect 41906 6526 41918 6578
rect 41970 6526 41982 6578
rect 54898 6526 54910 6578
rect 54962 6526 54974 6578
rect 69010 6526 69022 6578
rect 69074 6526 69086 6578
rect 78194 6526 78206 6578
rect 78258 6526 78270 6578
rect 98018 6526 98030 6578
rect 98082 6526 98094 6578
rect 36990 6514 37042 6526
rect 81790 6514 81842 6526
rect 1710 6466 1762 6478
rect 29374 6466 29426 6478
rect 27570 6414 27582 6466
rect 27634 6414 27646 6466
rect 1710 6402 1762 6414
rect 29374 6402 29426 6414
rect 37998 6466 38050 6478
rect 37998 6402 38050 6414
rect 45390 6466 45442 6478
rect 45390 6402 45442 6414
rect 59390 6466 59442 6478
rect 59390 6402 59442 6414
rect 74510 6466 74562 6478
rect 74510 6402 74562 6414
rect 74846 6466 74898 6478
rect 74846 6402 74898 6414
rect 75406 6466 75458 6478
rect 75406 6402 75458 6414
rect 81902 6466 81954 6478
rect 81902 6402 81954 6414
rect 82350 6466 82402 6478
rect 82350 6402 82402 6414
rect 1344 6298 98560 6332
rect 1344 6246 8896 6298
rect 8948 6246 9020 6298
rect 9072 6246 9144 6298
rect 9196 6246 9268 6298
rect 9320 6246 17896 6298
rect 17948 6246 18020 6298
rect 18072 6246 18144 6298
rect 18196 6246 18268 6298
rect 18320 6246 26896 6298
rect 26948 6246 27020 6298
rect 27072 6246 27144 6298
rect 27196 6246 27268 6298
rect 27320 6246 35896 6298
rect 35948 6246 36020 6298
rect 36072 6246 36144 6298
rect 36196 6246 36268 6298
rect 36320 6246 44896 6298
rect 44948 6246 45020 6298
rect 45072 6246 45144 6298
rect 45196 6246 45268 6298
rect 45320 6246 53896 6298
rect 53948 6246 54020 6298
rect 54072 6246 54144 6298
rect 54196 6246 54268 6298
rect 54320 6246 62896 6298
rect 62948 6246 63020 6298
rect 63072 6246 63144 6298
rect 63196 6246 63268 6298
rect 63320 6246 71896 6298
rect 71948 6246 72020 6298
rect 72072 6246 72144 6298
rect 72196 6246 72268 6298
rect 72320 6246 80896 6298
rect 80948 6246 81020 6298
rect 81072 6246 81144 6298
rect 81196 6246 81268 6298
rect 81320 6246 89896 6298
rect 89948 6246 90020 6298
rect 90072 6246 90144 6298
rect 90196 6246 90268 6298
rect 90320 6246 98560 6298
rect 1344 6212 98560 6246
rect 34862 6130 34914 6142
rect 34862 6066 34914 6078
rect 41022 6130 41074 6142
rect 41022 6066 41074 6078
rect 41694 6130 41746 6142
rect 41694 6066 41746 6078
rect 42142 6130 42194 6142
rect 42142 6066 42194 6078
rect 42590 6130 42642 6142
rect 42590 6066 42642 6078
rect 71262 6130 71314 6142
rect 71262 6066 71314 6078
rect 78094 6130 78146 6142
rect 78094 6066 78146 6078
rect 78542 6130 78594 6142
rect 78542 6066 78594 6078
rect 78990 6130 79042 6142
rect 78990 6066 79042 6078
rect 33518 6018 33570 6030
rect 40910 6018 40962 6030
rect 31042 5966 31054 6018
rect 31106 5966 31118 6018
rect 35634 5966 35646 6018
rect 35698 5966 35710 6018
rect 33518 5954 33570 5966
rect 40910 5954 40962 5966
rect 49982 6018 50034 6030
rect 63758 6018 63810 6030
rect 55346 5966 55358 6018
rect 55410 5966 55422 6018
rect 58818 5966 58830 6018
rect 58882 5966 58894 6018
rect 49982 5954 50034 5966
rect 63758 5954 63810 5966
rect 63870 6018 63922 6030
rect 70254 6018 70306 6030
rect 68786 5966 68798 6018
rect 68850 5966 68862 6018
rect 63870 5954 63922 5966
rect 70254 5954 70306 5966
rect 70814 6018 70866 6030
rect 72482 5966 72494 6018
rect 72546 5966 72558 6018
rect 83906 5966 83918 6018
rect 83970 5966 83982 6018
rect 90738 5966 90750 6018
rect 90802 5966 90814 6018
rect 70814 5954 70866 5966
rect 34190 5906 34242 5918
rect 1810 5854 1822 5906
rect 1874 5854 1886 5906
rect 27570 5854 27582 5906
rect 27634 5854 27646 5906
rect 33842 5854 33854 5906
rect 33906 5854 33918 5906
rect 34190 5842 34242 5854
rect 34750 5906 34802 5918
rect 49086 5906 49138 5918
rect 40114 5854 40126 5906
rect 40178 5854 40190 5906
rect 48178 5854 48190 5906
rect 48242 5854 48254 5906
rect 34750 5842 34802 5854
rect 49086 5842 49138 5854
rect 49310 5906 49362 5918
rect 49310 5842 49362 5854
rect 49870 5906 49922 5918
rect 62078 5906 62130 5918
rect 71710 5906 71762 5918
rect 50754 5854 50766 5906
rect 50818 5854 50830 5906
rect 57138 5854 57150 5906
rect 57202 5854 57214 5906
rect 62514 5854 62526 5906
rect 62578 5854 62590 5906
rect 62850 5854 62862 5906
rect 62914 5854 62926 5906
rect 64418 5854 64430 5906
rect 64482 5854 64494 5906
rect 71026 5854 71038 5906
rect 71090 5854 71102 5906
rect 76066 5854 76078 5906
rect 76130 5854 76142 5906
rect 80098 5854 80110 5906
rect 80162 5854 80174 5906
rect 88162 5854 88174 5906
rect 88226 5854 88238 5906
rect 49870 5842 49922 5854
rect 62078 5842 62130 5854
rect 71710 5842 71762 5854
rect 2270 5794 2322 5806
rect 2270 5730 2322 5742
rect 34526 5794 34578 5806
rect 50430 5794 50482 5806
rect 79438 5794 79490 5806
rect 45266 5742 45278 5794
rect 45330 5742 45342 5794
rect 62402 5742 62414 5794
rect 62466 5742 62478 5794
rect 70802 5742 70814 5794
rect 70866 5742 70878 5794
rect 34526 5730 34578 5742
rect 50430 5730 50482 5742
rect 79438 5730 79490 5742
rect 34302 5682 34354 5694
rect 34302 5618 34354 5630
rect 48974 5682 49026 5694
rect 48974 5618 49026 5630
rect 49422 5682 49474 5694
rect 49422 5618 49474 5630
rect 70366 5682 70418 5694
rect 70366 5618 70418 5630
rect 71598 5682 71650 5694
rect 71598 5618 71650 5630
rect 1344 5514 98560 5548
rect 1344 5462 4396 5514
rect 4448 5462 4520 5514
rect 4572 5462 4644 5514
rect 4696 5462 4768 5514
rect 4820 5462 13396 5514
rect 13448 5462 13520 5514
rect 13572 5462 13644 5514
rect 13696 5462 13768 5514
rect 13820 5462 22396 5514
rect 22448 5462 22520 5514
rect 22572 5462 22644 5514
rect 22696 5462 22768 5514
rect 22820 5462 31396 5514
rect 31448 5462 31520 5514
rect 31572 5462 31644 5514
rect 31696 5462 31768 5514
rect 31820 5462 40396 5514
rect 40448 5462 40520 5514
rect 40572 5462 40644 5514
rect 40696 5462 40768 5514
rect 40820 5462 49396 5514
rect 49448 5462 49520 5514
rect 49572 5462 49644 5514
rect 49696 5462 49768 5514
rect 49820 5462 58396 5514
rect 58448 5462 58520 5514
rect 58572 5462 58644 5514
rect 58696 5462 58768 5514
rect 58820 5462 67396 5514
rect 67448 5462 67520 5514
rect 67572 5462 67644 5514
rect 67696 5462 67768 5514
rect 67820 5462 76396 5514
rect 76448 5462 76520 5514
rect 76572 5462 76644 5514
rect 76696 5462 76768 5514
rect 76820 5462 85396 5514
rect 85448 5462 85520 5514
rect 85572 5462 85644 5514
rect 85696 5462 85768 5514
rect 85820 5462 94396 5514
rect 94448 5462 94520 5514
rect 94572 5462 94644 5514
rect 94696 5462 94768 5514
rect 94820 5462 98560 5514
rect 1344 5428 98560 5462
rect 30718 5346 30770 5358
rect 30718 5282 30770 5294
rect 37214 5346 37266 5358
rect 37214 5282 37266 5294
rect 58270 5346 58322 5358
rect 58270 5282 58322 5294
rect 59950 5346 60002 5358
rect 59950 5282 60002 5294
rect 67790 5346 67842 5358
rect 67790 5282 67842 5294
rect 74846 5346 74898 5358
rect 74846 5282 74898 5294
rect 1822 5234 1874 5246
rect 44942 5234 44994 5246
rect 73950 5234 74002 5246
rect 96574 5234 96626 5246
rect 26562 5182 26574 5234
rect 26626 5182 26638 5234
rect 34402 5182 34414 5234
rect 34466 5182 34478 5234
rect 42242 5182 42254 5234
rect 42306 5182 42318 5234
rect 46274 5182 46286 5234
rect 46338 5182 46350 5234
rect 51762 5182 51774 5234
rect 51826 5182 51838 5234
rect 54674 5182 54686 5234
rect 54738 5182 54750 5234
rect 60722 5182 60734 5234
rect 60786 5182 60798 5234
rect 70690 5182 70702 5234
rect 70754 5182 70766 5234
rect 79090 5182 79102 5234
rect 79154 5182 79166 5234
rect 87490 5182 87502 5234
rect 87554 5182 87566 5234
rect 1822 5170 1874 5182
rect 44942 5170 44994 5182
rect 73950 5170 74002 5182
rect 96574 5170 96626 5182
rect 37438 5122 37490 5134
rect 28466 5070 28478 5122
rect 28530 5070 28542 5122
rect 36418 5070 36430 5122
rect 36482 5070 36494 5122
rect 36978 5070 36990 5122
rect 37042 5070 37054 5122
rect 37438 5058 37490 5070
rect 37886 5122 37938 5134
rect 37886 5058 37938 5070
rect 37998 5122 38050 5134
rect 59166 5122 59218 5134
rect 42802 5070 42814 5122
rect 42866 5070 42878 5122
rect 45826 5070 45838 5122
rect 45890 5070 45902 5122
rect 46162 5070 46174 5122
rect 46226 5070 46238 5122
rect 48290 5070 48302 5122
rect 48354 5070 48366 5122
rect 57922 5070 57934 5122
rect 57986 5070 57998 5122
rect 37998 5058 38050 5070
rect 59166 5058 59218 5070
rect 59838 5122 59890 5134
rect 67342 5122 67394 5134
rect 96910 5122 96962 5134
rect 65426 5070 65438 5122
rect 65490 5070 65502 5122
rect 68338 5070 68350 5122
rect 68402 5070 68414 5122
rect 74386 5070 74398 5122
rect 74450 5070 74462 5122
rect 77074 5070 77086 5122
rect 77138 5070 77150 5122
rect 83234 5070 83246 5122
rect 83298 5070 83310 5122
rect 84242 5070 84254 5122
rect 84306 5070 84318 5122
rect 59838 5058 59890 5070
rect 67342 5058 67394 5070
rect 96910 5058 96962 5070
rect 97694 5122 97746 5134
rect 97694 5058 97746 5070
rect 59054 5010 59106 5022
rect 59614 5010 59666 5022
rect 59266 4958 59278 5010
rect 59330 4958 59342 5010
rect 82114 4958 82126 5010
rect 82178 4958 82190 5010
rect 59054 4946 59106 4958
rect 59614 4946 59666 4958
rect 37102 4898 37154 4910
rect 37102 4834 37154 4846
rect 38670 4898 38722 4910
rect 38670 4834 38722 4846
rect 46622 4898 46674 4910
rect 46622 4834 46674 4846
rect 75294 4898 75346 4910
rect 75294 4834 75346 4846
rect 1344 4730 98560 4764
rect 1344 4678 8896 4730
rect 8948 4678 9020 4730
rect 9072 4678 9144 4730
rect 9196 4678 9268 4730
rect 9320 4678 17896 4730
rect 17948 4678 18020 4730
rect 18072 4678 18144 4730
rect 18196 4678 18268 4730
rect 18320 4678 26896 4730
rect 26948 4678 27020 4730
rect 27072 4678 27144 4730
rect 27196 4678 27268 4730
rect 27320 4678 35896 4730
rect 35948 4678 36020 4730
rect 36072 4678 36144 4730
rect 36196 4678 36268 4730
rect 36320 4678 44896 4730
rect 44948 4678 45020 4730
rect 45072 4678 45144 4730
rect 45196 4678 45268 4730
rect 45320 4678 53896 4730
rect 53948 4678 54020 4730
rect 54072 4678 54144 4730
rect 54196 4678 54268 4730
rect 54320 4678 62896 4730
rect 62948 4678 63020 4730
rect 63072 4678 63144 4730
rect 63196 4678 63268 4730
rect 63320 4678 71896 4730
rect 71948 4678 72020 4730
rect 72072 4678 72144 4730
rect 72196 4678 72268 4730
rect 72320 4678 80896 4730
rect 80948 4678 81020 4730
rect 81072 4678 81144 4730
rect 81196 4678 81268 4730
rect 81320 4678 89896 4730
rect 89948 4678 90020 4730
rect 90072 4678 90144 4730
rect 90196 4678 90268 4730
rect 90320 4678 98560 4730
rect 1344 4644 98560 4678
rect 34526 4562 34578 4574
rect 34526 4498 34578 4510
rect 49870 4562 49922 4574
rect 49870 4498 49922 4510
rect 63198 4562 63250 4574
rect 63198 4498 63250 4510
rect 70142 4562 70194 4574
rect 70142 4498 70194 4510
rect 70926 4562 70978 4574
rect 70926 4498 70978 4510
rect 78430 4562 78482 4574
rect 96686 4562 96738 4574
rect 91186 4510 91198 4562
rect 91250 4510 91262 4562
rect 78430 4498 78482 4510
rect 96686 4498 96738 4510
rect 96910 4562 96962 4574
rect 96910 4498 96962 4510
rect 34078 4450 34130 4462
rect 41694 4450 41746 4462
rect 42254 4450 42306 4462
rect 49422 4450 49474 4462
rect 49982 4450 50034 4462
rect 62750 4450 62802 4462
rect 30146 4398 30158 4450
rect 30210 4398 30222 4450
rect 34402 4398 34414 4450
rect 34466 4398 34478 4450
rect 38322 4398 38334 4450
rect 38386 4398 38398 4450
rect 42018 4398 42030 4450
rect 42082 4398 42094 4450
rect 44146 4398 44158 4450
rect 44210 4398 44222 4450
rect 49746 4398 49758 4450
rect 49810 4398 49822 4450
rect 52770 4398 52782 4450
rect 52834 4398 52846 4450
rect 58706 4398 58718 4450
rect 58770 4398 58782 4450
rect 34078 4386 34130 4398
rect 41694 4386 41746 4398
rect 42254 4386 42306 4398
rect 49422 4386 49474 4398
rect 49982 4386 50034 4398
rect 62750 4386 62802 4398
rect 63534 4450 63586 4462
rect 71374 4450 71426 4462
rect 78318 4450 78370 4462
rect 65762 4398 65774 4450
rect 65826 4398 65838 4450
rect 75618 4398 75630 4450
rect 75682 4398 75694 4450
rect 82114 4398 82126 4450
rect 82178 4398 82190 4450
rect 63534 4386 63586 4398
rect 71374 4386 71426 4398
rect 78318 4386 78370 4398
rect 33854 4338 33906 4350
rect 31042 4286 31054 4338
rect 31106 4286 31118 4338
rect 33854 4274 33906 4286
rect 34638 4338 34690 4350
rect 41358 4338 41410 4350
rect 40226 4286 40238 4338
rect 40290 4286 40302 4338
rect 34638 4274 34690 4286
rect 41358 4274 41410 4286
rect 41470 4338 41522 4350
rect 49086 4338 49138 4350
rect 48178 4286 48190 4338
rect 48242 4286 48254 4338
rect 51314 4286 51326 4338
rect 51378 4286 51390 4338
rect 61842 4286 61854 4338
rect 61906 4286 61918 4338
rect 68898 4286 68910 4338
rect 68962 4286 68974 4338
rect 70018 4286 70030 4338
rect 70082 4286 70094 4338
rect 70690 4286 70702 4338
rect 70754 4286 70766 4338
rect 71026 4286 71038 4338
rect 71090 4286 71102 4338
rect 72818 4286 72830 4338
rect 72882 4286 72894 4338
rect 81554 4286 81566 4338
rect 81618 4286 81630 4338
rect 88050 4286 88062 4338
rect 88114 4286 88126 4338
rect 41470 4274 41522 4286
rect 49086 4274 49138 4286
rect 33406 4226 33458 4238
rect 62190 4226 62242 4238
rect 42354 4174 42366 4226
rect 42418 4174 42430 4226
rect 33406 4162 33458 4174
rect 62190 4162 62242 4174
rect 71710 4226 71762 4238
rect 71710 4162 71762 4174
rect 77982 4226 78034 4238
rect 77982 4162 78034 4174
rect 78878 4226 78930 4238
rect 78878 4162 78930 4174
rect 85934 4226 85986 4238
rect 85934 4162 85986 4174
rect 33742 4114 33794 4126
rect 33742 4050 33794 4062
rect 41022 4114 41074 4126
rect 41022 4050 41074 4062
rect 49198 4114 49250 4126
rect 49198 4050 49250 4062
rect 71598 4114 71650 4126
rect 71598 4050 71650 4062
rect 79438 4114 79490 4126
rect 79438 4050 79490 4062
rect 97694 4114 97746 4126
rect 97694 4050 97746 4062
rect 1344 3946 98560 3980
rect 1344 3894 4396 3946
rect 4448 3894 4520 3946
rect 4572 3894 4644 3946
rect 4696 3894 4768 3946
rect 4820 3894 13396 3946
rect 13448 3894 13520 3946
rect 13572 3894 13644 3946
rect 13696 3894 13768 3946
rect 13820 3894 22396 3946
rect 22448 3894 22520 3946
rect 22572 3894 22644 3946
rect 22696 3894 22768 3946
rect 22820 3894 31396 3946
rect 31448 3894 31520 3946
rect 31572 3894 31644 3946
rect 31696 3894 31768 3946
rect 31820 3894 40396 3946
rect 40448 3894 40520 3946
rect 40572 3894 40644 3946
rect 40696 3894 40768 3946
rect 40820 3894 49396 3946
rect 49448 3894 49520 3946
rect 49572 3894 49644 3946
rect 49696 3894 49768 3946
rect 49820 3894 58396 3946
rect 58448 3894 58520 3946
rect 58572 3894 58644 3946
rect 58696 3894 58768 3946
rect 58820 3894 67396 3946
rect 67448 3894 67520 3946
rect 67572 3894 67644 3946
rect 67696 3894 67768 3946
rect 67820 3894 76396 3946
rect 76448 3894 76520 3946
rect 76572 3894 76644 3946
rect 76696 3894 76768 3946
rect 76820 3894 85396 3946
rect 85448 3894 85520 3946
rect 85572 3894 85644 3946
rect 85696 3894 85768 3946
rect 85820 3894 94396 3946
rect 94448 3894 94520 3946
rect 94572 3894 94644 3946
rect 94696 3894 94768 3946
rect 94820 3894 98560 3946
rect 1344 3860 98560 3894
rect 34190 3778 34242 3790
rect 34190 3714 34242 3726
rect 34302 3778 34354 3790
rect 34302 3714 34354 3726
rect 34638 3778 34690 3790
rect 39230 3778 39282 3790
rect 37090 3726 37102 3778
rect 37154 3775 37166 3778
rect 38546 3775 38558 3778
rect 37154 3729 38558 3775
rect 37154 3726 37166 3729
rect 38546 3726 38558 3729
rect 38610 3726 38622 3778
rect 34638 3714 34690 3726
rect 39230 3714 39282 3726
rect 41022 3778 41074 3790
rect 41022 3714 41074 3726
rect 44046 3778 44098 3790
rect 44046 3714 44098 3726
rect 44830 3778 44882 3790
rect 44830 3714 44882 3726
rect 45166 3778 45218 3790
rect 45166 3714 45218 3726
rect 45278 3778 45330 3790
rect 45278 3714 45330 3726
rect 45950 3778 46002 3790
rect 45950 3714 46002 3726
rect 46846 3778 46898 3790
rect 46846 3714 46898 3726
rect 58270 3778 58322 3790
rect 58270 3714 58322 3726
rect 60846 3778 60898 3790
rect 60846 3714 60898 3726
rect 69582 3778 69634 3790
rect 69582 3714 69634 3726
rect 77982 3778 78034 3790
rect 77982 3714 78034 3726
rect 17838 3666 17890 3678
rect 31278 3666 31330 3678
rect 28802 3614 28814 3666
rect 28866 3614 28878 3666
rect 17838 3602 17890 3614
rect 31278 3602 31330 3614
rect 32510 3666 32562 3678
rect 32510 3602 32562 3614
rect 33070 3666 33122 3678
rect 35198 3666 35250 3678
rect 33394 3614 33406 3666
rect 33458 3614 33470 3666
rect 33070 3602 33122 3614
rect 35198 3602 35250 3614
rect 36542 3666 36594 3678
rect 36542 3602 36594 3614
rect 38782 3666 38834 3678
rect 38782 3602 38834 3614
rect 40910 3666 40962 3678
rect 44270 3666 44322 3678
rect 48526 3666 48578 3678
rect 51438 3666 51490 3678
rect 41906 3614 41918 3666
rect 41970 3614 41982 3666
rect 47730 3614 47742 3666
rect 47794 3614 47806 3666
rect 50306 3614 50318 3666
rect 50370 3614 50382 3666
rect 40910 3602 40962 3614
rect 44270 3602 44322 3614
rect 48526 3602 48578 3614
rect 51438 3602 51490 3614
rect 51886 3666 51938 3678
rect 51886 3602 51938 3614
rect 52334 3666 52386 3678
rect 57486 3666 57538 3678
rect 60734 3666 60786 3678
rect 55458 3614 55470 3666
rect 55522 3614 55534 3666
rect 59042 3614 59054 3666
rect 59106 3614 59118 3666
rect 52334 3602 52386 3614
rect 57486 3602 57538 3614
rect 60734 3602 60786 3614
rect 61742 3666 61794 3678
rect 61742 3602 61794 3614
rect 62750 3666 62802 3678
rect 62750 3602 62802 3614
rect 67454 3666 67506 3678
rect 67454 3602 67506 3614
rect 71038 3666 71090 3678
rect 71038 3602 71090 3614
rect 74286 3666 74338 3678
rect 74286 3602 74338 3614
rect 75518 3666 75570 3678
rect 82462 3666 82514 3678
rect 79986 3614 79998 3666
rect 80050 3614 80062 3666
rect 75518 3602 75570 3614
rect 82462 3602 82514 3614
rect 84702 3666 84754 3678
rect 96350 3666 96402 3678
rect 85698 3614 85710 3666
rect 85762 3614 85774 3666
rect 84702 3602 84754 3614
rect 96350 3602 96402 3614
rect 31726 3554 31778 3566
rect 34750 3554 34802 3566
rect 33282 3502 33294 3554
rect 33346 3502 33358 3554
rect 31726 3490 31778 3502
rect 34750 3490 34802 3502
rect 36094 3554 36146 3566
rect 36094 3490 36146 3502
rect 37438 3554 37490 3566
rect 37438 3490 37490 3502
rect 37886 3554 37938 3566
rect 37886 3490 37938 3502
rect 38334 3554 38386 3566
rect 38334 3490 38386 3502
rect 39118 3554 39170 3566
rect 39118 3490 39170 3502
rect 40350 3554 40402 3566
rect 41806 3554 41858 3566
rect 41570 3502 41582 3554
rect 41634 3502 41646 3554
rect 40350 3490 40402 3502
rect 41806 3490 41858 3502
rect 42478 3554 42530 3566
rect 42478 3490 42530 3502
rect 42926 3554 42978 3566
rect 42926 3490 42978 3502
rect 43486 3554 43538 3566
rect 43486 3490 43538 3502
rect 44494 3554 44546 3566
rect 44494 3490 44546 3502
rect 44942 3554 44994 3566
rect 49310 3554 49362 3566
rect 47954 3502 47966 3554
rect 48018 3502 48030 3554
rect 44942 3490 44994 3502
rect 49310 3490 49362 3502
rect 49422 3554 49474 3566
rect 50206 3554 50258 3566
rect 49970 3502 49982 3554
rect 50034 3502 50046 3554
rect 49422 3490 49474 3502
rect 50206 3490 50258 3502
rect 54574 3554 54626 3566
rect 54574 3490 54626 3502
rect 55022 3554 55074 3566
rect 55022 3490 55074 3502
rect 57822 3554 57874 3566
rect 57822 3490 57874 3502
rect 58158 3554 58210 3566
rect 60062 3554 60114 3566
rect 63198 3554 63250 3566
rect 59378 3502 59390 3554
rect 59442 3502 59454 3554
rect 60162 3502 60174 3554
rect 60226 3502 60238 3554
rect 61282 3502 61294 3554
rect 61346 3502 61358 3554
rect 58158 3490 58210 3502
rect 60062 3490 60114 3502
rect 63198 3490 63250 3502
rect 65998 3554 66050 3566
rect 82798 3554 82850 3566
rect 96910 3554 96962 3566
rect 66434 3502 66446 3554
rect 66498 3502 66510 3554
rect 71250 3502 71262 3554
rect 71314 3502 71326 3554
rect 77298 3502 77310 3554
rect 77362 3502 77374 3554
rect 78082 3502 78094 3554
rect 78146 3502 78158 3554
rect 80658 3502 80670 3554
rect 80722 3502 80734 3554
rect 86146 3502 86158 3554
rect 86210 3502 86222 3554
rect 94322 3502 94334 3554
rect 94386 3502 94398 3554
rect 65998 3490 66050 3502
rect 82798 3490 82850 3502
rect 96910 3490 96962 3502
rect 6078 3442 6130 3454
rect 6078 3378 6130 3390
rect 6302 3442 6354 3454
rect 6302 3378 6354 3390
rect 6638 3442 6690 3454
rect 6638 3378 6690 3390
rect 16494 3442 16546 3454
rect 16494 3378 16546 3390
rect 17278 3442 17330 3454
rect 17278 3378 17330 3390
rect 27918 3442 27970 3454
rect 27918 3378 27970 3390
rect 28366 3442 28418 3454
rect 33966 3442 34018 3454
rect 33618 3390 33630 3442
rect 33682 3390 33694 3442
rect 28366 3378 28418 3390
rect 33966 3378 34018 3390
rect 37102 3442 37154 3454
rect 37102 3378 37154 3390
rect 39790 3442 39842 3454
rect 39790 3378 39842 3390
rect 41246 3442 41298 3454
rect 41246 3378 41298 3390
rect 42590 3442 42642 3454
rect 46734 3442 46786 3454
rect 43810 3390 43822 3442
rect 43874 3390 43886 3442
rect 42590 3378 42642 3390
rect 46734 3378 46786 3390
rect 48862 3442 48914 3454
rect 48862 3378 48914 3390
rect 49758 3442 49810 3454
rect 49758 3378 49810 3390
rect 52670 3442 52722 3454
rect 52670 3378 52722 3390
rect 59950 3442 60002 3454
rect 59950 3378 60002 3390
rect 60510 3442 60562 3454
rect 60510 3378 60562 3390
rect 69694 3442 69746 3454
rect 69694 3378 69746 3390
rect 71822 3442 71874 3454
rect 71822 3378 71874 3390
rect 73278 3442 73330 3454
rect 73278 3378 73330 3390
rect 76750 3442 76802 3454
rect 76750 3378 76802 3390
rect 83246 3442 83298 3454
rect 83246 3378 83298 3390
rect 93886 3442 93938 3454
rect 93886 3378 93938 3390
rect 94110 3442 94162 3454
rect 94110 3378 94162 3390
rect 97694 3442 97746 3454
rect 97694 3378 97746 3390
rect 43038 3330 43090 3342
rect 46398 3330 46450 3342
rect 43922 3278 43934 3330
rect 43986 3278 43998 3330
rect 43038 3266 43090 3278
rect 46398 3266 46450 3278
rect 72718 3330 72770 3342
rect 72718 3266 72770 3278
rect 75854 3330 75906 3342
rect 75854 3266 75906 3278
rect 81902 3330 81954 3342
rect 81902 3266 81954 3278
rect 1344 3162 98560 3196
rect 1344 3110 8896 3162
rect 8948 3110 9020 3162
rect 9072 3110 9144 3162
rect 9196 3110 9268 3162
rect 9320 3110 17896 3162
rect 17948 3110 18020 3162
rect 18072 3110 18144 3162
rect 18196 3110 18268 3162
rect 18320 3110 26896 3162
rect 26948 3110 27020 3162
rect 27072 3110 27144 3162
rect 27196 3110 27268 3162
rect 27320 3110 35896 3162
rect 35948 3110 36020 3162
rect 36072 3110 36144 3162
rect 36196 3110 36268 3162
rect 36320 3110 44896 3162
rect 44948 3110 45020 3162
rect 45072 3110 45144 3162
rect 45196 3110 45268 3162
rect 45320 3110 53896 3162
rect 53948 3110 54020 3162
rect 54072 3110 54144 3162
rect 54196 3110 54268 3162
rect 54320 3110 62896 3162
rect 62948 3110 63020 3162
rect 63072 3110 63144 3162
rect 63196 3110 63268 3162
rect 63320 3110 71896 3162
rect 71948 3110 72020 3162
rect 72072 3110 72144 3162
rect 72196 3110 72268 3162
rect 72320 3110 80896 3162
rect 80948 3110 81020 3162
rect 81072 3110 81144 3162
rect 81196 3110 81268 3162
rect 81320 3110 89896 3162
rect 89948 3110 90020 3162
rect 90072 3110 90144 3162
rect 90196 3110 90268 3162
rect 90320 3110 98560 3162
rect 1344 3076 98560 3110
<< via1 >>
rect 6750 56590 6802 56642
rect 7310 56590 7362 56642
rect 43710 56590 43762 56642
rect 44382 56590 44434 56642
rect 56030 56590 56082 56642
rect 57038 56590 57090 56642
rect 80670 56590 80722 56642
rect 82238 56590 82290 56642
rect 92990 56590 93042 56642
rect 93998 56590 94050 56642
rect 8896 56422 8948 56474
rect 9020 56422 9072 56474
rect 9144 56422 9196 56474
rect 9268 56422 9320 56474
rect 17896 56422 17948 56474
rect 18020 56422 18072 56474
rect 18144 56422 18196 56474
rect 18268 56422 18320 56474
rect 26896 56422 26948 56474
rect 27020 56422 27072 56474
rect 27144 56422 27196 56474
rect 27268 56422 27320 56474
rect 35896 56422 35948 56474
rect 36020 56422 36072 56474
rect 36144 56422 36196 56474
rect 36268 56422 36320 56474
rect 44896 56422 44948 56474
rect 45020 56422 45072 56474
rect 45144 56422 45196 56474
rect 45268 56422 45320 56474
rect 53896 56422 53948 56474
rect 54020 56422 54072 56474
rect 54144 56422 54196 56474
rect 54268 56422 54320 56474
rect 62896 56422 62948 56474
rect 63020 56422 63072 56474
rect 63144 56422 63196 56474
rect 63268 56422 63320 56474
rect 71896 56422 71948 56474
rect 72020 56422 72072 56474
rect 72144 56422 72196 56474
rect 72268 56422 72320 56474
rect 80896 56422 80948 56474
rect 81020 56422 81072 56474
rect 81144 56422 81196 56474
rect 81268 56422 81320 56474
rect 89896 56422 89948 56474
rect 90020 56422 90072 56474
rect 90144 56422 90196 56474
rect 90268 56422 90320 56474
rect 32174 56254 32226 56306
rect 57038 56254 57090 56306
rect 93998 56254 94050 56306
rect 97694 56254 97746 56306
rect 2046 56142 2098 56194
rect 7310 56142 7362 56194
rect 1710 56030 1762 56082
rect 8206 56030 8258 56082
rect 20078 56030 20130 56082
rect 32846 56030 32898 56082
rect 43934 56030 43986 56082
rect 56254 56030 56306 56082
rect 68462 56030 68514 56082
rect 81678 56030 81730 56082
rect 93214 56030 93266 56082
rect 96350 56030 96402 56082
rect 96910 56030 96962 56082
rect 98142 56030 98194 56082
rect 2494 55918 2546 55970
rect 8766 55918 8818 55970
rect 19182 55918 19234 55970
rect 44382 55918 44434 55970
rect 69022 55918 69074 55970
rect 82238 55918 82290 55970
rect 95902 55918 95954 55970
rect 4396 55638 4448 55690
rect 4520 55638 4572 55690
rect 4644 55638 4696 55690
rect 4768 55638 4820 55690
rect 13396 55638 13448 55690
rect 13520 55638 13572 55690
rect 13644 55638 13696 55690
rect 13768 55638 13820 55690
rect 22396 55638 22448 55690
rect 22520 55638 22572 55690
rect 22644 55638 22696 55690
rect 22768 55638 22820 55690
rect 31396 55638 31448 55690
rect 31520 55638 31572 55690
rect 31644 55638 31696 55690
rect 31768 55638 31820 55690
rect 40396 55638 40448 55690
rect 40520 55638 40572 55690
rect 40644 55638 40696 55690
rect 40768 55638 40820 55690
rect 49396 55638 49448 55690
rect 49520 55638 49572 55690
rect 49644 55638 49696 55690
rect 49768 55638 49820 55690
rect 58396 55638 58448 55690
rect 58520 55638 58572 55690
rect 58644 55638 58696 55690
rect 58768 55638 58820 55690
rect 67396 55638 67448 55690
rect 67520 55638 67572 55690
rect 67644 55638 67696 55690
rect 67768 55638 67820 55690
rect 76396 55638 76448 55690
rect 76520 55638 76572 55690
rect 76644 55638 76696 55690
rect 76768 55638 76820 55690
rect 85396 55638 85448 55690
rect 85520 55638 85572 55690
rect 85644 55638 85696 55690
rect 85768 55638 85820 55690
rect 94396 55638 94448 55690
rect 94520 55638 94572 55690
rect 94644 55638 94696 55690
rect 94768 55638 94820 55690
rect 32062 55358 32114 55410
rect 36430 55358 36482 55410
rect 42590 55358 42642 55410
rect 48078 55358 48130 55410
rect 29262 55246 29314 55298
rect 33182 55246 33234 55298
rect 33630 55246 33682 55298
rect 37102 55246 37154 55298
rect 39790 55246 39842 55298
rect 43710 55246 43762 55298
rect 44270 55246 44322 55298
rect 45166 55246 45218 55298
rect 55806 55246 55858 55298
rect 66894 55246 66946 55298
rect 97022 55246 97074 55298
rect 1710 55134 1762 55186
rect 25454 55134 25506 55186
rect 25790 55134 25842 55186
rect 26126 55134 26178 55186
rect 26462 55134 26514 55186
rect 29934 55134 29986 55186
rect 32398 55134 32450 55186
rect 32734 55134 32786 55186
rect 34302 55134 34354 55186
rect 40462 55134 40514 55186
rect 42926 55134 42978 55186
rect 43262 55134 43314 55186
rect 45950 55134 46002 55186
rect 56030 55134 56082 55186
rect 58494 55134 58546 55186
rect 67118 55134 67170 55186
rect 68350 55134 68402 55186
rect 98030 55134 98082 55186
rect 2046 55022 2098 55074
rect 2494 55022 2546 55074
rect 48638 55022 48690 55074
rect 52222 55022 52274 55074
rect 52670 55022 52722 55074
rect 52782 55022 52834 55074
rect 52894 55022 52946 55074
rect 53118 55022 53170 55074
rect 57262 55022 57314 55074
rect 57486 55022 57538 55074
rect 57598 55022 57650 55074
rect 57710 55022 57762 55074
rect 57934 55022 57986 55074
rect 58382 55022 58434 55074
rect 68686 55022 68738 55074
rect 96574 55022 96626 55074
rect 8896 54854 8948 54906
rect 9020 54854 9072 54906
rect 9144 54854 9196 54906
rect 9268 54854 9320 54906
rect 17896 54854 17948 54906
rect 18020 54854 18072 54906
rect 18144 54854 18196 54906
rect 18268 54854 18320 54906
rect 26896 54854 26948 54906
rect 27020 54854 27072 54906
rect 27144 54854 27196 54906
rect 27268 54854 27320 54906
rect 35896 54854 35948 54906
rect 36020 54854 36072 54906
rect 36144 54854 36196 54906
rect 36268 54854 36320 54906
rect 44896 54854 44948 54906
rect 45020 54854 45072 54906
rect 45144 54854 45196 54906
rect 45268 54854 45320 54906
rect 53896 54854 53948 54906
rect 54020 54854 54072 54906
rect 54144 54854 54196 54906
rect 54268 54854 54320 54906
rect 62896 54854 62948 54906
rect 63020 54854 63072 54906
rect 63144 54854 63196 54906
rect 63268 54854 63320 54906
rect 71896 54854 71948 54906
rect 72020 54854 72072 54906
rect 72144 54854 72196 54906
rect 72268 54854 72320 54906
rect 80896 54854 80948 54906
rect 81020 54854 81072 54906
rect 81144 54854 81196 54906
rect 81268 54854 81320 54906
rect 89896 54854 89948 54906
rect 90020 54854 90072 54906
rect 90144 54854 90196 54906
rect 90268 54854 90320 54906
rect 40350 54686 40402 54738
rect 41246 54686 41298 54738
rect 41358 54686 41410 54738
rect 48862 54686 48914 54738
rect 49646 54686 49698 54738
rect 82126 54686 82178 54738
rect 44606 54574 44658 54626
rect 47742 54574 47794 54626
rect 47966 54574 48018 54626
rect 49758 54574 49810 54626
rect 51774 54574 51826 54626
rect 56814 54574 56866 54626
rect 57486 54574 57538 54626
rect 60510 54574 60562 54626
rect 40238 54462 40290 54514
rect 40910 54462 40962 54514
rect 41470 54462 41522 54514
rect 43262 54462 43314 54514
rect 44830 54462 44882 54514
rect 45166 54462 45218 54514
rect 47294 54462 47346 54514
rect 48750 54462 48802 54514
rect 48974 54462 49026 54514
rect 49422 54462 49474 54514
rect 50990 54462 51042 54514
rect 54350 54462 54402 54514
rect 55582 54462 55634 54514
rect 56030 54462 56082 54514
rect 56590 54462 56642 54514
rect 61294 54462 61346 54514
rect 81790 54462 81842 54514
rect 35198 54350 35250 54402
rect 36318 54350 36370 54402
rect 36766 54350 36818 54402
rect 39902 54350 39954 54402
rect 41918 54350 41970 54402
rect 44158 54350 44210 54402
rect 45502 54350 45554 54402
rect 45950 54350 46002 54402
rect 48078 54350 48130 54402
rect 50654 54350 50706 54402
rect 53902 54350 53954 54402
rect 57822 54350 57874 54402
rect 58382 54350 58434 54402
rect 61854 54350 61906 54402
rect 65774 54350 65826 54402
rect 81454 54350 81506 54402
rect 44942 54238 44994 54290
rect 47070 54238 47122 54290
rect 54238 54238 54290 54290
rect 4396 54070 4448 54122
rect 4520 54070 4572 54122
rect 4644 54070 4696 54122
rect 4768 54070 4820 54122
rect 13396 54070 13448 54122
rect 13520 54070 13572 54122
rect 13644 54070 13696 54122
rect 13768 54070 13820 54122
rect 22396 54070 22448 54122
rect 22520 54070 22572 54122
rect 22644 54070 22696 54122
rect 22768 54070 22820 54122
rect 31396 54070 31448 54122
rect 31520 54070 31572 54122
rect 31644 54070 31696 54122
rect 31768 54070 31820 54122
rect 40396 54070 40448 54122
rect 40520 54070 40572 54122
rect 40644 54070 40696 54122
rect 40768 54070 40820 54122
rect 49396 54070 49448 54122
rect 49520 54070 49572 54122
rect 49644 54070 49696 54122
rect 49768 54070 49820 54122
rect 58396 54070 58448 54122
rect 58520 54070 58572 54122
rect 58644 54070 58696 54122
rect 58768 54070 58820 54122
rect 67396 54070 67448 54122
rect 67520 54070 67572 54122
rect 67644 54070 67696 54122
rect 67768 54070 67820 54122
rect 76396 54070 76448 54122
rect 76520 54070 76572 54122
rect 76644 54070 76696 54122
rect 76768 54070 76820 54122
rect 85396 54070 85448 54122
rect 85520 54070 85572 54122
rect 85644 54070 85696 54122
rect 85768 54070 85820 54122
rect 94396 54070 94448 54122
rect 94520 54070 94572 54122
rect 94644 54070 94696 54122
rect 94768 54070 94820 54122
rect 59278 53902 59330 53954
rect 30046 53790 30098 53842
rect 34526 53790 34578 53842
rect 35310 53790 35362 53842
rect 36318 53790 36370 53842
rect 48750 53790 48802 53842
rect 59166 53790 59218 53842
rect 65326 53790 65378 53842
rect 72830 53790 72882 53842
rect 28478 53678 28530 53730
rect 29598 53678 29650 53730
rect 35086 53678 35138 53730
rect 35646 53678 35698 53730
rect 37214 53678 37266 53730
rect 38222 53678 38274 53730
rect 41358 53678 41410 53730
rect 41694 53678 41746 53730
rect 44942 53678 44994 53730
rect 46062 53678 46114 53730
rect 52782 53678 52834 53730
rect 56590 53678 56642 53730
rect 56814 53678 56866 53730
rect 57486 53678 57538 53730
rect 65214 53678 65266 53730
rect 65438 53678 65490 53730
rect 65998 53678 66050 53730
rect 66334 53678 66386 53730
rect 66558 53678 66610 53730
rect 66782 53678 66834 53730
rect 67118 53678 67170 53730
rect 69918 53678 69970 53730
rect 96910 53678 96962 53730
rect 1710 53566 1762 53618
rect 30830 53566 30882 53618
rect 35870 53566 35922 53618
rect 37326 53566 37378 53618
rect 38894 53566 38946 53618
rect 40798 53566 40850 53618
rect 42254 53566 42306 53618
rect 52894 53566 52946 53618
rect 56478 53566 56530 53618
rect 64878 53566 64930 53618
rect 66670 53566 66722 53618
rect 67230 53566 67282 53618
rect 70702 53566 70754 53618
rect 98030 53566 98082 53618
rect 2046 53454 2098 53506
rect 2494 53454 2546 53506
rect 29262 53454 29314 53506
rect 29934 53454 29986 53506
rect 30158 53454 30210 53506
rect 30718 53454 30770 53506
rect 31278 53454 31330 53506
rect 34414 53454 34466 53506
rect 34638 53454 34690 53506
rect 35422 53454 35474 53506
rect 36206 53454 36258 53506
rect 38334 53454 38386 53506
rect 41246 53454 41298 53506
rect 43822 53454 43874 53506
rect 44270 53454 44322 53506
rect 52110 53454 52162 53506
rect 56366 53454 56418 53506
rect 57262 53454 57314 53506
rect 57374 53454 57426 53506
rect 57934 53454 57986 53506
rect 59054 53454 59106 53506
rect 64542 53454 64594 53506
rect 65662 53454 65714 53506
rect 67678 53454 67730 53506
rect 69582 53454 69634 53506
rect 8896 53286 8948 53338
rect 9020 53286 9072 53338
rect 9144 53286 9196 53338
rect 9268 53286 9320 53338
rect 17896 53286 17948 53338
rect 18020 53286 18072 53338
rect 18144 53286 18196 53338
rect 18268 53286 18320 53338
rect 26896 53286 26948 53338
rect 27020 53286 27072 53338
rect 27144 53286 27196 53338
rect 27268 53286 27320 53338
rect 35896 53286 35948 53338
rect 36020 53286 36072 53338
rect 36144 53286 36196 53338
rect 36268 53286 36320 53338
rect 44896 53286 44948 53338
rect 45020 53286 45072 53338
rect 45144 53286 45196 53338
rect 45268 53286 45320 53338
rect 53896 53286 53948 53338
rect 54020 53286 54072 53338
rect 54144 53286 54196 53338
rect 54268 53286 54320 53338
rect 62896 53286 62948 53338
rect 63020 53286 63072 53338
rect 63144 53286 63196 53338
rect 63268 53286 63320 53338
rect 71896 53286 71948 53338
rect 72020 53286 72072 53338
rect 72144 53286 72196 53338
rect 72268 53286 72320 53338
rect 80896 53286 80948 53338
rect 81020 53286 81072 53338
rect 81144 53286 81196 53338
rect 81268 53286 81320 53338
rect 89896 53286 89948 53338
rect 90020 53286 90072 53338
rect 90144 53286 90196 53338
rect 90268 53286 90320 53338
rect 29038 53118 29090 53170
rect 33854 53118 33906 53170
rect 35534 53118 35586 53170
rect 35870 53118 35922 53170
rect 36990 53118 37042 53170
rect 39230 53118 39282 53170
rect 39454 53118 39506 53170
rect 48862 53118 48914 53170
rect 48974 53118 49026 53170
rect 51214 53118 51266 53170
rect 51662 53118 51714 53170
rect 60174 53118 60226 53170
rect 2046 53006 2098 53058
rect 27694 53006 27746 53058
rect 29598 53006 29650 53058
rect 29822 53006 29874 53058
rect 33742 53006 33794 53058
rect 35198 53006 35250 53058
rect 1710 52894 1762 52946
rect 27918 52894 27970 52946
rect 28142 52894 28194 52946
rect 28590 52894 28642 52946
rect 28814 52894 28866 52946
rect 35646 52950 35698 53002
rect 40910 53006 40962 53058
rect 45502 53006 45554 53058
rect 49758 53006 49810 53058
rect 50430 53006 50482 53058
rect 50766 53006 50818 53058
rect 58046 53006 58098 53058
rect 59502 53006 59554 53058
rect 65998 53006 66050 53058
rect 29150 52894 29202 52946
rect 30382 52894 30434 52946
rect 31278 52894 31330 52946
rect 34302 52894 34354 52946
rect 35310 52894 35362 52946
rect 36206 52894 36258 52946
rect 39678 52894 39730 52946
rect 41134 52894 41186 52946
rect 41358 52894 41410 52946
rect 41582 52894 41634 52946
rect 46622 52894 46674 52946
rect 49086 52894 49138 52946
rect 49422 52894 49474 52946
rect 50206 52894 50258 52946
rect 50990 52894 51042 52946
rect 55582 52894 55634 52946
rect 56926 52894 56978 52946
rect 58942 52894 58994 52946
rect 65214 52894 65266 52946
rect 68798 52894 68850 52946
rect 2494 52782 2546 52834
rect 28030 52782 28082 52834
rect 29710 52782 29762 52834
rect 30830 52782 30882 52834
rect 36542 52782 36594 52834
rect 38446 52782 38498 52834
rect 38894 52782 38946 52834
rect 39566 52782 39618 52834
rect 40126 52782 40178 52834
rect 41022 52782 41074 52834
rect 48190 52782 48242 52834
rect 50318 52782 50370 52834
rect 50878 52782 50930 52834
rect 52446 52782 52498 52834
rect 55134 52782 55186 52834
rect 56030 52782 56082 52834
rect 68126 52782 68178 52834
rect 28478 52670 28530 52722
rect 30046 52670 30098 52722
rect 49982 52670 50034 52722
rect 55022 52670 55074 52722
rect 55582 52670 55634 52722
rect 4396 52502 4448 52554
rect 4520 52502 4572 52554
rect 4644 52502 4696 52554
rect 4768 52502 4820 52554
rect 13396 52502 13448 52554
rect 13520 52502 13572 52554
rect 13644 52502 13696 52554
rect 13768 52502 13820 52554
rect 22396 52502 22448 52554
rect 22520 52502 22572 52554
rect 22644 52502 22696 52554
rect 22768 52502 22820 52554
rect 31396 52502 31448 52554
rect 31520 52502 31572 52554
rect 31644 52502 31696 52554
rect 31768 52502 31820 52554
rect 40396 52502 40448 52554
rect 40520 52502 40572 52554
rect 40644 52502 40696 52554
rect 40768 52502 40820 52554
rect 49396 52502 49448 52554
rect 49520 52502 49572 52554
rect 49644 52502 49696 52554
rect 49768 52502 49820 52554
rect 58396 52502 58448 52554
rect 58520 52502 58572 52554
rect 58644 52502 58696 52554
rect 58768 52502 58820 52554
rect 67396 52502 67448 52554
rect 67520 52502 67572 52554
rect 67644 52502 67696 52554
rect 67768 52502 67820 52554
rect 76396 52502 76448 52554
rect 76520 52502 76572 52554
rect 76644 52502 76696 52554
rect 76768 52502 76820 52554
rect 85396 52502 85448 52554
rect 85520 52502 85572 52554
rect 85644 52502 85696 52554
rect 85768 52502 85820 52554
rect 94396 52502 94448 52554
rect 94520 52502 94572 52554
rect 94644 52502 94696 52554
rect 94768 52502 94820 52554
rect 27918 52334 27970 52386
rect 28478 52334 28530 52386
rect 33294 52334 33346 52386
rect 41918 52334 41970 52386
rect 48750 52334 48802 52386
rect 49758 52334 49810 52386
rect 57822 52334 57874 52386
rect 58494 52334 58546 52386
rect 65998 52334 66050 52386
rect 22990 52222 23042 52274
rect 25118 52222 25170 52274
rect 28366 52222 28418 52274
rect 29262 52222 29314 52274
rect 30046 52222 30098 52274
rect 31726 52222 31778 52274
rect 32174 52222 32226 52274
rect 35758 52222 35810 52274
rect 45614 52222 45666 52274
rect 46734 52222 46786 52274
rect 47182 52222 47234 52274
rect 48302 52222 48354 52274
rect 48750 52222 48802 52274
rect 49198 52222 49250 52274
rect 50206 52222 50258 52274
rect 50766 52222 50818 52274
rect 51214 52222 51266 52274
rect 53342 52222 53394 52274
rect 53790 52222 53842 52274
rect 55694 52222 55746 52274
rect 58606 52222 58658 52274
rect 60510 52222 60562 52274
rect 62638 52222 62690 52274
rect 66110 52222 66162 52274
rect 66558 52222 66610 52274
rect 25902 52110 25954 52162
rect 26350 52110 26402 52162
rect 27582 52110 27634 52162
rect 28142 52110 28194 52162
rect 30158 52110 30210 52162
rect 31278 52110 31330 52162
rect 32958 52110 33010 52162
rect 33406 52110 33458 52162
rect 33742 52110 33794 52162
rect 34190 52110 34242 52162
rect 36206 52110 36258 52162
rect 43822 52110 43874 52162
rect 45950 52110 46002 52162
rect 46174 52110 46226 52162
rect 47742 52110 47794 52162
rect 49646 52110 49698 52162
rect 54350 52110 54402 52162
rect 55358 52110 55410 52162
rect 56590 52110 56642 52162
rect 56814 52110 56866 52162
rect 56926 52110 56978 52162
rect 57598 52110 57650 52162
rect 63422 52110 63474 52162
rect 63870 52110 63922 52162
rect 97694 52110 97746 52162
rect 26910 51998 26962 52050
rect 27806 51998 27858 52050
rect 29710 51998 29762 52050
rect 31166 51998 31218 52050
rect 49982 51998 50034 52050
rect 54462 51998 54514 52050
rect 56030 51998 56082 52050
rect 56366 51998 56418 52050
rect 57934 51998 57986 52050
rect 58158 51998 58210 52050
rect 27022 51886 27074 51938
rect 27134 51886 27186 51938
rect 32958 51886 33010 51938
rect 57150 51886 57202 51938
rect 96910 51886 96962 51938
rect 8896 51718 8948 51770
rect 9020 51718 9072 51770
rect 9144 51718 9196 51770
rect 9268 51718 9320 51770
rect 17896 51718 17948 51770
rect 18020 51718 18072 51770
rect 18144 51718 18196 51770
rect 18268 51718 18320 51770
rect 26896 51718 26948 51770
rect 27020 51718 27072 51770
rect 27144 51718 27196 51770
rect 27268 51718 27320 51770
rect 35896 51718 35948 51770
rect 36020 51718 36072 51770
rect 36144 51718 36196 51770
rect 36268 51718 36320 51770
rect 44896 51718 44948 51770
rect 45020 51718 45072 51770
rect 45144 51718 45196 51770
rect 45268 51718 45320 51770
rect 53896 51718 53948 51770
rect 54020 51718 54072 51770
rect 54144 51718 54196 51770
rect 54268 51718 54320 51770
rect 62896 51718 62948 51770
rect 63020 51718 63072 51770
rect 63144 51718 63196 51770
rect 63268 51718 63320 51770
rect 71896 51718 71948 51770
rect 72020 51718 72072 51770
rect 72144 51718 72196 51770
rect 72268 51718 72320 51770
rect 80896 51718 80948 51770
rect 81020 51718 81072 51770
rect 81144 51718 81196 51770
rect 81268 51718 81320 51770
rect 89896 51718 89948 51770
rect 90020 51718 90072 51770
rect 90144 51718 90196 51770
rect 90268 51718 90320 51770
rect 28814 51550 28866 51602
rect 37998 51550 38050 51602
rect 42702 51550 42754 51602
rect 43262 51550 43314 51602
rect 43710 51550 43762 51602
rect 44718 51550 44770 51602
rect 47854 51550 47906 51602
rect 50430 51550 50482 51602
rect 55806 51550 55858 51602
rect 57710 51550 57762 51602
rect 62078 51550 62130 51602
rect 90974 51550 91026 51602
rect 2046 51438 2098 51490
rect 11902 51438 11954 51490
rect 38670 51438 38722 51490
rect 40910 51438 40962 51490
rect 41022 51438 41074 51490
rect 41694 51438 41746 51490
rect 47070 51438 47122 51490
rect 70590 51438 70642 51490
rect 71038 51438 71090 51490
rect 71374 51438 71426 51490
rect 77086 51438 77138 51490
rect 1710 51326 1762 51378
rect 38446 51326 38498 51378
rect 39230 51326 39282 51378
rect 39678 51326 39730 51378
rect 41246 51326 41298 51378
rect 41470 51326 41522 51378
rect 42030 51326 42082 51378
rect 42254 51326 42306 51378
rect 44270 51326 44322 51378
rect 46174 51326 46226 51378
rect 46398 51326 46450 51378
rect 46734 51326 46786 51378
rect 47406 51326 47458 51378
rect 49982 51326 50034 51378
rect 62190 51326 62242 51378
rect 90750 51326 90802 51378
rect 2494 51214 2546 51266
rect 39790 51214 39842 51266
rect 40350 51214 40402 51266
rect 42814 51214 42866 51266
rect 55470 51214 55522 51266
rect 55694 51214 55746 51266
rect 57150 51214 57202 51266
rect 61742 51214 61794 51266
rect 76638 51214 76690 51266
rect 41582 51102 41634 51154
rect 57150 51102 57202 51154
rect 57486 51102 57538 51154
rect 4396 50934 4448 50986
rect 4520 50934 4572 50986
rect 4644 50934 4696 50986
rect 4768 50934 4820 50986
rect 13396 50934 13448 50986
rect 13520 50934 13572 50986
rect 13644 50934 13696 50986
rect 13768 50934 13820 50986
rect 22396 50934 22448 50986
rect 22520 50934 22572 50986
rect 22644 50934 22696 50986
rect 22768 50934 22820 50986
rect 31396 50934 31448 50986
rect 31520 50934 31572 50986
rect 31644 50934 31696 50986
rect 31768 50934 31820 50986
rect 40396 50934 40448 50986
rect 40520 50934 40572 50986
rect 40644 50934 40696 50986
rect 40768 50934 40820 50986
rect 49396 50934 49448 50986
rect 49520 50934 49572 50986
rect 49644 50934 49696 50986
rect 49768 50934 49820 50986
rect 58396 50934 58448 50986
rect 58520 50934 58572 50986
rect 58644 50934 58696 50986
rect 58768 50934 58820 50986
rect 67396 50934 67448 50986
rect 67520 50934 67572 50986
rect 67644 50934 67696 50986
rect 67768 50934 67820 50986
rect 76396 50934 76448 50986
rect 76520 50934 76572 50986
rect 76644 50934 76696 50986
rect 76768 50934 76820 50986
rect 85396 50934 85448 50986
rect 85520 50934 85572 50986
rect 85644 50934 85696 50986
rect 85768 50934 85820 50986
rect 94396 50934 94448 50986
rect 94520 50934 94572 50986
rect 94644 50934 94696 50986
rect 94768 50934 94820 50986
rect 27918 50766 27970 50818
rect 29374 50766 29426 50818
rect 32398 50766 32450 50818
rect 44270 50766 44322 50818
rect 49870 50766 49922 50818
rect 38558 50654 38610 50706
rect 39118 50654 39170 50706
rect 39566 50654 39618 50706
rect 55246 50654 55298 50706
rect 57374 50654 57426 50706
rect 58606 50654 58658 50706
rect 74286 50654 74338 50706
rect 16718 50542 16770 50594
rect 17278 50542 17330 50594
rect 29934 50542 29986 50594
rect 39902 50542 39954 50594
rect 40798 50542 40850 50594
rect 41246 50542 41298 50594
rect 45502 50542 45554 50594
rect 46174 50542 46226 50594
rect 46846 50542 46898 50594
rect 58046 50542 58098 50594
rect 60398 50542 60450 50594
rect 60958 50542 61010 50594
rect 70478 50542 70530 50594
rect 70926 50542 70978 50594
rect 76302 50542 76354 50594
rect 76974 50542 77026 50594
rect 77310 50542 77362 50594
rect 1710 50430 1762 50482
rect 2046 50430 2098 50482
rect 2494 50430 2546 50482
rect 16158 50430 16210 50482
rect 19630 50430 19682 50482
rect 20862 50430 20914 50482
rect 28030 50430 28082 50482
rect 29486 50430 29538 50482
rect 32286 50430 32338 50482
rect 32846 50430 32898 50482
rect 40462 50430 40514 50482
rect 46062 50430 46114 50482
rect 49086 50430 49138 50482
rect 63310 50430 63362 50482
rect 64094 50430 64146 50482
rect 64542 50430 64594 50482
rect 73166 50430 73218 50482
rect 73950 50430 74002 50482
rect 76526 50430 76578 50482
rect 79662 50430 79714 50482
rect 80446 50430 80498 50482
rect 96238 50430 96290 50482
rect 96574 50430 96626 50482
rect 5630 50318 5682 50370
rect 16494 50318 16546 50370
rect 20414 50318 20466 50370
rect 28478 50318 28530 50370
rect 43598 50318 43650 50370
rect 59950 50318 60002 50370
rect 65550 50318 65602 50370
rect 86830 50318 86882 50370
rect 8896 50150 8948 50202
rect 9020 50150 9072 50202
rect 9144 50150 9196 50202
rect 9268 50150 9320 50202
rect 17896 50150 17948 50202
rect 18020 50150 18072 50202
rect 18144 50150 18196 50202
rect 18268 50150 18320 50202
rect 26896 50150 26948 50202
rect 27020 50150 27072 50202
rect 27144 50150 27196 50202
rect 27268 50150 27320 50202
rect 35896 50150 35948 50202
rect 36020 50150 36072 50202
rect 36144 50150 36196 50202
rect 36268 50150 36320 50202
rect 44896 50150 44948 50202
rect 45020 50150 45072 50202
rect 45144 50150 45196 50202
rect 45268 50150 45320 50202
rect 53896 50150 53948 50202
rect 54020 50150 54072 50202
rect 54144 50150 54196 50202
rect 54268 50150 54320 50202
rect 62896 50150 62948 50202
rect 63020 50150 63072 50202
rect 63144 50150 63196 50202
rect 63268 50150 63320 50202
rect 71896 50150 71948 50202
rect 72020 50150 72072 50202
rect 72144 50150 72196 50202
rect 72268 50150 72320 50202
rect 80896 50150 80948 50202
rect 81020 50150 81072 50202
rect 81144 50150 81196 50202
rect 81268 50150 81320 50202
rect 89896 50150 89948 50202
rect 90020 50150 90072 50202
rect 90144 50150 90196 50202
rect 90268 50150 90320 50202
rect 8318 49982 8370 50034
rect 40350 49982 40402 50034
rect 60958 49982 61010 50034
rect 68126 49982 68178 50034
rect 69246 49982 69298 50034
rect 72382 49982 72434 50034
rect 75742 49982 75794 50034
rect 76862 49982 76914 50034
rect 1934 49870 1986 49922
rect 9550 49870 9602 49922
rect 10110 49870 10162 49922
rect 11342 49870 11394 49922
rect 14478 49870 14530 49922
rect 26238 49870 26290 49922
rect 29710 49870 29762 49922
rect 37662 49870 37714 49922
rect 51550 49870 51602 49922
rect 62302 49870 62354 49922
rect 62862 49870 62914 49922
rect 64990 49870 65042 49922
rect 72942 49870 72994 49922
rect 73502 49870 73554 49922
rect 77422 49870 77474 49922
rect 77758 49870 77810 49922
rect 86270 49870 86322 49922
rect 5518 49758 5570 49810
rect 5854 49758 5906 49810
rect 11678 49758 11730 49810
rect 12126 49758 12178 49810
rect 25566 49758 25618 49810
rect 29038 49758 29090 49810
rect 38446 49758 38498 49810
rect 42366 49758 42418 49810
rect 50430 49758 50482 49810
rect 50766 49758 50818 49810
rect 61294 49758 61346 49810
rect 61742 49758 61794 49810
rect 64766 49758 64818 49810
rect 65438 49758 65490 49810
rect 65774 49758 65826 49810
rect 77198 49758 77250 49810
rect 86046 49758 86098 49810
rect 96910 49758 96962 49810
rect 2494 49646 2546 49698
rect 28478 49646 28530 49698
rect 31950 49646 32002 49698
rect 32510 49646 32562 49698
rect 35534 49646 35586 49698
rect 39006 49646 39058 49698
rect 53790 49646 53842 49698
rect 60622 49646 60674 49698
rect 71262 49646 71314 49698
rect 71710 49646 71762 49698
rect 76190 49646 76242 49698
rect 92430 49646 92482 49698
rect 98030 49646 98082 49698
rect 8990 49534 9042 49586
rect 15262 49534 15314 49586
rect 62078 49534 62130 49586
rect 68910 49534 68962 49586
rect 72718 49534 72770 49586
rect 4396 49366 4448 49418
rect 4520 49366 4572 49418
rect 4644 49366 4696 49418
rect 4768 49366 4820 49418
rect 13396 49366 13448 49418
rect 13520 49366 13572 49418
rect 13644 49366 13696 49418
rect 13768 49366 13820 49418
rect 22396 49366 22448 49418
rect 22520 49366 22572 49418
rect 22644 49366 22696 49418
rect 22768 49366 22820 49418
rect 31396 49366 31448 49418
rect 31520 49366 31572 49418
rect 31644 49366 31696 49418
rect 31768 49366 31820 49418
rect 40396 49366 40448 49418
rect 40520 49366 40572 49418
rect 40644 49366 40696 49418
rect 40768 49366 40820 49418
rect 49396 49366 49448 49418
rect 49520 49366 49572 49418
rect 49644 49366 49696 49418
rect 49768 49366 49820 49418
rect 58396 49366 58448 49418
rect 58520 49366 58572 49418
rect 58644 49366 58696 49418
rect 58768 49366 58820 49418
rect 67396 49366 67448 49418
rect 67520 49366 67572 49418
rect 67644 49366 67696 49418
rect 67768 49366 67820 49418
rect 76396 49366 76448 49418
rect 76520 49366 76572 49418
rect 76644 49366 76696 49418
rect 76768 49366 76820 49418
rect 85396 49366 85448 49418
rect 85520 49366 85572 49418
rect 85644 49366 85696 49418
rect 85768 49366 85820 49418
rect 94396 49366 94448 49418
rect 94520 49366 94572 49418
rect 94644 49366 94696 49418
rect 94768 49366 94820 49418
rect 64766 49198 64818 49250
rect 86158 49198 86210 49250
rect 29262 49086 29314 49138
rect 32958 49086 33010 49138
rect 35086 49086 35138 49138
rect 35758 49086 35810 49138
rect 61294 49086 61346 49138
rect 63646 49086 63698 49138
rect 77646 49086 77698 49138
rect 79774 49086 79826 49138
rect 90526 49086 90578 49138
rect 8990 48974 9042 49026
rect 9326 48974 9378 49026
rect 32286 48974 32338 49026
rect 65102 48974 65154 49026
rect 72158 48974 72210 49026
rect 85150 48974 85202 49026
rect 85822 48974 85874 49026
rect 86718 48974 86770 49026
rect 87054 48974 87106 49026
rect 90190 48974 90242 49026
rect 92542 48974 92594 49026
rect 93102 48974 93154 49026
rect 1710 48862 1762 48914
rect 2382 48862 2434 48914
rect 3166 48862 3218 48914
rect 64206 48862 64258 48914
rect 65326 48862 65378 48914
rect 65886 48862 65938 48914
rect 71822 48862 71874 48914
rect 85038 48862 85090 48914
rect 92318 48862 92370 48914
rect 95454 48862 95506 48914
rect 2046 48750 2098 48802
rect 2718 48750 2770 48802
rect 11678 48750 11730 48802
rect 12462 48750 12514 48802
rect 14478 48750 14530 48802
rect 20750 48750 20802 48802
rect 55022 48750 55074 48802
rect 56366 48750 56418 48802
rect 73502 48750 73554 48802
rect 73950 48750 74002 48802
rect 80222 48750 80274 48802
rect 84702 48750 84754 48802
rect 89630 48750 89682 48802
rect 96238 48750 96290 48802
rect 8896 48582 8948 48634
rect 9020 48582 9072 48634
rect 9144 48582 9196 48634
rect 9268 48582 9320 48634
rect 17896 48582 17948 48634
rect 18020 48582 18072 48634
rect 18144 48582 18196 48634
rect 18268 48582 18320 48634
rect 26896 48582 26948 48634
rect 27020 48582 27072 48634
rect 27144 48582 27196 48634
rect 27268 48582 27320 48634
rect 35896 48582 35948 48634
rect 36020 48582 36072 48634
rect 36144 48582 36196 48634
rect 36268 48582 36320 48634
rect 44896 48582 44948 48634
rect 45020 48582 45072 48634
rect 45144 48582 45196 48634
rect 45268 48582 45320 48634
rect 53896 48582 53948 48634
rect 54020 48582 54072 48634
rect 54144 48582 54196 48634
rect 54268 48582 54320 48634
rect 62896 48582 62948 48634
rect 63020 48582 63072 48634
rect 63144 48582 63196 48634
rect 63268 48582 63320 48634
rect 71896 48582 71948 48634
rect 72020 48582 72072 48634
rect 72144 48582 72196 48634
rect 72268 48582 72320 48634
rect 80896 48582 80948 48634
rect 81020 48582 81072 48634
rect 81144 48582 81196 48634
rect 81268 48582 81320 48634
rect 89896 48582 89948 48634
rect 90020 48582 90072 48634
rect 90144 48582 90196 48634
rect 90268 48582 90320 48634
rect 4734 48414 4786 48466
rect 39902 48414 39954 48466
rect 41022 48414 41074 48466
rect 52334 48414 52386 48466
rect 53230 48414 53282 48466
rect 63870 48414 63922 48466
rect 65326 48414 65378 48466
rect 83134 48414 83186 48466
rect 96574 48414 96626 48466
rect 13582 48302 13634 48354
rect 14254 48302 14306 48354
rect 14926 48302 14978 48354
rect 19854 48302 19906 48354
rect 20414 48302 20466 48354
rect 43486 48302 43538 48354
rect 43934 48302 43986 48354
rect 48974 48302 49026 48354
rect 55694 48302 55746 48354
rect 57374 48302 57426 48354
rect 57822 48302 57874 48354
rect 64542 48302 64594 48354
rect 64878 48302 64930 48354
rect 65102 48302 65154 48354
rect 71038 48302 71090 48354
rect 71374 48302 71426 48354
rect 72942 48302 72994 48354
rect 73502 48302 73554 48354
rect 73950 48302 74002 48354
rect 74174 48302 74226 48354
rect 77198 48302 77250 48354
rect 77646 48302 77698 48354
rect 78318 48302 78370 48354
rect 83694 48302 83746 48354
rect 92542 48302 92594 48354
rect 1822 48190 1874 48242
rect 2158 48190 2210 48242
rect 14030 48190 14082 48242
rect 15038 48190 15090 48242
rect 15822 48190 15874 48242
rect 20302 48190 20354 48242
rect 36766 48190 36818 48242
rect 37326 48190 37378 48242
rect 44270 48190 44322 48242
rect 49198 48190 49250 48242
rect 49870 48190 49922 48242
rect 56030 48190 56082 48242
rect 56702 48190 56754 48242
rect 65550 48190 65602 48242
rect 71710 48190 71762 48242
rect 72382 48190 72434 48242
rect 72718 48190 72770 48242
rect 74398 48190 74450 48242
rect 74622 48190 74674 48242
rect 76414 48190 76466 48242
rect 76974 48190 77026 48242
rect 77422 48190 77474 48242
rect 78094 48190 78146 48242
rect 78878 48190 78930 48242
rect 80222 48190 80274 48242
rect 80558 48190 80610 48242
rect 91198 48190 91250 48242
rect 92318 48190 92370 48242
rect 93102 48190 93154 48242
rect 96238 48190 96290 48242
rect 96910 48190 96962 48242
rect 5630 48078 5682 48130
rect 16494 48078 16546 48130
rect 21086 48078 21138 48130
rect 22094 48078 22146 48130
rect 46398 48078 46450 48130
rect 58382 48078 58434 48130
rect 65214 48078 65266 48130
rect 74286 48078 74338 48130
rect 75966 48078 76018 48130
rect 77310 48078 77362 48130
rect 91646 48078 91698 48130
rect 98030 48078 98082 48130
rect 5294 47966 5346 48018
rect 15486 47966 15538 48018
rect 21422 47966 21474 48018
rect 40462 47966 40514 48018
rect 52894 47966 52946 48018
rect 57038 47966 57090 48018
rect 79214 47966 79266 48018
rect 93438 47966 93490 48018
rect 4396 47798 4448 47850
rect 4520 47798 4572 47850
rect 4644 47798 4696 47850
rect 4768 47798 4820 47850
rect 13396 47798 13448 47850
rect 13520 47798 13572 47850
rect 13644 47798 13696 47850
rect 13768 47798 13820 47850
rect 22396 47798 22448 47850
rect 22520 47798 22572 47850
rect 22644 47798 22696 47850
rect 22768 47798 22820 47850
rect 31396 47798 31448 47850
rect 31520 47798 31572 47850
rect 31644 47798 31696 47850
rect 31768 47798 31820 47850
rect 40396 47798 40448 47850
rect 40520 47798 40572 47850
rect 40644 47798 40696 47850
rect 40768 47798 40820 47850
rect 49396 47798 49448 47850
rect 49520 47798 49572 47850
rect 49644 47798 49696 47850
rect 49768 47798 49820 47850
rect 58396 47798 58448 47850
rect 58520 47798 58572 47850
rect 58644 47798 58696 47850
rect 58768 47798 58820 47850
rect 67396 47798 67448 47850
rect 67520 47798 67572 47850
rect 67644 47798 67696 47850
rect 67768 47798 67820 47850
rect 76396 47798 76448 47850
rect 76520 47798 76572 47850
rect 76644 47798 76696 47850
rect 76768 47798 76820 47850
rect 85396 47798 85448 47850
rect 85520 47798 85572 47850
rect 85644 47798 85696 47850
rect 85768 47798 85820 47850
rect 94396 47798 94448 47850
rect 94520 47798 94572 47850
rect 94644 47798 94696 47850
rect 94768 47798 94820 47850
rect 44942 47630 44994 47682
rect 74622 47630 74674 47682
rect 35758 47518 35810 47570
rect 38670 47518 38722 47570
rect 48750 47518 48802 47570
rect 54462 47518 54514 47570
rect 74958 47518 75010 47570
rect 77422 47518 77474 47570
rect 1822 47406 1874 47458
rect 10446 47406 10498 47458
rect 14142 47406 14194 47458
rect 14702 47406 14754 47458
rect 20526 47406 20578 47458
rect 21198 47406 21250 47458
rect 21758 47406 21810 47458
rect 33966 47406 34018 47458
rect 34638 47406 34690 47458
rect 43262 47406 43314 47458
rect 45278 47406 45330 47458
rect 45950 47406 46002 47458
rect 47406 47406 47458 47458
rect 47742 47406 47794 47458
rect 49198 47406 49250 47458
rect 54910 47406 54962 47458
rect 55358 47406 55410 47458
rect 71038 47406 71090 47458
rect 71486 47406 71538 47458
rect 79214 47406 79266 47458
rect 92654 47406 92706 47458
rect 2046 47294 2098 47346
rect 9662 47294 9714 47346
rect 10222 47294 10274 47346
rect 11342 47294 11394 47346
rect 20750 47294 20802 47346
rect 34750 47294 34802 47346
rect 36430 47294 36482 47346
rect 37326 47294 37378 47346
rect 37662 47294 37714 47346
rect 46062 47294 46114 47346
rect 46958 47294 47010 47346
rect 50542 47294 50594 47346
rect 50878 47294 50930 47346
rect 57598 47294 57650 47346
rect 79550 47294 79602 47346
rect 86718 47294 86770 47346
rect 87054 47294 87106 47346
rect 92878 47294 92930 47346
rect 2606 47182 2658 47234
rect 9102 47182 9154 47234
rect 10782 47182 10834 47234
rect 11790 47182 11842 47234
rect 17278 47182 17330 47234
rect 17838 47182 17890 47234
rect 18174 47182 18226 47234
rect 24110 47182 24162 47234
rect 24894 47182 24946 47234
rect 31166 47182 31218 47234
rect 33630 47182 33682 47234
rect 35310 47182 35362 47234
rect 43710 47182 43762 47234
rect 44270 47182 44322 47234
rect 47966 47182 48018 47234
rect 48190 47182 48242 47234
rect 58382 47182 58434 47234
rect 60734 47182 60786 47234
rect 74062 47182 74114 47234
rect 86382 47182 86434 47234
rect 8896 47014 8948 47066
rect 9020 47014 9072 47066
rect 9144 47014 9196 47066
rect 9268 47014 9320 47066
rect 17896 47014 17948 47066
rect 18020 47014 18072 47066
rect 18144 47014 18196 47066
rect 18268 47014 18320 47066
rect 26896 47014 26948 47066
rect 27020 47014 27072 47066
rect 27144 47014 27196 47066
rect 27268 47014 27320 47066
rect 35896 47014 35948 47066
rect 36020 47014 36072 47066
rect 36144 47014 36196 47066
rect 36268 47014 36320 47066
rect 44896 47014 44948 47066
rect 45020 47014 45072 47066
rect 45144 47014 45196 47066
rect 45268 47014 45320 47066
rect 53896 47014 53948 47066
rect 54020 47014 54072 47066
rect 54144 47014 54196 47066
rect 54268 47014 54320 47066
rect 62896 47014 62948 47066
rect 63020 47014 63072 47066
rect 63144 47014 63196 47066
rect 63268 47014 63320 47066
rect 71896 47014 71948 47066
rect 72020 47014 72072 47066
rect 72144 47014 72196 47066
rect 72268 47014 72320 47066
rect 80896 47014 80948 47066
rect 81020 47014 81072 47066
rect 81144 47014 81196 47066
rect 81268 47014 81320 47066
rect 89896 47014 89948 47066
rect 90020 47014 90072 47066
rect 90144 47014 90196 47066
rect 90268 47014 90320 47066
rect 5406 46846 5458 46898
rect 20974 46846 21026 46898
rect 28590 46846 28642 46898
rect 31614 46846 31666 46898
rect 38558 46846 38610 46898
rect 39118 46846 39170 46898
rect 43038 46846 43090 46898
rect 46958 46846 47010 46898
rect 51438 46846 51490 46898
rect 51886 46846 51938 46898
rect 85038 46846 85090 46898
rect 87278 46846 87330 46898
rect 96574 46846 96626 46898
rect 8654 46734 8706 46786
rect 8990 46734 9042 46786
rect 12350 46734 12402 46786
rect 30382 46734 30434 46786
rect 32174 46734 32226 46786
rect 32510 46734 32562 46786
rect 36766 46734 36818 46786
rect 37886 46734 37938 46786
rect 40014 46734 40066 46786
rect 46174 46734 46226 46786
rect 52446 46734 52498 46786
rect 53006 46734 53058 46786
rect 53566 46734 53618 46786
rect 57262 46734 57314 46786
rect 58382 46734 58434 46786
rect 61854 46734 61906 46786
rect 64990 46734 65042 46786
rect 65438 46734 65490 46786
rect 67566 46734 67618 46786
rect 73726 46734 73778 46786
rect 75294 46734 75346 46786
rect 76862 46734 76914 46786
rect 78430 46734 78482 46786
rect 86382 46734 86434 46786
rect 86718 46734 86770 46786
rect 92206 46734 92258 46786
rect 92542 46734 92594 46786
rect 1822 46622 1874 46674
rect 2494 46622 2546 46674
rect 2830 46622 2882 46674
rect 9550 46622 9602 46674
rect 9998 46622 10050 46674
rect 25678 46622 25730 46674
rect 26126 46622 26178 46674
rect 30606 46622 30658 46674
rect 33294 46622 33346 46674
rect 34750 46622 34802 46674
rect 34974 46622 35026 46674
rect 35646 46622 35698 46674
rect 38222 46622 38274 46674
rect 40238 46622 40290 46674
rect 43486 46622 43538 46674
rect 43934 46622 43986 46674
rect 55246 46622 55298 46674
rect 56590 46622 56642 46674
rect 58494 46622 58546 46674
rect 60062 46622 60114 46674
rect 60398 46622 60450 46674
rect 62190 46622 62242 46674
rect 65214 46622 65266 46674
rect 65774 46622 65826 46674
rect 66446 46622 66498 46674
rect 73950 46622 74002 46674
rect 74510 46622 74562 46674
rect 74958 46622 75010 46674
rect 77086 46622 77138 46674
rect 77646 46622 77698 46674
rect 78094 46622 78146 46674
rect 91870 46622 91922 46674
rect 96238 46622 96290 46674
rect 96910 46622 96962 46674
rect 29150 46510 29202 46562
rect 29822 46510 29874 46562
rect 31166 46510 31218 46562
rect 41022 46510 41074 46562
rect 54238 46510 54290 46562
rect 54686 46510 54738 46562
rect 55582 46510 55634 46562
rect 56030 46510 56082 46562
rect 58270 46510 58322 46562
rect 73390 46510 73442 46562
rect 76638 46510 76690 46562
rect 85486 46510 85538 46562
rect 98030 46510 98082 46562
rect 5966 46398 6018 46450
rect 13134 46398 13186 46450
rect 29486 46398 29538 46450
rect 39454 46398 39506 46450
rect 52222 46398 52274 46450
rect 54238 46398 54290 46450
rect 54686 46398 54738 46450
rect 55358 46398 55410 46450
rect 66782 46398 66834 46450
rect 86942 46398 86994 46450
rect 4396 46230 4448 46282
rect 4520 46230 4572 46282
rect 4644 46230 4696 46282
rect 4768 46230 4820 46282
rect 13396 46230 13448 46282
rect 13520 46230 13572 46282
rect 13644 46230 13696 46282
rect 13768 46230 13820 46282
rect 22396 46230 22448 46282
rect 22520 46230 22572 46282
rect 22644 46230 22696 46282
rect 22768 46230 22820 46282
rect 31396 46230 31448 46282
rect 31520 46230 31572 46282
rect 31644 46230 31696 46282
rect 31768 46230 31820 46282
rect 40396 46230 40448 46282
rect 40520 46230 40572 46282
rect 40644 46230 40696 46282
rect 40768 46230 40820 46282
rect 49396 46230 49448 46282
rect 49520 46230 49572 46282
rect 49644 46230 49696 46282
rect 49768 46230 49820 46282
rect 58396 46230 58448 46282
rect 58520 46230 58572 46282
rect 58644 46230 58696 46282
rect 58768 46230 58820 46282
rect 67396 46230 67448 46282
rect 67520 46230 67572 46282
rect 67644 46230 67696 46282
rect 67768 46230 67820 46282
rect 76396 46230 76448 46282
rect 76520 46230 76572 46282
rect 76644 46230 76696 46282
rect 76768 46230 76820 46282
rect 85396 46230 85448 46282
rect 85520 46230 85572 46282
rect 85644 46230 85696 46282
rect 85768 46230 85820 46282
rect 94396 46230 94448 46282
rect 94520 46230 94572 46282
rect 94644 46230 94696 46282
rect 94768 46230 94820 46282
rect 34526 46062 34578 46114
rect 73054 46062 73106 46114
rect 89630 46062 89682 46114
rect 14926 45950 14978 46002
rect 50318 45950 50370 46002
rect 54126 45950 54178 46002
rect 77982 45950 78034 46002
rect 79102 45950 79154 46002
rect 89966 45950 90018 46002
rect 27246 45838 27298 45890
rect 30942 45838 30994 45890
rect 31502 45838 31554 45890
rect 40686 45838 40738 45890
rect 47518 45838 47570 45890
rect 49198 45838 49250 45890
rect 55022 45838 55074 45890
rect 57710 45838 57762 45890
rect 58494 45838 58546 45890
rect 59950 45838 60002 45890
rect 60622 45838 60674 45890
rect 61070 45838 61122 45890
rect 64878 45838 64930 45890
rect 68238 45838 68290 45890
rect 68798 45838 68850 45890
rect 72718 45838 72770 45890
rect 72942 45838 72994 45890
rect 77086 45838 77138 45890
rect 77310 45838 77362 45890
rect 77646 45838 77698 45890
rect 79886 45838 79938 45890
rect 80446 45838 80498 45890
rect 86158 45838 86210 45890
rect 86494 45838 86546 45890
rect 91982 45838 92034 45890
rect 92542 45838 92594 45890
rect 1710 45726 1762 45778
rect 25678 45726 25730 45778
rect 26910 45726 26962 45778
rect 29262 45726 29314 45778
rect 30606 45726 30658 45778
rect 33742 45726 33794 45778
rect 38558 45726 38610 45778
rect 40238 45726 40290 45778
rect 48078 45726 48130 45778
rect 49086 45726 49138 45778
rect 55694 45726 55746 45778
rect 56814 45726 56866 45778
rect 64542 45726 64594 45778
rect 79326 45726 79378 45778
rect 82798 45726 82850 45778
rect 2046 45614 2098 45666
rect 2494 45614 2546 45666
rect 3166 45614 3218 45666
rect 21310 45614 21362 45666
rect 39006 45614 39058 45666
rect 39454 45614 39506 45666
rect 39902 45614 39954 45666
rect 54462 45614 54514 45666
rect 56926 45614 56978 45666
rect 63534 45614 63586 45666
rect 64094 45614 64146 45666
rect 64654 45614 64706 45666
rect 65326 45614 65378 45666
rect 67790 45614 67842 45666
rect 71374 45614 71426 45666
rect 71934 45614 71986 45666
rect 73054 45614 73106 45666
rect 77422 45614 77474 45666
rect 79662 45614 79714 45666
rect 83582 45614 83634 45666
rect 89070 45614 89122 45666
rect 91310 45614 91362 45666
rect 95006 45614 95058 45666
rect 95678 45614 95730 45666
rect 8896 45446 8948 45498
rect 9020 45446 9072 45498
rect 9144 45446 9196 45498
rect 9268 45446 9320 45498
rect 17896 45446 17948 45498
rect 18020 45446 18072 45498
rect 18144 45446 18196 45498
rect 18268 45446 18320 45498
rect 26896 45446 26948 45498
rect 27020 45446 27072 45498
rect 27144 45446 27196 45498
rect 27268 45446 27320 45498
rect 35896 45446 35948 45498
rect 36020 45446 36072 45498
rect 36144 45446 36196 45498
rect 36268 45446 36320 45498
rect 44896 45446 44948 45498
rect 45020 45446 45072 45498
rect 45144 45446 45196 45498
rect 45268 45446 45320 45498
rect 53896 45446 53948 45498
rect 54020 45446 54072 45498
rect 54144 45446 54196 45498
rect 54268 45446 54320 45498
rect 62896 45446 62948 45498
rect 63020 45446 63072 45498
rect 63144 45446 63196 45498
rect 63268 45446 63320 45498
rect 71896 45446 71948 45498
rect 72020 45446 72072 45498
rect 72144 45446 72196 45498
rect 72268 45446 72320 45498
rect 80896 45446 80948 45498
rect 81020 45446 81072 45498
rect 81144 45446 81196 45498
rect 81268 45446 81320 45498
rect 89896 45446 89948 45498
rect 90020 45446 90072 45498
rect 90144 45446 90196 45498
rect 90268 45446 90320 45498
rect 5742 45278 5794 45330
rect 20302 45278 20354 45330
rect 41022 45278 41074 45330
rect 44494 45278 44546 45330
rect 47294 45278 47346 45330
rect 54462 45278 54514 45330
rect 62414 45278 62466 45330
rect 64542 45278 64594 45330
rect 68574 45278 68626 45330
rect 78654 45278 78706 45330
rect 81006 45278 81058 45330
rect 91198 45278 91250 45330
rect 92878 45278 92930 45330
rect 2046 45166 2098 45218
rect 14254 45166 14306 45218
rect 14590 45166 14642 45218
rect 15486 45166 15538 45218
rect 19630 45166 19682 45218
rect 23438 45166 23490 45218
rect 37438 45166 37490 45218
rect 42030 45166 42082 45218
rect 43822 45166 43874 45218
rect 47518 45166 47570 45218
rect 50206 45166 50258 45218
rect 56926 45166 56978 45218
rect 61294 45166 61346 45218
rect 63310 45166 63362 45218
rect 71150 45166 71202 45218
rect 76750 45166 76802 45218
rect 77758 45166 77810 45218
rect 90638 45166 90690 45218
rect 91982 45166 92034 45218
rect 1710 45054 1762 45106
rect 3054 45054 3106 45106
rect 3390 45054 3442 45106
rect 14926 45054 14978 45106
rect 15374 45054 15426 45106
rect 16494 45054 16546 45106
rect 20078 45054 20130 45106
rect 20750 45054 20802 45106
rect 21086 45054 21138 45106
rect 37998 45054 38050 45106
rect 41358 45054 41410 45106
rect 42142 45054 42194 45106
rect 47630 45054 47682 45106
rect 48078 45054 48130 45106
rect 56590 45054 56642 45106
rect 62750 45054 62802 45106
rect 63534 45054 63586 45106
rect 68910 45054 68962 45106
rect 70142 45054 70194 45106
rect 70478 45054 70530 45106
rect 71262 45054 71314 45106
rect 77534 45054 77586 45106
rect 78318 45054 78370 45106
rect 91758 45054 91810 45106
rect 92542 45054 92594 45106
rect 2494 44942 2546 44994
rect 17614 44942 17666 44994
rect 40014 44942 40066 44994
rect 42702 44942 42754 44994
rect 51662 44942 51714 44994
rect 55918 44942 55970 44994
rect 61742 44942 61794 44994
rect 69470 44942 69522 44994
rect 73614 44942 73666 44994
rect 76302 44942 76354 44994
rect 6526 44830 6578 44882
rect 16158 44830 16210 44882
rect 24222 44830 24274 44882
rect 4396 44662 4448 44714
rect 4520 44662 4572 44714
rect 4644 44662 4696 44714
rect 4768 44662 4820 44714
rect 13396 44662 13448 44714
rect 13520 44662 13572 44714
rect 13644 44662 13696 44714
rect 13768 44662 13820 44714
rect 22396 44662 22448 44714
rect 22520 44662 22572 44714
rect 22644 44662 22696 44714
rect 22768 44662 22820 44714
rect 31396 44662 31448 44714
rect 31520 44662 31572 44714
rect 31644 44662 31696 44714
rect 31768 44662 31820 44714
rect 40396 44662 40448 44714
rect 40520 44662 40572 44714
rect 40644 44662 40696 44714
rect 40768 44662 40820 44714
rect 49396 44662 49448 44714
rect 49520 44662 49572 44714
rect 49644 44662 49696 44714
rect 49768 44662 49820 44714
rect 58396 44662 58448 44714
rect 58520 44662 58572 44714
rect 58644 44662 58696 44714
rect 58768 44662 58820 44714
rect 67396 44662 67448 44714
rect 67520 44662 67572 44714
rect 67644 44662 67696 44714
rect 67768 44662 67820 44714
rect 76396 44662 76448 44714
rect 76520 44662 76572 44714
rect 76644 44662 76696 44714
rect 76768 44662 76820 44714
rect 85396 44662 85448 44714
rect 85520 44662 85572 44714
rect 85644 44662 85696 44714
rect 85768 44662 85820 44714
rect 94396 44662 94448 44714
rect 94520 44662 94572 44714
rect 94644 44662 94696 44714
rect 94768 44662 94820 44714
rect 41470 44494 41522 44546
rect 45278 44494 45330 44546
rect 46398 44494 46450 44546
rect 46734 44494 46786 44546
rect 54910 44494 54962 44546
rect 56366 44494 56418 44546
rect 64430 44494 64482 44546
rect 74062 44494 74114 44546
rect 77982 44494 78034 44546
rect 22542 44382 22594 44434
rect 31054 44382 31106 44434
rect 35982 44382 36034 44434
rect 41806 44382 41858 44434
rect 49086 44382 49138 44434
rect 54126 44382 54178 44434
rect 63086 44382 63138 44434
rect 8766 44270 8818 44322
rect 9438 44270 9490 44322
rect 9774 44270 9826 44322
rect 10222 44270 10274 44322
rect 11566 44270 11618 44322
rect 14254 44270 14306 44322
rect 14814 44270 14866 44322
rect 21758 44270 21810 44322
rect 22206 44270 22258 44322
rect 34190 44270 34242 44322
rect 34862 44270 34914 44322
rect 37774 44270 37826 44322
rect 38446 44270 38498 44322
rect 45950 44270 46002 44322
rect 48078 44270 48130 44322
rect 51326 44270 51378 44322
rect 55470 44270 55522 44322
rect 56702 44270 56754 44322
rect 58494 44270 58546 44322
rect 69694 44270 69746 44322
rect 73614 44270 73666 44322
rect 73838 44270 73890 44322
rect 74510 44270 74562 44322
rect 75070 44270 75122 44322
rect 77310 44270 77362 44322
rect 96910 44270 96962 44322
rect 10334 44158 10386 44210
rect 14030 44158 14082 44210
rect 21422 44158 21474 44210
rect 34974 44158 35026 44210
rect 44270 44158 44322 44210
rect 44942 44158 44994 44210
rect 46062 44158 46114 44210
rect 47742 44158 47794 44210
rect 48638 44158 48690 44210
rect 49870 44158 49922 44210
rect 51998 44158 52050 44210
rect 54574 44158 54626 44210
rect 55694 44158 55746 44210
rect 56926 44158 56978 44210
rect 57486 44158 57538 44210
rect 64654 44158 64706 44210
rect 65214 44158 65266 44210
rect 74062 44158 74114 44210
rect 77422 44158 77474 44210
rect 78318 44158 78370 44210
rect 79774 44158 79826 44210
rect 95566 44158 95618 44210
rect 95902 44158 95954 44210
rect 96238 44158 96290 44210
rect 96574 44158 96626 44210
rect 98030 44158 98082 44210
rect 1822 44046 1874 44098
rect 2606 44046 2658 44098
rect 8318 44046 8370 44098
rect 8990 44046 9042 44098
rect 11118 44046 11170 44098
rect 17390 44046 17442 44098
rect 17950 44046 18002 44098
rect 20750 44046 20802 44098
rect 23102 44046 23154 44098
rect 33854 44046 33906 44098
rect 35534 44046 35586 44098
rect 40910 44046 40962 44098
rect 43934 44046 43986 44098
rect 46734 44046 46786 44098
rect 51662 44046 51714 44098
rect 52894 44046 52946 44098
rect 57934 44046 57986 44098
rect 63534 44046 63586 44098
rect 64094 44046 64146 44098
rect 73054 44046 73106 44098
rect 76638 44046 76690 44098
rect 80110 44046 80162 44098
rect 81118 44046 81170 44098
rect 8896 43878 8948 43930
rect 9020 43878 9072 43930
rect 9144 43878 9196 43930
rect 9268 43878 9320 43930
rect 17896 43878 17948 43930
rect 18020 43878 18072 43930
rect 18144 43878 18196 43930
rect 18268 43878 18320 43930
rect 26896 43878 26948 43930
rect 27020 43878 27072 43930
rect 27144 43878 27196 43930
rect 27268 43878 27320 43930
rect 35896 43878 35948 43930
rect 36020 43878 36072 43930
rect 36144 43878 36196 43930
rect 36268 43878 36320 43930
rect 44896 43878 44948 43930
rect 45020 43878 45072 43930
rect 45144 43878 45196 43930
rect 45268 43878 45320 43930
rect 53896 43878 53948 43930
rect 54020 43878 54072 43930
rect 54144 43878 54196 43930
rect 54268 43878 54320 43930
rect 62896 43878 62948 43930
rect 63020 43878 63072 43930
rect 63144 43878 63196 43930
rect 63268 43878 63320 43930
rect 71896 43878 71948 43930
rect 72020 43878 72072 43930
rect 72144 43878 72196 43930
rect 72268 43878 72320 43930
rect 80896 43878 80948 43930
rect 81020 43878 81072 43930
rect 81144 43878 81196 43930
rect 81268 43878 81320 43930
rect 89896 43878 89948 43930
rect 90020 43878 90072 43930
rect 90144 43878 90196 43930
rect 90268 43878 90320 43930
rect 5406 43710 5458 43762
rect 28590 43710 28642 43762
rect 38670 43710 38722 43762
rect 55582 43710 55634 43762
rect 60174 43710 60226 43762
rect 71262 43710 71314 43762
rect 75406 43710 75458 43762
rect 77086 43710 77138 43762
rect 2046 43598 2098 43650
rect 6750 43598 6802 43650
rect 7198 43598 7250 43650
rect 12350 43598 12402 43650
rect 13918 43598 13970 43650
rect 25342 43598 25394 43650
rect 30494 43598 30546 43650
rect 31726 43598 31778 43650
rect 33070 43598 33122 43650
rect 33406 43598 33458 43650
rect 37998 43598 38050 43650
rect 39678 43598 39730 43650
rect 43262 43598 43314 43650
rect 46398 43598 46450 43650
rect 47182 43598 47234 43650
rect 52782 43598 52834 43650
rect 53566 43598 53618 43650
rect 53902 43598 53954 43650
rect 56030 43598 56082 43650
rect 59390 43598 59442 43650
rect 62414 43598 62466 43650
rect 63086 43598 63138 43650
rect 63422 43598 63474 43650
rect 65998 43598 66050 43650
rect 69918 43598 69970 43650
rect 70366 43598 70418 43650
rect 71710 43598 71762 43650
rect 73502 43598 73554 43650
rect 76974 43598 77026 43650
rect 83694 43598 83746 43650
rect 84478 43598 84530 43650
rect 86606 43598 86658 43650
rect 91422 43598 91474 43650
rect 94558 43598 94610 43650
rect 1822 43486 1874 43538
rect 2494 43486 2546 43538
rect 2942 43486 2994 43538
rect 9438 43486 9490 43538
rect 10110 43486 10162 43538
rect 25566 43486 25618 43538
rect 26238 43486 26290 43538
rect 29262 43486 29314 43538
rect 29934 43486 29986 43538
rect 30606 43486 30658 43538
rect 34750 43486 34802 43538
rect 35198 43486 35250 43538
rect 35646 43486 35698 43538
rect 35870 43486 35922 43538
rect 38446 43486 38498 43538
rect 43598 43486 43650 43538
rect 44046 43486 44098 43538
rect 50094 43486 50146 43538
rect 50542 43486 50594 43538
rect 56702 43486 56754 43538
rect 57150 43486 57202 43538
rect 65438 43486 65490 43538
rect 65774 43486 65826 43538
rect 66334 43486 66386 43538
rect 67006 43486 67058 43538
rect 70702 43486 70754 43538
rect 72382 43486 72434 43538
rect 73166 43486 73218 43538
rect 75742 43486 75794 43538
rect 76638 43486 76690 43538
rect 77198 43486 77250 43538
rect 80782 43486 80834 43538
rect 81342 43486 81394 43538
rect 91646 43486 91698 43538
rect 92206 43486 92258 43538
rect 6302 43374 6354 43426
rect 31278 43374 31330 43426
rect 32510 43374 32562 43426
rect 39230 43374 39282 43426
rect 64542 43374 64594 43426
rect 64990 43374 65042 43426
rect 72718 43374 72770 43426
rect 74958 43374 75010 43426
rect 80558 43374 80610 43426
rect 90974 43374 91026 43426
rect 5966 43262 6018 43314
rect 13134 43262 13186 43314
rect 29598 43262 29650 43314
rect 66446 43262 66498 43314
rect 74958 43262 75010 43314
rect 75294 43262 75346 43314
rect 95342 43262 95394 43314
rect 4396 43094 4448 43146
rect 4520 43094 4572 43146
rect 4644 43094 4696 43146
rect 4768 43094 4820 43146
rect 13396 43094 13448 43146
rect 13520 43094 13572 43146
rect 13644 43094 13696 43146
rect 13768 43094 13820 43146
rect 22396 43094 22448 43146
rect 22520 43094 22572 43146
rect 22644 43094 22696 43146
rect 22768 43094 22820 43146
rect 31396 43094 31448 43146
rect 31520 43094 31572 43146
rect 31644 43094 31696 43146
rect 31768 43094 31820 43146
rect 40396 43094 40448 43146
rect 40520 43094 40572 43146
rect 40644 43094 40696 43146
rect 40768 43094 40820 43146
rect 49396 43094 49448 43146
rect 49520 43094 49572 43146
rect 49644 43094 49696 43146
rect 49768 43094 49820 43146
rect 58396 43094 58448 43146
rect 58520 43094 58572 43146
rect 58644 43094 58696 43146
rect 58768 43094 58820 43146
rect 67396 43094 67448 43146
rect 67520 43094 67572 43146
rect 67644 43094 67696 43146
rect 67768 43094 67820 43146
rect 76396 43094 76448 43146
rect 76520 43094 76572 43146
rect 76644 43094 76696 43146
rect 76768 43094 76820 43146
rect 85396 43094 85448 43146
rect 85520 43094 85572 43146
rect 85644 43094 85696 43146
rect 85768 43094 85820 43146
rect 94396 43094 94448 43146
rect 94520 43094 94572 43146
rect 94644 43094 94696 43146
rect 94768 43094 94820 43146
rect 35086 42926 35138 42978
rect 65774 42926 65826 42978
rect 73278 42926 73330 42978
rect 92766 42926 92818 42978
rect 29374 42814 29426 42866
rect 31166 42814 31218 42866
rect 61854 42814 61906 42866
rect 12686 42702 12738 42754
rect 13806 42702 13858 42754
rect 14366 42702 14418 42754
rect 18958 42702 19010 42754
rect 19518 42702 19570 42754
rect 20190 42702 20242 42754
rect 27246 42702 27298 42754
rect 31614 42702 31666 42754
rect 32062 42702 32114 42754
rect 62302 42702 62354 42754
rect 62750 42702 62802 42754
rect 69806 42702 69858 42754
rect 70254 42702 70306 42754
rect 86606 42702 86658 42754
rect 86942 42702 86994 42754
rect 90414 42702 90466 42754
rect 92318 42702 92370 42754
rect 96910 42702 96962 42754
rect 1710 42590 1762 42642
rect 13582 42590 13634 42642
rect 14702 42590 14754 42642
rect 19406 42590 19458 42642
rect 26910 42590 26962 42642
rect 34302 42590 34354 42642
rect 77758 42590 77810 42642
rect 91982 42590 92034 42642
rect 96238 42590 96290 42642
rect 96574 42590 96626 42642
rect 98030 42590 98082 42642
rect 2046 42478 2098 42530
rect 2494 42478 2546 42530
rect 2942 42478 2994 42530
rect 12238 42478 12290 42530
rect 12910 42478 12962 42530
rect 15262 42478 15314 42530
rect 20526 42478 20578 42530
rect 21310 42478 21362 42530
rect 21870 42478 21922 42530
rect 64990 42478 65042 42530
rect 69358 42478 69410 42530
rect 72494 42478 72546 42530
rect 75406 42478 75458 42530
rect 78094 42478 78146 42530
rect 89518 42478 89570 42530
rect 90078 42478 90130 42530
rect 90862 42478 90914 42530
rect 91422 42478 91474 42530
rect 93102 42478 93154 42530
rect 8896 42310 8948 42362
rect 9020 42310 9072 42362
rect 9144 42310 9196 42362
rect 9268 42310 9320 42362
rect 17896 42310 17948 42362
rect 18020 42310 18072 42362
rect 18144 42310 18196 42362
rect 18268 42310 18320 42362
rect 26896 42310 26948 42362
rect 27020 42310 27072 42362
rect 27144 42310 27196 42362
rect 27268 42310 27320 42362
rect 35896 42310 35948 42362
rect 36020 42310 36072 42362
rect 36144 42310 36196 42362
rect 36268 42310 36320 42362
rect 44896 42310 44948 42362
rect 45020 42310 45072 42362
rect 45144 42310 45196 42362
rect 45268 42310 45320 42362
rect 53896 42310 53948 42362
rect 54020 42310 54072 42362
rect 54144 42310 54196 42362
rect 54268 42310 54320 42362
rect 62896 42310 62948 42362
rect 63020 42310 63072 42362
rect 63144 42310 63196 42362
rect 63268 42310 63320 42362
rect 71896 42310 71948 42362
rect 72020 42310 72072 42362
rect 72144 42310 72196 42362
rect 72268 42310 72320 42362
rect 80896 42310 80948 42362
rect 81020 42310 81072 42362
rect 81144 42310 81196 42362
rect 81268 42310 81320 42362
rect 89896 42310 89948 42362
rect 90020 42310 90072 42362
rect 90144 42310 90196 42362
rect 90268 42310 90320 42362
rect 5742 42142 5794 42194
rect 16382 42142 16434 42194
rect 77534 42142 77586 42194
rect 86830 42142 86882 42194
rect 91982 42142 92034 42194
rect 20414 42030 20466 42082
rect 23550 42030 23602 42082
rect 24446 42030 24498 42082
rect 38558 42030 38610 42082
rect 39230 42030 39282 42082
rect 44046 42030 44098 42082
rect 49646 42030 49698 42082
rect 57598 42030 57650 42082
rect 58382 42030 58434 42082
rect 78206 42030 78258 42082
rect 78654 42030 78706 42082
rect 79102 42030 79154 42082
rect 88174 42030 88226 42082
rect 2830 41918 2882 41970
rect 3166 41918 3218 41970
rect 13246 41918 13298 41970
rect 13806 41918 13858 41970
rect 17502 41918 17554 41970
rect 19742 41918 19794 41970
rect 20190 41918 20242 41970
rect 20638 41918 20690 41970
rect 21198 41918 21250 41970
rect 39566 41918 39618 41970
rect 44494 41918 44546 41970
rect 54238 41918 54290 41970
rect 55582 41918 55634 41970
rect 57486 41918 57538 41970
rect 67790 41918 67842 41970
rect 76862 41918 76914 41970
rect 87166 41918 87218 41970
rect 88398 41918 88450 41970
rect 88846 41918 88898 41970
rect 89182 41918 89234 41970
rect 92318 41918 92370 41970
rect 2158 41806 2210 41858
rect 6638 41806 6690 41858
rect 50318 41806 50370 41858
rect 53342 41806 53394 41858
rect 53790 41806 53842 41858
rect 54686 41806 54738 41858
rect 56030 41806 56082 41858
rect 75966 41806 76018 41858
rect 76414 41806 76466 41858
rect 77870 41806 77922 41858
rect 6302 41694 6354 41746
rect 16942 41694 16994 41746
rect 56702 41694 56754 41746
rect 57038 41694 57090 41746
rect 4396 41526 4448 41578
rect 4520 41526 4572 41578
rect 4644 41526 4696 41578
rect 4768 41526 4820 41578
rect 13396 41526 13448 41578
rect 13520 41526 13572 41578
rect 13644 41526 13696 41578
rect 13768 41526 13820 41578
rect 22396 41526 22448 41578
rect 22520 41526 22572 41578
rect 22644 41526 22696 41578
rect 22768 41526 22820 41578
rect 31396 41526 31448 41578
rect 31520 41526 31572 41578
rect 31644 41526 31696 41578
rect 31768 41526 31820 41578
rect 40396 41526 40448 41578
rect 40520 41526 40572 41578
rect 40644 41526 40696 41578
rect 40768 41526 40820 41578
rect 49396 41526 49448 41578
rect 49520 41526 49572 41578
rect 49644 41526 49696 41578
rect 49768 41526 49820 41578
rect 58396 41526 58448 41578
rect 58520 41526 58572 41578
rect 58644 41526 58696 41578
rect 58768 41526 58820 41578
rect 67396 41526 67448 41578
rect 67520 41526 67572 41578
rect 67644 41526 67696 41578
rect 67768 41526 67820 41578
rect 76396 41526 76448 41578
rect 76520 41526 76572 41578
rect 76644 41526 76696 41578
rect 76768 41526 76820 41578
rect 85396 41526 85448 41578
rect 85520 41526 85572 41578
rect 85644 41526 85696 41578
rect 85768 41526 85820 41578
rect 94396 41526 94448 41578
rect 94520 41526 94572 41578
rect 94644 41526 94696 41578
rect 94768 41526 94820 41578
rect 53230 41358 53282 41410
rect 81566 41358 81618 41410
rect 33742 41246 33794 41298
rect 42366 41246 42418 41298
rect 76862 41246 76914 41298
rect 87614 41246 87666 41298
rect 34526 41134 34578 41186
rect 35310 41134 35362 41186
rect 35870 41134 35922 41186
rect 38558 41134 38610 41186
rect 39006 41134 39058 41186
rect 44046 41134 44098 41186
rect 44718 41134 44770 41186
rect 45278 41134 45330 41186
rect 48862 41134 48914 41186
rect 49534 41134 49586 41186
rect 54574 41134 54626 41186
rect 55694 41134 55746 41186
rect 56142 41134 56194 41186
rect 57038 41134 57090 41186
rect 58942 41134 58994 41186
rect 63982 41134 64034 41186
rect 64654 41134 64706 41186
rect 71038 41134 71090 41186
rect 71598 41134 71650 41186
rect 75070 41134 75122 41186
rect 76750 41134 76802 41186
rect 77982 41134 78034 41186
rect 78430 41134 78482 41186
rect 96910 41134 96962 41186
rect 1710 41022 1762 41074
rect 2382 41022 2434 41074
rect 8878 41022 8930 41074
rect 19070 41022 19122 41074
rect 35198 41022 35250 41074
rect 42030 41022 42082 41074
rect 44270 41022 44322 41074
rect 47630 41022 47682 41074
rect 48750 41022 48802 41074
rect 50990 41022 51042 41074
rect 52670 41022 52722 41074
rect 57822 41022 57874 41074
rect 63758 41022 63810 41074
rect 70814 41022 70866 41074
rect 74734 41022 74786 41074
rect 76302 41022 76354 41074
rect 76526 41022 76578 41074
rect 76862 41022 76914 41074
rect 96238 41022 96290 41074
rect 96574 41022 96626 41074
rect 98030 41022 98082 41074
rect 2046 40910 2098 40962
rect 2718 40910 2770 40962
rect 3166 40910 3218 40962
rect 5742 40910 5794 40962
rect 9326 40910 9378 40962
rect 25454 40910 25506 40962
rect 31502 40910 31554 40962
rect 33294 40910 33346 40962
rect 34190 40910 34242 40962
rect 41470 40910 41522 40962
rect 48414 40910 48466 40962
rect 48974 40910 49026 40962
rect 49982 40910 50034 40962
rect 50654 40910 50706 40962
rect 52222 40910 52274 40962
rect 59278 40910 59330 40962
rect 67006 40910 67058 40962
rect 67678 40910 67730 40962
rect 68574 40910 68626 40962
rect 74062 40910 74114 40962
rect 75630 40910 75682 40962
rect 77646 40910 77698 40962
rect 80894 40910 80946 40962
rect 82574 40910 82626 40962
rect 84590 40910 84642 40962
rect 8896 40742 8948 40794
rect 9020 40742 9072 40794
rect 9144 40742 9196 40794
rect 9268 40742 9320 40794
rect 17896 40742 17948 40794
rect 18020 40742 18072 40794
rect 18144 40742 18196 40794
rect 18268 40742 18320 40794
rect 26896 40742 26948 40794
rect 27020 40742 27072 40794
rect 27144 40742 27196 40794
rect 27268 40742 27320 40794
rect 35896 40742 35948 40794
rect 36020 40742 36072 40794
rect 36144 40742 36196 40794
rect 36268 40742 36320 40794
rect 44896 40742 44948 40794
rect 45020 40742 45072 40794
rect 45144 40742 45196 40794
rect 45268 40742 45320 40794
rect 53896 40742 53948 40794
rect 54020 40742 54072 40794
rect 54144 40742 54196 40794
rect 54268 40742 54320 40794
rect 62896 40742 62948 40794
rect 63020 40742 63072 40794
rect 63144 40742 63196 40794
rect 63268 40742 63320 40794
rect 71896 40742 71948 40794
rect 72020 40742 72072 40794
rect 72144 40742 72196 40794
rect 72268 40742 72320 40794
rect 80896 40742 80948 40794
rect 81020 40742 81072 40794
rect 81144 40742 81196 40794
rect 81268 40742 81320 40794
rect 89896 40742 89948 40794
rect 90020 40742 90072 40794
rect 90144 40742 90196 40794
rect 90268 40742 90320 40794
rect 4734 40574 4786 40626
rect 8318 40574 8370 40626
rect 12350 40574 12402 40626
rect 21982 40574 22034 40626
rect 22654 40574 22706 40626
rect 22990 40574 23042 40626
rect 28254 40574 28306 40626
rect 31390 40574 31442 40626
rect 39006 40574 39058 40626
rect 39902 40574 39954 40626
rect 41022 40574 41074 40626
rect 44830 40574 44882 40626
rect 46510 40574 46562 40626
rect 48862 40574 48914 40626
rect 52558 40574 52610 40626
rect 53678 40574 53730 40626
rect 55358 40574 55410 40626
rect 57822 40574 57874 40626
rect 60958 40574 61010 40626
rect 61742 40574 61794 40626
rect 65214 40574 65266 40626
rect 65998 40574 66050 40626
rect 72270 40574 72322 40626
rect 76302 40574 76354 40626
rect 85374 40574 85426 40626
rect 85934 40574 85986 40626
rect 90750 40574 90802 40626
rect 91422 40574 91474 40626
rect 94782 40574 94834 40626
rect 96574 40574 96626 40626
rect 16830 40462 16882 40514
rect 17614 40462 17666 40514
rect 30382 40462 30434 40514
rect 30942 40462 30994 40514
rect 33070 40462 33122 40514
rect 33406 40462 33458 40514
rect 37998 40462 38050 40514
rect 41582 40462 41634 40514
rect 42030 40462 42082 40514
rect 42702 40462 42754 40514
rect 45950 40462 46002 40514
rect 54574 40462 54626 40514
rect 57038 40462 57090 40514
rect 57374 40462 57426 40514
rect 67118 40462 67170 40514
rect 67454 40462 67506 40514
rect 68126 40462 68178 40514
rect 74174 40462 74226 40514
rect 76526 40462 76578 40514
rect 86270 40462 86322 40514
rect 1822 40350 1874 40402
rect 2158 40350 2210 40402
rect 5630 40350 5682 40402
rect 5966 40350 6018 40402
rect 9550 40350 9602 40402
rect 10110 40350 10162 40402
rect 13582 40350 13634 40402
rect 17502 40350 17554 40402
rect 18622 40350 18674 40402
rect 19182 40350 19234 40402
rect 19518 40350 19570 40402
rect 25454 40350 25506 40402
rect 25902 40350 25954 40402
rect 28926 40350 28978 40402
rect 29598 40350 29650 40402
rect 30158 40350 30210 40402
rect 34974 40350 35026 40402
rect 35422 40350 35474 40402
rect 35758 40350 35810 40402
rect 36094 40350 36146 40402
rect 38670 40350 38722 40402
rect 39454 40350 39506 40402
rect 45838 40350 45890 40402
rect 49422 40350 49474 40402
rect 50094 40350 50146 40402
rect 53118 40350 53170 40402
rect 54798 40350 54850 40402
rect 58158 40350 58210 40402
rect 58606 40350 58658 40402
rect 65550 40350 65602 40402
rect 66558 40350 66610 40402
rect 68238 40350 68290 40402
rect 68910 40350 68962 40402
rect 69358 40350 69410 40402
rect 71710 40350 71762 40402
rect 72606 40350 72658 40402
rect 73166 40350 73218 40402
rect 73950 40350 74002 40402
rect 76638 40350 76690 40402
rect 77422 40350 77474 40402
rect 77758 40350 77810 40402
rect 82462 40350 82514 40402
rect 82798 40350 82850 40402
rect 91198 40350 91250 40402
rect 91870 40350 91922 40402
rect 92206 40350 92258 40402
rect 95342 40350 95394 40402
rect 96238 40350 96290 40402
rect 18286 40238 18338 40290
rect 40350 40238 40402 40290
rect 44382 40238 44434 40290
rect 45166 40238 45218 40290
rect 54014 40238 54066 40290
rect 73502 40238 73554 40290
rect 78094 40238 78146 40290
rect 5294 40126 5346 40178
rect 9102 40126 9154 40178
rect 13134 40126 13186 40178
rect 29262 40126 29314 40178
rect 41358 40126 41410 40178
rect 66894 40126 66946 40178
rect 69694 40126 69746 40178
rect 4396 39958 4448 40010
rect 4520 39958 4572 40010
rect 4644 39958 4696 40010
rect 4768 39958 4820 40010
rect 13396 39958 13448 40010
rect 13520 39958 13572 40010
rect 13644 39958 13696 40010
rect 13768 39958 13820 40010
rect 22396 39958 22448 40010
rect 22520 39958 22572 40010
rect 22644 39958 22696 40010
rect 22768 39958 22820 40010
rect 31396 39958 31448 40010
rect 31520 39958 31572 40010
rect 31644 39958 31696 40010
rect 31768 39958 31820 40010
rect 40396 39958 40448 40010
rect 40520 39958 40572 40010
rect 40644 39958 40696 40010
rect 40768 39958 40820 40010
rect 49396 39958 49448 40010
rect 49520 39958 49572 40010
rect 49644 39958 49696 40010
rect 49768 39958 49820 40010
rect 58396 39958 58448 40010
rect 58520 39958 58572 40010
rect 58644 39958 58696 40010
rect 58768 39958 58820 40010
rect 67396 39958 67448 40010
rect 67520 39958 67572 40010
rect 67644 39958 67696 40010
rect 67768 39958 67820 40010
rect 76396 39958 76448 40010
rect 76520 39958 76572 40010
rect 76644 39958 76696 40010
rect 76768 39958 76820 40010
rect 85396 39958 85448 40010
rect 85520 39958 85572 40010
rect 85644 39958 85696 40010
rect 85768 39958 85820 40010
rect 94396 39958 94448 40010
rect 94520 39958 94572 40010
rect 94644 39958 94696 40010
rect 94768 39958 94820 40010
rect 12462 39790 12514 39842
rect 34862 39790 34914 39842
rect 9214 39678 9266 39730
rect 29262 39678 29314 39730
rect 30942 39678 30994 39730
rect 37662 39678 37714 39730
rect 48414 39678 48466 39730
rect 53230 39678 53282 39730
rect 53678 39678 53730 39730
rect 67230 39678 67282 39730
rect 67678 39678 67730 39730
rect 69022 39678 69074 39730
rect 82126 39678 82178 39730
rect 82574 39678 82626 39730
rect 90638 39678 90690 39730
rect 1822 39566 1874 39618
rect 11678 39566 11730 39618
rect 18398 39566 18450 39618
rect 26798 39566 26850 39618
rect 31166 39566 31218 39618
rect 31838 39566 31890 39618
rect 36542 39566 36594 39618
rect 37326 39566 37378 39618
rect 68350 39566 68402 39618
rect 68686 39566 68738 39618
rect 82462 39566 82514 39618
rect 83022 39566 83074 39618
rect 83918 39566 83970 39618
rect 84926 39566 84978 39618
rect 85038 39566 85090 39618
rect 85374 39566 85426 39618
rect 85598 39566 85650 39618
rect 86606 39566 86658 39618
rect 87166 39566 87218 39618
rect 96910 39566 96962 39618
rect 2382 39454 2434 39506
rect 5630 39454 5682 39506
rect 11902 39454 11954 39506
rect 12798 39454 12850 39506
rect 13470 39454 13522 39506
rect 19294 39454 19346 39506
rect 26574 39454 26626 39506
rect 36206 39454 36258 39506
rect 36990 39454 37042 39506
rect 37102 39454 37154 39506
rect 68462 39454 68514 39506
rect 84142 39454 84194 39506
rect 84254 39454 84306 39506
rect 84814 39454 84866 39506
rect 85934 39454 85986 39506
rect 86382 39454 86434 39506
rect 92094 39454 92146 39506
rect 98030 39454 98082 39506
rect 2046 39342 2098 39394
rect 11230 39342 11282 39394
rect 13806 39342 13858 39394
rect 14142 39342 14194 39394
rect 18622 39342 18674 39394
rect 34302 39342 34354 39394
rect 35870 39342 35922 39394
rect 36318 39342 36370 39394
rect 66110 39342 66162 39394
rect 72718 39342 72770 39394
rect 82686 39342 82738 39394
rect 83470 39342 83522 39394
rect 85822 39342 85874 39394
rect 89518 39342 89570 39394
rect 90302 39342 90354 39394
rect 8896 39174 8948 39226
rect 9020 39174 9072 39226
rect 9144 39174 9196 39226
rect 9268 39174 9320 39226
rect 17896 39174 17948 39226
rect 18020 39174 18072 39226
rect 18144 39174 18196 39226
rect 18268 39174 18320 39226
rect 26896 39174 26948 39226
rect 27020 39174 27072 39226
rect 27144 39174 27196 39226
rect 27268 39174 27320 39226
rect 35896 39174 35948 39226
rect 36020 39174 36072 39226
rect 36144 39174 36196 39226
rect 36268 39174 36320 39226
rect 44896 39174 44948 39226
rect 45020 39174 45072 39226
rect 45144 39174 45196 39226
rect 45268 39174 45320 39226
rect 53896 39174 53948 39226
rect 54020 39174 54072 39226
rect 54144 39174 54196 39226
rect 54268 39174 54320 39226
rect 62896 39174 62948 39226
rect 63020 39174 63072 39226
rect 63144 39174 63196 39226
rect 63268 39174 63320 39226
rect 71896 39174 71948 39226
rect 72020 39174 72072 39226
rect 72144 39174 72196 39226
rect 72268 39174 72320 39226
rect 80896 39174 80948 39226
rect 81020 39174 81072 39226
rect 81144 39174 81196 39226
rect 81268 39174 81320 39226
rect 89896 39174 89948 39226
rect 90020 39174 90072 39226
rect 90144 39174 90196 39226
rect 90268 39174 90320 39226
rect 16270 39006 16322 39058
rect 17502 39006 17554 39058
rect 21086 39006 21138 39058
rect 42142 39006 42194 39058
rect 44494 39006 44546 39058
rect 52894 39006 52946 39058
rect 66670 39006 66722 39058
rect 67118 39006 67170 39058
rect 67902 39006 67954 39058
rect 72494 39006 72546 39058
rect 72942 39006 72994 39058
rect 77310 39006 77362 39058
rect 77870 39006 77922 39058
rect 78542 39006 78594 39058
rect 84366 39006 84418 39058
rect 85262 39006 85314 39058
rect 89742 39006 89794 39058
rect 91982 39006 92034 39058
rect 2382 38894 2434 38946
rect 21646 38894 21698 38946
rect 38558 38894 38610 38946
rect 42590 38894 42642 38946
rect 43822 38894 43874 38946
rect 47742 38894 47794 38946
rect 47966 38894 48018 38946
rect 48078 38894 48130 38946
rect 49310 38894 49362 38946
rect 50542 38894 50594 38946
rect 53230 38894 53282 38946
rect 53902 38894 53954 38946
rect 58382 38894 58434 38946
rect 68014 38894 68066 38946
rect 76414 38894 76466 38946
rect 77534 38894 77586 38946
rect 78990 38894 79042 38946
rect 84702 38894 84754 38946
rect 90190 38894 90242 38946
rect 90974 38894 91026 38946
rect 91310 38894 91362 38946
rect 1822 38782 1874 38834
rect 13358 38782 13410 38834
rect 13806 38782 13858 38834
rect 48302 38782 48354 38834
rect 48750 38782 48802 38834
rect 51886 38782 51938 38834
rect 53566 38782 53618 38834
rect 60174 38782 60226 38834
rect 67790 38782 67842 38834
rect 68350 38782 68402 38834
rect 69022 38782 69074 38834
rect 74846 38782 74898 38834
rect 77198 38782 77250 38834
rect 91646 38782 91698 38834
rect 16830 38670 16882 38722
rect 28814 38670 28866 38722
rect 52446 38670 52498 38722
rect 76862 38670 76914 38722
rect 83694 38670 83746 38722
rect 85710 38670 85762 38722
rect 50094 38558 50146 38610
rect 75294 38558 75346 38610
rect 83694 38558 83746 38610
rect 84142 38558 84194 38610
rect 4396 38390 4448 38442
rect 4520 38390 4572 38442
rect 4644 38390 4696 38442
rect 4768 38390 4820 38442
rect 13396 38390 13448 38442
rect 13520 38390 13572 38442
rect 13644 38390 13696 38442
rect 13768 38390 13820 38442
rect 22396 38390 22448 38442
rect 22520 38390 22572 38442
rect 22644 38390 22696 38442
rect 22768 38390 22820 38442
rect 31396 38390 31448 38442
rect 31520 38390 31572 38442
rect 31644 38390 31696 38442
rect 31768 38390 31820 38442
rect 40396 38390 40448 38442
rect 40520 38390 40572 38442
rect 40644 38390 40696 38442
rect 40768 38390 40820 38442
rect 49396 38390 49448 38442
rect 49520 38390 49572 38442
rect 49644 38390 49696 38442
rect 49768 38390 49820 38442
rect 58396 38390 58448 38442
rect 58520 38390 58572 38442
rect 58644 38390 58696 38442
rect 58768 38390 58820 38442
rect 67396 38390 67448 38442
rect 67520 38390 67572 38442
rect 67644 38390 67696 38442
rect 67768 38390 67820 38442
rect 76396 38390 76448 38442
rect 76520 38390 76572 38442
rect 76644 38390 76696 38442
rect 76768 38390 76820 38442
rect 85396 38390 85448 38442
rect 85520 38390 85572 38442
rect 85644 38390 85696 38442
rect 85768 38390 85820 38442
rect 94396 38390 94448 38442
rect 94520 38390 94572 38442
rect 94644 38390 94696 38442
rect 94768 38390 94820 38442
rect 42030 38222 42082 38274
rect 45278 38222 45330 38274
rect 46398 38222 46450 38274
rect 46734 38222 46786 38274
rect 60958 38222 61010 38274
rect 76078 38222 76130 38274
rect 33406 38110 33458 38162
rect 51550 38110 51602 38162
rect 56702 38110 56754 38162
rect 67678 38110 67730 38162
rect 68798 38110 68850 38162
rect 75406 38110 75458 38162
rect 87166 38110 87218 38162
rect 20526 37998 20578 38050
rect 21534 37998 21586 38050
rect 21870 37998 21922 38050
rect 27694 37998 27746 38050
rect 28366 37998 28418 38050
rect 34302 37998 34354 38050
rect 35086 37998 35138 38050
rect 38558 37998 38610 38050
rect 39006 37998 39058 38050
rect 42366 37998 42418 38050
rect 45950 37998 46002 38050
rect 48190 37998 48242 38050
rect 49758 37998 49810 38050
rect 52670 37998 52722 38050
rect 53230 37998 53282 38050
rect 63310 37998 63362 38050
rect 63982 37998 64034 38050
rect 68574 37998 68626 38050
rect 72494 37998 72546 38050
rect 73166 37998 73218 38050
rect 73502 37998 73554 38050
rect 73950 37998 74002 38050
rect 76190 37998 76242 38050
rect 76974 37998 77026 38050
rect 77422 37998 77474 38050
rect 78318 37998 78370 38050
rect 78878 37998 78930 38050
rect 79326 37998 79378 38050
rect 84926 37998 84978 38050
rect 85150 37998 85202 38050
rect 87502 37998 87554 38050
rect 1710 37886 1762 37938
rect 20750 37886 20802 37938
rect 28478 37886 28530 37938
rect 32958 37886 33010 37938
rect 34862 37886 34914 37938
rect 36990 37886 37042 37938
rect 43374 37886 43426 37938
rect 44270 37886 44322 37938
rect 44942 37886 44994 37938
rect 46062 37886 46114 37938
rect 48974 37886 49026 37938
rect 49982 37886 50034 37938
rect 59278 37886 59330 37938
rect 60622 37886 60674 37938
rect 61182 37886 61234 37938
rect 61742 37886 61794 37938
rect 63086 37886 63138 37938
rect 68350 37886 68402 37938
rect 74286 37886 74338 37938
rect 76302 37886 76354 37938
rect 78542 37886 78594 37938
rect 81678 37886 81730 37938
rect 85486 37886 85538 37938
rect 96238 37886 96290 37938
rect 96574 37886 96626 37938
rect 2046 37774 2098 37826
rect 2494 37774 2546 37826
rect 5966 37774 6018 37826
rect 24222 37774 24274 37826
rect 25006 37774 25058 37826
rect 26350 37774 26402 37826
rect 27358 37774 27410 37826
rect 29598 37774 29650 37826
rect 30046 37774 30098 37826
rect 33966 37774 34018 37826
rect 35646 37774 35698 37826
rect 37102 37774 37154 37826
rect 37326 37774 37378 37826
rect 41470 37774 41522 37826
rect 43934 37774 43986 37826
rect 46622 37774 46674 37826
rect 55806 37774 55858 37826
rect 56366 37774 56418 37826
rect 58942 37774 58994 37826
rect 59950 37774 60002 37826
rect 66446 37774 66498 37826
rect 67006 37774 67058 37826
rect 67230 37774 67282 37826
rect 68798 37774 68850 37826
rect 68910 37774 68962 37826
rect 71934 37774 71986 37826
rect 72718 37774 72770 37826
rect 74958 37774 75010 37826
rect 82462 37774 82514 37826
rect 83470 37774 83522 37826
rect 84254 37774 84306 37826
rect 84366 37774 84418 37826
rect 84478 37774 84530 37826
rect 85374 37774 85426 37826
rect 85934 37774 85986 37826
rect 88062 37774 88114 37826
rect 8896 37606 8948 37658
rect 9020 37606 9072 37658
rect 9144 37606 9196 37658
rect 9268 37606 9320 37658
rect 17896 37606 17948 37658
rect 18020 37606 18072 37658
rect 18144 37606 18196 37658
rect 18268 37606 18320 37658
rect 26896 37606 26948 37658
rect 27020 37606 27072 37658
rect 27144 37606 27196 37658
rect 27268 37606 27320 37658
rect 35896 37606 35948 37658
rect 36020 37606 36072 37658
rect 36144 37606 36196 37658
rect 36268 37606 36320 37658
rect 44896 37606 44948 37658
rect 45020 37606 45072 37658
rect 45144 37606 45196 37658
rect 45268 37606 45320 37658
rect 53896 37606 53948 37658
rect 54020 37606 54072 37658
rect 54144 37606 54196 37658
rect 54268 37606 54320 37658
rect 62896 37606 62948 37658
rect 63020 37606 63072 37658
rect 63144 37606 63196 37658
rect 63268 37606 63320 37658
rect 71896 37606 71948 37658
rect 72020 37606 72072 37658
rect 72144 37606 72196 37658
rect 72268 37606 72320 37658
rect 80896 37606 80948 37658
rect 81020 37606 81072 37658
rect 81144 37606 81196 37658
rect 81268 37606 81320 37658
rect 89896 37606 89948 37658
rect 90020 37606 90072 37658
rect 90144 37606 90196 37658
rect 90268 37606 90320 37658
rect 18398 37438 18450 37490
rect 20190 37438 20242 37490
rect 21646 37438 21698 37490
rect 29150 37438 29202 37490
rect 38558 37438 38610 37490
rect 39454 37438 39506 37490
rect 40462 37438 40514 37490
rect 47182 37438 47234 37490
rect 49870 37438 49922 37490
rect 52110 37438 52162 37490
rect 53678 37438 53730 37490
rect 55358 37438 55410 37490
rect 57934 37438 57986 37490
rect 60958 37438 61010 37490
rect 61742 37438 61794 37490
rect 63870 37438 63922 37490
rect 64430 37438 64482 37490
rect 67790 37438 67842 37490
rect 68238 37438 68290 37490
rect 75294 37438 75346 37490
rect 75854 37438 75906 37490
rect 76862 37438 76914 37490
rect 78654 37438 78706 37490
rect 86830 37438 86882 37490
rect 88062 37438 88114 37490
rect 96462 37438 96514 37490
rect 5070 37326 5122 37378
rect 5854 37326 5906 37378
rect 6078 37326 6130 37378
rect 8318 37326 8370 37378
rect 8654 37326 8706 37378
rect 8990 37326 9042 37378
rect 9662 37326 9714 37378
rect 10222 37326 10274 37378
rect 10558 37326 10610 37378
rect 15262 37326 15314 37378
rect 20638 37326 20690 37378
rect 31726 37326 31778 37378
rect 33070 37326 33122 37378
rect 33406 37326 33458 37378
rect 36878 37326 36930 37378
rect 37998 37326 38050 37378
rect 41918 37326 41970 37378
rect 43374 37326 43426 37378
rect 46398 37326 46450 37378
rect 50654 37326 50706 37378
rect 54238 37326 54290 37378
rect 54574 37326 54626 37378
rect 66334 37326 66386 37378
rect 77646 37326 77698 37378
rect 90414 37326 90466 37378
rect 2382 37214 2434 37266
rect 2718 37214 2770 37266
rect 6526 37214 6578 37266
rect 15598 37214 15650 37266
rect 20526 37214 20578 37266
rect 21310 37214 21362 37266
rect 26238 37214 26290 37266
rect 26686 37214 26738 37266
rect 29710 37214 29762 37266
rect 29934 37214 29986 37266
rect 34862 37214 34914 37266
rect 35086 37214 35138 37266
rect 35758 37214 35810 37266
rect 38334 37214 38386 37266
rect 39790 37214 39842 37266
rect 41022 37214 41074 37266
rect 41358 37214 41410 37266
rect 42030 37214 42082 37266
rect 43598 37214 43650 37266
rect 44046 37214 44098 37266
rect 50206 37214 50258 37266
rect 50430 37214 50482 37266
rect 51550 37214 51602 37266
rect 58158 37214 58210 37266
rect 58718 37214 58770 37266
rect 64766 37214 64818 37266
rect 65214 37214 65266 37266
rect 65550 37214 65602 37266
rect 66110 37214 66162 37266
rect 72382 37214 72434 37266
rect 72718 37214 72770 37266
rect 77534 37214 77586 37266
rect 78318 37214 78370 37266
rect 83918 37214 83970 37266
rect 84366 37214 84418 37266
rect 96126 37214 96178 37266
rect 96910 37214 96962 37266
rect 1822 37102 1874 37154
rect 7086 37102 7138 37154
rect 11342 37102 11394 37154
rect 11902 37102 11954 37154
rect 19630 37102 19682 37154
rect 39118 37102 39170 37154
rect 42702 37102 42754 37154
rect 48974 37102 49026 37154
rect 49422 37102 49474 37154
rect 51214 37102 51266 37154
rect 54014 37102 54066 37154
rect 66894 37102 66946 37154
rect 76190 37102 76242 37154
rect 98030 37102 98082 37154
rect 9998 36990 10050 37042
rect 30942 36990 30994 37042
rect 87502 36990 87554 37042
rect 4396 36822 4448 36874
rect 4520 36822 4572 36874
rect 4644 36822 4696 36874
rect 4768 36822 4820 36874
rect 13396 36822 13448 36874
rect 13520 36822 13572 36874
rect 13644 36822 13696 36874
rect 13768 36822 13820 36874
rect 22396 36822 22448 36874
rect 22520 36822 22572 36874
rect 22644 36822 22696 36874
rect 22768 36822 22820 36874
rect 31396 36822 31448 36874
rect 31520 36822 31572 36874
rect 31644 36822 31696 36874
rect 31768 36822 31820 36874
rect 40396 36822 40448 36874
rect 40520 36822 40572 36874
rect 40644 36822 40696 36874
rect 40768 36822 40820 36874
rect 49396 36822 49448 36874
rect 49520 36822 49572 36874
rect 49644 36822 49696 36874
rect 49768 36822 49820 36874
rect 58396 36822 58448 36874
rect 58520 36822 58572 36874
rect 58644 36822 58696 36874
rect 58768 36822 58820 36874
rect 67396 36822 67448 36874
rect 67520 36822 67572 36874
rect 67644 36822 67696 36874
rect 67768 36822 67820 36874
rect 76396 36822 76448 36874
rect 76520 36822 76572 36874
rect 76644 36822 76696 36874
rect 76768 36822 76820 36874
rect 85396 36822 85448 36874
rect 85520 36822 85572 36874
rect 85644 36822 85696 36874
rect 85768 36822 85820 36874
rect 94396 36822 94448 36874
rect 94520 36822 94572 36874
rect 94644 36822 94696 36874
rect 94768 36822 94820 36874
rect 18958 36654 19010 36706
rect 35086 36654 35138 36706
rect 53342 36654 53394 36706
rect 3278 36542 3330 36594
rect 7310 36542 7362 36594
rect 46958 36542 47010 36594
rect 50878 36542 50930 36594
rect 51998 36542 52050 36594
rect 56814 36542 56866 36594
rect 64878 36542 64930 36594
rect 67454 36542 67506 36594
rect 68798 36542 68850 36594
rect 77198 36542 77250 36594
rect 1710 36430 1762 36482
rect 6750 36430 6802 36482
rect 8654 36430 8706 36482
rect 9214 36430 9266 36482
rect 12350 36430 12402 36482
rect 14814 36430 14866 36482
rect 15374 36430 15426 36482
rect 19742 36430 19794 36482
rect 27470 36430 27522 36482
rect 31614 36430 31666 36482
rect 32062 36430 32114 36482
rect 37326 36430 37378 36482
rect 47742 36430 47794 36482
rect 51550 36430 51602 36482
rect 52782 36430 52834 36482
rect 53006 36430 53058 36482
rect 53230 36430 53282 36482
rect 69470 36430 69522 36482
rect 92206 36430 92258 36482
rect 92430 36430 92482 36482
rect 14590 36318 14642 36370
rect 17726 36318 17778 36370
rect 18510 36318 18562 36370
rect 27134 36318 27186 36370
rect 36990 36318 37042 36370
rect 37102 36318 37154 36370
rect 37662 36318 37714 36370
rect 46734 36318 46786 36370
rect 53454 36318 53506 36370
rect 67790 36318 67842 36370
rect 69582 36318 69634 36370
rect 90526 36318 90578 36370
rect 96238 36318 96290 36370
rect 96574 36318 96626 36370
rect 2046 36206 2098 36258
rect 2718 36206 2770 36258
rect 6302 36206 6354 36258
rect 8430 36206 8482 36258
rect 11566 36206 11618 36258
rect 21310 36206 21362 36258
rect 29822 36206 29874 36258
rect 31166 36206 31218 36258
rect 34302 36206 34354 36258
rect 38894 36206 38946 36258
rect 45950 36206 46002 36258
rect 46398 36206 46450 36258
rect 48414 36206 48466 36258
rect 48974 36206 49026 36258
rect 53902 36206 53954 36258
rect 68462 36206 68514 36258
rect 78990 36206 79042 36258
rect 90862 36206 90914 36258
rect 91310 36206 91362 36258
rect 91870 36206 91922 36258
rect 8896 36038 8948 36090
rect 9020 36038 9072 36090
rect 9144 36038 9196 36090
rect 9268 36038 9320 36090
rect 17896 36038 17948 36090
rect 18020 36038 18072 36090
rect 18144 36038 18196 36090
rect 18268 36038 18320 36090
rect 26896 36038 26948 36090
rect 27020 36038 27072 36090
rect 27144 36038 27196 36090
rect 27268 36038 27320 36090
rect 35896 36038 35948 36090
rect 36020 36038 36072 36090
rect 36144 36038 36196 36090
rect 36268 36038 36320 36090
rect 44896 36038 44948 36090
rect 45020 36038 45072 36090
rect 45144 36038 45196 36090
rect 45268 36038 45320 36090
rect 53896 36038 53948 36090
rect 54020 36038 54072 36090
rect 54144 36038 54196 36090
rect 54268 36038 54320 36090
rect 62896 36038 62948 36090
rect 63020 36038 63072 36090
rect 63144 36038 63196 36090
rect 63268 36038 63320 36090
rect 71896 36038 71948 36090
rect 72020 36038 72072 36090
rect 72144 36038 72196 36090
rect 72268 36038 72320 36090
rect 80896 36038 80948 36090
rect 81020 36038 81072 36090
rect 81144 36038 81196 36090
rect 81268 36038 81320 36090
rect 89896 36038 89948 36090
rect 90020 36038 90072 36090
rect 90144 36038 90196 36090
rect 90268 36038 90320 36090
rect 5630 35870 5682 35922
rect 6638 35870 6690 35922
rect 16494 35870 16546 35922
rect 17502 35870 17554 35922
rect 18622 35870 18674 35922
rect 19742 35870 19794 35922
rect 36766 35870 36818 35922
rect 37326 35870 37378 35922
rect 38670 35870 38722 35922
rect 39118 35870 39170 35922
rect 52446 35870 52498 35922
rect 57150 35870 57202 35922
rect 57374 35870 57426 35922
rect 2046 35758 2098 35810
rect 15486 35758 15538 35810
rect 20302 35758 20354 35810
rect 22094 35758 22146 35810
rect 39566 35758 39618 35810
rect 46510 35758 46562 35810
rect 47742 35758 47794 35810
rect 49758 35758 49810 35810
rect 53342 35758 53394 35810
rect 53566 35758 53618 35810
rect 62974 35758 63026 35810
rect 68350 35814 68402 35866
rect 77982 35870 78034 35922
rect 78206 35870 78258 35922
rect 78430 35870 78482 35922
rect 84254 35870 84306 35922
rect 84590 35870 84642 35922
rect 89854 35870 89906 35922
rect 92990 35870 93042 35922
rect 93774 35870 93826 35922
rect 68686 35758 68738 35810
rect 72382 35758 72434 35810
rect 79102 35758 79154 35810
rect 80222 35758 80274 35810
rect 85486 35758 85538 35810
rect 89294 35758 89346 35810
rect 1710 35646 1762 35698
rect 2718 35646 2770 35698
rect 3054 35646 3106 35698
rect 6190 35646 6242 35698
rect 15374 35646 15426 35698
rect 16158 35646 16210 35698
rect 20190 35646 20242 35698
rect 21310 35646 21362 35698
rect 21758 35646 21810 35698
rect 36654 35646 36706 35698
rect 39006 35646 39058 35698
rect 39342 35646 39394 35698
rect 47182 35646 47234 35698
rect 48974 35646 49026 35698
rect 53118 35646 53170 35698
rect 53790 35646 53842 35698
rect 56030 35646 56082 35698
rect 57150 35646 57202 35698
rect 57598 35646 57650 35698
rect 57822 35646 57874 35698
rect 62638 35646 62690 35698
rect 68126 35646 68178 35698
rect 78878 35646 78930 35698
rect 79998 35646 80050 35698
rect 80334 35646 80386 35698
rect 84702 35646 84754 35698
rect 84814 35646 84866 35698
rect 85262 35646 85314 35698
rect 86046 35646 86098 35698
rect 90302 35646 90354 35698
rect 90750 35646 90802 35698
rect 96910 35646 96962 35698
rect 14926 35534 14978 35586
rect 36206 35534 36258 35586
rect 45054 35534 45106 35586
rect 45390 35534 45442 35586
rect 45502 35534 45554 35586
rect 20974 35422 21026 35474
rect 36766 35422 36818 35474
rect 45950 35534 46002 35586
rect 56702 35534 56754 35586
rect 78318 35534 78370 35586
rect 80782 35534 80834 35586
rect 89070 35534 89122 35586
rect 45950 35422 46002 35474
rect 46286 35422 46338 35474
rect 46622 35422 46674 35474
rect 54126 35422 54178 35474
rect 89518 35422 89570 35474
rect 97694 35422 97746 35474
rect 4396 35254 4448 35306
rect 4520 35254 4572 35306
rect 4644 35254 4696 35306
rect 4768 35254 4820 35306
rect 13396 35254 13448 35306
rect 13520 35254 13572 35306
rect 13644 35254 13696 35306
rect 13768 35254 13820 35306
rect 22396 35254 22448 35306
rect 22520 35254 22572 35306
rect 22644 35254 22696 35306
rect 22768 35254 22820 35306
rect 31396 35254 31448 35306
rect 31520 35254 31572 35306
rect 31644 35254 31696 35306
rect 31768 35254 31820 35306
rect 40396 35254 40448 35306
rect 40520 35254 40572 35306
rect 40644 35254 40696 35306
rect 40768 35254 40820 35306
rect 49396 35254 49448 35306
rect 49520 35254 49572 35306
rect 49644 35254 49696 35306
rect 49768 35254 49820 35306
rect 58396 35254 58448 35306
rect 58520 35254 58572 35306
rect 58644 35254 58696 35306
rect 58768 35254 58820 35306
rect 67396 35254 67448 35306
rect 67520 35254 67572 35306
rect 67644 35254 67696 35306
rect 67768 35254 67820 35306
rect 76396 35254 76448 35306
rect 76520 35254 76572 35306
rect 76644 35254 76696 35306
rect 76768 35254 76820 35306
rect 85396 35254 85448 35306
rect 85520 35254 85572 35306
rect 85644 35254 85696 35306
rect 85768 35254 85820 35306
rect 94396 35254 94448 35306
rect 94520 35254 94572 35306
rect 94644 35254 94696 35306
rect 94768 35254 94820 35306
rect 44046 35086 44098 35138
rect 52782 35086 52834 35138
rect 71934 35086 71986 35138
rect 81566 35086 81618 35138
rect 20750 34974 20802 35026
rect 35310 34974 35362 35026
rect 39006 34974 39058 35026
rect 51662 34974 51714 35026
rect 52110 34974 52162 35026
rect 89966 34974 90018 35026
rect 5518 34862 5570 34914
rect 6078 34862 6130 34914
rect 21198 34862 21250 34914
rect 21870 34862 21922 34914
rect 35870 34862 35922 34914
rect 38670 34862 38722 34914
rect 39118 34862 39170 34914
rect 45502 34862 45554 34914
rect 46062 34862 46114 34914
rect 47294 34862 47346 34914
rect 51102 34862 51154 34914
rect 52558 34862 52610 34914
rect 55246 34862 55298 34914
rect 55806 34862 55858 34914
rect 58942 34862 58994 34914
rect 61630 34862 61682 34914
rect 61966 34862 62018 34914
rect 68462 34862 68514 34914
rect 68910 34862 68962 34914
rect 72158 34862 72210 34914
rect 72718 34862 72770 34914
rect 78094 34862 78146 34914
rect 78430 34862 78482 34914
rect 84590 34862 84642 34914
rect 85038 34862 85090 34914
rect 1710 34750 1762 34802
rect 5070 34750 5122 34802
rect 24894 34750 24946 34802
rect 35758 34750 35810 34802
rect 36990 34750 37042 34802
rect 40798 34750 40850 34802
rect 43038 34750 43090 34802
rect 44942 34750 44994 34802
rect 46846 34750 46898 34802
rect 48414 34750 48466 34802
rect 49870 34750 49922 34802
rect 53118 34750 53170 34802
rect 55022 34750 55074 34802
rect 65438 34750 65490 34802
rect 77646 34750 77698 34802
rect 80782 34750 80834 34802
rect 88174 34750 88226 34802
rect 96238 34750 96290 34802
rect 96574 34750 96626 34802
rect 2046 34638 2098 34690
rect 2382 34638 2434 34690
rect 2942 34638 2994 34690
rect 8654 34638 8706 34690
rect 9214 34638 9266 34690
rect 11342 34638 11394 34690
rect 24222 34638 24274 34690
rect 26238 34638 26290 34690
rect 27470 34638 27522 34690
rect 35534 34638 35586 34690
rect 36430 34638 36482 34690
rect 41246 34638 41298 34690
rect 46958 34638 47010 34690
rect 50318 34638 50370 34690
rect 52894 34638 52946 34690
rect 54686 34638 54738 34690
rect 58158 34638 58210 34690
rect 67902 34638 67954 34690
rect 71150 34638 71202 34690
rect 75182 34638 75234 34690
rect 75742 34638 75794 34690
rect 76414 34638 76466 34690
rect 84366 34638 84418 34690
rect 87390 34638 87442 34690
rect 8896 34470 8948 34522
rect 9020 34470 9072 34522
rect 9144 34470 9196 34522
rect 9268 34470 9320 34522
rect 17896 34470 17948 34522
rect 18020 34470 18072 34522
rect 18144 34470 18196 34522
rect 18268 34470 18320 34522
rect 26896 34470 26948 34522
rect 27020 34470 27072 34522
rect 27144 34470 27196 34522
rect 27268 34470 27320 34522
rect 35896 34470 35948 34522
rect 36020 34470 36072 34522
rect 36144 34470 36196 34522
rect 36268 34470 36320 34522
rect 44896 34470 44948 34522
rect 45020 34470 45072 34522
rect 45144 34470 45196 34522
rect 45268 34470 45320 34522
rect 53896 34470 53948 34522
rect 54020 34470 54072 34522
rect 54144 34470 54196 34522
rect 54268 34470 54320 34522
rect 62896 34470 62948 34522
rect 63020 34470 63072 34522
rect 63144 34470 63196 34522
rect 63268 34470 63320 34522
rect 71896 34470 71948 34522
rect 72020 34470 72072 34522
rect 72144 34470 72196 34522
rect 72268 34470 72320 34522
rect 80896 34470 80948 34522
rect 81020 34470 81072 34522
rect 81144 34470 81196 34522
rect 81268 34470 81320 34522
rect 89896 34470 89948 34522
rect 90020 34470 90072 34522
rect 90144 34470 90196 34522
rect 90268 34470 90320 34522
rect 4734 34302 4786 34354
rect 30158 34302 30210 34354
rect 37102 34302 37154 34354
rect 38670 34302 38722 34354
rect 39566 34302 39618 34354
rect 41022 34302 41074 34354
rect 41470 34302 41522 34354
rect 46286 34302 46338 34354
rect 47966 34302 48018 34354
rect 50430 34302 50482 34354
rect 50990 34302 51042 34354
rect 51550 34302 51602 34354
rect 55694 34302 55746 34354
rect 61630 34302 61682 34354
rect 62190 34302 62242 34354
rect 64654 34302 64706 34354
rect 72494 34302 72546 34354
rect 72830 34302 72882 34354
rect 74510 34302 74562 34354
rect 85374 34302 85426 34354
rect 85822 34302 85874 34354
rect 14030 34190 14082 34242
rect 20862 34190 20914 34242
rect 30942 34190 30994 34242
rect 32510 34190 32562 34242
rect 35870 34190 35922 34242
rect 40238 34190 40290 34242
rect 47518 34190 47570 34242
rect 52670 34190 52722 34242
rect 55358 34190 55410 34242
rect 57374 34190 57426 34242
rect 57710 34190 57762 34242
rect 63086 34190 63138 34242
rect 63758 34190 63810 34242
rect 76190 34190 76242 34242
rect 76526 34190 76578 34242
rect 85934 34190 85986 34242
rect 1822 34078 1874 34130
rect 2270 34078 2322 34130
rect 11342 34078 11394 34130
rect 11790 34078 11842 34130
rect 27358 34078 27410 34130
rect 27806 34078 27858 34130
rect 32958 34078 33010 34130
rect 33518 34078 33570 34130
rect 39006 34078 39058 34130
rect 39342 34078 39394 34130
rect 39790 34078 39842 34130
rect 40126 34078 40178 34130
rect 46846 34078 46898 34130
rect 47294 34078 47346 34130
rect 47406 34078 47458 34130
rect 49310 34078 49362 34130
rect 49758 34078 49810 34130
rect 50094 34078 50146 34130
rect 52334 34078 52386 34130
rect 56030 34078 56082 34130
rect 56814 34078 56866 34130
rect 62974 34078 63026 34130
rect 64318 34078 64370 34130
rect 64654 34078 64706 34130
rect 64878 34078 64930 34130
rect 65438 34078 65490 34130
rect 72718 34078 72770 34130
rect 72942 34078 72994 34130
rect 73390 34078 73442 34130
rect 74286 34078 74338 34130
rect 74622 34078 74674 34130
rect 96574 34078 96626 34130
rect 97022 34078 97074 34130
rect 5294 33966 5346 34018
rect 5630 33966 5682 34018
rect 27022 33966 27074 34018
rect 31390 33966 31442 34018
rect 32174 33966 32226 34018
rect 38222 33966 38274 34018
rect 39454 33966 39506 34018
rect 44606 33966 44658 34018
rect 45278 33966 45330 34018
rect 48862 33966 48914 34018
rect 61070 33966 61122 34018
rect 73726 33966 73778 34018
rect 75070 33966 75122 34018
rect 14814 33854 14866 33906
rect 57150 33854 57202 33906
rect 62526 33854 62578 33906
rect 85822 33854 85874 33906
rect 97694 33854 97746 33906
rect 4396 33686 4448 33738
rect 4520 33686 4572 33738
rect 4644 33686 4696 33738
rect 4768 33686 4820 33738
rect 13396 33686 13448 33738
rect 13520 33686 13572 33738
rect 13644 33686 13696 33738
rect 13768 33686 13820 33738
rect 22396 33686 22448 33738
rect 22520 33686 22572 33738
rect 22644 33686 22696 33738
rect 22768 33686 22820 33738
rect 31396 33686 31448 33738
rect 31520 33686 31572 33738
rect 31644 33686 31696 33738
rect 31768 33686 31820 33738
rect 40396 33686 40448 33738
rect 40520 33686 40572 33738
rect 40644 33686 40696 33738
rect 40768 33686 40820 33738
rect 49396 33686 49448 33738
rect 49520 33686 49572 33738
rect 49644 33686 49696 33738
rect 49768 33686 49820 33738
rect 58396 33686 58448 33738
rect 58520 33686 58572 33738
rect 58644 33686 58696 33738
rect 58768 33686 58820 33738
rect 67396 33686 67448 33738
rect 67520 33686 67572 33738
rect 67644 33686 67696 33738
rect 67768 33686 67820 33738
rect 76396 33686 76448 33738
rect 76520 33686 76572 33738
rect 76644 33686 76696 33738
rect 76768 33686 76820 33738
rect 85396 33686 85448 33738
rect 85520 33686 85572 33738
rect 85644 33686 85696 33738
rect 85768 33686 85820 33738
rect 94396 33686 94448 33738
rect 94520 33686 94572 33738
rect 94644 33686 94696 33738
rect 94768 33686 94820 33738
rect 45502 33518 45554 33570
rect 14590 33406 14642 33458
rect 19070 33406 19122 33458
rect 45950 33406 46002 33458
rect 53230 33406 53282 33458
rect 60846 33406 60898 33458
rect 67006 33406 67058 33458
rect 15038 33294 15090 33346
rect 15822 33294 15874 33346
rect 16718 33294 16770 33346
rect 19630 33294 19682 33346
rect 20302 33294 20354 33346
rect 20638 33294 20690 33346
rect 21534 33294 21586 33346
rect 38894 33294 38946 33346
rect 39342 33294 39394 33346
rect 44270 33294 44322 33346
rect 45054 33294 45106 33346
rect 45166 33294 45218 33346
rect 45390 33294 45442 33346
rect 48526 33294 48578 33346
rect 48862 33294 48914 33346
rect 61854 33294 61906 33346
rect 63198 33294 63250 33346
rect 63534 33294 63586 33346
rect 1710 33182 1762 33234
rect 2494 33182 2546 33234
rect 15150 33182 15202 33234
rect 19518 33182 19570 33234
rect 43934 33182 43986 33234
rect 47406 33182 47458 33234
rect 49422 33182 49474 33234
rect 62078 33182 62130 33234
rect 62526 33182 62578 33234
rect 2046 33070 2098 33122
rect 8878 33070 8930 33122
rect 16158 33070 16210 33122
rect 21310 33070 21362 33122
rect 32510 33070 32562 33122
rect 38558 33070 38610 33122
rect 41806 33070 41858 33122
rect 42366 33070 42418 33122
rect 44046 33070 44098 33122
rect 46398 33070 46450 33122
rect 50430 33070 50482 33122
rect 56366 33070 56418 33122
rect 61518 33070 61570 33122
rect 66110 33070 66162 33122
rect 66670 33070 66722 33122
rect 8896 32902 8948 32954
rect 9020 32902 9072 32954
rect 9144 32902 9196 32954
rect 9268 32902 9320 32954
rect 17896 32902 17948 32954
rect 18020 32902 18072 32954
rect 18144 32902 18196 32954
rect 18268 32902 18320 32954
rect 26896 32902 26948 32954
rect 27020 32902 27072 32954
rect 27144 32902 27196 32954
rect 27268 32902 27320 32954
rect 35896 32902 35948 32954
rect 36020 32902 36072 32954
rect 36144 32902 36196 32954
rect 36268 32902 36320 32954
rect 44896 32902 44948 32954
rect 45020 32902 45072 32954
rect 45144 32902 45196 32954
rect 45268 32902 45320 32954
rect 53896 32902 53948 32954
rect 54020 32902 54072 32954
rect 54144 32902 54196 32954
rect 54268 32902 54320 32954
rect 62896 32902 62948 32954
rect 63020 32902 63072 32954
rect 63144 32902 63196 32954
rect 63268 32902 63320 32954
rect 71896 32902 71948 32954
rect 72020 32902 72072 32954
rect 72144 32902 72196 32954
rect 72268 32902 72320 32954
rect 80896 32902 80948 32954
rect 81020 32902 81072 32954
rect 81144 32902 81196 32954
rect 81268 32902 81320 32954
rect 89896 32902 89948 32954
rect 90020 32902 90072 32954
rect 90144 32902 90196 32954
rect 90268 32902 90320 32954
rect 13134 32734 13186 32786
rect 29038 32734 29090 32786
rect 38894 32734 38946 32786
rect 41022 32734 41074 32786
rect 41470 32734 41522 32786
rect 46174 32734 46226 32786
rect 47854 32734 47906 32786
rect 48302 32734 48354 32786
rect 52558 32734 52610 32786
rect 53118 32734 53170 32786
rect 55246 32734 55298 32786
rect 55694 32734 55746 32786
rect 59838 32734 59890 32786
rect 60734 32734 60786 32786
rect 61182 32734 61234 32786
rect 63758 32734 63810 32786
rect 2046 32622 2098 32674
rect 8542 32622 8594 32674
rect 12350 32622 12402 32674
rect 14814 32622 14866 32674
rect 15150 32622 15202 32674
rect 15486 32622 15538 32674
rect 20302 32622 20354 32674
rect 23438 32622 23490 32674
rect 29710 32622 29762 32674
rect 35982 32622 36034 32674
rect 39230 32622 39282 32674
rect 44046 32622 44098 32674
rect 46398 32622 46450 32674
rect 49198 32622 49250 32674
rect 54574 32622 54626 32674
rect 56030 32622 56082 32674
rect 57262 32622 57314 32674
rect 57822 32622 57874 32674
rect 61406 32622 61458 32674
rect 63310 32622 63362 32674
rect 1710 32510 1762 32562
rect 9102 32510 9154 32562
rect 9550 32510 9602 32562
rect 9998 32510 10050 32562
rect 20526 32510 20578 32562
rect 21198 32510 21250 32562
rect 26126 32510 26178 32562
rect 26462 32510 26514 32562
rect 35870 32510 35922 32562
rect 36206 32510 36258 32562
rect 39342 32510 39394 32562
rect 39678 32510 39730 32562
rect 39902 32510 39954 32562
rect 40238 32510 40290 32562
rect 43822 32510 43874 32562
rect 45726 32510 45778 32562
rect 46510 32510 46562 32562
rect 49422 32510 49474 32562
rect 50094 32510 50146 32562
rect 53790 32510 53842 32562
rect 54462 32510 54514 32562
rect 57038 32510 57090 32562
rect 61742 32510 61794 32562
rect 62526 32510 62578 32562
rect 62974 32510 63026 32562
rect 2494 32398 2546 32450
rect 25790 32398 25842 32450
rect 30158 32398 30210 32450
rect 38446 32398 38498 32450
rect 44606 32398 44658 32450
rect 60286 32398 60338 32450
rect 63086 32398 63138 32450
rect 64878 32398 64930 32450
rect 24222 32286 24274 32338
rect 53454 32286 53506 32338
rect 56702 32286 56754 32338
rect 4396 32118 4448 32170
rect 4520 32118 4572 32170
rect 4644 32118 4696 32170
rect 4768 32118 4820 32170
rect 13396 32118 13448 32170
rect 13520 32118 13572 32170
rect 13644 32118 13696 32170
rect 13768 32118 13820 32170
rect 22396 32118 22448 32170
rect 22520 32118 22572 32170
rect 22644 32118 22696 32170
rect 22768 32118 22820 32170
rect 31396 32118 31448 32170
rect 31520 32118 31572 32170
rect 31644 32118 31696 32170
rect 31768 32118 31820 32170
rect 40396 32118 40448 32170
rect 40520 32118 40572 32170
rect 40644 32118 40696 32170
rect 40768 32118 40820 32170
rect 49396 32118 49448 32170
rect 49520 32118 49572 32170
rect 49644 32118 49696 32170
rect 49768 32118 49820 32170
rect 58396 32118 58448 32170
rect 58520 32118 58572 32170
rect 58644 32118 58696 32170
rect 58768 32118 58820 32170
rect 67396 32118 67448 32170
rect 67520 32118 67572 32170
rect 67644 32118 67696 32170
rect 67768 32118 67820 32170
rect 76396 32118 76448 32170
rect 76520 32118 76572 32170
rect 76644 32118 76696 32170
rect 76768 32118 76820 32170
rect 85396 32118 85448 32170
rect 85520 32118 85572 32170
rect 85644 32118 85696 32170
rect 85768 32118 85820 32170
rect 94396 32118 94448 32170
rect 94520 32118 94572 32170
rect 94644 32118 94696 32170
rect 94768 32118 94820 32170
rect 42366 31950 42418 32002
rect 43374 31950 43426 32002
rect 64094 31950 64146 32002
rect 9214 31838 9266 31890
rect 38894 31838 38946 31890
rect 42926 31838 42978 31890
rect 45838 31838 45890 31890
rect 53118 31838 53170 31890
rect 64430 31838 64482 31890
rect 68574 31838 68626 31890
rect 5518 31726 5570 31778
rect 6078 31726 6130 31778
rect 14590 31726 14642 31778
rect 14926 31726 14978 31778
rect 27134 31726 27186 31778
rect 36206 31726 36258 31778
rect 39230 31726 39282 31778
rect 41470 31726 41522 31778
rect 43598 31726 43650 31778
rect 44046 31726 44098 31778
rect 44830 31726 44882 31778
rect 46510 31726 46562 31778
rect 51214 31726 51266 31778
rect 56142 31726 56194 31778
rect 60398 31726 60450 31778
rect 61070 31726 61122 31778
rect 65774 31726 65826 31778
rect 69246 31726 69298 31778
rect 69806 31726 69858 31778
rect 96910 31726 96962 31778
rect 1710 31614 1762 31666
rect 5070 31614 5122 31666
rect 18062 31614 18114 31666
rect 35870 31614 35922 31666
rect 36318 31614 36370 31666
rect 36542 31614 36594 31666
rect 40686 31614 40738 31666
rect 41582 31614 41634 31666
rect 45390 31614 45442 31666
rect 50878 31614 50930 31666
rect 59950 31614 60002 31666
rect 65102 31614 65154 31666
rect 69022 31614 69074 31666
rect 72942 31614 72994 31666
rect 74062 31614 74114 31666
rect 98030 31614 98082 31666
rect 2046 31502 2098 31554
rect 2382 31502 2434 31554
rect 2942 31502 2994 31554
rect 8654 31502 8706 31554
rect 17502 31502 17554 31554
rect 18398 31502 18450 31554
rect 26798 31502 26850 31554
rect 27470 31502 27522 31554
rect 30046 31502 30098 31554
rect 32734 31502 32786 31554
rect 38446 31502 38498 31554
rect 55806 31502 55858 31554
rect 56478 31502 56530 31554
rect 63534 31502 63586 31554
rect 65214 31502 65266 31554
rect 65326 31502 65378 31554
rect 65998 31502 66050 31554
rect 66558 31502 66610 31554
rect 72158 31502 72210 31554
rect 74398 31502 74450 31554
rect 96686 31502 96738 31554
rect 8896 31334 8948 31386
rect 9020 31334 9072 31386
rect 9144 31334 9196 31386
rect 9268 31334 9320 31386
rect 17896 31334 17948 31386
rect 18020 31334 18072 31386
rect 18144 31334 18196 31386
rect 18268 31334 18320 31386
rect 26896 31334 26948 31386
rect 27020 31334 27072 31386
rect 27144 31334 27196 31386
rect 27268 31334 27320 31386
rect 35896 31334 35948 31386
rect 36020 31334 36072 31386
rect 36144 31334 36196 31386
rect 36268 31334 36320 31386
rect 44896 31334 44948 31386
rect 45020 31334 45072 31386
rect 45144 31334 45196 31386
rect 45268 31334 45320 31386
rect 53896 31334 53948 31386
rect 54020 31334 54072 31386
rect 54144 31334 54196 31386
rect 54268 31334 54320 31386
rect 62896 31334 62948 31386
rect 63020 31334 63072 31386
rect 63144 31334 63196 31386
rect 63268 31334 63320 31386
rect 71896 31334 71948 31386
rect 72020 31334 72072 31386
rect 72144 31334 72196 31386
rect 72268 31334 72320 31386
rect 80896 31334 80948 31386
rect 81020 31334 81072 31386
rect 81144 31334 81196 31386
rect 81268 31334 81320 31386
rect 89896 31334 89948 31386
rect 90020 31334 90072 31386
rect 90144 31334 90196 31386
rect 90268 31334 90320 31386
rect 4734 31166 4786 31218
rect 19966 31166 20018 31218
rect 29374 31166 29426 31218
rect 30606 31166 30658 31218
rect 38894 31166 38946 31218
rect 39790 31166 39842 31218
rect 42702 31166 42754 31218
rect 61182 31166 61234 31218
rect 67902 31166 67954 31218
rect 68910 31166 68962 31218
rect 69806 31166 69858 31218
rect 69918 31166 69970 31218
rect 70702 31166 70754 31218
rect 72382 31166 72434 31218
rect 72942 31166 72994 31218
rect 20862 31054 20914 31106
rect 23998 31054 24050 31106
rect 31054 31054 31106 31106
rect 35870 31054 35922 31106
rect 43822 31054 43874 31106
rect 45054 31054 45106 31106
rect 46846 31054 46898 31106
rect 69470 31054 69522 31106
rect 69694 31054 69746 31106
rect 1822 30942 1874 30994
rect 2158 30942 2210 30994
rect 20414 30942 20466 30994
rect 21086 30942 21138 30994
rect 21646 30942 21698 30994
rect 26462 30942 26514 30994
rect 26798 30942 26850 30994
rect 30942 30942 30994 30994
rect 32958 30942 33010 30994
rect 33518 30942 33570 30994
rect 39678 30942 39730 30994
rect 40014 30942 40066 30994
rect 44046 30942 44098 30994
rect 46398 30942 46450 30994
rect 47182 30942 47234 30994
rect 61518 30942 61570 30994
rect 65102 30942 65154 30994
rect 65438 30942 65490 30994
rect 70366 30942 70418 30994
rect 72494 30942 72546 30994
rect 14702 30830 14754 30882
rect 31726 30830 31778 30882
rect 39454 30830 39506 30882
rect 44494 30830 44546 30882
rect 46958 30830 47010 30882
rect 5294 30718 5346 30770
rect 24782 30718 24834 30770
rect 29934 30718 29986 30770
rect 32062 30718 32114 30770
rect 36654 30718 36706 30770
rect 39230 30718 39282 30770
rect 39454 30718 39506 30770
rect 68574 30718 68626 30770
rect 72382 30718 72434 30770
rect 4396 30550 4448 30602
rect 4520 30550 4572 30602
rect 4644 30550 4696 30602
rect 4768 30550 4820 30602
rect 13396 30550 13448 30602
rect 13520 30550 13572 30602
rect 13644 30550 13696 30602
rect 13768 30550 13820 30602
rect 22396 30550 22448 30602
rect 22520 30550 22572 30602
rect 22644 30550 22696 30602
rect 22768 30550 22820 30602
rect 31396 30550 31448 30602
rect 31520 30550 31572 30602
rect 31644 30550 31696 30602
rect 31768 30550 31820 30602
rect 40396 30550 40448 30602
rect 40520 30550 40572 30602
rect 40644 30550 40696 30602
rect 40768 30550 40820 30602
rect 49396 30550 49448 30602
rect 49520 30550 49572 30602
rect 49644 30550 49696 30602
rect 49768 30550 49820 30602
rect 58396 30550 58448 30602
rect 58520 30550 58572 30602
rect 58644 30550 58696 30602
rect 58768 30550 58820 30602
rect 67396 30550 67448 30602
rect 67520 30550 67572 30602
rect 67644 30550 67696 30602
rect 67768 30550 67820 30602
rect 76396 30550 76448 30602
rect 76520 30550 76572 30602
rect 76644 30550 76696 30602
rect 76768 30550 76820 30602
rect 85396 30550 85448 30602
rect 85520 30550 85572 30602
rect 85644 30550 85696 30602
rect 85768 30550 85820 30602
rect 94396 30550 94448 30602
rect 94520 30550 94572 30602
rect 94644 30550 94696 30602
rect 94768 30550 94820 30602
rect 27918 30382 27970 30434
rect 28254 30382 28306 30434
rect 15934 30270 15986 30322
rect 43038 30270 43090 30322
rect 85150 30270 85202 30322
rect 8878 30158 8930 30210
rect 9438 30158 9490 30210
rect 15150 30158 15202 30210
rect 26238 30158 26290 30210
rect 27246 30158 27298 30210
rect 30270 30158 30322 30210
rect 31838 30158 31890 30210
rect 32734 30158 32786 30210
rect 42142 30158 42194 30210
rect 44158 30158 44210 30210
rect 45054 30158 45106 30210
rect 47070 30158 47122 30210
rect 49758 30158 49810 30210
rect 52670 30158 52722 30210
rect 66446 30158 66498 30210
rect 72494 30158 72546 30210
rect 83470 30158 83522 30210
rect 84478 30158 84530 30210
rect 96910 30158 96962 30210
rect 1710 30046 1762 30098
rect 8654 30046 8706 30098
rect 14702 30046 14754 30098
rect 15374 30046 15426 30098
rect 16270 30046 16322 30098
rect 27134 30046 27186 30098
rect 32062 30046 32114 30098
rect 36990 30046 37042 30098
rect 37102 30046 37154 30098
rect 41582 30046 41634 30098
rect 43598 30046 43650 30098
rect 45614 30046 45666 30098
rect 47630 30046 47682 30098
rect 49198 30046 49250 30098
rect 66670 30046 66722 30098
rect 66782 30046 66834 30098
rect 67230 30046 67282 30098
rect 72830 30046 72882 30098
rect 96686 30046 96738 30098
rect 98030 30046 98082 30098
rect 2046 29934 2098 29986
rect 2494 29934 2546 29986
rect 12014 29934 12066 29986
rect 12574 29934 12626 29986
rect 13918 29934 13970 29986
rect 14366 29934 14418 29986
rect 16830 29934 16882 29986
rect 26686 29934 26738 29986
rect 33182 29934 33234 29986
rect 37326 29934 37378 29986
rect 46734 29934 46786 29986
rect 49310 29934 49362 29986
rect 50206 29934 50258 29986
rect 52110 29934 52162 29986
rect 59054 29934 59106 29986
rect 8896 29766 8948 29818
rect 9020 29766 9072 29818
rect 9144 29766 9196 29818
rect 9268 29766 9320 29818
rect 17896 29766 17948 29818
rect 18020 29766 18072 29818
rect 18144 29766 18196 29818
rect 18268 29766 18320 29818
rect 26896 29766 26948 29818
rect 27020 29766 27072 29818
rect 27144 29766 27196 29818
rect 27268 29766 27320 29818
rect 35896 29766 35948 29818
rect 36020 29766 36072 29818
rect 36144 29766 36196 29818
rect 36268 29766 36320 29818
rect 44896 29766 44948 29818
rect 45020 29766 45072 29818
rect 45144 29766 45196 29818
rect 45268 29766 45320 29818
rect 53896 29766 53948 29818
rect 54020 29766 54072 29818
rect 54144 29766 54196 29818
rect 54268 29766 54320 29818
rect 62896 29766 62948 29818
rect 63020 29766 63072 29818
rect 63144 29766 63196 29818
rect 63268 29766 63320 29818
rect 71896 29766 71948 29818
rect 72020 29766 72072 29818
rect 72144 29766 72196 29818
rect 72268 29766 72320 29818
rect 80896 29766 80948 29818
rect 81020 29766 81072 29818
rect 81144 29766 81196 29818
rect 81268 29766 81320 29818
rect 89896 29766 89948 29818
rect 90020 29766 90072 29818
rect 90144 29766 90196 29818
rect 90268 29766 90320 29818
rect 5070 29598 5122 29650
rect 21534 29598 21586 29650
rect 22430 29598 22482 29650
rect 39342 29598 39394 29650
rect 39790 29598 39842 29650
rect 44046 29598 44098 29650
rect 44494 29598 44546 29650
rect 46174 29598 46226 29650
rect 46286 29598 46338 29650
rect 53118 29598 53170 29650
rect 68798 29598 68850 29650
rect 69694 29598 69746 29650
rect 1934 29486 1986 29538
rect 16158 29486 16210 29538
rect 18174 29486 18226 29538
rect 38782 29486 38834 29538
rect 43150 29486 43202 29538
rect 44158 29486 44210 29538
rect 54238 29486 54290 29538
rect 56030 29486 56082 29538
rect 56926 29486 56978 29538
rect 57598 29486 57650 29538
rect 2158 29374 2210 29426
rect 2718 29374 2770 29426
rect 13470 29374 13522 29426
rect 13918 29374 13970 29426
rect 17726 29374 17778 29426
rect 18398 29374 18450 29426
rect 18958 29374 19010 29426
rect 42478 29374 42530 29426
rect 43262 29374 43314 29426
rect 44718 29374 44770 29426
rect 45502 29374 45554 29426
rect 45838 29374 45890 29426
rect 46062 29374 46114 29426
rect 46398 29374 46450 29426
rect 46958 29374 47010 29426
rect 50206 29374 50258 29426
rect 50542 29374 50594 29426
rect 56814 29374 56866 29426
rect 57150 29374 57202 29426
rect 68574 29374 68626 29426
rect 69246 29374 69298 29426
rect 75854 29374 75906 29426
rect 13022 29262 13074 29314
rect 68350 29262 68402 29314
rect 68686 29262 68738 29314
rect 5854 29150 5906 29202
rect 16942 29150 16994 29202
rect 22094 29150 22146 29202
rect 42142 29150 42194 29202
rect 44046 29150 44098 29202
rect 53678 29150 53730 29202
rect 4396 28982 4448 29034
rect 4520 28982 4572 29034
rect 4644 28982 4696 29034
rect 4768 28982 4820 29034
rect 13396 28982 13448 29034
rect 13520 28982 13572 29034
rect 13644 28982 13696 29034
rect 13768 28982 13820 29034
rect 22396 28982 22448 29034
rect 22520 28982 22572 29034
rect 22644 28982 22696 29034
rect 22768 28982 22820 29034
rect 31396 28982 31448 29034
rect 31520 28982 31572 29034
rect 31644 28982 31696 29034
rect 31768 28982 31820 29034
rect 40396 28982 40448 29034
rect 40520 28982 40572 29034
rect 40644 28982 40696 29034
rect 40768 28982 40820 29034
rect 49396 28982 49448 29034
rect 49520 28982 49572 29034
rect 49644 28982 49696 29034
rect 49768 28982 49820 29034
rect 58396 28982 58448 29034
rect 58520 28982 58572 29034
rect 58644 28982 58696 29034
rect 58768 28982 58820 29034
rect 67396 28982 67448 29034
rect 67520 28982 67572 29034
rect 67644 28982 67696 29034
rect 67768 28982 67820 29034
rect 76396 28982 76448 29034
rect 76520 28982 76572 29034
rect 76644 28982 76696 29034
rect 76768 28982 76820 29034
rect 85396 28982 85448 29034
rect 85520 28982 85572 29034
rect 85644 28982 85696 29034
rect 85768 28982 85820 29034
rect 94396 28982 94448 29034
rect 94520 28982 94572 29034
rect 94644 28982 94696 29034
rect 94768 28982 94820 29034
rect 45054 28814 45106 28866
rect 54910 28814 54962 28866
rect 58942 28814 58994 28866
rect 61182 28814 61234 28866
rect 61742 28814 61794 28866
rect 75406 28814 75458 28866
rect 2494 28702 2546 28754
rect 24222 28702 24274 28754
rect 25902 28702 25954 28754
rect 46510 28702 46562 28754
rect 60734 28702 60786 28754
rect 67342 28702 67394 28754
rect 76750 28702 76802 28754
rect 1710 28590 1762 28642
rect 13806 28590 13858 28642
rect 25454 28590 25506 28642
rect 26238 28590 26290 28642
rect 26798 28590 26850 28642
rect 29262 28590 29314 28642
rect 41694 28590 41746 28642
rect 44382 28590 44434 28642
rect 45838 28590 45890 28642
rect 46846 28590 46898 28642
rect 47406 28590 47458 28642
rect 47742 28590 47794 28642
rect 55358 28590 55410 28642
rect 55806 28590 55858 28642
rect 62302 28590 62354 28642
rect 63198 28590 63250 28642
rect 63646 28590 63698 28642
rect 64430 28590 64482 28642
rect 68238 28590 68290 28642
rect 68798 28590 68850 28642
rect 71934 28590 71986 28642
rect 72382 28590 72434 28642
rect 77422 28590 77474 28642
rect 96574 28590 96626 28642
rect 97022 28590 97074 28642
rect 97694 28590 97746 28642
rect 2046 28478 2098 28530
rect 25230 28478 25282 28530
rect 30270 28478 30322 28530
rect 30606 28478 30658 28530
rect 55022 28478 55074 28530
rect 61070 28478 61122 28530
rect 61182 28478 61234 28530
rect 7422 28366 7474 28418
rect 24670 28366 24722 28418
rect 30942 28366 30994 28418
rect 35422 28366 35474 28418
rect 41358 28366 41410 28418
rect 48078 28366 48130 28418
rect 48526 28366 48578 28418
rect 54574 28366 54626 28418
rect 61630 28422 61682 28474
rect 61742 28478 61794 28530
rect 62974 28478 63026 28530
rect 67790 28478 67842 28530
rect 71150 28478 71202 28530
rect 72718 28478 72770 28530
rect 74174 28478 74226 28530
rect 74398 28478 74450 28530
rect 54910 28366 54962 28418
rect 58158 28366 58210 28418
rect 63086 28366 63138 28418
rect 63870 28366 63922 28418
rect 77758 28366 77810 28418
rect 8896 28198 8948 28250
rect 9020 28198 9072 28250
rect 9144 28198 9196 28250
rect 9268 28198 9320 28250
rect 17896 28198 17948 28250
rect 18020 28198 18072 28250
rect 18144 28198 18196 28250
rect 18268 28198 18320 28250
rect 26896 28198 26948 28250
rect 27020 28198 27072 28250
rect 27144 28198 27196 28250
rect 27268 28198 27320 28250
rect 35896 28198 35948 28250
rect 36020 28198 36072 28250
rect 36144 28198 36196 28250
rect 36268 28198 36320 28250
rect 44896 28198 44948 28250
rect 45020 28198 45072 28250
rect 45144 28198 45196 28250
rect 45268 28198 45320 28250
rect 53896 28198 53948 28250
rect 54020 28198 54072 28250
rect 54144 28198 54196 28250
rect 54268 28198 54320 28250
rect 62896 28198 62948 28250
rect 63020 28198 63072 28250
rect 63144 28198 63196 28250
rect 63268 28198 63320 28250
rect 71896 28198 71948 28250
rect 72020 28198 72072 28250
rect 72144 28198 72196 28250
rect 72268 28198 72320 28250
rect 80896 28198 80948 28250
rect 81020 28198 81072 28250
rect 81144 28198 81196 28250
rect 81268 28198 81320 28250
rect 89896 28198 89948 28250
rect 90020 28198 90072 28250
rect 90144 28198 90196 28250
rect 90268 28198 90320 28250
rect 5070 28030 5122 28082
rect 14478 28030 14530 28082
rect 28254 28030 28306 28082
rect 32062 28030 32114 28082
rect 33182 28030 33234 28082
rect 39902 28030 39954 28082
rect 43934 28030 43986 28082
rect 44494 28030 44546 28082
rect 51774 28030 51826 28082
rect 52894 28030 52946 28082
rect 55022 28030 55074 28082
rect 59614 28030 59666 28082
rect 66222 28030 66274 28082
rect 70478 28030 70530 28082
rect 70702 28030 70754 28082
rect 75742 28030 75794 28082
rect 1934 27918 1986 27970
rect 12462 27918 12514 27970
rect 14142 27918 14194 27970
rect 24670 27918 24722 27970
rect 34862 27918 34914 27970
rect 37998 27918 38050 27970
rect 40350 27918 40402 27970
rect 60174 27918 60226 27970
rect 65662 27918 65714 27970
rect 70814 27918 70866 27970
rect 71262 27918 71314 27970
rect 78878 27918 78930 27970
rect 2158 27806 2210 27858
rect 2718 27806 2770 27858
rect 6078 27806 6130 27858
rect 12238 27806 12290 27858
rect 13022 27806 13074 27858
rect 13358 27806 13410 27858
rect 13806 27806 13858 27858
rect 24446 27806 24498 27858
rect 25118 27806 25170 27858
rect 25678 27806 25730 27858
rect 29150 27806 29202 27858
rect 29598 27806 29650 27858
rect 35310 27806 35362 27858
rect 35646 27806 35698 27858
rect 40798 27806 40850 27858
rect 41358 27806 41410 27858
rect 46398 27806 46450 27858
rect 48638 27806 48690 27858
rect 49198 27806 49250 27858
rect 52446 27806 52498 27858
rect 56478 27806 56530 27858
rect 57150 27806 57202 27858
rect 65774 27806 65826 27858
rect 73614 27806 73666 27858
rect 76190 27806 76242 27858
rect 76526 27806 76578 27858
rect 6750 27694 6802 27746
rect 11790 27694 11842 27746
rect 45726 27694 45778 27746
rect 46846 27694 46898 27746
rect 56030 27694 56082 27746
rect 73166 27694 73218 27746
rect 74622 27694 74674 27746
rect 5854 27582 5906 27634
rect 28814 27582 28866 27634
rect 32622 27582 32674 27634
rect 38782 27582 38834 27634
rect 65662 27582 65714 27634
rect 79662 27582 79714 27634
rect 4396 27414 4448 27466
rect 4520 27414 4572 27466
rect 4644 27414 4696 27466
rect 4768 27414 4820 27466
rect 13396 27414 13448 27466
rect 13520 27414 13572 27466
rect 13644 27414 13696 27466
rect 13768 27414 13820 27466
rect 22396 27414 22448 27466
rect 22520 27414 22572 27466
rect 22644 27414 22696 27466
rect 22768 27414 22820 27466
rect 31396 27414 31448 27466
rect 31520 27414 31572 27466
rect 31644 27414 31696 27466
rect 31768 27414 31820 27466
rect 40396 27414 40448 27466
rect 40520 27414 40572 27466
rect 40644 27414 40696 27466
rect 40768 27414 40820 27466
rect 49396 27414 49448 27466
rect 49520 27414 49572 27466
rect 49644 27414 49696 27466
rect 49768 27414 49820 27466
rect 58396 27414 58448 27466
rect 58520 27414 58572 27466
rect 58644 27414 58696 27466
rect 58768 27414 58820 27466
rect 67396 27414 67448 27466
rect 67520 27414 67572 27466
rect 67644 27414 67696 27466
rect 67768 27414 67820 27466
rect 76396 27414 76448 27466
rect 76520 27414 76572 27466
rect 76644 27414 76696 27466
rect 76768 27414 76820 27466
rect 85396 27414 85448 27466
rect 85520 27414 85572 27466
rect 85644 27414 85696 27466
rect 85768 27414 85820 27466
rect 94396 27414 94448 27466
rect 94520 27414 94572 27466
rect 94644 27414 94696 27466
rect 94768 27414 94820 27466
rect 17390 27246 17442 27298
rect 31502 27246 31554 27298
rect 37326 27246 37378 27298
rect 56926 27246 56978 27298
rect 57262 27246 57314 27298
rect 57934 27246 57986 27298
rect 66222 27246 66274 27298
rect 17726 27134 17778 27186
rect 20750 27134 20802 27186
rect 29486 27134 29538 27186
rect 29934 27134 29986 27186
rect 32062 27134 32114 27186
rect 37550 27134 37602 27186
rect 38110 27134 38162 27186
rect 53678 27134 53730 27186
rect 59950 27134 60002 27186
rect 73838 27134 73890 27186
rect 76414 27134 76466 27186
rect 96574 27134 96626 27186
rect 1710 27022 1762 27074
rect 2606 27022 2658 27074
rect 7310 27022 7362 27074
rect 7646 27022 7698 27074
rect 13918 27022 13970 27074
rect 14254 27022 14306 27074
rect 21758 27022 21810 27074
rect 30382 27022 30434 27074
rect 31166 27022 31218 27074
rect 35422 27022 35474 27074
rect 57822 27022 57874 27074
rect 60846 27022 60898 27074
rect 61070 27022 61122 27074
rect 61630 27022 61682 27074
rect 62750 27022 62802 27074
rect 63086 27022 63138 27074
rect 67230 27022 67282 27074
rect 74286 27022 74338 27074
rect 76302 27022 76354 27074
rect 76974 27022 77026 27074
rect 77310 27022 77362 27074
rect 96910 27022 96962 27074
rect 2046 26910 2098 26962
rect 3166 26910 3218 26962
rect 5742 26910 5794 26962
rect 9998 26910 10050 26962
rect 16606 26910 16658 26962
rect 21982 26910 22034 26962
rect 22318 26910 22370 26962
rect 30494 26910 30546 26962
rect 35646 26910 35698 26962
rect 57934 26910 57986 26962
rect 60510 26910 60562 26962
rect 60622 26910 60674 26962
rect 61182 26910 61234 26962
rect 61742 26910 61794 26962
rect 61966 26910 62018 26962
rect 62302 26910 62354 26962
rect 65438 26910 65490 26962
rect 67566 26910 67618 26962
rect 75294 26910 75346 26962
rect 77534 26910 77586 26962
rect 77646 26910 77698 26962
rect 78094 26910 78146 26962
rect 97694 26910 97746 26962
rect 2382 26798 2434 26850
rect 10782 26798 10834 26850
rect 19742 26798 19794 26850
rect 21422 26798 21474 26850
rect 23102 26798 23154 26850
rect 36990 26798 37042 26850
rect 54238 26798 54290 26850
rect 57038 26798 57090 26850
rect 61406 26798 61458 26850
rect 76526 26798 76578 26850
rect 8896 26630 8948 26682
rect 9020 26630 9072 26682
rect 9144 26630 9196 26682
rect 9268 26630 9320 26682
rect 17896 26630 17948 26682
rect 18020 26630 18072 26682
rect 18144 26630 18196 26682
rect 18268 26630 18320 26682
rect 26896 26630 26948 26682
rect 27020 26630 27072 26682
rect 27144 26630 27196 26682
rect 27268 26630 27320 26682
rect 35896 26630 35948 26682
rect 36020 26630 36072 26682
rect 36144 26630 36196 26682
rect 36268 26630 36320 26682
rect 44896 26630 44948 26682
rect 45020 26630 45072 26682
rect 45144 26630 45196 26682
rect 45268 26630 45320 26682
rect 53896 26630 53948 26682
rect 54020 26630 54072 26682
rect 54144 26630 54196 26682
rect 54268 26630 54320 26682
rect 62896 26630 62948 26682
rect 63020 26630 63072 26682
rect 63144 26630 63196 26682
rect 63268 26630 63320 26682
rect 71896 26630 71948 26682
rect 72020 26630 72072 26682
rect 72144 26630 72196 26682
rect 72268 26630 72320 26682
rect 80896 26630 80948 26682
rect 81020 26630 81072 26682
rect 81144 26630 81196 26682
rect 81268 26630 81320 26682
rect 89896 26630 89948 26682
rect 90020 26630 90072 26682
rect 90144 26630 90196 26682
rect 90268 26630 90320 26682
rect 2494 26462 2546 26514
rect 11454 26462 11506 26514
rect 12014 26462 12066 26514
rect 19182 26462 19234 26514
rect 22318 26462 22370 26514
rect 23102 26462 23154 26514
rect 53006 26462 53058 26514
rect 53566 26462 53618 26514
rect 57598 26462 57650 26514
rect 59614 26462 59666 26514
rect 60062 26462 60114 26514
rect 60846 26462 60898 26514
rect 67118 26462 67170 26514
rect 72494 26462 72546 26514
rect 74734 26462 74786 26514
rect 1934 26350 1986 26402
rect 5294 26350 5346 26402
rect 26686 26350 26738 26402
rect 49646 26350 49698 26402
rect 53790 26350 53842 26402
rect 58494 26350 58546 26402
rect 59950 26350 60002 26402
rect 66670 26350 66722 26402
rect 67342 26350 67394 26402
rect 68126 26350 68178 26402
rect 72718 26350 72770 26402
rect 73502 26350 73554 26402
rect 77086 26350 77138 26402
rect 84254 26350 84306 26402
rect 19630 26238 19682 26290
rect 20078 26238 20130 26290
rect 26462 26238 26514 26290
rect 49870 26238 49922 26290
rect 50430 26238 50482 26290
rect 57038 26238 57090 26290
rect 57934 26238 57986 26290
rect 62302 26238 62354 26290
rect 67790 26238 67842 26290
rect 73166 26238 73218 26290
rect 75070 26238 75122 26290
rect 84030 26238 84082 26290
rect 10894 26126 10946 26178
rect 54798 26126 54850 26178
rect 67230 26126 67282 26178
rect 72606 26126 72658 26178
rect 75742 26126 75794 26178
rect 77982 26126 78034 26178
rect 60062 26014 60114 26066
rect 4396 25846 4448 25898
rect 4520 25846 4572 25898
rect 4644 25846 4696 25898
rect 4768 25846 4820 25898
rect 13396 25846 13448 25898
rect 13520 25846 13572 25898
rect 13644 25846 13696 25898
rect 13768 25846 13820 25898
rect 22396 25846 22448 25898
rect 22520 25846 22572 25898
rect 22644 25846 22696 25898
rect 22768 25846 22820 25898
rect 31396 25846 31448 25898
rect 31520 25846 31572 25898
rect 31644 25846 31696 25898
rect 31768 25846 31820 25898
rect 40396 25846 40448 25898
rect 40520 25846 40572 25898
rect 40644 25846 40696 25898
rect 40768 25846 40820 25898
rect 49396 25846 49448 25898
rect 49520 25846 49572 25898
rect 49644 25846 49696 25898
rect 49768 25846 49820 25898
rect 58396 25846 58448 25898
rect 58520 25846 58572 25898
rect 58644 25846 58696 25898
rect 58768 25846 58820 25898
rect 67396 25846 67448 25898
rect 67520 25846 67572 25898
rect 67644 25846 67696 25898
rect 67768 25846 67820 25898
rect 76396 25846 76448 25898
rect 76520 25846 76572 25898
rect 76644 25846 76696 25898
rect 76768 25846 76820 25898
rect 85396 25846 85448 25898
rect 85520 25846 85572 25898
rect 85644 25846 85696 25898
rect 85768 25846 85820 25898
rect 94396 25846 94448 25898
rect 94520 25846 94572 25898
rect 94644 25846 94696 25898
rect 94768 25846 94820 25898
rect 27246 25678 27298 25730
rect 35422 25678 35474 25730
rect 48414 25678 48466 25730
rect 57710 25678 57762 25730
rect 76078 25678 76130 25730
rect 76750 25678 76802 25730
rect 77086 25678 77138 25730
rect 25230 25566 25282 25618
rect 25678 25566 25730 25618
rect 53454 25566 53506 25618
rect 58046 25566 58098 25618
rect 65774 25566 65826 25618
rect 69358 25566 69410 25618
rect 76750 25566 76802 25618
rect 5518 25454 5570 25506
rect 6078 25454 6130 25506
rect 9214 25454 9266 25506
rect 11342 25454 11394 25506
rect 20638 25454 20690 25506
rect 26238 25454 26290 25506
rect 26910 25454 26962 25506
rect 34862 25454 34914 25506
rect 35086 25454 35138 25506
rect 38894 25454 38946 25506
rect 43150 25454 43202 25506
rect 43374 25454 43426 25506
rect 44718 25454 44770 25506
rect 45278 25454 45330 25506
rect 54238 25454 54290 25506
rect 54574 25454 54626 25506
rect 62302 25454 62354 25506
rect 62974 25454 63026 25506
rect 64990 25454 65042 25506
rect 65326 25454 65378 25506
rect 68574 25454 68626 25506
rect 68910 25454 68962 25506
rect 72046 25454 72098 25506
rect 72606 25454 72658 25506
rect 76302 25454 76354 25506
rect 77310 25454 77362 25506
rect 77422 25454 77474 25506
rect 77534 25454 77586 25506
rect 77870 25454 77922 25506
rect 78430 25454 78482 25506
rect 78766 25454 78818 25506
rect 1710 25342 1762 25394
rect 2046 25342 2098 25394
rect 2494 25342 2546 25394
rect 8430 25342 8482 25394
rect 10558 25342 10610 25394
rect 11118 25342 11170 25394
rect 12350 25342 12402 25394
rect 20302 25342 20354 25394
rect 26126 25342 26178 25394
rect 33070 25342 33122 25394
rect 43038 25342 43090 25394
rect 43822 25342 43874 25394
rect 44270 25342 44322 25394
rect 71822 25342 71874 25394
rect 81118 25342 81170 25394
rect 9550 25230 9602 25282
rect 11678 25230 11730 25282
rect 12686 25230 12738 25282
rect 27694 25230 27746 25282
rect 28254 25230 28306 25282
rect 33406 25230 33458 25282
rect 34078 25230 34130 25282
rect 34526 25230 34578 25282
rect 39118 25230 39170 25282
rect 39454 25230 39506 25282
rect 42702 25230 42754 25282
rect 47630 25230 47682 25282
rect 57150 25230 57202 25282
rect 61854 25230 61906 25282
rect 62414 25230 62466 25282
rect 62526 25230 62578 25282
rect 63310 25230 63362 25282
rect 65214 25230 65266 25282
rect 68798 25230 68850 25282
rect 75070 25230 75122 25282
rect 75742 25230 75794 25282
rect 81902 25230 81954 25282
rect 8896 25062 8948 25114
rect 9020 25062 9072 25114
rect 9144 25062 9196 25114
rect 9268 25062 9320 25114
rect 17896 25062 17948 25114
rect 18020 25062 18072 25114
rect 18144 25062 18196 25114
rect 18268 25062 18320 25114
rect 26896 25062 26948 25114
rect 27020 25062 27072 25114
rect 27144 25062 27196 25114
rect 27268 25062 27320 25114
rect 35896 25062 35948 25114
rect 36020 25062 36072 25114
rect 36144 25062 36196 25114
rect 36268 25062 36320 25114
rect 44896 25062 44948 25114
rect 45020 25062 45072 25114
rect 45144 25062 45196 25114
rect 45268 25062 45320 25114
rect 53896 25062 53948 25114
rect 54020 25062 54072 25114
rect 54144 25062 54196 25114
rect 54268 25062 54320 25114
rect 62896 25062 62948 25114
rect 63020 25062 63072 25114
rect 63144 25062 63196 25114
rect 63268 25062 63320 25114
rect 71896 25062 71948 25114
rect 72020 25062 72072 25114
rect 72144 25062 72196 25114
rect 72268 25062 72320 25114
rect 80896 25062 80948 25114
rect 81020 25062 81072 25114
rect 81144 25062 81196 25114
rect 81268 25062 81320 25114
rect 89896 25062 89948 25114
rect 90020 25062 90072 25114
rect 90144 25062 90196 25114
rect 90268 25062 90320 25114
rect 4734 24894 4786 24946
rect 5294 24894 5346 24946
rect 10334 24894 10386 24946
rect 11902 24894 11954 24946
rect 29374 24894 29426 24946
rect 30158 24894 30210 24946
rect 32062 24894 32114 24946
rect 39566 24894 39618 24946
rect 43038 24894 43090 24946
rect 43374 24894 43426 24946
rect 44270 24894 44322 24946
rect 60174 24894 60226 24946
rect 60622 24894 60674 24946
rect 66334 24894 66386 24946
rect 70254 24894 70306 24946
rect 74174 24894 74226 24946
rect 75070 24894 75122 24946
rect 76974 24894 77026 24946
rect 77758 24894 77810 24946
rect 77870 24894 77922 24946
rect 78094 24894 78146 24946
rect 78542 24894 78594 24946
rect 10894 24782 10946 24834
rect 12462 24782 12514 24834
rect 15598 24782 15650 24834
rect 16606 24782 16658 24834
rect 30494 24782 30546 24834
rect 32510 24782 32562 24834
rect 35870 24782 35922 24834
rect 37550 24782 37602 24834
rect 38558 24782 38610 24834
rect 60510 24782 60562 24834
rect 69470 24782 69522 24834
rect 74398 24782 74450 24834
rect 74510 24782 74562 24834
rect 83134 24782 83186 24834
rect 83470 24782 83522 24834
rect 1822 24670 1874 24722
rect 2270 24670 2322 24722
rect 5630 24670 5682 24722
rect 9774 24670 9826 24722
rect 11678 24670 11730 24722
rect 12686 24670 12738 24722
rect 13246 24670 13298 24722
rect 26462 24670 26514 24722
rect 27022 24670 27074 24722
rect 32958 24670 33010 24722
rect 33630 24670 33682 24722
rect 36654 24670 36706 24722
rect 38446 24670 38498 24722
rect 43486 24670 43538 24722
rect 66670 24670 66722 24722
rect 67230 24670 67282 24722
rect 78206 24670 78258 24722
rect 96910 24670 96962 24722
rect 38110 24558 38162 24610
rect 40238 24558 40290 24610
rect 98030 24558 98082 24610
rect 16382 24446 16434 24498
rect 39230 24446 39282 24498
rect 60622 24446 60674 24498
rect 4396 24278 4448 24330
rect 4520 24278 4572 24330
rect 4644 24278 4696 24330
rect 4768 24278 4820 24330
rect 13396 24278 13448 24330
rect 13520 24278 13572 24330
rect 13644 24278 13696 24330
rect 13768 24278 13820 24330
rect 22396 24278 22448 24330
rect 22520 24278 22572 24330
rect 22644 24278 22696 24330
rect 22768 24278 22820 24330
rect 31396 24278 31448 24330
rect 31520 24278 31572 24330
rect 31644 24278 31696 24330
rect 31768 24278 31820 24330
rect 40396 24278 40448 24330
rect 40520 24278 40572 24330
rect 40644 24278 40696 24330
rect 40768 24278 40820 24330
rect 49396 24278 49448 24330
rect 49520 24278 49572 24330
rect 49644 24278 49696 24330
rect 49768 24278 49820 24330
rect 58396 24278 58448 24330
rect 58520 24278 58572 24330
rect 58644 24278 58696 24330
rect 58768 24278 58820 24330
rect 67396 24278 67448 24330
rect 67520 24278 67572 24330
rect 67644 24278 67696 24330
rect 67768 24278 67820 24330
rect 76396 24278 76448 24330
rect 76520 24278 76572 24330
rect 76644 24278 76696 24330
rect 76768 24278 76820 24330
rect 85396 24278 85448 24330
rect 85520 24278 85572 24330
rect 85644 24278 85696 24330
rect 85768 24278 85820 24330
rect 94396 24278 94448 24330
rect 94520 24278 94572 24330
rect 94644 24278 94696 24330
rect 94768 24278 94820 24330
rect 33854 24110 33906 24162
rect 34190 24110 34242 24162
rect 3614 23998 3666 24050
rect 11230 23998 11282 24050
rect 19630 23998 19682 24050
rect 20302 23998 20354 24050
rect 34750 23998 34802 24050
rect 59390 23998 59442 24050
rect 1710 23886 1762 23938
rect 10894 23886 10946 23938
rect 15822 23886 15874 23938
rect 16158 23886 16210 23938
rect 21534 23886 21586 23938
rect 22206 23886 22258 23938
rect 38894 23886 38946 23938
rect 39230 23886 39282 23938
rect 60510 23886 60562 23938
rect 61742 23886 61794 23938
rect 62190 23886 62242 23938
rect 71150 23886 71202 23938
rect 76302 23886 76354 23938
rect 2382 23774 2434 23826
rect 10446 23774 10498 23826
rect 21422 23774 21474 23826
rect 32622 23774 32674 23826
rect 33070 23774 33122 23826
rect 33518 23774 33570 23826
rect 59726 23774 59778 23826
rect 59838 23774 59890 23826
rect 61070 23774 61122 23826
rect 61182 23774 61234 23826
rect 2046 23662 2098 23714
rect 2718 23662 2770 23714
rect 3166 23662 3218 23714
rect 12462 23662 12514 23714
rect 18734 23662 18786 23714
rect 19294 23662 19346 23714
rect 20638 23662 20690 23714
rect 22542 23662 22594 23714
rect 23102 23662 23154 23714
rect 26910 23662 26962 23714
rect 32174 23662 32226 23714
rect 38446 23662 38498 23714
rect 41582 23662 41634 23714
rect 42366 23662 42418 23714
rect 60062 23662 60114 23714
rect 60622 23662 60674 23714
rect 60846 23662 60898 23714
rect 61406 23662 61458 23714
rect 64654 23662 64706 23714
rect 65214 23662 65266 23714
rect 65550 23662 65602 23714
rect 71486 23662 71538 23714
rect 76638 23662 76690 23714
rect 8896 23494 8948 23546
rect 9020 23494 9072 23546
rect 9144 23494 9196 23546
rect 9268 23494 9320 23546
rect 17896 23494 17948 23546
rect 18020 23494 18072 23546
rect 18144 23494 18196 23546
rect 18268 23494 18320 23546
rect 26896 23494 26948 23546
rect 27020 23494 27072 23546
rect 27144 23494 27196 23546
rect 27268 23494 27320 23546
rect 35896 23494 35948 23546
rect 36020 23494 36072 23546
rect 36144 23494 36196 23546
rect 36268 23494 36320 23546
rect 44896 23494 44948 23546
rect 45020 23494 45072 23546
rect 45144 23494 45196 23546
rect 45268 23494 45320 23546
rect 53896 23494 53948 23546
rect 54020 23494 54072 23546
rect 54144 23494 54196 23546
rect 54268 23494 54320 23546
rect 62896 23494 62948 23546
rect 63020 23494 63072 23546
rect 63144 23494 63196 23546
rect 63268 23494 63320 23546
rect 71896 23494 71948 23546
rect 72020 23494 72072 23546
rect 72144 23494 72196 23546
rect 72268 23494 72320 23546
rect 80896 23494 80948 23546
rect 81020 23494 81072 23546
rect 81144 23494 81196 23546
rect 81268 23494 81320 23546
rect 89896 23494 89948 23546
rect 90020 23494 90072 23546
rect 90144 23494 90196 23546
rect 90268 23494 90320 23546
rect 4734 23326 4786 23378
rect 6078 23326 6130 23378
rect 10110 23326 10162 23378
rect 26350 23326 26402 23378
rect 29486 23326 29538 23378
rect 30606 23326 30658 23378
rect 60286 23326 60338 23378
rect 60846 23326 60898 23378
rect 62302 23326 62354 23378
rect 62526 23326 62578 23378
rect 63310 23326 63362 23378
rect 65998 23326 66050 23378
rect 69806 23326 69858 23378
rect 73502 23326 73554 23378
rect 77422 23326 77474 23378
rect 77982 23326 78034 23378
rect 81006 23326 81058 23378
rect 82238 23326 82290 23378
rect 96574 23326 96626 23378
rect 5294 23214 5346 23266
rect 5630 23214 5682 23266
rect 10222 23214 10274 23266
rect 20302 23214 20354 23266
rect 23438 23214 23490 23266
rect 46062 23214 46114 23266
rect 66334 23214 66386 23266
rect 66670 23214 66722 23266
rect 72942 23214 72994 23266
rect 73726 23214 73778 23266
rect 74510 23214 74562 23266
rect 77758 23214 77810 23266
rect 78654 23214 78706 23266
rect 85710 23214 85762 23266
rect 1822 23102 1874 23154
rect 2270 23102 2322 23154
rect 10894 23102 10946 23154
rect 20638 23102 20690 23154
rect 21198 23102 21250 23154
rect 24222 23102 24274 23154
rect 26574 23102 26626 23154
rect 27134 23102 27186 23154
rect 45166 23102 45218 23154
rect 45950 23102 46002 23154
rect 46286 23102 46338 23154
rect 62974 23102 63026 23154
rect 67118 23102 67170 23154
rect 67566 23102 67618 23154
rect 74174 23102 74226 23154
rect 78430 23102 78482 23154
rect 82014 23102 82066 23154
rect 82126 23102 82178 23154
rect 82686 23102 82738 23154
rect 83022 23102 83074 23154
rect 83358 23102 83410 23154
rect 96910 23102 96962 23154
rect 45614 22990 45666 23042
rect 62414 22990 62466 23042
rect 73614 22990 73666 23042
rect 77870 22990 77922 23042
rect 81454 22990 81506 23042
rect 98030 22990 98082 23042
rect 30270 22878 30322 22930
rect 70590 22878 70642 22930
rect 86494 22878 86546 22930
rect 4396 22710 4448 22762
rect 4520 22710 4572 22762
rect 4644 22710 4696 22762
rect 4768 22710 4820 22762
rect 13396 22710 13448 22762
rect 13520 22710 13572 22762
rect 13644 22710 13696 22762
rect 13768 22710 13820 22762
rect 22396 22710 22448 22762
rect 22520 22710 22572 22762
rect 22644 22710 22696 22762
rect 22768 22710 22820 22762
rect 31396 22710 31448 22762
rect 31520 22710 31572 22762
rect 31644 22710 31696 22762
rect 31768 22710 31820 22762
rect 40396 22710 40448 22762
rect 40520 22710 40572 22762
rect 40644 22710 40696 22762
rect 40768 22710 40820 22762
rect 49396 22710 49448 22762
rect 49520 22710 49572 22762
rect 49644 22710 49696 22762
rect 49768 22710 49820 22762
rect 58396 22710 58448 22762
rect 58520 22710 58572 22762
rect 58644 22710 58696 22762
rect 58768 22710 58820 22762
rect 67396 22710 67448 22762
rect 67520 22710 67572 22762
rect 67644 22710 67696 22762
rect 67768 22710 67820 22762
rect 76396 22710 76448 22762
rect 76520 22710 76572 22762
rect 76644 22710 76696 22762
rect 76768 22710 76820 22762
rect 85396 22710 85448 22762
rect 85520 22710 85572 22762
rect 85644 22710 85696 22762
rect 85768 22710 85820 22762
rect 94396 22710 94448 22762
rect 94520 22710 94572 22762
rect 94644 22710 94696 22762
rect 94768 22710 94820 22762
rect 9214 22542 9266 22594
rect 65662 22542 65714 22594
rect 9550 22430 9602 22482
rect 38110 22430 38162 22482
rect 68462 22430 68514 22482
rect 69918 22430 69970 22482
rect 76302 22430 76354 22482
rect 77758 22430 77810 22482
rect 5630 22318 5682 22370
rect 6078 22318 6130 22370
rect 10894 22318 10946 22370
rect 21646 22318 21698 22370
rect 33630 22318 33682 22370
rect 38558 22318 38610 22370
rect 39342 22318 39394 22370
rect 64318 22318 64370 22370
rect 64654 22318 64706 22370
rect 68350 22318 68402 22370
rect 68574 22318 68626 22370
rect 68910 22318 68962 22370
rect 69134 22318 69186 22370
rect 72158 22318 72210 22370
rect 72718 22318 72770 22370
rect 78206 22318 78258 22370
rect 78542 22318 78594 22370
rect 82574 22318 82626 22370
rect 84926 22318 84978 22370
rect 1710 22206 1762 22258
rect 2382 22206 2434 22258
rect 8430 22206 8482 22258
rect 10782 22206 10834 22258
rect 21310 22206 21362 22258
rect 27806 22206 27858 22258
rect 28590 22206 28642 22258
rect 38670 22206 38722 22258
rect 67118 22206 67170 22258
rect 69358 22206 69410 22258
rect 69470 22206 69522 22258
rect 83134 22206 83186 22258
rect 84590 22206 84642 22258
rect 84814 22206 84866 22258
rect 2046 22094 2098 22146
rect 2942 22094 2994 22146
rect 11678 22094 11730 22146
rect 14590 22094 14642 22146
rect 14926 22094 14978 22146
rect 29150 22094 29202 22146
rect 29710 22094 29762 22146
rect 33854 22094 33906 22146
rect 34190 22094 34242 22146
rect 39678 22094 39730 22146
rect 40126 22094 40178 22146
rect 61854 22094 61906 22146
rect 70366 22094 70418 22146
rect 75070 22094 75122 22146
rect 75742 22094 75794 22146
rect 80894 22094 80946 22146
rect 81678 22094 81730 22146
rect 84366 22094 84418 22146
rect 8896 21926 8948 21978
rect 9020 21926 9072 21978
rect 9144 21926 9196 21978
rect 9268 21926 9320 21978
rect 17896 21926 17948 21978
rect 18020 21926 18072 21978
rect 18144 21926 18196 21978
rect 18268 21926 18320 21978
rect 26896 21926 26948 21978
rect 27020 21926 27072 21978
rect 27144 21926 27196 21978
rect 27268 21926 27320 21978
rect 35896 21926 35948 21978
rect 36020 21926 36072 21978
rect 36144 21926 36196 21978
rect 36268 21926 36320 21978
rect 44896 21926 44948 21978
rect 45020 21926 45072 21978
rect 45144 21926 45196 21978
rect 45268 21926 45320 21978
rect 53896 21926 53948 21978
rect 54020 21926 54072 21978
rect 54144 21926 54196 21978
rect 54268 21926 54320 21978
rect 62896 21926 62948 21978
rect 63020 21926 63072 21978
rect 63144 21926 63196 21978
rect 63268 21926 63320 21978
rect 71896 21926 71948 21978
rect 72020 21926 72072 21978
rect 72144 21926 72196 21978
rect 72268 21926 72320 21978
rect 80896 21926 80948 21978
rect 81020 21926 81072 21978
rect 81144 21926 81196 21978
rect 81268 21926 81320 21978
rect 89896 21926 89948 21978
rect 90020 21926 90072 21978
rect 90144 21926 90196 21978
rect 90268 21926 90320 21978
rect 8990 21758 9042 21810
rect 13022 21758 13074 21810
rect 31950 21758 32002 21810
rect 43374 21758 43426 21810
rect 43822 21758 43874 21810
rect 64318 21758 64370 21810
rect 74958 21758 75010 21810
rect 80222 21758 80274 21810
rect 96574 21758 96626 21810
rect 2046 21646 2098 21698
rect 9886 21646 9938 21698
rect 13806 21646 13858 21698
rect 14590 21646 14642 21698
rect 15150 21646 15202 21698
rect 15598 21646 15650 21698
rect 25230 21646 25282 21698
rect 36206 21646 36258 21698
rect 39342 21646 39394 21698
rect 64542 21646 64594 21698
rect 64654 21646 64706 21698
rect 65102 21646 65154 21698
rect 75182 21646 75234 21698
rect 80446 21646 80498 21698
rect 87054 21646 87106 21698
rect 87390 21646 87442 21698
rect 1710 21534 1762 21586
rect 6414 21534 6466 21586
rect 10110 21534 10162 21586
rect 10670 21534 10722 21586
rect 14366 21534 14418 21586
rect 16158 21534 16210 21586
rect 17838 21534 17890 21586
rect 27358 21534 27410 21586
rect 29038 21534 29090 21586
rect 29374 21534 29426 21586
rect 33406 21534 33458 21586
rect 33854 21534 33906 21586
rect 39118 21534 39170 21586
rect 43710 21534 43762 21586
rect 75294 21534 75346 21586
rect 80558 21534 80610 21586
rect 81006 21534 81058 21586
rect 96910 21534 96962 21586
rect 2494 21422 2546 21474
rect 6862 21422 6914 21474
rect 16830 21422 16882 21474
rect 17502 21422 17554 21474
rect 18734 21422 18786 21474
rect 26574 21422 26626 21474
rect 27022 21422 27074 21474
rect 28366 21422 28418 21474
rect 75742 21422 75794 21474
rect 98030 21422 98082 21474
rect 5854 21310 5906 21362
rect 15822 21310 15874 21362
rect 32510 21310 32562 21362
rect 36990 21310 37042 21362
rect 43822 21310 43874 21362
rect 4396 21142 4448 21194
rect 4520 21142 4572 21194
rect 4644 21142 4696 21194
rect 4768 21142 4820 21194
rect 13396 21142 13448 21194
rect 13520 21142 13572 21194
rect 13644 21142 13696 21194
rect 13768 21142 13820 21194
rect 22396 21142 22448 21194
rect 22520 21142 22572 21194
rect 22644 21142 22696 21194
rect 22768 21142 22820 21194
rect 31396 21142 31448 21194
rect 31520 21142 31572 21194
rect 31644 21142 31696 21194
rect 31768 21142 31820 21194
rect 40396 21142 40448 21194
rect 40520 21142 40572 21194
rect 40644 21142 40696 21194
rect 40768 21142 40820 21194
rect 49396 21142 49448 21194
rect 49520 21142 49572 21194
rect 49644 21142 49696 21194
rect 49768 21142 49820 21194
rect 58396 21142 58448 21194
rect 58520 21142 58572 21194
rect 58644 21142 58696 21194
rect 58768 21142 58820 21194
rect 67396 21142 67448 21194
rect 67520 21142 67572 21194
rect 67644 21142 67696 21194
rect 67768 21142 67820 21194
rect 76396 21142 76448 21194
rect 76520 21142 76572 21194
rect 76644 21142 76696 21194
rect 76768 21142 76820 21194
rect 85396 21142 85448 21194
rect 85520 21142 85572 21194
rect 85644 21142 85696 21194
rect 85768 21142 85820 21194
rect 94396 21142 94448 21194
rect 94520 21142 94572 21194
rect 94644 21142 94696 21194
rect 94768 21142 94820 21194
rect 9886 20974 9938 21026
rect 30158 20974 30210 21026
rect 34750 20974 34802 21026
rect 42926 20974 42978 21026
rect 65214 20974 65266 21026
rect 74846 20974 74898 21026
rect 4286 20862 4338 20914
rect 18398 20862 18450 20914
rect 18734 20862 18786 20914
rect 32622 20862 32674 20914
rect 33070 20862 33122 20914
rect 39006 20862 39058 20914
rect 43486 20862 43538 20914
rect 55470 20862 55522 20914
rect 56702 20862 56754 20914
rect 65550 20862 65602 20914
rect 73726 20862 73778 20914
rect 80670 20862 80722 20914
rect 84366 20862 84418 20914
rect 4622 20750 4674 20802
rect 6190 20750 6242 20802
rect 6750 20750 6802 20802
rect 14926 20750 14978 20802
rect 15262 20750 15314 20802
rect 22990 20750 23042 20802
rect 24222 20750 24274 20802
rect 25118 20750 25170 20802
rect 25566 20750 25618 20802
rect 28590 20750 28642 20802
rect 29150 20750 29202 20802
rect 33742 20750 33794 20802
rect 34414 20750 34466 20802
rect 39230 20750 39282 20802
rect 39790 20750 39842 20802
rect 43822 20750 43874 20802
rect 56030 20750 56082 20802
rect 56366 20750 56418 20802
rect 61742 20750 61794 20802
rect 62190 20750 62242 20802
rect 72046 20750 72098 20802
rect 72718 20750 72770 20802
rect 74174 20750 74226 20802
rect 84926 20750 84978 20802
rect 85598 20750 85650 20802
rect 5070 20638 5122 20690
rect 5966 20638 6018 20690
rect 9102 20638 9154 20690
rect 23438 20638 23490 20690
rect 23998 20638 24050 20690
rect 27806 20638 27858 20690
rect 33630 20638 33682 20690
rect 42142 20638 42194 20690
rect 43934 20638 43986 20690
rect 56142 20638 56194 20690
rect 1934 20526 1986 20578
rect 17838 20526 17890 20578
rect 19070 20526 19122 20578
rect 24558 20526 24610 20578
rect 44158 20526 44210 20578
rect 64654 20526 64706 20578
rect 72158 20526 72210 20578
rect 72270 20526 72322 20578
rect 73054 20526 73106 20578
rect 76302 20526 76354 20578
rect 85038 20526 85090 20578
rect 85150 20526 85202 20578
rect 8896 20358 8948 20410
rect 9020 20358 9072 20410
rect 9144 20358 9196 20410
rect 9268 20358 9320 20410
rect 17896 20358 17948 20410
rect 18020 20358 18072 20410
rect 18144 20358 18196 20410
rect 18268 20358 18320 20410
rect 26896 20358 26948 20410
rect 27020 20358 27072 20410
rect 27144 20358 27196 20410
rect 27268 20358 27320 20410
rect 35896 20358 35948 20410
rect 36020 20358 36072 20410
rect 36144 20358 36196 20410
rect 36268 20358 36320 20410
rect 44896 20358 44948 20410
rect 45020 20358 45072 20410
rect 45144 20358 45196 20410
rect 45268 20358 45320 20410
rect 53896 20358 53948 20410
rect 54020 20358 54072 20410
rect 54144 20358 54196 20410
rect 54268 20358 54320 20410
rect 62896 20358 62948 20410
rect 63020 20358 63072 20410
rect 63144 20358 63196 20410
rect 63268 20358 63320 20410
rect 71896 20358 71948 20410
rect 72020 20358 72072 20410
rect 72144 20358 72196 20410
rect 72268 20358 72320 20410
rect 80896 20358 80948 20410
rect 81020 20358 81072 20410
rect 81144 20358 81196 20410
rect 81268 20358 81320 20410
rect 89896 20358 89948 20410
rect 90020 20358 90072 20410
rect 90144 20358 90196 20410
rect 90268 20358 90320 20410
rect 18174 20190 18226 20242
rect 21758 20190 21810 20242
rect 25566 20190 25618 20242
rect 28926 20190 28978 20242
rect 73166 20190 73218 20242
rect 75518 20190 75570 20242
rect 76302 20190 76354 20242
rect 81230 20190 81282 20242
rect 81902 20190 81954 20242
rect 86046 20190 86098 20242
rect 4510 20078 4562 20130
rect 5294 20078 5346 20130
rect 22430 20078 22482 20130
rect 28478 20078 28530 20130
rect 29374 20078 29426 20130
rect 39902 20078 39954 20130
rect 40126 20078 40178 20130
rect 40238 20078 40290 20130
rect 65886 20078 65938 20130
rect 66222 20078 66274 20130
rect 71038 20078 71090 20130
rect 73390 20078 73442 20130
rect 73502 20078 73554 20130
rect 75070 20078 75122 20130
rect 75966 20078 76018 20130
rect 78094 20078 78146 20130
rect 78206 20078 78258 20130
rect 78766 20078 78818 20130
rect 82910 20078 82962 20130
rect 83246 20078 83298 20130
rect 83358 20078 83410 20130
rect 85598 20078 85650 20130
rect 85822 20078 85874 20130
rect 1822 19966 1874 20018
rect 2158 19966 2210 20018
rect 5742 19966 5794 20018
rect 18958 19966 19010 20018
rect 19294 19966 19346 20018
rect 25342 19966 25394 20018
rect 40462 19966 40514 20018
rect 76526 19966 76578 20018
rect 76974 19966 77026 20018
rect 81006 19966 81058 20018
rect 81678 19966 81730 20018
rect 83022 19966 83074 20018
rect 85486 19966 85538 20018
rect 6078 19854 6130 19906
rect 7310 19854 7362 19906
rect 18510 19854 18562 19906
rect 73054 19854 73106 19906
rect 76414 19854 76466 19906
rect 77422 19854 77474 19906
rect 80446 19854 80498 19906
rect 81118 19854 81170 19906
rect 84702 19854 84754 19906
rect 85262 19854 85314 19906
rect 74510 19742 74562 19794
rect 78094 19742 78146 19794
rect 4396 19574 4448 19626
rect 4520 19574 4572 19626
rect 4644 19574 4696 19626
rect 4768 19574 4820 19626
rect 13396 19574 13448 19626
rect 13520 19574 13572 19626
rect 13644 19574 13696 19626
rect 13768 19574 13820 19626
rect 22396 19574 22448 19626
rect 22520 19574 22572 19626
rect 22644 19574 22696 19626
rect 22768 19574 22820 19626
rect 31396 19574 31448 19626
rect 31520 19574 31572 19626
rect 31644 19574 31696 19626
rect 31768 19574 31820 19626
rect 40396 19574 40448 19626
rect 40520 19574 40572 19626
rect 40644 19574 40696 19626
rect 40768 19574 40820 19626
rect 49396 19574 49448 19626
rect 49520 19574 49572 19626
rect 49644 19574 49696 19626
rect 49768 19574 49820 19626
rect 58396 19574 58448 19626
rect 58520 19574 58572 19626
rect 58644 19574 58696 19626
rect 58768 19574 58820 19626
rect 67396 19574 67448 19626
rect 67520 19574 67572 19626
rect 67644 19574 67696 19626
rect 67768 19574 67820 19626
rect 76396 19574 76448 19626
rect 76520 19574 76572 19626
rect 76644 19574 76696 19626
rect 76768 19574 76820 19626
rect 85396 19574 85448 19626
rect 85520 19574 85572 19626
rect 85644 19574 85696 19626
rect 85768 19574 85820 19626
rect 94396 19574 94448 19626
rect 94520 19574 94572 19626
rect 94644 19574 94696 19626
rect 94768 19574 94820 19626
rect 74398 19406 74450 19458
rect 79774 19406 79826 19458
rect 89070 19406 89122 19458
rect 3166 19294 3218 19346
rect 6078 19294 6130 19346
rect 6526 19294 6578 19346
rect 74734 19294 74786 19346
rect 75630 19294 75682 19346
rect 1710 19182 1762 19234
rect 40014 19182 40066 19234
rect 44270 19182 44322 19234
rect 70926 19182 70978 19234
rect 71374 19182 71426 19234
rect 76078 19182 76130 19234
rect 76638 19182 76690 19234
rect 80110 19182 80162 19234
rect 80558 19182 80610 19234
rect 85598 19182 85650 19234
rect 86046 19182 86098 19234
rect 96910 19182 96962 19234
rect 2382 19070 2434 19122
rect 2718 19070 2770 19122
rect 42030 19070 42082 19122
rect 96686 19070 96738 19122
rect 98030 19070 98082 19122
rect 2046 18958 2098 19010
rect 73838 18958 73890 19010
rect 79214 18958 79266 19010
rect 82798 18958 82850 19010
rect 83582 18958 83634 19010
rect 85150 18958 85202 19010
rect 88286 18958 88338 19010
rect 8896 18790 8948 18842
rect 9020 18790 9072 18842
rect 9144 18790 9196 18842
rect 9268 18790 9320 18842
rect 17896 18790 17948 18842
rect 18020 18790 18072 18842
rect 18144 18790 18196 18842
rect 18268 18790 18320 18842
rect 26896 18790 26948 18842
rect 27020 18790 27072 18842
rect 27144 18790 27196 18842
rect 27268 18790 27320 18842
rect 35896 18790 35948 18842
rect 36020 18790 36072 18842
rect 36144 18790 36196 18842
rect 36268 18790 36320 18842
rect 44896 18790 44948 18842
rect 45020 18790 45072 18842
rect 45144 18790 45196 18842
rect 45268 18790 45320 18842
rect 53896 18790 53948 18842
rect 54020 18790 54072 18842
rect 54144 18790 54196 18842
rect 54268 18790 54320 18842
rect 62896 18790 62948 18842
rect 63020 18790 63072 18842
rect 63144 18790 63196 18842
rect 63268 18790 63320 18842
rect 71896 18790 71948 18842
rect 72020 18790 72072 18842
rect 72144 18790 72196 18842
rect 72268 18790 72320 18842
rect 80896 18790 80948 18842
rect 81020 18790 81072 18842
rect 81144 18790 81196 18842
rect 81268 18790 81320 18842
rect 89896 18790 89948 18842
rect 90020 18790 90072 18842
rect 90144 18790 90196 18842
rect 90268 18790 90320 18842
rect 79662 18622 79714 18674
rect 75182 18510 75234 18562
rect 75518 18510 75570 18562
rect 80222 18510 80274 18562
rect 80558 18510 80610 18562
rect 89966 18510 90018 18562
rect 90302 18510 90354 18562
rect 2158 18398 2210 18450
rect 4396 18006 4448 18058
rect 4520 18006 4572 18058
rect 4644 18006 4696 18058
rect 4768 18006 4820 18058
rect 13396 18006 13448 18058
rect 13520 18006 13572 18058
rect 13644 18006 13696 18058
rect 13768 18006 13820 18058
rect 22396 18006 22448 18058
rect 22520 18006 22572 18058
rect 22644 18006 22696 18058
rect 22768 18006 22820 18058
rect 31396 18006 31448 18058
rect 31520 18006 31572 18058
rect 31644 18006 31696 18058
rect 31768 18006 31820 18058
rect 40396 18006 40448 18058
rect 40520 18006 40572 18058
rect 40644 18006 40696 18058
rect 40768 18006 40820 18058
rect 49396 18006 49448 18058
rect 49520 18006 49572 18058
rect 49644 18006 49696 18058
rect 49768 18006 49820 18058
rect 58396 18006 58448 18058
rect 58520 18006 58572 18058
rect 58644 18006 58696 18058
rect 58768 18006 58820 18058
rect 67396 18006 67448 18058
rect 67520 18006 67572 18058
rect 67644 18006 67696 18058
rect 67768 18006 67820 18058
rect 76396 18006 76448 18058
rect 76520 18006 76572 18058
rect 76644 18006 76696 18058
rect 76768 18006 76820 18058
rect 85396 18006 85448 18058
rect 85520 18006 85572 18058
rect 85644 18006 85696 18058
rect 85768 18006 85820 18058
rect 94396 18006 94448 18058
rect 94520 18006 94572 18058
rect 94644 18006 94696 18058
rect 94768 18006 94820 18058
rect 85710 17614 85762 17666
rect 96910 17614 96962 17666
rect 1710 17502 1762 17554
rect 2046 17502 2098 17554
rect 2494 17502 2546 17554
rect 98030 17502 98082 17554
rect 86046 17390 86098 17442
rect 96686 17390 96738 17442
rect 8896 17222 8948 17274
rect 9020 17222 9072 17274
rect 9144 17222 9196 17274
rect 9268 17222 9320 17274
rect 17896 17222 17948 17274
rect 18020 17222 18072 17274
rect 18144 17222 18196 17274
rect 18268 17222 18320 17274
rect 26896 17222 26948 17274
rect 27020 17222 27072 17274
rect 27144 17222 27196 17274
rect 27268 17222 27320 17274
rect 35896 17222 35948 17274
rect 36020 17222 36072 17274
rect 36144 17222 36196 17274
rect 36268 17222 36320 17274
rect 44896 17222 44948 17274
rect 45020 17222 45072 17274
rect 45144 17222 45196 17274
rect 45268 17222 45320 17274
rect 53896 17222 53948 17274
rect 54020 17222 54072 17274
rect 54144 17222 54196 17274
rect 54268 17222 54320 17274
rect 62896 17222 62948 17274
rect 63020 17222 63072 17274
rect 63144 17222 63196 17274
rect 63268 17222 63320 17274
rect 71896 17222 71948 17274
rect 72020 17222 72072 17274
rect 72144 17222 72196 17274
rect 72268 17222 72320 17274
rect 80896 17222 80948 17274
rect 81020 17222 81072 17274
rect 81144 17222 81196 17274
rect 81268 17222 81320 17274
rect 89896 17222 89948 17274
rect 90020 17222 90072 17274
rect 90144 17222 90196 17274
rect 90268 17222 90320 17274
rect 2046 17054 2098 17106
rect 1710 16830 1762 16882
rect 2494 16830 2546 16882
rect 4396 16438 4448 16490
rect 4520 16438 4572 16490
rect 4644 16438 4696 16490
rect 4768 16438 4820 16490
rect 13396 16438 13448 16490
rect 13520 16438 13572 16490
rect 13644 16438 13696 16490
rect 13768 16438 13820 16490
rect 22396 16438 22448 16490
rect 22520 16438 22572 16490
rect 22644 16438 22696 16490
rect 22768 16438 22820 16490
rect 31396 16438 31448 16490
rect 31520 16438 31572 16490
rect 31644 16438 31696 16490
rect 31768 16438 31820 16490
rect 40396 16438 40448 16490
rect 40520 16438 40572 16490
rect 40644 16438 40696 16490
rect 40768 16438 40820 16490
rect 49396 16438 49448 16490
rect 49520 16438 49572 16490
rect 49644 16438 49696 16490
rect 49768 16438 49820 16490
rect 58396 16438 58448 16490
rect 58520 16438 58572 16490
rect 58644 16438 58696 16490
rect 58768 16438 58820 16490
rect 67396 16438 67448 16490
rect 67520 16438 67572 16490
rect 67644 16438 67696 16490
rect 67768 16438 67820 16490
rect 76396 16438 76448 16490
rect 76520 16438 76572 16490
rect 76644 16438 76696 16490
rect 76768 16438 76820 16490
rect 85396 16438 85448 16490
rect 85520 16438 85572 16490
rect 85644 16438 85696 16490
rect 85768 16438 85820 16490
rect 94396 16438 94448 16490
rect 94520 16438 94572 16490
rect 94644 16438 94696 16490
rect 94768 16438 94820 16490
rect 96686 16046 96738 16098
rect 96910 16046 96962 16098
rect 98030 15934 98082 15986
rect 8896 15654 8948 15706
rect 9020 15654 9072 15706
rect 9144 15654 9196 15706
rect 9268 15654 9320 15706
rect 17896 15654 17948 15706
rect 18020 15654 18072 15706
rect 18144 15654 18196 15706
rect 18268 15654 18320 15706
rect 26896 15654 26948 15706
rect 27020 15654 27072 15706
rect 27144 15654 27196 15706
rect 27268 15654 27320 15706
rect 35896 15654 35948 15706
rect 36020 15654 36072 15706
rect 36144 15654 36196 15706
rect 36268 15654 36320 15706
rect 44896 15654 44948 15706
rect 45020 15654 45072 15706
rect 45144 15654 45196 15706
rect 45268 15654 45320 15706
rect 53896 15654 53948 15706
rect 54020 15654 54072 15706
rect 54144 15654 54196 15706
rect 54268 15654 54320 15706
rect 62896 15654 62948 15706
rect 63020 15654 63072 15706
rect 63144 15654 63196 15706
rect 63268 15654 63320 15706
rect 71896 15654 71948 15706
rect 72020 15654 72072 15706
rect 72144 15654 72196 15706
rect 72268 15654 72320 15706
rect 80896 15654 80948 15706
rect 81020 15654 81072 15706
rect 81144 15654 81196 15706
rect 81268 15654 81320 15706
rect 89896 15654 89948 15706
rect 90020 15654 90072 15706
rect 90144 15654 90196 15706
rect 90268 15654 90320 15706
rect 42254 15374 42306 15426
rect 44606 15374 44658 15426
rect 41694 15262 41746 15314
rect 43038 15262 43090 15314
rect 44830 15262 44882 15314
rect 41134 15150 41186 15202
rect 43934 15150 43986 15202
rect 79662 15150 79714 15202
rect 80334 15150 80386 15202
rect 82798 15150 82850 15202
rect 4396 14870 4448 14922
rect 4520 14870 4572 14922
rect 4644 14870 4696 14922
rect 4768 14870 4820 14922
rect 13396 14870 13448 14922
rect 13520 14870 13572 14922
rect 13644 14870 13696 14922
rect 13768 14870 13820 14922
rect 22396 14870 22448 14922
rect 22520 14870 22572 14922
rect 22644 14870 22696 14922
rect 22768 14870 22820 14922
rect 31396 14870 31448 14922
rect 31520 14870 31572 14922
rect 31644 14870 31696 14922
rect 31768 14870 31820 14922
rect 40396 14870 40448 14922
rect 40520 14870 40572 14922
rect 40644 14870 40696 14922
rect 40768 14870 40820 14922
rect 49396 14870 49448 14922
rect 49520 14870 49572 14922
rect 49644 14870 49696 14922
rect 49768 14870 49820 14922
rect 58396 14870 58448 14922
rect 58520 14870 58572 14922
rect 58644 14870 58696 14922
rect 58768 14870 58820 14922
rect 67396 14870 67448 14922
rect 67520 14870 67572 14922
rect 67644 14870 67696 14922
rect 67768 14870 67820 14922
rect 76396 14870 76448 14922
rect 76520 14870 76572 14922
rect 76644 14870 76696 14922
rect 76768 14870 76820 14922
rect 85396 14870 85448 14922
rect 85520 14870 85572 14922
rect 85644 14870 85696 14922
rect 85768 14870 85820 14922
rect 94396 14870 94448 14922
rect 94520 14870 94572 14922
rect 94644 14870 94696 14922
rect 94768 14870 94820 14922
rect 46622 14590 46674 14642
rect 21422 14478 21474 14530
rect 44942 14478 44994 14530
rect 45390 14478 45442 14530
rect 46734 14478 46786 14530
rect 47070 14478 47122 14530
rect 70030 14478 70082 14530
rect 71710 14478 71762 14530
rect 74174 14478 74226 14530
rect 78430 14478 78482 14530
rect 80558 14478 80610 14530
rect 81902 14478 81954 14530
rect 82798 14478 82850 14530
rect 96910 14478 96962 14530
rect 70590 14366 70642 14418
rect 74174 14366 74226 14418
rect 78318 14366 78370 14418
rect 81678 14366 81730 14418
rect 83134 14366 83186 14418
rect 98030 14366 98082 14418
rect 20750 14254 20802 14306
rect 27694 14254 27746 14306
rect 44270 14254 44322 14306
rect 73950 14254 74002 14306
rect 74622 14254 74674 14306
rect 75070 14254 75122 14306
rect 82238 14254 82290 14306
rect 8896 14086 8948 14138
rect 9020 14086 9072 14138
rect 9144 14086 9196 14138
rect 9268 14086 9320 14138
rect 17896 14086 17948 14138
rect 18020 14086 18072 14138
rect 18144 14086 18196 14138
rect 18268 14086 18320 14138
rect 26896 14086 26948 14138
rect 27020 14086 27072 14138
rect 27144 14086 27196 14138
rect 27268 14086 27320 14138
rect 35896 14086 35948 14138
rect 36020 14086 36072 14138
rect 36144 14086 36196 14138
rect 36268 14086 36320 14138
rect 44896 14086 44948 14138
rect 45020 14086 45072 14138
rect 45144 14086 45196 14138
rect 45268 14086 45320 14138
rect 53896 14086 53948 14138
rect 54020 14086 54072 14138
rect 54144 14086 54196 14138
rect 54268 14086 54320 14138
rect 62896 14086 62948 14138
rect 63020 14086 63072 14138
rect 63144 14086 63196 14138
rect 63268 14086 63320 14138
rect 71896 14086 71948 14138
rect 72020 14086 72072 14138
rect 72144 14086 72196 14138
rect 72268 14086 72320 14138
rect 80896 14086 80948 14138
rect 81020 14086 81072 14138
rect 81144 14086 81196 14138
rect 81268 14086 81320 14138
rect 89896 14086 89948 14138
rect 90020 14086 90072 14138
rect 90144 14086 90196 14138
rect 90268 14086 90320 14138
rect 2046 13918 2098 13970
rect 55582 13918 55634 13970
rect 55134 13806 55186 13858
rect 59054 13806 59106 13858
rect 61854 13806 61906 13858
rect 72270 13806 72322 13858
rect 72606 13806 72658 13858
rect 80222 13806 80274 13858
rect 1710 13694 1762 13746
rect 34862 13694 34914 13746
rect 43150 13694 43202 13746
rect 51662 13694 51714 13746
rect 52110 13694 52162 13746
rect 53006 13694 53058 13746
rect 53454 13694 53506 13746
rect 54574 13694 54626 13746
rect 58830 13694 58882 13746
rect 60510 13694 60562 13746
rect 61966 13694 62018 13746
rect 74062 13694 74114 13746
rect 75518 13694 75570 13746
rect 76974 13694 77026 13746
rect 77310 13694 77362 13746
rect 77982 13694 78034 13746
rect 80110 13694 80162 13746
rect 81790 13694 81842 13746
rect 82798 13694 82850 13746
rect 83582 13694 83634 13746
rect 2494 13582 2546 13634
rect 37214 13582 37266 13634
rect 44270 13582 44322 13634
rect 51214 13582 51266 13634
rect 52334 13582 52386 13634
rect 61070 13582 61122 13634
rect 75406 13582 75458 13634
rect 78878 13582 78930 13634
rect 79326 13582 79378 13634
rect 82686 13582 82738 13634
rect 4396 13302 4448 13354
rect 4520 13302 4572 13354
rect 4644 13302 4696 13354
rect 4768 13302 4820 13354
rect 13396 13302 13448 13354
rect 13520 13302 13572 13354
rect 13644 13302 13696 13354
rect 13768 13302 13820 13354
rect 22396 13302 22448 13354
rect 22520 13302 22572 13354
rect 22644 13302 22696 13354
rect 22768 13302 22820 13354
rect 31396 13302 31448 13354
rect 31520 13302 31572 13354
rect 31644 13302 31696 13354
rect 31768 13302 31820 13354
rect 40396 13302 40448 13354
rect 40520 13302 40572 13354
rect 40644 13302 40696 13354
rect 40768 13302 40820 13354
rect 49396 13302 49448 13354
rect 49520 13302 49572 13354
rect 49644 13302 49696 13354
rect 49768 13302 49820 13354
rect 58396 13302 58448 13354
rect 58520 13302 58572 13354
rect 58644 13302 58696 13354
rect 58768 13302 58820 13354
rect 67396 13302 67448 13354
rect 67520 13302 67572 13354
rect 67644 13302 67696 13354
rect 67768 13302 67820 13354
rect 76396 13302 76448 13354
rect 76520 13302 76572 13354
rect 76644 13302 76696 13354
rect 76768 13302 76820 13354
rect 85396 13302 85448 13354
rect 85520 13302 85572 13354
rect 85644 13302 85696 13354
rect 85768 13302 85820 13354
rect 94396 13302 94448 13354
rect 94520 13302 94572 13354
rect 94644 13302 94696 13354
rect 94768 13302 94820 13354
rect 45390 13022 45442 13074
rect 80446 13022 80498 13074
rect 37214 12910 37266 12962
rect 46958 12910 47010 12962
rect 48078 12910 48130 12962
rect 50094 12910 50146 12962
rect 66110 12910 66162 12962
rect 73838 12910 73890 12962
rect 82238 12910 82290 12962
rect 41470 12798 41522 12850
rect 47182 12798 47234 12850
rect 49534 12798 49586 12850
rect 61070 12798 61122 12850
rect 69694 12798 69746 12850
rect 47854 12686 47906 12738
rect 50878 12686 50930 12738
rect 51326 12686 51378 12738
rect 66558 12686 66610 12738
rect 74286 12686 74338 12738
rect 8896 12518 8948 12570
rect 9020 12518 9072 12570
rect 9144 12518 9196 12570
rect 9268 12518 9320 12570
rect 17896 12518 17948 12570
rect 18020 12518 18072 12570
rect 18144 12518 18196 12570
rect 18268 12518 18320 12570
rect 26896 12518 26948 12570
rect 27020 12518 27072 12570
rect 27144 12518 27196 12570
rect 27268 12518 27320 12570
rect 35896 12518 35948 12570
rect 36020 12518 36072 12570
rect 36144 12518 36196 12570
rect 36268 12518 36320 12570
rect 44896 12518 44948 12570
rect 45020 12518 45072 12570
rect 45144 12518 45196 12570
rect 45268 12518 45320 12570
rect 53896 12518 53948 12570
rect 54020 12518 54072 12570
rect 54144 12518 54196 12570
rect 54268 12518 54320 12570
rect 62896 12518 62948 12570
rect 63020 12518 63072 12570
rect 63144 12518 63196 12570
rect 63268 12518 63320 12570
rect 71896 12518 71948 12570
rect 72020 12518 72072 12570
rect 72144 12518 72196 12570
rect 72268 12518 72320 12570
rect 80896 12518 80948 12570
rect 81020 12518 81072 12570
rect 81144 12518 81196 12570
rect 81268 12518 81320 12570
rect 89896 12518 89948 12570
rect 90020 12518 90072 12570
rect 90144 12518 90196 12570
rect 90268 12518 90320 12570
rect 2046 12238 2098 12290
rect 48862 12238 48914 12290
rect 52782 12238 52834 12290
rect 60398 12238 60450 12290
rect 68462 12238 68514 12290
rect 71710 12238 71762 12290
rect 96574 12238 96626 12290
rect 1710 12126 1762 12178
rect 40014 12126 40066 12178
rect 42702 12126 42754 12178
rect 48750 12126 48802 12178
rect 51102 12126 51154 12178
rect 52446 12126 52498 12178
rect 63758 12126 63810 12178
rect 67902 12126 67954 12178
rect 69694 12126 69746 12178
rect 71486 12126 71538 12178
rect 76078 12126 76130 12178
rect 80110 12126 80162 12178
rect 81342 12126 81394 12178
rect 82574 12126 82626 12178
rect 83470 12126 83522 12178
rect 96910 12126 96962 12178
rect 2494 12014 2546 12066
rect 36878 12014 36930 12066
rect 44382 12014 44434 12066
rect 48190 12014 48242 12066
rect 51326 12014 51378 12066
rect 70142 12014 70194 12066
rect 72494 12014 72546 12066
rect 78878 12014 78930 12066
rect 79326 12014 79378 12066
rect 83806 12014 83858 12066
rect 98030 12014 98082 12066
rect 83918 11902 83970 11954
rect 4396 11734 4448 11786
rect 4520 11734 4572 11786
rect 4644 11734 4696 11786
rect 4768 11734 4820 11786
rect 13396 11734 13448 11786
rect 13520 11734 13572 11786
rect 13644 11734 13696 11786
rect 13768 11734 13820 11786
rect 22396 11734 22448 11786
rect 22520 11734 22572 11786
rect 22644 11734 22696 11786
rect 22768 11734 22820 11786
rect 31396 11734 31448 11786
rect 31520 11734 31572 11786
rect 31644 11734 31696 11786
rect 31768 11734 31820 11786
rect 40396 11734 40448 11786
rect 40520 11734 40572 11786
rect 40644 11734 40696 11786
rect 40768 11734 40820 11786
rect 49396 11734 49448 11786
rect 49520 11734 49572 11786
rect 49644 11734 49696 11786
rect 49768 11734 49820 11786
rect 58396 11734 58448 11786
rect 58520 11734 58572 11786
rect 58644 11734 58696 11786
rect 58768 11734 58820 11786
rect 67396 11734 67448 11786
rect 67520 11734 67572 11786
rect 67644 11734 67696 11786
rect 67768 11734 67820 11786
rect 76396 11734 76448 11786
rect 76520 11734 76572 11786
rect 76644 11734 76696 11786
rect 76768 11734 76820 11786
rect 85396 11734 85448 11786
rect 85520 11734 85572 11786
rect 85644 11734 85696 11786
rect 85768 11734 85820 11786
rect 94396 11734 94448 11786
rect 94520 11734 94572 11786
rect 94644 11734 94696 11786
rect 94768 11734 94820 11786
rect 67566 11566 67618 11618
rect 62190 11454 62242 11506
rect 71150 11454 71202 11506
rect 31166 11342 31218 11394
rect 39006 11342 39058 11394
rect 46398 11342 46450 11394
rect 56142 11342 56194 11394
rect 58158 11342 58210 11394
rect 59390 11342 59442 11394
rect 63646 11342 63698 11394
rect 73614 11342 73666 11394
rect 81902 11342 81954 11394
rect 1710 11230 1762 11282
rect 33966 11230 34018 11282
rect 41022 11230 41074 11282
rect 47070 11230 47122 11282
rect 56702 11230 56754 11282
rect 58046 11230 58098 11282
rect 59166 11230 59218 11282
rect 2046 11118 2098 11170
rect 2494 11118 2546 11170
rect 60622 11118 60674 11170
rect 61070 11118 61122 11170
rect 78206 11118 78258 11170
rect 8896 10950 8948 11002
rect 9020 10950 9072 11002
rect 9144 10950 9196 11002
rect 9268 10950 9320 11002
rect 17896 10950 17948 11002
rect 18020 10950 18072 11002
rect 18144 10950 18196 11002
rect 18268 10950 18320 11002
rect 26896 10950 26948 11002
rect 27020 10950 27072 11002
rect 27144 10950 27196 11002
rect 27268 10950 27320 11002
rect 35896 10950 35948 11002
rect 36020 10950 36072 11002
rect 36144 10950 36196 11002
rect 36268 10950 36320 11002
rect 44896 10950 44948 11002
rect 45020 10950 45072 11002
rect 45144 10950 45196 11002
rect 45268 10950 45320 11002
rect 53896 10950 53948 11002
rect 54020 10950 54072 11002
rect 54144 10950 54196 11002
rect 54268 10950 54320 11002
rect 62896 10950 62948 11002
rect 63020 10950 63072 11002
rect 63144 10950 63196 11002
rect 63268 10950 63320 11002
rect 71896 10950 71948 11002
rect 72020 10950 72072 11002
rect 72144 10950 72196 11002
rect 72268 10950 72320 11002
rect 80896 10950 80948 11002
rect 81020 10950 81072 11002
rect 81144 10950 81196 11002
rect 81268 10950 81320 11002
rect 89896 10950 89948 11002
rect 90020 10950 90072 11002
rect 90144 10950 90196 11002
rect 90268 10950 90320 11002
rect 65550 10782 65602 10834
rect 76078 10670 76130 10722
rect 77870 10670 77922 10722
rect 78206 10670 78258 10722
rect 96686 10670 96738 10722
rect 35310 10558 35362 10610
rect 47182 10558 47234 10610
rect 53230 10558 53282 10610
rect 59950 10558 60002 10610
rect 69694 10558 69746 10610
rect 72606 10558 72658 10610
rect 81566 10558 81618 10610
rect 96910 10558 96962 10610
rect 38110 10446 38162 10498
rect 43710 10446 43762 10498
rect 50430 10446 50482 10498
rect 63534 10446 63586 10498
rect 85150 10446 85202 10498
rect 98030 10446 98082 10498
rect 4396 10166 4448 10218
rect 4520 10166 4572 10218
rect 4644 10166 4696 10218
rect 4768 10166 4820 10218
rect 13396 10166 13448 10218
rect 13520 10166 13572 10218
rect 13644 10166 13696 10218
rect 13768 10166 13820 10218
rect 22396 10166 22448 10218
rect 22520 10166 22572 10218
rect 22644 10166 22696 10218
rect 22768 10166 22820 10218
rect 31396 10166 31448 10218
rect 31520 10166 31572 10218
rect 31644 10166 31696 10218
rect 31768 10166 31820 10218
rect 40396 10166 40448 10218
rect 40520 10166 40572 10218
rect 40644 10166 40696 10218
rect 40768 10166 40820 10218
rect 49396 10166 49448 10218
rect 49520 10166 49572 10218
rect 49644 10166 49696 10218
rect 49768 10166 49820 10218
rect 58396 10166 58448 10218
rect 58520 10166 58572 10218
rect 58644 10166 58696 10218
rect 58768 10166 58820 10218
rect 67396 10166 67448 10218
rect 67520 10166 67572 10218
rect 67644 10166 67696 10218
rect 67768 10166 67820 10218
rect 76396 10166 76448 10218
rect 76520 10166 76572 10218
rect 76644 10166 76696 10218
rect 76768 10166 76820 10218
rect 85396 10166 85448 10218
rect 85520 10166 85572 10218
rect 85644 10166 85696 10218
rect 85768 10166 85820 10218
rect 94396 10166 94448 10218
rect 94520 10166 94572 10218
rect 94644 10166 94696 10218
rect 94768 10166 94820 10218
rect 45054 9886 45106 9938
rect 46062 9886 46114 9938
rect 54686 9886 54738 9938
rect 35422 9774 35474 9826
rect 39006 9774 39058 9826
rect 47070 9774 47122 9826
rect 52782 9774 52834 9826
rect 64318 9774 64370 9826
rect 75070 9774 75122 9826
rect 81454 9774 81506 9826
rect 88958 9774 89010 9826
rect 1710 9662 1762 9714
rect 2494 9662 2546 9714
rect 31950 9662 32002 9714
rect 41022 9662 41074 9714
rect 48974 9662 49026 9714
rect 62414 9662 62466 9714
rect 70702 9662 70754 9714
rect 77310 9662 77362 9714
rect 84366 9662 84418 9714
rect 2046 9550 2098 9602
rect 45166 9550 45218 9602
rect 45950 9550 46002 9602
rect 8896 9382 8948 9434
rect 9020 9382 9072 9434
rect 9144 9382 9196 9434
rect 9268 9382 9320 9434
rect 17896 9382 17948 9434
rect 18020 9382 18072 9434
rect 18144 9382 18196 9434
rect 18268 9382 18320 9434
rect 26896 9382 26948 9434
rect 27020 9382 27072 9434
rect 27144 9382 27196 9434
rect 27268 9382 27320 9434
rect 35896 9382 35948 9434
rect 36020 9382 36072 9434
rect 36144 9382 36196 9434
rect 36268 9382 36320 9434
rect 44896 9382 44948 9434
rect 45020 9382 45072 9434
rect 45144 9382 45196 9434
rect 45268 9382 45320 9434
rect 53896 9382 53948 9434
rect 54020 9382 54072 9434
rect 54144 9382 54196 9434
rect 54268 9382 54320 9434
rect 62896 9382 62948 9434
rect 63020 9382 63072 9434
rect 63144 9382 63196 9434
rect 63268 9382 63320 9434
rect 71896 9382 71948 9434
rect 72020 9382 72072 9434
rect 72144 9382 72196 9434
rect 72268 9382 72320 9434
rect 80896 9382 80948 9434
rect 81020 9382 81072 9434
rect 81144 9382 81196 9434
rect 81268 9382 81320 9434
rect 89896 9382 89948 9434
rect 90020 9382 90072 9434
rect 90144 9382 90196 9434
rect 90268 9382 90320 9434
rect 96686 9214 96738 9266
rect 96910 9214 96962 9266
rect 48862 9102 48914 9154
rect 49198 9102 49250 9154
rect 80670 9102 80722 9154
rect 31838 8990 31890 9042
rect 35534 8990 35586 9042
rect 43150 8990 43202 9042
rect 50206 8990 50258 9042
rect 50542 8990 50594 9042
rect 63086 8990 63138 9042
rect 68910 8990 68962 9042
rect 76078 8990 76130 9042
rect 84030 8990 84082 9042
rect 30158 8878 30210 8930
rect 34526 8878 34578 8930
rect 37214 8878 37266 8930
rect 42702 8878 42754 8930
rect 45950 8878 46002 8930
rect 49758 8878 49810 8930
rect 54574 8878 54626 8930
rect 59838 8878 59890 8930
rect 65550 8878 65602 8930
rect 72494 8878 72546 8930
rect 48750 8766 48802 8818
rect 50094 8766 50146 8818
rect 97694 8766 97746 8818
rect 4396 8598 4448 8650
rect 4520 8598 4572 8650
rect 4644 8598 4696 8650
rect 4768 8598 4820 8650
rect 13396 8598 13448 8650
rect 13520 8598 13572 8650
rect 13644 8598 13696 8650
rect 13768 8598 13820 8650
rect 22396 8598 22448 8650
rect 22520 8598 22572 8650
rect 22644 8598 22696 8650
rect 22768 8598 22820 8650
rect 31396 8598 31448 8650
rect 31520 8598 31572 8650
rect 31644 8598 31696 8650
rect 31768 8598 31820 8650
rect 40396 8598 40448 8650
rect 40520 8598 40572 8650
rect 40644 8598 40696 8650
rect 40768 8598 40820 8650
rect 49396 8598 49448 8650
rect 49520 8598 49572 8650
rect 49644 8598 49696 8650
rect 49768 8598 49820 8650
rect 58396 8598 58448 8650
rect 58520 8598 58572 8650
rect 58644 8598 58696 8650
rect 58768 8598 58820 8650
rect 67396 8598 67448 8650
rect 67520 8598 67572 8650
rect 67644 8598 67696 8650
rect 67768 8598 67820 8650
rect 76396 8598 76448 8650
rect 76520 8598 76572 8650
rect 76644 8598 76696 8650
rect 76768 8598 76820 8650
rect 85396 8598 85448 8650
rect 85520 8598 85572 8650
rect 85644 8598 85696 8650
rect 85768 8598 85820 8650
rect 94396 8598 94448 8650
rect 94520 8598 94572 8650
rect 94644 8598 94696 8650
rect 94768 8598 94820 8650
rect 45726 8318 45778 8370
rect 58830 8318 58882 8370
rect 81454 8318 81506 8370
rect 81790 8318 81842 8370
rect 36430 8206 36482 8258
rect 40014 8206 40066 8258
rect 45390 8206 45442 8258
rect 45838 8206 45890 8258
rect 46286 8206 46338 8258
rect 51886 8206 51938 8258
rect 52670 8206 52722 8258
rect 58942 8206 58994 8258
rect 59166 8206 59218 8258
rect 61966 8206 62018 8258
rect 69022 8206 69074 8258
rect 81454 8206 81506 8258
rect 88062 8206 88114 8258
rect 34302 8094 34354 8146
rect 44046 8094 44098 8146
rect 44830 8094 44882 8146
rect 48638 8094 48690 8146
rect 54686 8094 54738 8146
rect 63870 8094 63922 8146
rect 71374 8094 71426 8146
rect 76414 8094 76466 8146
rect 86158 8094 86210 8146
rect 58830 7982 58882 8034
rect 66222 7982 66274 8034
rect 81902 7982 81954 8034
rect 8896 7814 8948 7866
rect 9020 7814 9072 7866
rect 9144 7814 9196 7866
rect 9268 7814 9320 7866
rect 17896 7814 17948 7866
rect 18020 7814 18072 7866
rect 18144 7814 18196 7866
rect 18268 7814 18320 7866
rect 26896 7814 26948 7866
rect 27020 7814 27072 7866
rect 27144 7814 27196 7866
rect 27268 7814 27320 7866
rect 35896 7814 35948 7866
rect 36020 7814 36072 7866
rect 36144 7814 36196 7866
rect 36268 7814 36320 7866
rect 44896 7814 44948 7866
rect 45020 7814 45072 7866
rect 45144 7814 45196 7866
rect 45268 7814 45320 7866
rect 53896 7814 53948 7866
rect 54020 7814 54072 7866
rect 54144 7814 54196 7866
rect 54268 7814 54320 7866
rect 62896 7814 62948 7866
rect 63020 7814 63072 7866
rect 63144 7814 63196 7866
rect 63268 7814 63320 7866
rect 71896 7814 71948 7866
rect 72020 7814 72072 7866
rect 72144 7814 72196 7866
rect 72268 7814 72320 7866
rect 80896 7814 80948 7866
rect 81020 7814 81072 7866
rect 81144 7814 81196 7866
rect 81268 7814 81320 7866
rect 89896 7814 89948 7866
rect 90020 7814 90072 7866
rect 90144 7814 90196 7866
rect 90268 7814 90320 7866
rect 42478 7646 42530 7698
rect 48974 7646 49026 7698
rect 49870 7646 49922 7698
rect 30046 7534 30098 7586
rect 33518 7534 33570 7586
rect 34302 7534 34354 7586
rect 34638 7534 34690 7586
rect 41246 7534 41298 7586
rect 59278 7534 59330 7586
rect 62190 7534 62242 7586
rect 66446 7534 66498 7586
rect 90862 7534 90914 7586
rect 32510 7422 32562 7474
rect 40126 7422 40178 7474
rect 42142 7422 42194 7474
rect 42478 7422 42530 7474
rect 42926 7422 42978 7474
rect 50318 7422 50370 7474
rect 51998 7422 52050 7474
rect 56590 7422 56642 7474
rect 64654 7422 64706 7474
rect 71038 7422 71090 7474
rect 71374 7422 71426 7474
rect 77198 7422 77250 7474
rect 78318 7422 78370 7474
rect 84030 7422 84082 7474
rect 87950 7422 88002 7474
rect 1822 7310 1874 7362
rect 38334 7310 38386 7362
rect 45390 7310 45442 7362
rect 53790 7310 53842 7362
rect 70366 7310 70418 7362
rect 74062 7310 74114 7362
rect 77982 7310 78034 7362
rect 81566 7310 81618 7362
rect 34190 7198 34242 7250
rect 34750 7198 34802 7250
rect 41694 7198 41746 7250
rect 42366 7198 42418 7250
rect 71150 7198 71202 7250
rect 71486 7198 71538 7250
rect 4396 7030 4448 7082
rect 4520 7030 4572 7082
rect 4644 7030 4696 7082
rect 4768 7030 4820 7082
rect 13396 7030 13448 7082
rect 13520 7030 13572 7082
rect 13644 7030 13696 7082
rect 13768 7030 13820 7082
rect 22396 7030 22448 7082
rect 22520 7030 22572 7082
rect 22644 7030 22696 7082
rect 22768 7030 22820 7082
rect 31396 7030 31448 7082
rect 31520 7030 31572 7082
rect 31644 7030 31696 7082
rect 31768 7030 31820 7082
rect 40396 7030 40448 7082
rect 40520 7030 40572 7082
rect 40644 7030 40696 7082
rect 40768 7030 40820 7082
rect 49396 7030 49448 7082
rect 49520 7030 49572 7082
rect 49644 7030 49696 7082
rect 49768 7030 49820 7082
rect 58396 7030 58448 7082
rect 58520 7030 58572 7082
rect 58644 7030 58696 7082
rect 58768 7030 58820 7082
rect 67396 7030 67448 7082
rect 67520 7030 67572 7082
rect 67644 7030 67696 7082
rect 67768 7030 67820 7082
rect 76396 7030 76448 7082
rect 76520 7030 76572 7082
rect 76644 7030 76696 7082
rect 76768 7030 76820 7082
rect 85396 7030 85448 7082
rect 85520 7030 85572 7082
rect 85644 7030 85696 7082
rect 85768 7030 85820 7082
rect 94396 7030 94448 7082
rect 94520 7030 94572 7082
rect 94644 7030 94696 7082
rect 94768 7030 94820 7082
rect 37102 6862 37154 6914
rect 37326 6862 37378 6914
rect 37438 6862 37490 6914
rect 59278 6862 59330 6914
rect 59502 6862 59554 6914
rect 59726 6862 59778 6914
rect 46286 6750 46338 6802
rect 51886 6750 51938 6802
rect 64318 6750 64370 6802
rect 87950 6750 88002 6802
rect 2270 6638 2322 6690
rect 25118 6638 25170 6690
rect 25902 6638 25954 6690
rect 26798 6638 26850 6690
rect 28366 6638 28418 6690
rect 35646 6638 35698 6690
rect 44270 6638 44322 6690
rect 45614 6638 45666 6690
rect 46062 6638 46114 6690
rect 47854 6638 47906 6690
rect 54350 6638 54402 6690
rect 59838 6638 59890 6690
rect 60510 6638 60562 6690
rect 72718 6638 72770 6690
rect 73950 6638 74002 6690
rect 74062 6638 74114 6690
rect 76190 6638 76242 6690
rect 84030 6638 84082 6690
rect 96686 6638 96738 6690
rect 96910 6638 96962 6690
rect 27918 6526 27970 6578
rect 34414 6526 34466 6578
rect 36990 6526 37042 6578
rect 41918 6526 41970 6578
rect 54910 6526 54962 6578
rect 69022 6526 69074 6578
rect 78206 6526 78258 6578
rect 81790 6526 81842 6578
rect 98030 6526 98082 6578
rect 1710 6414 1762 6466
rect 27582 6414 27634 6466
rect 29374 6414 29426 6466
rect 37998 6414 38050 6466
rect 45390 6414 45442 6466
rect 59390 6414 59442 6466
rect 74510 6414 74562 6466
rect 74846 6414 74898 6466
rect 75406 6414 75458 6466
rect 81902 6414 81954 6466
rect 82350 6414 82402 6466
rect 8896 6246 8948 6298
rect 9020 6246 9072 6298
rect 9144 6246 9196 6298
rect 9268 6246 9320 6298
rect 17896 6246 17948 6298
rect 18020 6246 18072 6298
rect 18144 6246 18196 6298
rect 18268 6246 18320 6298
rect 26896 6246 26948 6298
rect 27020 6246 27072 6298
rect 27144 6246 27196 6298
rect 27268 6246 27320 6298
rect 35896 6246 35948 6298
rect 36020 6246 36072 6298
rect 36144 6246 36196 6298
rect 36268 6246 36320 6298
rect 44896 6246 44948 6298
rect 45020 6246 45072 6298
rect 45144 6246 45196 6298
rect 45268 6246 45320 6298
rect 53896 6246 53948 6298
rect 54020 6246 54072 6298
rect 54144 6246 54196 6298
rect 54268 6246 54320 6298
rect 62896 6246 62948 6298
rect 63020 6246 63072 6298
rect 63144 6246 63196 6298
rect 63268 6246 63320 6298
rect 71896 6246 71948 6298
rect 72020 6246 72072 6298
rect 72144 6246 72196 6298
rect 72268 6246 72320 6298
rect 80896 6246 80948 6298
rect 81020 6246 81072 6298
rect 81144 6246 81196 6298
rect 81268 6246 81320 6298
rect 89896 6246 89948 6298
rect 90020 6246 90072 6298
rect 90144 6246 90196 6298
rect 90268 6246 90320 6298
rect 34862 6078 34914 6130
rect 41022 6078 41074 6130
rect 41694 6078 41746 6130
rect 42142 6078 42194 6130
rect 42590 6078 42642 6130
rect 71262 6078 71314 6130
rect 78094 6078 78146 6130
rect 78542 6078 78594 6130
rect 78990 6078 79042 6130
rect 31054 5966 31106 6018
rect 33518 5966 33570 6018
rect 35646 5966 35698 6018
rect 40910 5966 40962 6018
rect 49982 5966 50034 6018
rect 55358 5966 55410 6018
rect 58830 5966 58882 6018
rect 63758 5966 63810 6018
rect 63870 5966 63922 6018
rect 68798 5966 68850 6018
rect 70254 5966 70306 6018
rect 70814 5966 70866 6018
rect 72494 5966 72546 6018
rect 83918 5966 83970 6018
rect 90750 5966 90802 6018
rect 1822 5854 1874 5906
rect 27582 5854 27634 5906
rect 33854 5854 33906 5906
rect 34190 5854 34242 5906
rect 34750 5854 34802 5906
rect 40126 5854 40178 5906
rect 48190 5854 48242 5906
rect 49086 5854 49138 5906
rect 49310 5854 49362 5906
rect 49870 5854 49922 5906
rect 50766 5854 50818 5906
rect 57150 5854 57202 5906
rect 62078 5854 62130 5906
rect 62526 5854 62578 5906
rect 62862 5854 62914 5906
rect 64430 5854 64482 5906
rect 71038 5854 71090 5906
rect 71710 5854 71762 5906
rect 76078 5854 76130 5906
rect 80110 5854 80162 5906
rect 88174 5854 88226 5906
rect 2270 5742 2322 5794
rect 34526 5742 34578 5794
rect 45278 5742 45330 5794
rect 50430 5742 50482 5794
rect 62414 5742 62466 5794
rect 70814 5742 70866 5794
rect 79438 5742 79490 5794
rect 34302 5630 34354 5682
rect 48974 5630 49026 5682
rect 49422 5630 49474 5682
rect 70366 5630 70418 5682
rect 71598 5630 71650 5682
rect 4396 5462 4448 5514
rect 4520 5462 4572 5514
rect 4644 5462 4696 5514
rect 4768 5462 4820 5514
rect 13396 5462 13448 5514
rect 13520 5462 13572 5514
rect 13644 5462 13696 5514
rect 13768 5462 13820 5514
rect 22396 5462 22448 5514
rect 22520 5462 22572 5514
rect 22644 5462 22696 5514
rect 22768 5462 22820 5514
rect 31396 5462 31448 5514
rect 31520 5462 31572 5514
rect 31644 5462 31696 5514
rect 31768 5462 31820 5514
rect 40396 5462 40448 5514
rect 40520 5462 40572 5514
rect 40644 5462 40696 5514
rect 40768 5462 40820 5514
rect 49396 5462 49448 5514
rect 49520 5462 49572 5514
rect 49644 5462 49696 5514
rect 49768 5462 49820 5514
rect 58396 5462 58448 5514
rect 58520 5462 58572 5514
rect 58644 5462 58696 5514
rect 58768 5462 58820 5514
rect 67396 5462 67448 5514
rect 67520 5462 67572 5514
rect 67644 5462 67696 5514
rect 67768 5462 67820 5514
rect 76396 5462 76448 5514
rect 76520 5462 76572 5514
rect 76644 5462 76696 5514
rect 76768 5462 76820 5514
rect 85396 5462 85448 5514
rect 85520 5462 85572 5514
rect 85644 5462 85696 5514
rect 85768 5462 85820 5514
rect 94396 5462 94448 5514
rect 94520 5462 94572 5514
rect 94644 5462 94696 5514
rect 94768 5462 94820 5514
rect 30718 5294 30770 5346
rect 37214 5294 37266 5346
rect 58270 5294 58322 5346
rect 59950 5294 60002 5346
rect 67790 5294 67842 5346
rect 74846 5294 74898 5346
rect 1822 5182 1874 5234
rect 26574 5182 26626 5234
rect 34414 5182 34466 5234
rect 42254 5182 42306 5234
rect 44942 5182 44994 5234
rect 46286 5182 46338 5234
rect 51774 5182 51826 5234
rect 54686 5182 54738 5234
rect 60734 5182 60786 5234
rect 70702 5182 70754 5234
rect 73950 5182 74002 5234
rect 79102 5182 79154 5234
rect 87502 5182 87554 5234
rect 96574 5182 96626 5234
rect 28478 5070 28530 5122
rect 36430 5070 36482 5122
rect 36990 5070 37042 5122
rect 37438 5070 37490 5122
rect 37886 5070 37938 5122
rect 37998 5070 38050 5122
rect 42814 5070 42866 5122
rect 45838 5070 45890 5122
rect 46174 5070 46226 5122
rect 48302 5070 48354 5122
rect 57934 5070 57986 5122
rect 59166 5070 59218 5122
rect 59838 5070 59890 5122
rect 65438 5070 65490 5122
rect 67342 5070 67394 5122
rect 68350 5070 68402 5122
rect 74398 5070 74450 5122
rect 77086 5070 77138 5122
rect 83246 5070 83298 5122
rect 84254 5070 84306 5122
rect 96910 5070 96962 5122
rect 97694 5070 97746 5122
rect 59054 4958 59106 5010
rect 59278 4958 59330 5010
rect 59614 4958 59666 5010
rect 82126 4958 82178 5010
rect 37102 4846 37154 4898
rect 38670 4846 38722 4898
rect 46622 4846 46674 4898
rect 75294 4846 75346 4898
rect 8896 4678 8948 4730
rect 9020 4678 9072 4730
rect 9144 4678 9196 4730
rect 9268 4678 9320 4730
rect 17896 4678 17948 4730
rect 18020 4678 18072 4730
rect 18144 4678 18196 4730
rect 18268 4678 18320 4730
rect 26896 4678 26948 4730
rect 27020 4678 27072 4730
rect 27144 4678 27196 4730
rect 27268 4678 27320 4730
rect 35896 4678 35948 4730
rect 36020 4678 36072 4730
rect 36144 4678 36196 4730
rect 36268 4678 36320 4730
rect 44896 4678 44948 4730
rect 45020 4678 45072 4730
rect 45144 4678 45196 4730
rect 45268 4678 45320 4730
rect 53896 4678 53948 4730
rect 54020 4678 54072 4730
rect 54144 4678 54196 4730
rect 54268 4678 54320 4730
rect 62896 4678 62948 4730
rect 63020 4678 63072 4730
rect 63144 4678 63196 4730
rect 63268 4678 63320 4730
rect 71896 4678 71948 4730
rect 72020 4678 72072 4730
rect 72144 4678 72196 4730
rect 72268 4678 72320 4730
rect 80896 4678 80948 4730
rect 81020 4678 81072 4730
rect 81144 4678 81196 4730
rect 81268 4678 81320 4730
rect 89896 4678 89948 4730
rect 90020 4678 90072 4730
rect 90144 4678 90196 4730
rect 90268 4678 90320 4730
rect 34526 4510 34578 4562
rect 49870 4510 49922 4562
rect 63198 4510 63250 4562
rect 70142 4510 70194 4562
rect 70926 4510 70978 4562
rect 78430 4510 78482 4562
rect 91198 4510 91250 4562
rect 96686 4510 96738 4562
rect 96910 4510 96962 4562
rect 30158 4398 30210 4450
rect 34078 4398 34130 4450
rect 34414 4398 34466 4450
rect 38334 4398 38386 4450
rect 41694 4398 41746 4450
rect 42030 4398 42082 4450
rect 42254 4398 42306 4450
rect 44158 4398 44210 4450
rect 49422 4398 49474 4450
rect 49758 4398 49810 4450
rect 49982 4398 50034 4450
rect 52782 4398 52834 4450
rect 58718 4398 58770 4450
rect 62750 4398 62802 4450
rect 63534 4398 63586 4450
rect 65774 4398 65826 4450
rect 71374 4398 71426 4450
rect 75630 4398 75682 4450
rect 78318 4398 78370 4450
rect 82126 4398 82178 4450
rect 31054 4286 31106 4338
rect 33854 4286 33906 4338
rect 34638 4286 34690 4338
rect 40238 4286 40290 4338
rect 41358 4286 41410 4338
rect 41470 4286 41522 4338
rect 48190 4286 48242 4338
rect 49086 4286 49138 4338
rect 51326 4286 51378 4338
rect 61854 4286 61906 4338
rect 68910 4286 68962 4338
rect 70030 4286 70082 4338
rect 70702 4286 70754 4338
rect 71038 4286 71090 4338
rect 72830 4286 72882 4338
rect 81566 4286 81618 4338
rect 88062 4286 88114 4338
rect 33406 4174 33458 4226
rect 42366 4174 42418 4226
rect 62190 4174 62242 4226
rect 71710 4174 71762 4226
rect 77982 4174 78034 4226
rect 78878 4174 78930 4226
rect 85934 4174 85986 4226
rect 33742 4062 33794 4114
rect 41022 4062 41074 4114
rect 49198 4062 49250 4114
rect 71598 4062 71650 4114
rect 79438 4062 79490 4114
rect 97694 4062 97746 4114
rect 4396 3894 4448 3946
rect 4520 3894 4572 3946
rect 4644 3894 4696 3946
rect 4768 3894 4820 3946
rect 13396 3894 13448 3946
rect 13520 3894 13572 3946
rect 13644 3894 13696 3946
rect 13768 3894 13820 3946
rect 22396 3894 22448 3946
rect 22520 3894 22572 3946
rect 22644 3894 22696 3946
rect 22768 3894 22820 3946
rect 31396 3894 31448 3946
rect 31520 3894 31572 3946
rect 31644 3894 31696 3946
rect 31768 3894 31820 3946
rect 40396 3894 40448 3946
rect 40520 3894 40572 3946
rect 40644 3894 40696 3946
rect 40768 3894 40820 3946
rect 49396 3894 49448 3946
rect 49520 3894 49572 3946
rect 49644 3894 49696 3946
rect 49768 3894 49820 3946
rect 58396 3894 58448 3946
rect 58520 3894 58572 3946
rect 58644 3894 58696 3946
rect 58768 3894 58820 3946
rect 67396 3894 67448 3946
rect 67520 3894 67572 3946
rect 67644 3894 67696 3946
rect 67768 3894 67820 3946
rect 76396 3894 76448 3946
rect 76520 3894 76572 3946
rect 76644 3894 76696 3946
rect 76768 3894 76820 3946
rect 85396 3894 85448 3946
rect 85520 3894 85572 3946
rect 85644 3894 85696 3946
rect 85768 3894 85820 3946
rect 94396 3894 94448 3946
rect 94520 3894 94572 3946
rect 94644 3894 94696 3946
rect 94768 3894 94820 3946
rect 34190 3726 34242 3778
rect 34302 3726 34354 3778
rect 34638 3726 34690 3778
rect 37102 3726 37154 3778
rect 38558 3726 38610 3778
rect 39230 3726 39282 3778
rect 41022 3726 41074 3778
rect 44046 3726 44098 3778
rect 44830 3726 44882 3778
rect 45166 3726 45218 3778
rect 45278 3726 45330 3778
rect 45950 3726 46002 3778
rect 46846 3726 46898 3778
rect 58270 3726 58322 3778
rect 60846 3726 60898 3778
rect 69582 3726 69634 3778
rect 77982 3726 78034 3778
rect 17838 3614 17890 3666
rect 28814 3614 28866 3666
rect 31278 3614 31330 3666
rect 32510 3614 32562 3666
rect 33070 3614 33122 3666
rect 33406 3614 33458 3666
rect 35198 3614 35250 3666
rect 36542 3614 36594 3666
rect 38782 3614 38834 3666
rect 40910 3614 40962 3666
rect 41918 3614 41970 3666
rect 44270 3614 44322 3666
rect 47742 3614 47794 3666
rect 48526 3614 48578 3666
rect 50318 3614 50370 3666
rect 51438 3614 51490 3666
rect 51886 3614 51938 3666
rect 52334 3614 52386 3666
rect 55470 3614 55522 3666
rect 57486 3614 57538 3666
rect 59054 3614 59106 3666
rect 60734 3614 60786 3666
rect 61742 3614 61794 3666
rect 62750 3614 62802 3666
rect 67454 3614 67506 3666
rect 71038 3614 71090 3666
rect 74286 3614 74338 3666
rect 75518 3614 75570 3666
rect 79998 3614 80050 3666
rect 82462 3614 82514 3666
rect 84702 3614 84754 3666
rect 85710 3614 85762 3666
rect 96350 3614 96402 3666
rect 31726 3502 31778 3554
rect 33294 3502 33346 3554
rect 34750 3502 34802 3554
rect 36094 3502 36146 3554
rect 37438 3502 37490 3554
rect 37886 3502 37938 3554
rect 38334 3502 38386 3554
rect 39118 3502 39170 3554
rect 40350 3502 40402 3554
rect 41582 3502 41634 3554
rect 41806 3502 41858 3554
rect 42478 3502 42530 3554
rect 42926 3502 42978 3554
rect 43486 3502 43538 3554
rect 44494 3502 44546 3554
rect 44942 3502 44994 3554
rect 47966 3502 48018 3554
rect 49310 3502 49362 3554
rect 49422 3502 49474 3554
rect 49982 3502 50034 3554
rect 50206 3502 50258 3554
rect 54574 3502 54626 3554
rect 55022 3502 55074 3554
rect 57822 3502 57874 3554
rect 58158 3502 58210 3554
rect 59390 3502 59442 3554
rect 60062 3502 60114 3554
rect 60174 3502 60226 3554
rect 61294 3502 61346 3554
rect 63198 3502 63250 3554
rect 65998 3502 66050 3554
rect 66446 3502 66498 3554
rect 71262 3502 71314 3554
rect 77310 3502 77362 3554
rect 78094 3502 78146 3554
rect 80670 3502 80722 3554
rect 82798 3502 82850 3554
rect 86158 3502 86210 3554
rect 94334 3502 94386 3554
rect 96910 3502 96962 3554
rect 6078 3390 6130 3442
rect 6302 3390 6354 3442
rect 6638 3390 6690 3442
rect 16494 3390 16546 3442
rect 17278 3390 17330 3442
rect 27918 3390 27970 3442
rect 28366 3390 28418 3442
rect 33630 3390 33682 3442
rect 33966 3390 34018 3442
rect 37102 3390 37154 3442
rect 39790 3390 39842 3442
rect 41246 3390 41298 3442
rect 42590 3390 42642 3442
rect 43822 3390 43874 3442
rect 46734 3390 46786 3442
rect 48862 3390 48914 3442
rect 49758 3390 49810 3442
rect 52670 3390 52722 3442
rect 59950 3390 60002 3442
rect 60510 3390 60562 3442
rect 69694 3390 69746 3442
rect 71822 3390 71874 3442
rect 73278 3390 73330 3442
rect 76750 3390 76802 3442
rect 83246 3390 83298 3442
rect 93886 3390 93938 3442
rect 94110 3390 94162 3442
rect 97694 3390 97746 3442
rect 43038 3278 43090 3330
rect 43934 3278 43986 3330
rect 46398 3278 46450 3330
rect 72718 3278 72770 3330
rect 75854 3278 75906 3330
rect 81902 3278 81954 3330
rect 8896 3110 8948 3162
rect 9020 3110 9072 3162
rect 9144 3110 9196 3162
rect 9268 3110 9320 3162
rect 17896 3110 17948 3162
rect 18020 3110 18072 3162
rect 18144 3110 18196 3162
rect 18268 3110 18320 3162
rect 26896 3110 26948 3162
rect 27020 3110 27072 3162
rect 27144 3110 27196 3162
rect 27268 3110 27320 3162
rect 35896 3110 35948 3162
rect 36020 3110 36072 3162
rect 36144 3110 36196 3162
rect 36268 3110 36320 3162
rect 44896 3110 44948 3162
rect 45020 3110 45072 3162
rect 45144 3110 45196 3162
rect 45268 3110 45320 3162
rect 53896 3110 53948 3162
rect 54020 3110 54072 3162
rect 54144 3110 54196 3162
rect 54268 3110 54320 3162
rect 62896 3110 62948 3162
rect 63020 3110 63072 3162
rect 63144 3110 63196 3162
rect 63268 3110 63320 3162
rect 71896 3110 71948 3162
rect 72020 3110 72072 3162
rect 72144 3110 72196 3162
rect 72268 3110 72320 3162
rect 80896 3110 80948 3162
rect 81020 3110 81072 3162
rect 81144 3110 81196 3162
rect 81268 3110 81320 3162
rect 89896 3110 89948 3162
rect 90020 3110 90072 3162
rect 90144 3110 90196 3162
rect 90268 3110 90320 3162
<< metal2 >>
rect 6720 59200 6832 60000
rect 19040 59200 19152 60000
rect 31360 59200 31472 60000
rect 43680 59200 43792 60000
rect 56000 59200 56112 60000
rect 68320 59200 68432 60000
rect 80640 59200 80752 60000
rect 92960 59200 93072 60000
rect 6748 56642 6804 59200
rect 6748 56590 6750 56642
rect 6802 56590 6804 56642
rect 6748 56578 6804 56590
rect 7308 56642 7364 56654
rect 7308 56590 7310 56642
rect 7362 56590 7364 56642
rect 2044 56196 2100 56206
rect 2044 56102 2100 56140
rect 7308 56194 7364 56590
rect 8768 56476 9448 56486
rect 8824 56420 8872 56476
rect 8928 56474 8976 56476
rect 9032 56474 9080 56476
rect 8948 56422 8976 56474
rect 9072 56422 9080 56474
rect 8928 56420 8976 56422
rect 9032 56420 9080 56422
rect 9136 56474 9184 56476
rect 9240 56474 9288 56476
rect 9136 56422 9144 56474
rect 9240 56422 9268 56474
rect 9136 56420 9184 56422
rect 9240 56420 9288 56422
rect 9344 56420 9392 56476
rect 8768 56410 9448 56420
rect 17768 56476 18448 56486
rect 17824 56420 17872 56476
rect 17928 56474 17976 56476
rect 18032 56474 18080 56476
rect 17948 56422 17976 56474
rect 18072 56422 18080 56474
rect 17928 56420 17976 56422
rect 18032 56420 18080 56422
rect 18136 56474 18184 56476
rect 18240 56474 18288 56476
rect 18136 56422 18144 56474
rect 18240 56422 18268 56474
rect 18136 56420 18184 56422
rect 18240 56420 18288 56422
rect 18344 56420 18392 56476
rect 17768 56410 18448 56420
rect 7308 56142 7310 56194
rect 7362 56142 7364 56194
rect 7308 56130 7364 56142
rect 12124 56196 12180 56206
rect 1708 56082 1764 56094
rect 1708 56030 1710 56082
rect 1762 56030 1764 56082
rect 1708 55636 1764 56030
rect 8204 56082 8260 56094
rect 8204 56030 8206 56082
rect 8258 56030 8260 56082
rect 1708 55570 1764 55580
rect 2492 55970 2548 55982
rect 2492 55918 2494 55970
rect 2546 55918 2548 55970
rect 2492 55636 2548 55918
rect 8204 55972 8260 56030
rect 8204 55906 8260 55916
rect 8764 55972 8820 55982
rect 8764 55878 8820 55916
rect 4268 55692 4948 55702
rect 4324 55636 4372 55692
rect 4428 55690 4476 55692
rect 4532 55690 4580 55692
rect 4448 55638 4476 55690
rect 4572 55638 4580 55690
rect 4428 55636 4476 55638
rect 4532 55636 4580 55638
rect 4636 55690 4684 55692
rect 4740 55690 4788 55692
rect 4636 55638 4644 55690
rect 4740 55638 4768 55690
rect 4636 55636 4684 55638
rect 4740 55636 4788 55638
rect 4844 55636 4892 55692
rect 4268 55626 4948 55636
rect 2492 55570 2548 55580
rect 1708 55186 1764 55198
rect 1708 55134 1710 55186
rect 1762 55134 1764 55186
rect 1708 55076 1764 55134
rect 1708 54516 1764 55020
rect 1708 54450 1764 54460
rect 2044 55074 2100 55086
rect 2044 55022 2046 55074
rect 2098 55022 2100 55074
rect 2044 53732 2100 55022
rect 2492 55076 2548 55086
rect 2492 54982 2548 55020
rect 8768 54908 9448 54918
rect 8824 54852 8872 54908
rect 8928 54906 8976 54908
rect 9032 54906 9080 54908
rect 8948 54854 8976 54906
rect 9072 54854 9080 54906
rect 8928 54852 8976 54854
rect 9032 54852 9080 54854
rect 9136 54906 9184 54908
rect 9240 54906 9288 54908
rect 9136 54854 9144 54906
rect 9240 54854 9268 54906
rect 9136 54852 9184 54854
rect 9240 54852 9288 54854
rect 9344 54852 9392 54908
rect 8768 54842 9448 54852
rect 4268 54124 4948 54134
rect 4324 54068 4372 54124
rect 4428 54122 4476 54124
rect 4532 54122 4580 54124
rect 4448 54070 4476 54122
rect 4572 54070 4580 54122
rect 4428 54068 4476 54070
rect 4532 54068 4580 54070
rect 4636 54122 4684 54124
rect 4740 54122 4788 54124
rect 4636 54070 4644 54122
rect 4740 54070 4768 54122
rect 4636 54068 4684 54070
rect 4740 54068 4788 54070
rect 4844 54068 4892 54124
rect 4268 54058 4948 54068
rect 1820 53676 2100 53732
rect 1708 53618 1764 53630
rect 1708 53566 1710 53618
rect 1762 53566 1764 53618
rect 1708 53396 1764 53566
rect 1708 53330 1764 53340
rect 1708 52946 1764 52958
rect 1708 52894 1710 52946
rect 1762 52894 1764 52946
rect 1708 52836 1764 52894
rect 1708 52276 1764 52780
rect 1708 52210 1764 52220
rect 1708 51378 1764 51390
rect 1708 51326 1710 51378
rect 1762 51326 1764 51378
rect 1708 51156 1764 51326
rect 1708 51090 1764 51100
rect 1708 50482 1764 50494
rect 1708 50430 1710 50482
rect 1762 50430 1764 50482
rect 1708 50036 1764 50430
rect 1820 50148 1876 53676
rect 2044 53508 2100 53518
rect 1932 53506 2100 53508
rect 1932 53454 2046 53506
rect 2098 53454 2100 53506
rect 1932 53452 2100 53454
rect 1932 50484 1988 53452
rect 2044 53442 2100 53452
rect 2492 53506 2548 53518
rect 2492 53454 2494 53506
rect 2546 53454 2548 53506
rect 2492 53396 2548 53454
rect 2492 53330 2548 53340
rect 8768 53340 9448 53350
rect 8824 53284 8872 53340
rect 8928 53338 8976 53340
rect 9032 53338 9080 53340
rect 8948 53286 8976 53338
rect 9072 53286 9080 53338
rect 8928 53284 8976 53286
rect 9032 53284 9080 53286
rect 9136 53338 9184 53340
rect 9240 53338 9288 53340
rect 9136 53286 9144 53338
rect 9240 53286 9268 53338
rect 9136 53284 9184 53286
rect 9240 53284 9288 53286
rect 9344 53284 9392 53340
rect 8768 53274 9448 53284
rect 2044 53058 2100 53070
rect 2044 53006 2046 53058
rect 2098 53006 2100 53058
rect 2044 51716 2100 53006
rect 2492 52836 2548 52846
rect 2492 52742 2548 52780
rect 4268 52556 4948 52566
rect 4324 52500 4372 52556
rect 4428 52554 4476 52556
rect 4532 52554 4580 52556
rect 4448 52502 4476 52554
rect 4572 52502 4580 52554
rect 4428 52500 4476 52502
rect 4532 52500 4580 52502
rect 4636 52554 4684 52556
rect 4740 52554 4788 52556
rect 4636 52502 4644 52554
rect 4740 52502 4768 52554
rect 4636 52500 4684 52502
rect 4740 52500 4788 52502
rect 4844 52500 4892 52556
rect 4268 52490 4948 52500
rect 8768 51772 9448 51782
rect 2044 51650 2100 51660
rect 5852 51716 5908 51726
rect 8824 51716 8872 51772
rect 8928 51770 8976 51772
rect 9032 51770 9080 51772
rect 8948 51718 8976 51770
rect 9072 51718 9080 51770
rect 8928 51716 8976 51718
rect 9032 51716 9080 51718
rect 9136 51770 9184 51772
rect 9240 51770 9288 51772
rect 9136 51718 9144 51770
rect 9240 51718 9268 51770
rect 9136 51716 9184 51718
rect 9240 51716 9288 51718
rect 9344 51716 9392 51772
rect 8768 51706 9448 51716
rect 2044 51492 2100 51502
rect 2044 51490 2324 51492
rect 2044 51438 2046 51490
rect 2098 51438 2324 51490
rect 2044 51436 2324 51438
rect 2044 51426 2100 51436
rect 1932 50418 1988 50428
rect 2044 50482 2100 50494
rect 2044 50430 2046 50482
rect 2098 50430 2100 50482
rect 2044 50372 2100 50430
rect 2044 50306 2100 50316
rect 1820 50092 2212 50148
rect 1708 49970 1764 49980
rect 1932 49924 1988 49934
rect 1820 49922 1988 49924
rect 1820 49870 1934 49922
rect 1986 49870 1988 49922
rect 1820 49868 1988 49870
rect 1708 48914 1764 48926
rect 1708 48862 1710 48914
rect 1762 48862 1764 48914
rect 1708 48692 1764 48862
rect 1708 47796 1764 48636
rect 1820 48242 1876 49868
rect 1932 49858 1988 49868
rect 1820 48190 1822 48242
rect 1874 48190 1876 48242
rect 1820 48178 1876 48190
rect 2044 48802 2100 48814
rect 2044 48750 2046 48802
rect 2098 48750 2100 48802
rect 1708 47730 1764 47740
rect 2044 47572 2100 48750
rect 2156 48242 2212 50092
rect 2268 49028 2324 51436
rect 2492 51266 2548 51278
rect 2492 51214 2494 51266
rect 2546 51214 2548 51266
rect 2492 51156 2548 51214
rect 2492 51090 2548 51100
rect 4268 50988 4948 50998
rect 4324 50932 4372 50988
rect 4428 50986 4476 50988
rect 4532 50986 4580 50988
rect 4448 50934 4476 50986
rect 4572 50934 4580 50986
rect 4428 50932 4476 50934
rect 4532 50932 4580 50934
rect 4636 50986 4684 50988
rect 4740 50986 4788 50988
rect 4636 50934 4644 50986
rect 4740 50934 4768 50986
rect 4636 50932 4684 50934
rect 4740 50932 4788 50934
rect 4844 50932 4892 50988
rect 4268 50922 4948 50932
rect 2492 50482 2548 50494
rect 2492 50430 2494 50482
rect 2546 50430 2548 50482
rect 2492 50036 2548 50430
rect 2492 49970 2548 49980
rect 2828 50372 2884 50382
rect 2268 48962 2324 48972
rect 2492 49698 2548 49710
rect 2492 49646 2494 49698
rect 2546 49646 2548 49698
rect 2380 48916 2436 48926
rect 2380 48822 2436 48860
rect 2492 48692 2548 49646
rect 2492 48626 2548 48636
rect 2716 48802 2772 48814
rect 2716 48750 2718 48802
rect 2770 48750 2772 48802
rect 2156 48190 2158 48242
rect 2210 48190 2212 48242
rect 2156 48178 2212 48190
rect 2044 47516 2436 47572
rect 1820 47458 1876 47470
rect 1820 47406 1822 47458
rect 1874 47406 1876 47458
rect 1820 46676 1876 47406
rect 2044 47348 2100 47358
rect 2044 47254 2100 47292
rect 1820 46582 1876 46620
rect 1708 45778 1764 45790
rect 1708 45726 1710 45778
rect 1762 45726 1764 45778
rect 1708 45556 1764 45726
rect 2044 45668 2100 45678
rect 2044 45666 2212 45668
rect 2044 45614 2046 45666
rect 2098 45614 2212 45666
rect 2044 45612 2212 45614
rect 2044 45602 2100 45612
rect 1708 45490 1764 45500
rect 2044 45220 2100 45230
rect 1932 45218 2100 45220
rect 1932 45166 2046 45218
rect 2098 45166 2100 45218
rect 1932 45164 2100 45166
rect 1708 45106 1764 45118
rect 1708 45054 1710 45106
rect 1762 45054 1764 45106
rect 1708 44996 1764 45054
rect 1708 44436 1764 44940
rect 1708 44370 1764 44380
rect 1820 44098 1876 44110
rect 1820 44046 1822 44098
rect 1874 44046 1876 44098
rect 1820 43538 1876 44046
rect 1820 43486 1822 43538
rect 1874 43486 1876 43538
rect 1820 43316 1876 43486
rect 1820 43250 1876 43260
rect 1708 42642 1764 42654
rect 1708 42590 1710 42642
rect 1762 42590 1764 42642
rect 1708 42196 1764 42590
rect 1708 42130 1764 42140
rect 1708 41074 1764 41086
rect 1708 41022 1710 41074
rect 1762 41022 1764 41074
rect 1708 39956 1764 41022
rect 1708 39890 1764 39900
rect 1820 40402 1876 40414
rect 1820 40350 1822 40402
rect 1874 40350 1876 40402
rect 1820 39844 1876 40350
rect 1932 40404 1988 45164
rect 2044 45154 2100 45164
rect 2044 43650 2100 43662
rect 2044 43598 2046 43650
rect 2098 43598 2100 43650
rect 2044 42868 2100 43598
rect 2156 43092 2212 45612
rect 2380 44772 2436 47516
rect 2604 47236 2660 47246
rect 2492 47234 2660 47236
rect 2492 47182 2606 47234
rect 2658 47182 2660 47234
rect 2492 47180 2660 47182
rect 2492 46674 2548 47180
rect 2604 47170 2660 47180
rect 2492 46622 2494 46674
rect 2546 46622 2548 46674
rect 2492 46610 2548 46622
rect 2492 45666 2548 45678
rect 2492 45614 2494 45666
rect 2546 45614 2548 45666
rect 2492 45556 2548 45614
rect 2492 45490 2548 45500
rect 2716 45108 2772 48750
rect 2828 46674 2884 50316
rect 5628 50370 5684 50382
rect 5628 50318 5630 50370
rect 5682 50318 5684 50370
rect 5516 49812 5572 49822
rect 5628 49812 5684 50318
rect 5516 49810 5684 49812
rect 5516 49758 5518 49810
rect 5570 49758 5684 49810
rect 5516 49756 5684 49758
rect 5852 49810 5908 51660
rect 11900 51492 11956 51502
rect 11676 51490 11956 51492
rect 11676 51438 11902 51490
rect 11954 51438 11956 51490
rect 11676 51436 11956 51438
rect 8768 50204 9448 50214
rect 8824 50148 8872 50204
rect 8928 50202 8976 50204
rect 9032 50202 9080 50204
rect 8948 50150 8976 50202
rect 9072 50150 9080 50202
rect 8928 50148 8976 50150
rect 9032 50148 9080 50150
rect 9136 50202 9184 50204
rect 9240 50202 9288 50204
rect 9136 50150 9144 50202
rect 9240 50150 9268 50202
rect 9136 50148 9184 50150
rect 9240 50148 9288 50150
rect 9344 50148 9392 50204
rect 8768 50138 9448 50148
rect 5852 49758 5854 49810
rect 5906 49758 5908 49810
rect 5516 49746 5572 49756
rect 5852 49746 5908 49758
rect 8316 50034 8372 50046
rect 8316 49982 8318 50034
rect 8370 49982 8372 50034
rect 8316 49700 8372 49982
rect 9548 49924 9604 49934
rect 8316 49634 8372 49644
rect 9100 49922 9604 49924
rect 9100 49870 9550 49922
rect 9602 49870 9604 49922
rect 9100 49868 9604 49870
rect 5852 49588 5908 49598
rect 8988 49588 9044 49598
rect 4268 49420 4948 49430
rect 4324 49364 4372 49420
rect 4428 49418 4476 49420
rect 4532 49418 4580 49420
rect 4448 49366 4476 49418
rect 4572 49366 4580 49418
rect 4428 49364 4476 49366
rect 4532 49364 4580 49366
rect 4636 49418 4684 49420
rect 4740 49418 4788 49420
rect 4636 49366 4644 49418
rect 4740 49366 4768 49418
rect 4636 49364 4684 49366
rect 4740 49364 4788 49366
rect 4844 49364 4892 49420
rect 4268 49354 4948 49364
rect 3164 48916 3220 48926
rect 3164 48822 3220 48860
rect 4732 48466 4788 48478
rect 4732 48414 4734 48466
rect 4786 48414 4788 48466
rect 4732 48132 4788 48414
rect 4732 48066 4788 48076
rect 5628 48132 5684 48142
rect 5292 48020 5348 48030
rect 5292 47926 5348 47964
rect 5628 47908 5684 48076
rect 5852 47908 5908 49532
rect 4268 47852 4948 47862
rect 5628 47852 5908 47908
rect 4324 47796 4372 47852
rect 4428 47850 4476 47852
rect 4532 47850 4580 47852
rect 4448 47798 4476 47850
rect 4572 47798 4580 47850
rect 4428 47796 4476 47798
rect 4532 47796 4580 47798
rect 4636 47850 4684 47852
rect 4740 47850 4788 47852
rect 4636 47798 4644 47850
rect 4740 47798 4768 47850
rect 4636 47796 4684 47798
rect 4740 47796 4788 47798
rect 4844 47796 4892 47852
rect 4268 47786 4948 47796
rect 5404 46900 5460 46910
rect 5404 46898 5796 46900
rect 5404 46846 5406 46898
rect 5458 46846 5796 46898
rect 5404 46844 5796 46846
rect 5404 46834 5460 46844
rect 2828 46622 2830 46674
rect 2882 46622 2884 46674
rect 2828 46610 2884 46622
rect 4268 46284 4948 46294
rect 4324 46228 4372 46284
rect 4428 46282 4476 46284
rect 4532 46282 4580 46284
rect 4448 46230 4476 46282
rect 4572 46230 4580 46282
rect 4428 46228 4476 46230
rect 4532 46228 4580 46230
rect 4636 46282 4684 46284
rect 4740 46282 4788 46284
rect 4636 46230 4644 46282
rect 4740 46230 4768 46282
rect 4636 46228 4684 46230
rect 4740 46228 4788 46230
rect 4844 46228 4892 46284
rect 4268 46218 4948 46228
rect 3164 45668 3220 45678
rect 2716 45042 2772 45052
rect 3052 45666 3220 45668
rect 3052 45614 3166 45666
rect 3218 45614 3220 45666
rect 3052 45612 3220 45614
rect 3052 45106 3108 45612
rect 3164 45602 3220 45612
rect 5740 45330 5796 46844
rect 5740 45278 5742 45330
rect 5794 45278 5796 45330
rect 3052 45054 3054 45106
rect 3106 45054 3108 45106
rect 3052 45042 3108 45054
rect 3388 45108 3444 45118
rect 3388 45014 3444 45052
rect 2492 44996 2548 45006
rect 2492 44902 2548 44940
rect 2380 44716 2996 44772
rect 2604 44098 2660 44110
rect 2604 44046 2606 44098
rect 2658 44046 2660 44098
rect 2492 43540 2548 43550
rect 2604 43540 2660 44046
rect 2492 43538 2660 43540
rect 2492 43486 2494 43538
rect 2546 43486 2660 43538
rect 2492 43484 2660 43486
rect 2940 43538 2996 44716
rect 4268 44716 4948 44726
rect 4324 44660 4372 44716
rect 4428 44714 4476 44716
rect 4532 44714 4580 44716
rect 4448 44662 4476 44714
rect 4572 44662 4580 44714
rect 4428 44660 4476 44662
rect 4532 44660 4580 44662
rect 4636 44714 4684 44716
rect 4740 44714 4788 44716
rect 4636 44662 4644 44714
rect 4740 44662 4768 44714
rect 4636 44660 4684 44662
rect 4740 44660 4788 44662
rect 4844 44660 4892 44716
rect 4268 44650 4948 44660
rect 5404 43764 5460 43774
rect 5740 43764 5796 45278
rect 5404 43762 5796 43764
rect 5404 43710 5406 43762
rect 5458 43710 5796 43762
rect 5404 43708 5796 43710
rect 5404 43698 5460 43708
rect 5740 43652 5796 43708
rect 5740 43586 5796 43596
rect 2940 43486 2942 43538
rect 2994 43486 2996 43538
rect 2492 43474 2548 43484
rect 2940 43474 2996 43486
rect 4268 43148 4948 43158
rect 4324 43092 4372 43148
rect 4428 43146 4476 43148
rect 4532 43146 4580 43148
rect 4448 43094 4476 43146
rect 4572 43094 4580 43146
rect 4428 43092 4476 43094
rect 4532 43092 4580 43094
rect 4636 43146 4684 43148
rect 4740 43146 4788 43148
rect 4636 43094 4644 43146
rect 4740 43094 4768 43146
rect 4636 43092 4684 43094
rect 4740 43092 4788 43094
rect 4844 43092 4892 43148
rect 2156 43036 3108 43092
rect 4268 43082 4948 43092
rect 2044 42812 2660 42868
rect 2044 42530 2100 42542
rect 2044 42478 2046 42530
rect 2098 42478 2100 42530
rect 2044 41412 2100 42478
rect 2492 42530 2548 42542
rect 2492 42478 2494 42530
rect 2546 42478 2548 42530
rect 2492 42196 2548 42478
rect 2492 42130 2548 42140
rect 2044 41346 2100 41356
rect 2156 41858 2212 41870
rect 2156 41806 2158 41858
rect 2210 41806 2212 41858
rect 2156 41076 2212 41806
rect 2380 41076 2436 41086
rect 2156 41020 2380 41076
rect 2380 40982 2436 41020
rect 2044 40962 2100 40974
rect 2044 40910 2046 40962
rect 2098 40910 2100 40962
rect 2044 40628 2100 40910
rect 2044 40572 2548 40628
rect 2156 40404 2212 40414
rect 1932 40402 2212 40404
rect 1932 40350 2158 40402
rect 2210 40350 2212 40402
rect 1932 40348 2212 40350
rect 2156 40338 2212 40348
rect 1820 39788 2436 39844
rect 1820 39618 1876 39630
rect 1820 39566 1822 39618
rect 1874 39566 1876 39618
rect 1820 38836 1876 39566
rect 2380 39506 2436 39788
rect 2380 39454 2382 39506
rect 2434 39454 2436 39506
rect 2380 39442 2436 39454
rect 2044 39396 2100 39406
rect 2044 39302 2100 39340
rect 2492 39284 2548 40572
rect 1820 38742 1876 38780
rect 2268 39228 2548 39284
rect 1708 37938 1764 37950
rect 1708 37886 1710 37938
rect 1762 37886 1764 37938
rect 1708 37716 1764 37886
rect 2044 37828 2100 37838
rect 1708 37650 1764 37660
rect 1932 37826 2100 37828
rect 1932 37774 2046 37826
rect 2098 37774 2100 37826
rect 1932 37772 2100 37774
rect 1820 37154 1876 37166
rect 1820 37102 1822 37154
rect 1874 37102 1876 37154
rect 1708 36596 1764 36606
rect 1708 36482 1764 36540
rect 1708 36430 1710 36482
rect 1762 36430 1764 36482
rect 1708 36418 1764 36430
rect 1708 35700 1764 35710
rect 1820 35700 1876 37102
rect 1708 35698 1876 35700
rect 1708 35646 1710 35698
rect 1762 35646 1876 35698
rect 1708 35644 1876 35646
rect 1708 35476 1764 35644
rect 1708 35410 1764 35420
rect 1708 34802 1764 34814
rect 1708 34750 1710 34802
rect 1762 34750 1764 34802
rect 1708 34356 1764 34750
rect 1708 34290 1764 34300
rect 1820 34468 1876 34478
rect 1932 34468 1988 37772
rect 2044 37762 2100 37772
rect 2044 36260 2100 36270
rect 2044 36258 2212 36260
rect 2044 36206 2046 36258
rect 2098 36206 2212 36258
rect 2044 36204 2212 36206
rect 2044 36194 2100 36204
rect 2044 35812 2100 35822
rect 2044 35718 2100 35756
rect 2156 34916 2212 36204
rect 2156 34850 2212 34860
rect 2044 34692 2100 34702
rect 2044 34598 2100 34636
rect 1932 34412 2100 34468
rect 1820 34130 1876 34412
rect 1820 34078 1822 34130
rect 1874 34078 1876 34130
rect 1820 34066 1876 34078
rect 2044 33348 2100 34412
rect 2268 34130 2324 39228
rect 2380 38946 2436 38958
rect 2380 38894 2382 38946
rect 2434 38894 2436 38946
rect 2380 37266 2436 38894
rect 2492 37826 2548 37838
rect 2492 37774 2494 37826
rect 2546 37774 2548 37826
rect 2492 37716 2548 37774
rect 2492 37650 2548 37660
rect 2380 37214 2382 37266
rect 2434 37214 2436 37266
rect 2380 37202 2436 37214
rect 2604 37268 2660 42812
rect 2940 42532 2996 42542
rect 2828 42530 2996 42532
rect 2828 42478 2942 42530
rect 2994 42478 2996 42530
rect 2828 42476 2996 42478
rect 2828 41970 2884 42476
rect 2940 42466 2996 42476
rect 2828 41918 2830 41970
rect 2882 41918 2884 41970
rect 2828 41906 2884 41918
rect 3052 41972 3108 43036
rect 5740 42196 5796 42206
rect 5852 42196 5908 47852
rect 8540 49586 9044 49588
rect 8540 49534 8990 49586
rect 9042 49534 9044 49586
rect 8540 49532 9044 49534
rect 8540 46900 8596 49532
rect 8988 49522 9044 49532
rect 8988 49028 9044 49038
rect 9100 49028 9156 49868
rect 9548 49858 9604 49868
rect 10108 49924 10164 49934
rect 10108 49830 10164 49868
rect 11340 49924 11396 49934
rect 11340 49830 11396 49868
rect 11676 49810 11732 51436
rect 11900 51426 11956 51436
rect 11676 49758 11678 49810
rect 11730 49758 11732 49810
rect 11676 49746 11732 49758
rect 12124 49810 12180 56140
rect 19068 55972 19124 59200
rect 26768 56476 27448 56486
rect 26824 56420 26872 56476
rect 26928 56474 26976 56476
rect 27032 56474 27080 56476
rect 26948 56422 26976 56474
rect 27072 56422 27080 56474
rect 26928 56420 26976 56422
rect 27032 56420 27080 56422
rect 27136 56474 27184 56476
rect 27240 56474 27288 56476
rect 27136 56422 27144 56474
rect 27240 56422 27268 56474
rect 27136 56420 27184 56422
rect 27240 56420 27288 56422
rect 27344 56420 27392 56476
rect 26768 56410 27448 56420
rect 31388 56308 31444 59200
rect 43708 56642 43764 59200
rect 43708 56590 43710 56642
rect 43762 56590 43764 56642
rect 43708 56578 43764 56590
rect 44380 56642 44436 56654
rect 44380 56590 44382 56642
rect 44434 56590 44436 56642
rect 35768 56476 36448 56486
rect 35824 56420 35872 56476
rect 35928 56474 35976 56476
rect 36032 56474 36080 56476
rect 35948 56422 35976 56474
rect 36072 56422 36080 56474
rect 35928 56420 35976 56422
rect 36032 56420 36080 56422
rect 36136 56474 36184 56476
rect 36240 56474 36288 56476
rect 36136 56422 36144 56474
rect 36240 56422 36268 56474
rect 36136 56420 36184 56422
rect 36240 56420 36288 56422
rect 36344 56420 36392 56476
rect 35768 56410 36448 56420
rect 31388 56242 31444 56252
rect 32172 56308 32228 56318
rect 32172 56214 32228 56252
rect 20076 56084 20132 56094
rect 20076 55990 20132 56028
rect 25452 56084 25508 56094
rect 32844 56084 32900 56094
rect 43932 56084 43988 56094
rect 19180 55972 19236 55982
rect 19068 55970 19236 55972
rect 19068 55918 19182 55970
rect 19234 55918 19236 55970
rect 19068 55916 19236 55918
rect 19180 55906 19236 55916
rect 13268 55692 13948 55702
rect 13324 55636 13372 55692
rect 13428 55690 13476 55692
rect 13532 55690 13580 55692
rect 13448 55638 13476 55690
rect 13572 55638 13580 55690
rect 13428 55636 13476 55638
rect 13532 55636 13580 55638
rect 13636 55690 13684 55692
rect 13740 55690 13788 55692
rect 13636 55638 13644 55690
rect 13740 55638 13768 55690
rect 13636 55636 13684 55638
rect 13740 55636 13788 55638
rect 13844 55636 13892 55692
rect 13268 55626 13948 55636
rect 22268 55692 22948 55702
rect 22324 55636 22372 55692
rect 22428 55690 22476 55692
rect 22532 55690 22580 55692
rect 22448 55638 22476 55690
rect 22572 55638 22580 55690
rect 22428 55636 22476 55638
rect 22532 55636 22580 55638
rect 22636 55690 22684 55692
rect 22740 55690 22788 55692
rect 22636 55638 22644 55690
rect 22740 55638 22768 55690
rect 22636 55636 22684 55638
rect 22740 55636 22788 55638
rect 22844 55636 22892 55692
rect 22268 55626 22948 55636
rect 25452 55186 25508 56028
rect 32396 56082 32900 56084
rect 32396 56030 32846 56082
rect 32898 56030 32900 56082
rect 32396 56028 32900 56030
rect 26124 55972 26180 55982
rect 25452 55134 25454 55186
rect 25506 55134 25508 55186
rect 25452 55122 25508 55134
rect 25788 55186 25844 55198
rect 25788 55134 25790 55186
rect 25842 55134 25844 55186
rect 17768 54908 18448 54918
rect 17824 54852 17872 54908
rect 17928 54906 17976 54908
rect 18032 54906 18080 54908
rect 17948 54854 17976 54906
rect 18072 54854 18080 54906
rect 17928 54852 17976 54854
rect 18032 54852 18080 54854
rect 18136 54906 18184 54908
rect 18240 54906 18288 54908
rect 18136 54854 18144 54906
rect 18240 54854 18268 54906
rect 18136 54852 18184 54854
rect 18240 54852 18288 54854
rect 18344 54852 18392 54908
rect 17768 54842 18448 54852
rect 13268 54124 13948 54134
rect 13324 54068 13372 54124
rect 13428 54122 13476 54124
rect 13532 54122 13580 54124
rect 13448 54070 13476 54122
rect 13572 54070 13580 54122
rect 13428 54068 13476 54070
rect 13532 54068 13580 54070
rect 13636 54122 13684 54124
rect 13740 54122 13788 54124
rect 13636 54070 13644 54122
rect 13740 54070 13768 54122
rect 13636 54068 13684 54070
rect 13740 54068 13788 54070
rect 13844 54068 13892 54124
rect 13268 54058 13948 54068
rect 22268 54124 22948 54134
rect 22324 54068 22372 54124
rect 22428 54122 22476 54124
rect 22532 54122 22580 54124
rect 22448 54070 22476 54122
rect 22572 54070 22580 54122
rect 22428 54068 22476 54070
rect 22532 54068 22580 54070
rect 22636 54122 22684 54124
rect 22740 54122 22788 54124
rect 22636 54070 22644 54122
rect 22740 54070 22768 54122
rect 22636 54068 22684 54070
rect 22740 54068 22788 54070
rect 22844 54068 22892 54124
rect 22268 54058 22948 54068
rect 17768 53340 18448 53350
rect 17824 53284 17872 53340
rect 17928 53338 17976 53340
rect 18032 53338 18080 53340
rect 17948 53286 17976 53338
rect 18072 53286 18080 53338
rect 17928 53284 17976 53286
rect 18032 53284 18080 53286
rect 18136 53338 18184 53340
rect 18240 53338 18288 53340
rect 18136 53286 18144 53338
rect 18240 53286 18268 53338
rect 18136 53284 18184 53286
rect 18240 53284 18288 53286
rect 18344 53284 18392 53340
rect 17768 53274 18448 53284
rect 25788 53060 25844 55134
rect 26124 55186 26180 55916
rect 31268 55692 31948 55702
rect 31324 55636 31372 55692
rect 31428 55690 31476 55692
rect 31532 55690 31580 55692
rect 31448 55638 31476 55690
rect 31572 55638 31580 55690
rect 31428 55636 31476 55638
rect 31532 55636 31580 55638
rect 31636 55690 31684 55692
rect 31740 55690 31788 55692
rect 31636 55638 31644 55690
rect 31740 55638 31768 55690
rect 31636 55636 31684 55638
rect 31740 55636 31788 55638
rect 31844 55636 31892 55692
rect 31268 55626 31948 55636
rect 32060 55410 32116 55422
rect 32060 55358 32062 55410
rect 32114 55358 32116 55410
rect 29260 55300 29316 55310
rect 29260 55206 29316 55244
rect 26124 55134 26126 55186
rect 26178 55134 26180 55186
rect 26124 55122 26180 55134
rect 26460 55188 26516 55198
rect 29932 55188 29988 55198
rect 26460 55186 26628 55188
rect 26460 55134 26462 55186
rect 26514 55134 26628 55186
rect 26460 55132 26628 55134
rect 26460 55122 26516 55132
rect 26572 53172 26628 55132
rect 29932 55186 30100 55188
rect 29932 55134 29934 55186
rect 29986 55134 30100 55186
rect 29932 55132 30100 55134
rect 29932 55122 29988 55132
rect 26768 54908 27448 54918
rect 26824 54852 26872 54908
rect 26928 54906 26976 54908
rect 27032 54906 27080 54908
rect 26948 54854 26976 54906
rect 27072 54854 27080 54906
rect 26928 54852 26976 54854
rect 27032 54852 27080 54854
rect 27136 54906 27184 54908
rect 27240 54906 27288 54908
rect 27136 54854 27144 54906
rect 27240 54854 27268 54906
rect 27136 54852 27184 54854
rect 27240 54852 27288 54854
rect 27344 54852 27392 54908
rect 26768 54842 27448 54852
rect 28476 53956 28532 53966
rect 28476 53732 28532 53900
rect 30044 53842 30100 55132
rect 31268 54124 31948 54134
rect 31324 54068 31372 54124
rect 31428 54122 31476 54124
rect 31532 54122 31580 54124
rect 31448 54070 31476 54122
rect 31572 54070 31580 54122
rect 31428 54068 31476 54070
rect 31532 54068 31580 54070
rect 31636 54122 31684 54124
rect 31740 54122 31788 54124
rect 31636 54070 31644 54122
rect 31740 54070 31768 54122
rect 31636 54068 31684 54070
rect 31740 54068 31788 54070
rect 31844 54068 31892 54124
rect 31268 54058 31948 54068
rect 30044 53790 30046 53842
rect 30098 53790 30100 53842
rect 30044 53778 30100 53790
rect 28252 53730 28532 53732
rect 28252 53678 28478 53730
rect 28530 53678 28532 53730
rect 28252 53676 28532 53678
rect 26768 53340 27448 53350
rect 26824 53284 26872 53340
rect 26928 53338 26976 53340
rect 27032 53338 27080 53340
rect 26948 53286 26976 53338
rect 27072 53286 27080 53338
rect 26928 53284 26976 53286
rect 27032 53284 27080 53286
rect 27136 53338 27184 53340
rect 27240 53338 27288 53340
rect 27136 53286 27144 53338
rect 27240 53286 27268 53338
rect 27136 53284 27184 53286
rect 27240 53284 27288 53286
rect 27344 53284 27392 53340
rect 26768 53274 27448 53284
rect 26572 53116 27188 53172
rect 25788 52994 25844 53004
rect 25116 52836 25172 52846
rect 13268 52556 13948 52566
rect 13324 52500 13372 52556
rect 13428 52554 13476 52556
rect 13532 52554 13580 52556
rect 13448 52502 13476 52554
rect 13572 52502 13580 52554
rect 13428 52500 13476 52502
rect 13532 52500 13580 52502
rect 13636 52554 13684 52556
rect 13740 52554 13788 52556
rect 13636 52502 13644 52554
rect 13740 52502 13768 52554
rect 13636 52500 13684 52502
rect 13740 52500 13788 52502
rect 13844 52500 13892 52556
rect 13268 52490 13948 52500
rect 22268 52556 22948 52566
rect 22324 52500 22372 52556
rect 22428 52554 22476 52556
rect 22532 52554 22580 52556
rect 22448 52502 22476 52554
rect 22572 52502 22580 52554
rect 22428 52500 22476 52502
rect 22532 52500 22580 52502
rect 22636 52554 22684 52556
rect 22740 52554 22788 52556
rect 22636 52502 22644 52554
rect 22740 52502 22768 52554
rect 22636 52500 22684 52502
rect 22740 52500 22788 52502
rect 22844 52500 22892 52556
rect 22268 52490 22948 52500
rect 22988 52276 23044 52286
rect 22988 52182 23044 52220
rect 25116 52274 25172 52780
rect 25116 52222 25118 52274
rect 25170 52222 25172 52274
rect 25116 52210 25172 52222
rect 25900 52164 25956 52174
rect 26348 52164 26404 52174
rect 25900 52162 26404 52164
rect 25900 52110 25902 52162
rect 25954 52110 26350 52162
rect 26402 52110 26404 52162
rect 25900 52108 26404 52110
rect 25900 52098 25956 52108
rect 26236 51940 26292 51950
rect 17768 51772 18448 51782
rect 17824 51716 17872 51772
rect 17928 51770 17976 51772
rect 18032 51770 18080 51772
rect 17948 51718 17976 51770
rect 18072 51718 18080 51770
rect 17928 51716 17976 51718
rect 18032 51716 18080 51718
rect 18136 51770 18184 51772
rect 18240 51770 18288 51772
rect 18136 51718 18144 51770
rect 18240 51718 18268 51770
rect 18136 51716 18184 51718
rect 18240 51716 18288 51718
rect 18344 51716 18392 51772
rect 17768 51706 18448 51716
rect 13268 50988 13948 50998
rect 13324 50932 13372 50988
rect 13428 50986 13476 50988
rect 13532 50986 13580 50988
rect 13448 50934 13476 50986
rect 13572 50934 13580 50986
rect 13428 50932 13476 50934
rect 13532 50932 13580 50934
rect 13636 50986 13684 50988
rect 13740 50986 13788 50988
rect 13636 50934 13644 50986
rect 13740 50934 13768 50986
rect 13636 50932 13684 50934
rect 13740 50932 13788 50934
rect 13844 50932 13892 50988
rect 13268 50922 13948 50932
rect 22268 50988 22948 50998
rect 22324 50932 22372 50988
rect 22428 50986 22476 50988
rect 22532 50986 22580 50988
rect 22448 50934 22476 50986
rect 22572 50934 22580 50986
rect 22428 50932 22476 50934
rect 22532 50932 22580 50934
rect 22636 50986 22684 50988
rect 22740 50986 22788 50988
rect 22636 50934 22644 50986
rect 22740 50934 22768 50986
rect 22636 50932 22684 50934
rect 22740 50932 22788 50934
rect 22844 50932 22892 50988
rect 22268 50922 22948 50932
rect 16716 50596 16772 50606
rect 16492 50594 16772 50596
rect 16492 50542 16718 50594
rect 16770 50542 16772 50594
rect 16492 50540 16772 50542
rect 16156 50484 16212 50494
rect 16156 50390 16212 50428
rect 16492 50370 16548 50540
rect 16716 50530 16772 50540
rect 17276 50594 17332 50606
rect 17276 50542 17278 50594
rect 17330 50542 17332 50594
rect 17276 50484 17332 50542
rect 17276 50418 17332 50428
rect 19628 50484 19684 50494
rect 19628 50390 19684 50428
rect 20524 50484 20580 50494
rect 16492 50318 16494 50370
rect 16546 50318 16548 50370
rect 16492 50306 16548 50318
rect 20412 50370 20468 50382
rect 20412 50318 20414 50370
rect 20466 50318 20468 50370
rect 17768 50204 18448 50214
rect 17824 50148 17872 50204
rect 17928 50202 17976 50204
rect 18032 50202 18080 50204
rect 17948 50150 17976 50202
rect 18072 50150 18080 50202
rect 17928 50148 17976 50150
rect 18032 50148 18080 50150
rect 18136 50202 18184 50204
rect 18240 50202 18288 50204
rect 18136 50150 18144 50202
rect 18240 50150 18268 50202
rect 18136 50148 18184 50150
rect 18240 50148 18288 50150
rect 18344 50148 18392 50204
rect 17768 50138 18448 50148
rect 14476 49924 14532 49934
rect 14476 49830 14532 49868
rect 12124 49758 12126 49810
rect 12178 49758 12180 49810
rect 12124 49746 12180 49758
rect 15260 49588 15316 49598
rect 15260 49586 15652 49588
rect 15260 49534 15262 49586
rect 15314 49534 15652 49586
rect 15260 49532 15652 49534
rect 15260 49522 15316 49532
rect 13268 49420 13948 49430
rect 13324 49364 13372 49420
rect 13428 49418 13476 49420
rect 13532 49418 13580 49420
rect 13448 49366 13476 49418
rect 13572 49366 13580 49418
rect 13428 49364 13476 49366
rect 13532 49364 13580 49366
rect 13636 49418 13684 49420
rect 13740 49418 13788 49420
rect 13636 49366 13644 49418
rect 13740 49366 13768 49418
rect 13636 49364 13684 49366
rect 13740 49364 13788 49366
rect 13844 49364 13892 49420
rect 13268 49354 13948 49364
rect 8988 49026 9156 49028
rect 8988 48974 8990 49026
rect 9042 48974 9156 49026
rect 8988 48972 9156 48974
rect 9324 49028 9380 49038
rect 8988 48962 9044 48972
rect 9324 48934 9380 48972
rect 11676 48802 11732 48814
rect 11676 48750 11678 48802
rect 11730 48750 11732 48802
rect 8768 48636 9448 48646
rect 8824 48580 8872 48636
rect 8928 48634 8976 48636
rect 9032 48634 9080 48636
rect 8948 48582 8976 48634
rect 9072 48582 9080 48634
rect 8928 48580 8976 48582
rect 9032 48580 9080 48582
rect 9136 48634 9184 48636
rect 9240 48634 9288 48636
rect 9136 48582 9144 48634
rect 9240 48582 9268 48634
rect 9136 48580 9184 48582
rect 9240 48580 9288 48582
rect 9344 48580 9392 48636
rect 8768 48570 9448 48580
rect 9660 48020 9716 48030
rect 9660 47346 9716 47964
rect 9660 47294 9662 47346
rect 9714 47294 9716 47346
rect 9660 47282 9716 47294
rect 10108 47460 10164 47470
rect 8764 47236 8820 47246
rect 8540 46834 8596 46844
rect 8652 47180 8764 47236
rect 8652 46786 8708 47180
rect 8764 47170 8820 47180
rect 9100 47236 9156 47246
rect 9100 47234 9604 47236
rect 9100 47182 9102 47234
rect 9154 47182 9604 47234
rect 9100 47180 9604 47182
rect 9100 47170 9156 47180
rect 8768 47068 9448 47078
rect 8824 47012 8872 47068
rect 8928 47066 8976 47068
rect 9032 47066 9080 47068
rect 8948 47014 8976 47066
rect 9072 47014 9080 47066
rect 8928 47012 8976 47014
rect 9032 47012 9080 47014
rect 9136 47066 9184 47068
rect 9240 47066 9288 47068
rect 9136 47014 9144 47066
rect 9240 47014 9268 47066
rect 9136 47012 9184 47014
rect 9240 47012 9288 47014
rect 9344 47012 9392 47068
rect 8768 47002 9448 47012
rect 8652 46734 8654 46786
rect 8706 46734 8708 46786
rect 8652 46722 8708 46734
rect 8988 46786 9044 46798
rect 8988 46734 8990 46786
rect 9042 46734 9044 46786
rect 8988 46676 9044 46734
rect 8988 46610 9044 46620
rect 9548 46674 9604 47180
rect 9548 46622 9550 46674
rect 9602 46622 9604 46674
rect 9548 46610 9604 46622
rect 9996 46676 10052 46686
rect 9996 46582 10052 46620
rect 5964 46450 6020 46462
rect 5964 46398 5966 46450
rect 6018 46398 6020 46450
rect 5964 45220 6020 46398
rect 8768 45500 9448 45510
rect 8824 45444 8872 45500
rect 8928 45498 8976 45500
rect 9032 45498 9080 45500
rect 8948 45446 8976 45498
rect 9072 45446 9080 45498
rect 8928 45444 8976 45446
rect 9032 45444 9080 45446
rect 9136 45498 9184 45500
rect 9240 45498 9288 45500
rect 9136 45446 9144 45498
rect 9240 45446 9268 45498
rect 9136 45444 9184 45446
rect 9240 45444 9288 45446
rect 9344 45444 9392 45500
rect 8768 45434 9448 45444
rect 5964 45154 6020 45164
rect 6524 44882 6580 44894
rect 6524 44830 6526 44882
rect 6578 44830 6580 44882
rect 6524 44548 6580 44830
rect 6524 44482 6580 44492
rect 8764 44324 8820 44334
rect 9436 44324 9492 44334
rect 8764 44322 9492 44324
rect 8764 44270 8766 44322
rect 8818 44270 9438 44322
rect 9490 44270 9492 44322
rect 8764 44268 9492 44270
rect 8764 44258 8820 44268
rect 9436 44258 9492 44268
rect 9772 44324 9828 44334
rect 10108 44324 10164 47404
rect 10444 47460 10500 47470
rect 10444 47366 10500 47404
rect 9772 44230 9828 44268
rect 9996 44268 10164 44324
rect 10220 47348 10276 47358
rect 10220 44322 10276 47292
rect 11340 47348 11396 47358
rect 11340 47254 11396 47292
rect 10780 47236 10836 47246
rect 10780 47142 10836 47180
rect 10220 44270 10222 44322
rect 10274 44270 10276 44322
rect 7196 44212 7252 44222
rect 6300 43652 6356 43662
rect 6300 43426 6356 43596
rect 6300 43374 6302 43426
rect 6354 43374 6356 43426
rect 6300 43362 6356 43374
rect 6748 43652 6804 43662
rect 7196 43652 7252 44156
rect 8316 44098 8372 44110
rect 8316 44046 8318 44098
rect 8370 44046 8372 44098
rect 8316 43764 8372 44046
rect 8988 44100 9044 44138
rect 8988 44034 9044 44044
rect 9772 44100 9828 44110
rect 8768 43932 9448 43942
rect 8824 43876 8872 43932
rect 8928 43930 8976 43932
rect 9032 43930 9080 43932
rect 8948 43878 8976 43930
rect 9072 43878 9080 43930
rect 8928 43876 8976 43878
rect 9032 43876 9080 43878
rect 9136 43930 9184 43932
rect 9240 43930 9288 43932
rect 9136 43878 9144 43930
rect 9240 43878 9268 43930
rect 9136 43876 9184 43878
rect 9240 43876 9288 43878
rect 9344 43876 9392 43932
rect 8768 43866 9448 43876
rect 8316 43698 8372 43708
rect 9436 43764 9492 43774
rect 6748 43650 7252 43652
rect 6748 43598 6750 43650
rect 6802 43598 7198 43650
rect 7250 43598 7252 43650
rect 6748 43596 7252 43598
rect 5964 43316 6020 43326
rect 5964 43222 6020 43260
rect 6188 42196 6244 42206
rect 5740 42194 5908 42196
rect 5740 42142 5742 42194
rect 5794 42142 5908 42194
rect 5740 42140 5908 42142
rect 6076 42140 6188 42196
rect 3164 41972 3220 41982
rect 3052 41970 3220 41972
rect 3052 41918 3166 41970
rect 3218 41918 3220 41970
rect 3052 41916 3220 41918
rect 3164 41906 3220 41916
rect 4268 41580 4948 41590
rect 4324 41524 4372 41580
rect 4428 41578 4476 41580
rect 4532 41578 4580 41580
rect 4448 41526 4476 41578
rect 4572 41526 4580 41578
rect 4428 41524 4476 41526
rect 4532 41524 4580 41526
rect 4636 41578 4684 41580
rect 4740 41578 4788 41580
rect 4636 41526 4644 41578
rect 4740 41526 4768 41578
rect 4636 41524 4684 41526
rect 4740 41524 4788 41526
rect 4844 41524 4892 41580
rect 4268 41514 4948 41524
rect 2716 40964 2772 40974
rect 2716 40962 2884 40964
rect 2716 40910 2718 40962
rect 2770 40910 2884 40962
rect 2716 40908 2884 40910
rect 2716 40898 2772 40908
rect 2716 37268 2772 37278
rect 2604 37266 2772 37268
rect 2604 37214 2718 37266
rect 2770 37214 2772 37266
rect 2604 37212 2772 37214
rect 2716 37202 2772 37212
rect 2716 36258 2772 36270
rect 2716 36206 2718 36258
rect 2770 36206 2772 36258
rect 2380 35812 2436 35822
rect 2436 35756 2660 35812
rect 2380 35746 2436 35756
rect 2380 34690 2436 34702
rect 2380 34638 2382 34690
rect 2434 34638 2436 34690
rect 2380 34468 2436 34638
rect 2380 34402 2436 34412
rect 2268 34078 2270 34130
rect 2322 34078 2324 34130
rect 2268 34066 2324 34078
rect 2044 33292 2212 33348
rect 1708 33236 1764 33246
rect 1708 33142 1764 33180
rect 2044 33124 2100 33134
rect 1820 33122 2100 33124
rect 1820 33070 2046 33122
rect 2098 33070 2100 33122
rect 1820 33068 2100 33070
rect 1708 32562 1764 32574
rect 1708 32510 1710 32562
rect 1762 32510 1764 32562
rect 1708 32116 1764 32510
rect 1708 32050 1764 32060
rect 1820 32004 1876 33068
rect 2044 33058 2100 33068
rect 2156 32900 2212 33292
rect 2492 33236 2548 33246
rect 2492 33142 2548 33180
rect 1820 31938 1876 31948
rect 1932 32844 2212 32900
rect 1708 31666 1764 31678
rect 1708 31614 1710 31666
rect 1762 31614 1764 31666
rect 1708 31556 1764 31614
rect 1708 30996 1764 31500
rect 1708 30930 1764 30940
rect 1820 31220 1876 31230
rect 1820 30994 1876 31164
rect 1820 30942 1822 30994
rect 1874 30942 1876 30994
rect 1820 30930 1876 30942
rect 1932 30996 1988 32844
rect 2044 32674 2100 32686
rect 2044 32622 2046 32674
rect 2098 32622 2100 32674
rect 2044 31892 2100 32622
rect 2492 32450 2548 32462
rect 2492 32398 2494 32450
rect 2546 32398 2548 32450
rect 2492 32116 2548 32398
rect 2492 32050 2548 32060
rect 2044 31836 2324 31892
rect 2268 31780 2324 31836
rect 2604 31780 2660 35756
rect 2716 35698 2772 36206
rect 2716 35646 2718 35698
rect 2770 35646 2772 35698
rect 2716 35634 2772 35646
rect 2828 35700 2884 40908
rect 3164 40962 3220 40974
rect 3164 40910 3166 40962
rect 3218 40910 3220 40962
rect 3164 39956 3220 40910
rect 5740 40964 5796 42140
rect 5964 41412 6020 41422
rect 5740 40962 5908 40964
rect 5740 40910 5742 40962
rect 5794 40910 5908 40962
rect 5740 40908 5908 40910
rect 5740 40898 5796 40908
rect 4732 40628 4788 40638
rect 4732 40534 4788 40572
rect 5852 40628 5908 40908
rect 5628 40402 5684 40414
rect 5628 40350 5630 40402
rect 5682 40350 5684 40402
rect 5292 40178 5348 40190
rect 5292 40126 5294 40178
rect 5346 40126 5348 40178
rect 4268 40012 4948 40022
rect 4324 39956 4372 40012
rect 4428 40010 4476 40012
rect 4532 40010 4580 40012
rect 4448 39958 4476 40010
rect 4572 39958 4580 40010
rect 4428 39956 4476 39958
rect 4532 39956 4580 39958
rect 4636 40010 4684 40012
rect 4740 40010 4788 40012
rect 4636 39958 4644 40010
rect 4740 39958 4768 40010
rect 4636 39956 4684 39958
rect 4740 39956 4788 39958
rect 4844 39956 4892 40012
rect 4268 39946 4948 39956
rect 3164 39890 3220 39900
rect 4268 38444 4948 38454
rect 4324 38388 4372 38444
rect 4428 38442 4476 38444
rect 4532 38442 4580 38444
rect 4448 38390 4476 38442
rect 4572 38390 4580 38442
rect 4428 38388 4476 38390
rect 4532 38388 4580 38390
rect 4636 38442 4684 38444
rect 4740 38442 4788 38444
rect 4636 38390 4644 38442
rect 4740 38390 4768 38442
rect 4636 38388 4684 38390
rect 4740 38388 4788 38390
rect 4844 38388 4892 38444
rect 4268 38378 4948 38388
rect 5292 37828 5348 40126
rect 5628 39506 5684 40350
rect 5628 39454 5630 39506
rect 5682 39454 5684 39506
rect 5628 39442 5684 39454
rect 5852 37828 5908 40572
rect 5964 40402 6020 41356
rect 5964 40350 5966 40402
rect 6018 40350 6020 40402
rect 5964 40338 6020 40350
rect 5964 37828 6020 37838
rect 5852 37826 6020 37828
rect 5852 37774 5966 37826
rect 6018 37774 6020 37826
rect 5852 37772 6020 37774
rect 5292 37762 5348 37772
rect 5068 37378 5124 37390
rect 5068 37326 5070 37378
rect 5122 37326 5124 37378
rect 4268 36876 4948 36886
rect 4324 36820 4372 36876
rect 4428 36874 4476 36876
rect 4532 36874 4580 36876
rect 4448 36822 4476 36874
rect 4572 36822 4580 36874
rect 4428 36820 4476 36822
rect 4532 36820 4580 36822
rect 4636 36874 4684 36876
rect 4740 36874 4788 36876
rect 4636 36822 4644 36874
rect 4740 36822 4768 36874
rect 4636 36820 4684 36822
rect 4740 36820 4788 36822
rect 4844 36820 4892 36876
rect 4268 36810 4948 36820
rect 3276 36596 3332 36606
rect 3276 36502 3332 36540
rect 5068 36260 5124 37326
rect 5852 37380 5908 37390
rect 5852 37286 5908 37324
rect 5068 36194 5124 36204
rect 5628 36260 5684 36270
rect 5628 35922 5684 36204
rect 5964 36260 6020 37772
rect 6076 37378 6132 42140
rect 6188 42130 6244 42140
rect 6748 42196 6804 43596
rect 7196 43558 7252 43596
rect 9436 43538 9492 43708
rect 9772 43708 9828 44044
rect 9996 43876 10052 44268
rect 10220 43988 10276 44270
rect 10332 46900 10388 46910
rect 10332 44210 10388 46844
rect 11676 46788 11732 48750
rect 12460 48804 12516 48814
rect 14476 48804 14532 48814
rect 12460 48710 12516 48748
rect 14140 48802 14532 48804
rect 14140 48750 14478 48802
rect 14530 48750 14532 48802
rect 14140 48748 14532 48750
rect 13580 48356 13636 48366
rect 13580 48262 13636 48300
rect 14028 48244 14084 48254
rect 14028 48150 14084 48188
rect 13268 47852 13948 47862
rect 13324 47796 13372 47852
rect 13428 47850 13476 47852
rect 13532 47850 13580 47852
rect 13448 47798 13476 47850
rect 13572 47798 13580 47850
rect 13428 47796 13476 47798
rect 13532 47796 13580 47798
rect 13636 47850 13684 47852
rect 13740 47850 13788 47852
rect 13636 47798 13644 47850
rect 13740 47798 13768 47850
rect 13636 47796 13684 47798
rect 13740 47796 13788 47798
rect 13844 47796 13892 47852
rect 13268 47786 13948 47796
rect 14140 47458 14196 48748
rect 14476 48738 14532 48748
rect 14924 48804 14980 48814
rect 14140 47406 14142 47458
rect 14194 47406 14196 47458
rect 14140 47394 14196 47406
rect 14252 48354 14308 48366
rect 14252 48302 14254 48354
rect 14306 48302 14308 48354
rect 14252 47460 14308 48302
rect 14924 48354 14980 48748
rect 14924 48302 14926 48354
rect 14978 48302 14980 48354
rect 14924 48290 14980 48302
rect 15036 48356 15092 48366
rect 15036 48242 15092 48300
rect 15036 48190 15038 48242
rect 15090 48190 15092 48242
rect 14700 47460 14756 47470
rect 14252 47458 14756 47460
rect 14252 47406 14702 47458
rect 14754 47406 14756 47458
rect 14252 47404 14756 47406
rect 14700 47394 14756 47404
rect 11788 47236 11844 47246
rect 11788 47142 11844 47180
rect 13132 47236 13188 47246
rect 12348 46788 12404 46798
rect 11676 46786 12404 46788
rect 11676 46734 12350 46786
rect 12402 46734 12404 46786
rect 11676 46732 12404 46734
rect 11564 44324 11620 44334
rect 11564 44230 11620 44268
rect 10332 44158 10334 44210
rect 10386 44158 10388 44210
rect 10332 44146 10388 44158
rect 11116 44098 11172 44110
rect 11116 44046 11118 44098
rect 11170 44046 11172 44098
rect 10220 43932 10500 43988
rect 9996 43820 10276 43876
rect 9772 43652 10164 43708
rect 9436 43486 9438 43538
rect 9490 43486 9492 43538
rect 9436 43474 9492 43486
rect 10108 43538 10164 43652
rect 10108 43486 10110 43538
rect 10162 43486 10164 43538
rect 10108 43474 10164 43486
rect 8768 42364 9448 42374
rect 8824 42308 8872 42364
rect 8928 42362 8976 42364
rect 9032 42362 9080 42364
rect 8948 42310 8976 42362
rect 9072 42310 9080 42362
rect 8928 42308 8976 42310
rect 9032 42308 9080 42310
rect 9136 42362 9184 42364
rect 9240 42362 9288 42364
rect 9136 42310 9144 42362
rect 9240 42310 9268 42362
rect 9136 42308 9184 42310
rect 9240 42308 9288 42310
rect 9344 42308 9392 42364
rect 8768 42298 9448 42308
rect 6748 42130 6804 42140
rect 6636 41858 6692 41870
rect 6636 41806 6638 41858
rect 6690 41806 6692 41858
rect 6300 41748 6356 41758
rect 6300 41654 6356 41692
rect 6636 40628 6692 41806
rect 8876 41132 9604 41188
rect 8876 41074 8932 41132
rect 8876 41022 8878 41074
rect 8930 41022 8932 41074
rect 8876 41010 8932 41022
rect 9324 40964 9380 41002
rect 9324 40898 9380 40908
rect 8768 40796 9448 40806
rect 8824 40740 8872 40796
rect 8928 40794 8976 40796
rect 9032 40794 9080 40796
rect 8948 40742 8976 40794
rect 9072 40742 9080 40794
rect 8928 40740 8976 40742
rect 9032 40740 9080 40742
rect 9136 40794 9184 40796
rect 9240 40794 9288 40796
rect 9136 40742 9144 40794
rect 9240 40742 9268 40794
rect 9136 40740 9184 40742
rect 9240 40740 9288 40742
rect 9344 40740 9392 40796
rect 8768 40730 9448 40740
rect 6636 40562 6692 40572
rect 8316 40628 8372 40638
rect 8316 40534 8372 40572
rect 9548 40402 9604 41132
rect 9548 40350 9550 40402
rect 9602 40350 9604 40402
rect 9548 40338 9604 40350
rect 9660 40964 9716 40974
rect 9100 40178 9156 40190
rect 9660 40180 9716 40908
rect 10108 40404 10164 40414
rect 10220 40404 10276 43820
rect 10444 43708 10500 43932
rect 11116 43708 11172 44046
rect 10108 40402 10276 40404
rect 10108 40350 10110 40402
rect 10162 40350 10276 40402
rect 10108 40348 10276 40350
rect 10332 43652 11172 43708
rect 12348 43652 12404 46732
rect 13132 46450 13188 47180
rect 13132 46398 13134 46450
rect 13186 46398 13188 46450
rect 13132 46004 13188 46398
rect 13268 46284 13948 46294
rect 13324 46228 13372 46284
rect 13428 46282 13476 46284
rect 13532 46282 13580 46284
rect 13448 46230 13476 46282
rect 13572 46230 13580 46282
rect 13428 46228 13476 46230
rect 13532 46228 13580 46230
rect 13636 46282 13684 46284
rect 13740 46282 13788 46284
rect 13636 46230 13644 46282
rect 13740 46230 13768 46282
rect 13636 46228 13684 46230
rect 13740 46228 13788 46230
rect 13844 46228 13892 46284
rect 13268 46218 13948 46228
rect 13244 46004 13300 46014
rect 13132 45948 13244 46004
rect 13244 45938 13300 45948
rect 14924 46004 14980 46014
rect 15036 46004 15092 48190
rect 15484 48020 15540 48030
rect 15484 47926 15540 47964
rect 14924 46002 15092 46004
rect 14924 45950 14926 46002
rect 14978 45950 15092 46002
rect 14924 45948 15092 45950
rect 14924 45938 14980 45948
rect 14252 45218 14308 45230
rect 14252 45166 14254 45218
rect 14306 45166 14308 45218
rect 13268 44716 13948 44726
rect 13324 44660 13372 44716
rect 13428 44714 13476 44716
rect 13532 44714 13580 44716
rect 13448 44662 13476 44714
rect 13572 44662 13580 44714
rect 13428 44660 13476 44662
rect 13532 44660 13580 44662
rect 13636 44714 13684 44716
rect 13740 44714 13788 44716
rect 13636 44662 13644 44714
rect 13740 44662 13768 44714
rect 13636 44660 13684 44662
rect 13740 44660 13788 44662
rect 13844 44660 13892 44716
rect 13268 44650 13948 44660
rect 10332 42532 10388 43652
rect 12348 43558 12404 43596
rect 13132 44324 13188 44334
rect 13132 43314 13188 44268
rect 14252 44322 14308 45166
rect 14252 44270 14254 44322
rect 14306 44270 14308 44322
rect 14252 44258 14308 44270
rect 14588 45218 14644 45230
rect 14588 45166 14590 45218
rect 14642 45166 14644 45218
rect 14588 44324 14644 45166
rect 14924 45108 14980 45118
rect 15036 45108 15092 45948
rect 15484 45220 15540 45230
rect 15484 45126 15540 45164
rect 15372 45108 15428 45118
rect 15036 45106 15428 45108
rect 15036 45054 15374 45106
rect 15426 45054 15428 45106
rect 15036 45052 15428 45054
rect 14924 45014 14980 45052
rect 14812 44324 14868 44334
rect 14588 44322 14868 44324
rect 14588 44270 14814 44322
rect 14866 44270 14868 44322
rect 14588 44268 14868 44270
rect 14812 44258 14868 44268
rect 14028 44212 14084 44222
rect 14028 44118 14084 44156
rect 13916 43652 13972 43662
rect 13916 43650 14084 43652
rect 13916 43598 13918 43650
rect 13970 43598 14084 43650
rect 13916 43596 14084 43598
rect 13916 43586 13972 43596
rect 13132 43262 13134 43314
rect 13186 43262 13188 43314
rect 12684 42754 12740 42766
rect 12684 42702 12686 42754
rect 12738 42702 12740 42754
rect 12684 42644 12740 42702
rect 12684 42578 12740 42588
rect 10108 40338 10164 40348
rect 9100 40126 9102 40178
rect 9154 40126 9156 40178
rect 9100 39620 9156 40126
rect 9212 40124 9716 40180
rect 9212 39730 9268 40124
rect 9212 39678 9214 39730
rect 9266 39678 9268 39730
rect 9212 39666 9268 39678
rect 9100 39554 9156 39564
rect 8768 39228 9448 39238
rect 8824 39172 8872 39228
rect 8928 39226 8976 39228
rect 9032 39226 9080 39228
rect 8948 39174 8976 39226
rect 9072 39174 9080 39226
rect 8928 39172 8976 39174
rect 9032 39172 9080 39174
rect 9136 39226 9184 39228
rect 9240 39226 9288 39228
rect 9136 39174 9144 39226
rect 9240 39174 9268 39226
rect 9136 39172 9184 39174
rect 9240 39172 9288 39174
rect 9344 39172 9392 39228
rect 8768 39162 9448 39172
rect 8768 37660 9448 37670
rect 8824 37604 8872 37660
rect 8928 37658 8976 37660
rect 9032 37658 9080 37660
rect 8948 37606 8976 37658
rect 9072 37606 9080 37658
rect 8928 37604 8976 37606
rect 9032 37604 9080 37606
rect 9136 37658 9184 37660
rect 9240 37658 9288 37660
rect 9136 37606 9144 37658
rect 9240 37606 9268 37658
rect 9136 37604 9184 37606
rect 9240 37604 9288 37606
rect 9344 37604 9392 37660
rect 8768 37594 9448 37604
rect 6076 37326 6078 37378
rect 6130 37326 6132 37378
rect 6076 37044 6132 37326
rect 7308 37492 7364 37502
rect 6076 36978 6132 36988
rect 6524 37266 6580 37278
rect 6524 37214 6526 37266
rect 6578 37214 6580 37266
rect 6524 37156 6580 37214
rect 7084 37156 7140 37166
rect 6524 37154 7140 37156
rect 6524 37102 7086 37154
rect 7138 37102 7140 37154
rect 6524 37100 7140 37102
rect 5964 36194 6020 36204
rect 6300 36260 6356 36270
rect 6300 36166 6356 36204
rect 5628 35870 5630 35922
rect 5682 35870 5684 35922
rect 5628 35858 5684 35870
rect 3052 35700 3108 35710
rect 2828 35698 3108 35700
rect 2828 35646 3054 35698
rect 3106 35646 3108 35698
rect 2828 35644 3108 35646
rect 3052 35634 3108 35644
rect 6188 35700 6244 35710
rect 6188 35606 6244 35644
rect 4268 35308 4948 35318
rect 4324 35252 4372 35308
rect 4428 35306 4476 35308
rect 4532 35306 4580 35308
rect 4448 35254 4476 35306
rect 4572 35254 4580 35306
rect 4428 35252 4476 35254
rect 4532 35252 4580 35254
rect 4636 35306 4684 35308
rect 4740 35306 4788 35308
rect 4636 35254 4644 35306
rect 4740 35254 4768 35306
rect 4636 35252 4684 35254
rect 4740 35252 4788 35254
rect 4844 35252 4892 35308
rect 4268 35242 4948 35252
rect 5516 34916 5572 34926
rect 5068 34914 5572 34916
rect 5068 34862 5518 34914
rect 5570 34862 5572 34914
rect 5068 34860 5572 34862
rect 5068 34802 5124 34860
rect 5516 34850 5572 34860
rect 6076 34916 6132 34926
rect 6076 34822 6132 34860
rect 5068 34750 5070 34802
rect 5122 34750 5124 34802
rect 5068 34738 5124 34750
rect 2268 31724 2548 31780
rect 2044 31612 2212 31668
rect 2044 31554 2100 31612
rect 2044 31502 2046 31554
rect 2098 31502 2100 31554
rect 2044 31490 2100 31502
rect 2156 31444 2212 31612
rect 2380 31554 2436 31566
rect 2380 31502 2382 31554
rect 2434 31502 2436 31554
rect 2156 31388 2324 31444
rect 2156 30996 2212 31006
rect 1932 30994 2212 30996
rect 1932 30942 2158 30994
rect 2210 30942 2212 30994
rect 1932 30940 2212 30942
rect 2156 30930 2212 30940
rect 1708 30098 1764 30110
rect 1708 30046 1710 30098
rect 1762 30046 1764 30098
rect 1708 29876 1764 30046
rect 1708 29810 1764 29820
rect 2044 29986 2100 29998
rect 2044 29934 2046 29986
rect 2098 29934 2100 29986
rect 2044 29652 2100 29934
rect 2268 29764 2324 31388
rect 2380 31220 2436 31502
rect 2380 31154 2436 31164
rect 2492 30212 2548 31724
rect 2604 31714 2660 31724
rect 2716 34692 2772 34702
rect 2604 30212 2660 30222
rect 2492 30156 2604 30212
rect 2604 30146 2660 30156
rect 2492 29986 2548 29998
rect 2492 29934 2494 29986
rect 2546 29934 2548 29986
rect 2492 29876 2548 29934
rect 2492 29810 2548 29820
rect 2268 29708 2436 29764
rect 2044 29596 2324 29652
rect 1932 29538 1988 29550
rect 1932 29486 1934 29538
rect 1986 29486 1988 29538
rect 1932 29428 1988 29486
rect 2156 29428 2212 29438
rect 1932 29426 2212 29428
rect 1932 29374 2158 29426
rect 2210 29374 2212 29426
rect 1932 29372 2212 29374
rect 2156 29362 2212 29372
rect 1708 28756 1764 28766
rect 1708 28642 1764 28700
rect 1708 28590 1710 28642
rect 1762 28590 1764 28642
rect 1708 28578 1764 28590
rect 2044 28644 2100 28654
rect 2044 28530 2100 28588
rect 2044 28478 2046 28530
rect 2098 28478 2100 28530
rect 2044 28466 2100 28478
rect 1932 27970 1988 27982
rect 1932 27918 1934 27970
rect 1986 27918 1988 27970
rect 1932 27860 1988 27918
rect 2156 27860 2212 27870
rect 1932 27858 2212 27860
rect 1932 27806 2158 27858
rect 2210 27806 2212 27858
rect 1932 27804 2212 27806
rect 2268 27860 2324 29596
rect 2380 29428 2436 29708
rect 2380 29362 2436 29372
rect 2716 29426 2772 34636
rect 2940 34690 2996 34702
rect 2940 34638 2942 34690
rect 2994 34638 2996 34690
rect 2940 34356 2996 34638
rect 2940 34290 2996 34300
rect 4732 34354 4788 34366
rect 4732 34302 4734 34354
rect 4786 34302 4788 34354
rect 4732 34244 4788 34302
rect 4732 34178 4788 34188
rect 5628 34244 5684 34254
rect 5292 34020 5348 34030
rect 5292 33926 5348 33964
rect 5628 34018 5684 34188
rect 5628 33966 5630 34018
rect 5682 33966 5684 34018
rect 4268 33740 4948 33750
rect 4324 33684 4372 33740
rect 4428 33738 4476 33740
rect 4532 33738 4580 33740
rect 4448 33686 4476 33738
rect 4572 33686 4580 33738
rect 4428 33684 4476 33686
rect 4532 33684 4580 33686
rect 4636 33738 4684 33740
rect 4740 33738 4788 33740
rect 4636 33686 4644 33738
rect 4740 33686 4768 33738
rect 4636 33684 4684 33686
rect 4740 33684 4788 33686
rect 4844 33684 4892 33740
rect 4268 33674 4948 33684
rect 5628 32564 5684 33966
rect 5628 32498 5684 32508
rect 4268 32172 4948 32182
rect 4324 32116 4372 32172
rect 4428 32170 4476 32172
rect 4532 32170 4580 32172
rect 4448 32118 4476 32170
rect 4572 32118 4580 32170
rect 4428 32116 4476 32118
rect 4532 32116 4580 32118
rect 4636 32170 4684 32172
rect 4740 32170 4788 32172
rect 4636 32118 4644 32170
rect 4740 32118 4768 32170
rect 4636 32116 4684 32118
rect 4740 32116 4788 32118
rect 4844 32116 4892 32172
rect 4268 32106 4948 32116
rect 6524 31948 6580 37100
rect 7084 37090 7140 37100
rect 6748 36932 6804 36942
rect 6748 36596 6804 36876
rect 7308 36596 7364 37436
rect 8316 37380 8372 37390
rect 8652 37380 8708 37390
rect 8316 37378 8484 37380
rect 8316 37326 8318 37378
rect 8370 37326 8484 37378
rect 8316 37324 8484 37326
rect 8316 37314 8372 37324
rect 6748 36594 7364 36596
rect 6748 36542 7310 36594
rect 7362 36542 7364 36594
rect 6748 36540 7364 36542
rect 6748 36482 6804 36540
rect 7308 36530 7364 36540
rect 6748 36430 6750 36482
rect 6802 36430 6804 36482
rect 6748 36418 6804 36430
rect 8428 36484 8484 37324
rect 8652 37286 8708 37324
rect 8988 37378 9044 37390
rect 8988 37326 8990 37378
rect 9042 37326 9044 37378
rect 8652 36484 8708 36494
rect 8428 36482 8708 36484
rect 8428 36430 8654 36482
rect 8706 36430 8708 36482
rect 8428 36428 8708 36430
rect 8988 36484 9044 37326
rect 9660 37380 9716 37390
rect 10220 37380 10276 37390
rect 9660 37286 9716 37324
rect 10108 37378 10276 37380
rect 10108 37326 10222 37378
rect 10274 37326 10276 37378
rect 10108 37324 10276 37326
rect 9996 37044 10052 37054
rect 9996 36950 10052 36988
rect 10108 36932 10164 37324
rect 10220 37314 10276 37324
rect 9212 36484 9268 36494
rect 8988 36482 9268 36484
rect 8988 36430 9214 36482
rect 9266 36430 9268 36482
rect 8988 36428 9268 36430
rect 8652 36418 8708 36428
rect 9212 36418 9268 36428
rect 6636 36260 6692 36270
rect 6636 35922 6692 36204
rect 8428 36260 8484 36270
rect 8428 36166 8484 36204
rect 8768 36092 9448 36102
rect 8824 36036 8872 36092
rect 8928 36090 8976 36092
rect 9032 36090 9080 36092
rect 8948 36038 8976 36090
rect 9072 36038 9080 36090
rect 8928 36036 8976 36038
rect 9032 36036 9080 36038
rect 9136 36090 9184 36092
rect 9240 36090 9288 36092
rect 9136 36038 9144 36090
rect 9240 36038 9268 36090
rect 9136 36036 9184 36038
rect 9240 36036 9288 36038
rect 9344 36036 9392 36092
rect 8768 36026 9448 36036
rect 6636 35870 6638 35922
rect 6690 35870 6692 35922
rect 6636 35858 6692 35870
rect 8652 34690 8708 34702
rect 8652 34638 8654 34690
rect 8706 34638 8708 34690
rect 8652 33684 8708 34638
rect 9212 34692 9268 34702
rect 9212 34690 9604 34692
rect 9212 34638 9214 34690
rect 9266 34638 9604 34690
rect 9212 34636 9604 34638
rect 9212 34626 9268 34636
rect 8768 34524 9448 34534
rect 8824 34468 8872 34524
rect 8928 34522 8976 34524
rect 9032 34522 9080 34524
rect 8948 34470 8976 34522
rect 9072 34470 9080 34522
rect 8928 34468 8976 34470
rect 9032 34468 9080 34470
rect 9136 34522 9184 34524
rect 9240 34522 9288 34524
rect 9136 34470 9144 34522
rect 9240 34470 9268 34522
rect 9136 34468 9184 34470
rect 9240 34468 9288 34470
rect 9344 34468 9392 34524
rect 8768 34458 9448 34468
rect 8540 32676 8596 32686
rect 8540 31948 8596 32620
rect 3276 31892 3332 31902
rect 2940 31556 2996 31566
rect 2940 31462 2996 31500
rect 3276 30884 3332 31836
rect 6300 31892 6580 31948
rect 8428 31892 8596 31948
rect 5516 31780 5572 31790
rect 5068 31778 5572 31780
rect 5068 31726 5518 31778
rect 5570 31726 5572 31778
rect 5068 31724 5572 31726
rect 5068 31666 5124 31724
rect 5516 31714 5572 31724
rect 6076 31780 6132 31790
rect 6076 31686 6132 31724
rect 5068 31614 5070 31666
rect 5122 31614 5124 31666
rect 5068 31602 5124 31614
rect 4732 31220 4788 31230
rect 4732 31218 5124 31220
rect 4732 31166 4734 31218
rect 4786 31166 5124 31218
rect 4732 31164 5124 31166
rect 4732 31154 4788 31164
rect 3276 30818 3332 30828
rect 4268 30604 4948 30614
rect 4324 30548 4372 30604
rect 4428 30602 4476 30604
rect 4532 30602 4580 30604
rect 4448 30550 4476 30602
rect 4572 30550 4580 30602
rect 4428 30548 4476 30550
rect 4532 30548 4580 30550
rect 4636 30602 4684 30604
rect 4740 30602 4788 30604
rect 4636 30550 4644 30602
rect 4740 30550 4768 30602
rect 4636 30548 4684 30550
rect 4740 30548 4788 30550
rect 4844 30548 4892 30604
rect 4268 30538 4948 30548
rect 2716 29374 2718 29426
rect 2770 29374 2772 29426
rect 2716 29362 2772 29374
rect 5068 29650 5124 31164
rect 5068 29598 5070 29650
rect 5122 29598 5124 29650
rect 4268 29036 4948 29046
rect 4324 28980 4372 29036
rect 4428 29034 4476 29036
rect 4532 29034 4580 29036
rect 4448 28982 4476 29034
rect 4572 28982 4580 29034
rect 4428 28980 4476 28982
rect 4532 28980 4580 28982
rect 4636 29034 4684 29036
rect 4740 29034 4788 29036
rect 4636 28982 4644 29034
rect 4740 28982 4768 29034
rect 4636 28980 4684 28982
rect 4740 28980 4788 28982
rect 4844 28980 4892 29036
rect 4268 28970 4948 28980
rect 2492 28756 2548 28766
rect 2492 28662 2548 28700
rect 5068 28084 5124 29598
rect 5292 30770 5348 30782
rect 5292 30718 5294 30770
rect 5346 30718 5348 30770
rect 5292 29652 5348 30718
rect 5292 29586 5348 29596
rect 6076 29316 6132 29326
rect 6300 29316 6356 31892
rect 6132 29260 6356 29316
rect 5852 29204 5908 29214
rect 5068 27990 5124 28028
rect 5628 29202 5908 29204
rect 5628 29150 5854 29202
rect 5906 29150 5908 29202
rect 5628 29148 5908 29150
rect 2716 27860 2772 27870
rect 2268 27858 2772 27860
rect 2268 27806 2718 27858
rect 2770 27806 2772 27858
rect 2268 27804 2772 27806
rect 2156 27794 2212 27804
rect 2716 27794 2772 27804
rect 1708 27636 1764 27646
rect 1708 27076 1764 27580
rect 4268 27468 4948 27478
rect 4324 27412 4372 27468
rect 4428 27466 4476 27468
rect 4532 27466 4580 27468
rect 4448 27414 4476 27466
rect 4572 27414 4580 27466
rect 4428 27412 4476 27414
rect 4532 27412 4580 27414
rect 4636 27466 4684 27468
rect 4740 27466 4788 27468
rect 4636 27414 4644 27466
rect 4740 27414 4768 27466
rect 4636 27412 4684 27414
rect 4740 27412 4788 27414
rect 4844 27412 4892 27468
rect 4268 27402 4948 27412
rect 5628 27300 5684 29148
rect 5852 29138 5908 29148
rect 6076 27860 6132 29260
rect 7644 28644 7700 28654
rect 7420 28420 7476 28430
rect 7308 28418 7476 28420
rect 7308 28366 7422 28418
rect 7474 28366 7476 28418
rect 7308 28364 7476 28366
rect 5628 27234 5684 27244
rect 5740 27858 6132 27860
rect 5740 27806 6078 27858
rect 6130 27806 6132 27858
rect 5740 27804 6132 27806
rect 1708 26982 1764 27020
rect 2492 27076 2548 27086
rect 2044 26964 2100 26974
rect 2044 26962 2212 26964
rect 2044 26910 2046 26962
rect 2098 26910 2212 26962
rect 2044 26908 2212 26910
rect 2044 26898 2100 26908
rect 1932 26402 1988 26414
rect 1932 26350 1934 26402
rect 1986 26350 1988 26402
rect 1708 25396 1764 25406
rect 1708 25302 1764 25340
rect 1820 24724 1876 24734
rect 1932 24724 1988 26350
rect 2044 25732 2100 25742
rect 2044 25394 2100 25676
rect 2156 25508 2212 26908
rect 2380 26852 2436 26862
rect 2156 25442 2212 25452
rect 2268 26850 2436 26852
rect 2268 26798 2382 26850
rect 2434 26798 2436 26850
rect 2268 26796 2436 26798
rect 2044 25342 2046 25394
rect 2098 25342 2100 25394
rect 2044 25330 2100 25342
rect 1820 24722 1988 24724
rect 1820 24670 1822 24722
rect 1874 24670 1988 24722
rect 1820 24668 1988 24670
rect 2268 24722 2324 26796
rect 2380 26786 2436 26796
rect 2492 26514 2548 27020
rect 2492 26462 2494 26514
rect 2546 26462 2548 26514
rect 2492 26450 2548 26462
rect 2604 27074 2660 27086
rect 2604 27022 2606 27074
rect 2658 27022 2660 27074
rect 2604 26964 2660 27022
rect 3164 26964 3220 26974
rect 2604 26962 3220 26964
rect 2604 26910 3166 26962
rect 3218 26910 3220 26962
rect 2604 26908 3220 26910
rect 2604 26516 2660 26908
rect 3164 26898 3220 26908
rect 5740 26962 5796 27804
rect 6076 27794 6132 27804
rect 6748 28084 6804 28094
rect 6748 27746 6804 28028
rect 6748 27694 6750 27746
rect 6802 27694 6804 27746
rect 6748 27682 6804 27694
rect 5740 26910 5742 26962
rect 5794 26910 5796 26962
rect 2604 26450 2660 26460
rect 5292 26402 5348 26414
rect 5292 26350 5294 26402
rect 5346 26350 5348 26402
rect 4268 25900 4948 25910
rect 4324 25844 4372 25900
rect 4428 25898 4476 25900
rect 4532 25898 4580 25900
rect 4448 25846 4476 25898
rect 4572 25846 4580 25898
rect 4428 25844 4476 25846
rect 4532 25844 4580 25846
rect 4636 25898 4684 25900
rect 4740 25898 4788 25900
rect 4636 25846 4644 25898
rect 4740 25846 4768 25898
rect 4636 25844 4684 25846
rect 4740 25844 4788 25846
rect 4844 25844 4892 25900
rect 4268 25834 4948 25844
rect 5292 25508 5348 26350
rect 5516 25508 5572 25518
rect 5292 25506 5572 25508
rect 5292 25454 5518 25506
rect 5570 25454 5572 25506
rect 5292 25452 5572 25454
rect 5516 25442 5572 25452
rect 2492 25396 2548 25406
rect 5740 25396 5796 26910
rect 5852 27634 5908 27646
rect 5852 27582 5854 27634
rect 5906 27582 5908 27634
rect 5852 25620 5908 27582
rect 7308 27074 7364 28364
rect 7420 28354 7476 28364
rect 7308 27022 7310 27074
rect 7362 27022 7364 27074
rect 7308 27010 7364 27022
rect 7644 27074 7700 28588
rect 7644 27022 7646 27074
rect 7698 27022 7700 27074
rect 7644 27010 7700 27022
rect 5852 25554 5908 25564
rect 6076 25508 6132 25518
rect 6076 25414 6132 25452
rect 5740 25340 5908 25396
rect 2492 25302 2548 25340
rect 4732 24946 4788 24958
rect 4732 24894 4734 24946
rect 4786 24894 4788 24946
rect 4732 24836 4788 24894
rect 5292 24948 5348 24958
rect 5292 24854 5348 24892
rect 4732 24770 4788 24780
rect 5068 24836 5124 24846
rect 5740 24836 5796 24846
rect 2268 24670 2270 24722
rect 2322 24670 2324 24722
rect 1820 24658 1876 24668
rect 2268 24658 2324 24670
rect 4268 24332 4948 24342
rect 1708 24276 1764 24286
rect 1708 23938 1764 24220
rect 3612 24276 3668 24286
rect 4324 24276 4372 24332
rect 4428 24330 4476 24332
rect 4532 24330 4580 24332
rect 4448 24278 4476 24330
rect 4572 24278 4580 24330
rect 4428 24276 4476 24278
rect 4532 24276 4580 24278
rect 4636 24330 4684 24332
rect 4740 24330 4788 24332
rect 4636 24278 4644 24330
rect 4740 24278 4768 24330
rect 4636 24276 4684 24278
rect 4740 24276 4788 24278
rect 4844 24276 4892 24332
rect 4268 24266 4948 24276
rect 3612 24050 3668 24220
rect 3612 23998 3614 24050
rect 3666 23998 3668 24050
rect 3612 23986 3668 23998
rect 1708 23886 1710 23938
rect 1762 23886 1764 23938
rect 1708 23874 1764 23886
rect 2380 23826 2436 23838
rect 2380 23774 2382 23826
rect 2434 23774 2436 23826
rect 2044 23714 2100 23726
rect 2044 23662 2046 23714
rect 2098 23662 2100 23714
rect 2044 23380 2100 23662
rect 2380 23548 2436 23774
rect 2044 23314 2100 23324
rect 2156 23492 2436 23548
rect 1820 23154 1876 23166
rect 1820 23102 1822 23154
rect 1874 23102 1876 23154
rect 1820 22708 1876 23102
rect 2156 23156 2212 23492
rect 2380 23416 2436 23436
rect 2716 23714 2772 23726
rect 2716 23662 2718 23714
rect 2770 23662 2772 23714
rect 2156 23090 2212 23100
rect 2268 23156 2324 23166
rect 2268 23154 2660 23156
rect 2268 23102 2270 23154
rect 2322 23102 2660 23154
rect 2268 23100 2660 23102
rect 2268 23090 2324 23100
rect 1820 22652 2212 22708
rect 1708 22258 1764 22270
rect 1708 22206 1710 22258
rect 1762 22206 1764 22258
rect 1708 22036 1764 22206
rect 2156 22260 2212 22652
rect 2380 22260 2436 22270
rect 2156 22258 2436 22260
rect 2156 22206 2382 22258
rect 2434 22206 2436 22258
rect 2156 22204 2436 22206
rect 2380 22194 2436 22204
rect 2044 22148 2100 22158
rect 1708 21970 1764 21980
rect 1932 22146 2100 22148
rect 1932 22094 2046 22146
rect 2098 22094 2100 22146
rect 1932 22092 2100 22094
rect 1708 21586 1764 21598
rect 1708 21534 1710 21586
rect 1762 21534 1764 21586
rect 1708 21476 1764 21534
rect 1932 21588 1988 22092
rect 2044 22082 2100 22092
rect 2044 21700 2100 21710
rect 2044 21698 2436 21700
rect 2044 21646 2046 21698
rect 2098 21646 2436 21698
rect 2044 21644 2436 21646
rect 2044 21634 2100 21644
rect 1932 21522 1988 21532
rect 1708 20916 1764 21420
rect 1708 20850 1764 20860
rect 2044 20804 2100 20814
rect 1932 20578 1988 20590
rect 1932 20526 1934 20578
rect 1986 20526 1988 20578
rect 1820 20020 1876 20030
rect 1932 20020 1988 20526
rect 1820 20018 1988 20020
rect 1820 19966 1822 20018
rect 1874 19966 1988 20018
rect 1820 19964 1988 19966
rect 1820 19954 1876 19964
rect 1708 19796 1764 19806
rect 1708 19348 1764 19740
rect 1708 19234 1764 19292
rect 2044 19236 2100 20748
rect 1708 19182 1710 19234
rect 1762 19182 1764 19234
rect 1708 19170 1764 19182
rect 1932 19180 2100 19236
rect 2156 20018 2212 20030
rect 2156 19966 2158 20018
rect 2210 19966 2212 20018
rect 1708 17556 1764 17566
rect 1708 17462 1764 17500
rect 1932 17108 1988 19180
rect 2044 19012 2100 19022
rect 2044 18918 2100 18956
rect 2156 18676 2212 19966
rect 2380 19460 2436 21644
rect 2492 21476 2548 21486
rect 2492 21382 2548 21420
rect 2604 21252 2660 23100
rect 2716 21476 2772 23662
rect 3164 23714 3220 23726
rect 3164 23662 3166 23714
rect 3218 23662 3220 23714
rect 3164 23492 3220 23662
rect 5068 23492 5124 24780
rect 5628 24780 5740 24836
rect 5628 24722 5684 24780
rect 5740 24770 5796 24780
rect 5628 24670 5630 24722
rect 5682 24670 5684 24722
rect 5628 24658 5684 24670
rect 5852 24612 5908 25340
rect 8428 25394 8484 31892
rect 8652 31554 8708 33628
rect 9548 33348 9604 34636
rect 9548 33282 9604 33292
rect 10108 33460 10164 36876
rect 8876 33124 8932 33134
rect 8876 33122 9604 33124
rect 8876 33070 8878 33122
rect 8930 33070 9604 33122
rect 8876 33068 9604 33070
rect 8876 33058 8932 33068
rect 8768 32956 9448 32966
rect 8824 32900 8872 32956
rect 8928 32954 8976 32956
rect 9032 32954 9080 32956
rect 8948 32902 8976 32954
rect 9072 32902 9080 32954
rect 8928 32900 8976 32902
rect 9032 32900 9080 32902
rect 9136 32954 9184 32956
rect 9240 32954 9288 32956
rect 9136 32902 9144 32954
rect 9240 32902 9268 32954
rect 9136 32900 9184 32902
rect 9240 32900 9288 32902
rect 9344 32900 9392 32956
rect 8768 32890 9448 32900
rect 9100 32564 9156 32574
rect 9100 32470 9156 32508
rect 9548 32562 9604 33068
rect 9548 32510 9550 32562
rect 9602 32510 9604 32562
rect 9548 32498 9604 32510
rect 9996 32564 10052 32574
rect 9996 31948 10052 32508
rect 9212 31892 9268 31902
rect 9212 31798 9268 31836
rect 9884 31892 10052 31948
rect 8652 31502 8654 31554
rect 8706 31502 8708 31554
rect 8652 31490 8708 31502
rect 8768 31388 9448 31398
rect 8824 31332 8872 31388
rect 8928 31386 8976 31388
rect 9032 31386 9080 31388
rect 8948 31334 8976 31386
rect 9072 31334 9080 31386
rect 8928 31332 8976 31334
rect 9032 31332 9080 31334
rect 9136 31386 9184 31388
rect 9240 31386 9288 31388
rect 9136 31334 9144 31386
rect 9240 31334 9268 31386
rect 9136 31332 9184 31334
rect 9240 31332 9288 31334
rect 9344 31332 9392 31388
rect 8768 31322 9448 31332
rect 8876 30212 8932 30222
rect 8652 30210 8932 30212
rect 8652 30158 8878 30210
rect 8930 30158 8932 30210
rect 8652 30156 8932 30158
rect 8652 30098 8708 30156
rect 8876 30146 8932 30156
rect 9436 30212 9492 30222
rect 9436 30118 9492 30156
rect 8652 30046 8654 30098
rect 8706 30046 8708 30098
rect 8652 30034 8708 30046
rect 8768 29820 9448 29830
rect 8824 29764 8872 29820
rect 8928 29818 8976 29820
rect 9032 29818 9080 29820
rect 8948 29766 8976 29818
rect 9072 29766 9080 29818
rect 8928 29764 8976 29766
rect 9032 29764 9080 29766
rect 9136 29818 9184 29820
rect 9240 29818 9288 29820
rect 9136 29766 9144 29818
rect 9240 29766 9268 29818
rect 9136 29764 9184 29766
rect 9240 29764 9288 29766
rect 9344 29764 9392 29820
rect 8768 29754 9448 29764
rect 8768 28252 9448 28262
rect 8824 28196 8872 28252
rect 8928 28250 8976 28252
rect 9032 28250 9080 28252
rect 8948 28198 8976 28250
rect 9072 28198 9080 28250
rect 8928 28196 8976 28198
rect 9032 28196 9080 28198
rect 9136 28250 9184 28252
rect 9240 28250 9288 28252
rect 9136 28198 9144 28250
rect 9240 28198 9268 28250
rect 9136 28196 9184 28198
rect 9240 28196 9288 28198
rect 9344 28196 9392 28252
rect 8768 28186 9448 28196
rect 8768 26684 9448 26694
rect 8824 26628 8872 26684
rect 8928 26682 8976 26684
rect 9032 26682 9080 26684
rect 8948 26630 8976 26682
rect 9072 26630 9080 26682
rect 8928 26628 8976 26630
rect 9032 26628 9080 26630
rect 9136 26682 9184 26684
rect 9240 26682 9288 26684
rect 9136 26630 9144 26682
rect 9240 26630 9268 26682
rect 9136 26628 9184 26630
rect 9240 26628 9288 26630
rect 9344 26628 9392 26684
rect 8768 26618 9448 26628
rect 9212 25508 9268 25518
rect 9212 25506 9716 25508
rect 9212 25454 9214 25506
rect 9266 25454 9716 25506
rect 9212 25452 9716 25454
rect 9212 25442 9268 25452
rect 8428 25342 8430 25394
rect 8482 25342 8484 25394
rect 8428 25284 8484 25342
rect 9548 25284 9604 25294
rect 8428 25282 9604 25284
rect 8428 25230 9550 25282
rect 9602 25230 9604 25282
rect 8428 25228 9604 25230
rect 3164 23426 3220 23436
rect 4732 23436 5124 23492
rect 5740 24556 5908 24612
rect 6076 24836 6132 24846
rect 4732 23378 4788 23436
rect 4732 23326 4734 23378
rect 4786 23326 4788 23378
rect 4732 23314 4788 23326
rect 5292 23268 5348 23278
rect 5292 23174 5348 23212
rect 5628 23266 5684 23278
rect 5628 23214 5630 23266
rect 5682 23214 5684 23266
rect 4268 22764 4948 22774
rect 4324 22708 4372 22764
rect 4428 22762 4476 22764
rect 4532 22762 4580 22764
rect 4448 22710 4476 22762
rect 4572 22710 4580 22762
rect 4428 22708 4476 22710
rect 4532 22708 4580 22710
rect 4636 22762 4684 22764
rect 4740 22762 4788 22764
rect 4636 22710 4644 22762
rect 4740 22710 4768 22762
rect 4636 22708 4684 22710
rect 4740 22708 4788 22710
rect 4844 22708 4892 22764
rect 4268 22698 4948 22708
rect 2716 21410 2772 21420
rect 2828 22372 2884 22382
rect 2380 19394 2436 19404
rect 2492 21196 2660 21252
rect 2380 19124 2436 19134
rect 2492 19124 2548 21196
rect 2380 19122 2548 19124
rect 2380 19070 2382 19122
rect 2434 19070 2548 19122
rect 2380 19068 2548 19070
rect 2716 19122 2772 19134
rect 2716 19070 2718 19122
rect 2770 19070 2772 19122
rect 2380 19058 2436 19068
rect 2044 18620 2212 18676
rect 2268 18676 2324 18686
rect 2044 17554 2100 18620
rect 2156 18452 2212 18462
rect 2268 18452 2324 18620
rect 2716 18676 2772 19070
rect 2828 19012 2884 22316
rect 5628 22370 5684 23214
rect 5628 22318 5630 22370
rect 5682 22318 5684 22370
rect 5628 22306 5684 22318
rect 2940 22146 2996 22158
rect 2940 22094 2942 22146
rect 2994 22094 2996 22146
rect 2940 22036 2996 22094
rect 2940 21970 2996 21980
rect 4268 21196 4948 21206
rect 4324 21140 4372 21196
rect 4428 21194 4476 21196
rect 4532 21194 4580 21196
rect 4448 21142 4476 21194
rect 4572 21142 4580 21194
rect 4428 21140 4476 21142
rect 4532 21140 4580 21142
rect 4636 21194 4684 21196
rect 4740 21194 4788 21196
rect 4636 21142 4644 21194
rect 4740 21142 4768 21194
rect 4636 21140 4684 21142
rect 4740 21140 4788 21142
rect 4844 21140 4892 21196
rect 4268 21130 4948 21140
rect 4620 21028 4676 21038
rect 4284 20916 4340 20926
rect 4620 20916 4676 20972
rect 4284 20914 4676 20916
rect 4284 20862 4286 20914
rect 4338 20862 4676 20914
rect 4284 20860 4676 20862
rect 4284 20850 4340 20860
rect 4620 20802 4676 20860
rect 4620 20750 4622 20802
rect 4674 20750 4676 20802
rect 4620 20738 4676 20750
rect 5068 20690 5124 20702
rect 5068 20638 5070 20690
rect 5122 20638 5124 20690
rect 4508 20130 4564 20142
rect 4508 20078 4510 20130
rect 4562 20078 4564 20130
rect 4508 20020 4564 20078
rect 4508 19954 4564 19964
rect 5068 19908 5124 20638
rect 5292 20132 5348 20142
rect 5292 20038 5348 20076
rect 5068 19842 5124 19852
rect 5740 20018 5796 24556
rect 6076 23380 6132 24780
rect 8428 24836 8484 25228
rect 9548 25218 9604 25228
rect 8768 25116 9448 25126
rect 8824 25060 8872 25116
rect 8928 25114 8976 25116
rect 9032 25114 9080 25116
rect 8948 25062 8976 25114
rect 9072 25062 9080 25114
rect 8928 25060 8976 25062
rect 9032 25060 9080 25062
rect 9136 25114 9184 25116
rect 9240 25114 9288 25116
rect 9136 25062 9144 25114
rect 9240 25062 9268 25114
rect 9136 25060 9184 25062
rect 9240 25060 9288 25062
rect 9344 25060 9392 25116
rect 8768 25050 9448 25060
rect 6076 23378 6356 23380
rect 6076 23326 6078 23378
rect 6130 23326 6356 23378
rect 6076 23324 6356 23326
rect 6076 23314 6132 23324
rect 6076 22372 6132 22382
rect 6076 22278 6132 22316
rect 5852 21362 5908 21374
rect 5852 21310 5854 21362
rect 5906 21310 5908 21362
rect 5852 21028 5908 21310
rect 5852 20962 5908 20972
rect 6188 20804 6244 20814
rect 5964 20802 6244 20804
rect 5964 20750 6190 20802
rect 6242 20750 6244 20802
rect 5964 20748 6244 20750
rect 5964 20690 6020 20748
rect 6188 20738 6244 20748
rect 5964 20638 5966 20690
rect 6018 20638 6020 20690
rect 5964 20626 6020 20638
rect 6300 20188 6356 23324
rect 8428 22484 8484 24780
rect 9660 23828 9716 25452
rect 9660 23762 9716 23772
rect 9772 24722 9828 24734
rect 9772 24670 9774 24722
rect 9826 24670 9828 24722
rect 9772 23604 9828 24670
rect 8768 23548 9448 23558
rect 8824 23492 8872 23548
rect 8928 23546 8976 23548
rect 9032 23546 9080 23548
rect 8948 23494 8976 23546
rect 9072 23494 9080 23546
rect 8928 23492 8976 23494
rect 9032 23492 9080 23494
rect 9136 23546 9184 23548
rect 9240 23546 9288 23548
rect 9136 23494 9144 23546
rect 9240 23494 9268 23546
rect 9136 23492 9184 23494
rect 9240 23492 9288 23494
rect 9344 23492 9392 23548
rect 8768 23482 9448 23492
rect 9548 23548 9828 23604
rect 9548 23380 9604 23548
rect 9884 23492 9940 31892
rect 9996 29988 10052 29998
rect 9996 27972 10052 29932
rect 9996 26962 10052 27916
rect 9996 26910 9998 26962
rect 10050 26910 10052 26962
rect 9996 26898 10052 26910
rect 9212 23324 9604 23380
rect 9660 23436 9940 23492
rect 9212 22594 9268 23324
rect 9212 22542 9214 22594
rect 9266 22542 9268 22594
rect 9212 22530 9268 22542
rect 8428 22260 8484 22428
rect 9548 22484 9604 22494
rect 9548 22390 9604 22428
rect 8428 22258 8708 22260
rect 8428 22206 8430 22258
rect 8482 22206 8708 22258
rect 8428 22204 8708 22206
rect 8428 22194 8484 22204
rect 8652 21812 8708 22204
rect 8768 21980 9448 21990
rect 8824 21924 8872 21980
rect 8928 21978 8976 21980
rect 9032 21978 9080 21980
rect 8948 21926 8976 21978
rect 9072 21926 9080 21978
rect 8928 21924 8976 21926
rect 9032 21924 9080 21926
rect 9136 21978 9184 21980
rect 9240 21978 9288 21980
rect 9136 21926 9144 21978
rect 9240 21926 9268 21978
rect 9136 21924 9184 21926
rect 9240 21924 9288 21926
rect 9344 21924 9392 21980
rect 8768 21914 9448 21924
rect 8988 21812 9044 21822
rect 9100 21812 9156 21822
rect 8652 21810 9100 21812
rect 8652 21758 8990 21810
rect 9042 21758 9100 21810
rect 8652 21756 9100 21758
rect 8988 21746 9044 21756
rect 6412 21586 6468 21598
rect 6412 21534 6414 21586
rect 6466 21534 6468 21586
rect 6412 21476 6468 21534
rect 6860 21476 6916 21486
rect 6412 21474 6916 21476
rect 6412 21422 6862 21474
rect 6914 21422 6916 21474
rect 6412 21420 6916 21422
rect 6748 20804 6804 20814
rect 6748 20710 6804 20748
rect 6860 20188 6916 21420
rect 9100 20690 9156 21756
rect 9100 20638 9102 20690
rect 9154 20638 9156 20690
rect 9100 20626 9156 20638
rect 8768 20412 9448 20422
rect 8824 20356 8872 20412
rect 8928 20410 8976 20412
rect 9032 20410 9080 20412
rect 8948 20358 8976 20410
rect 9072 20358 9080 20410
rect 8928 20356 8976 20358
rect 9032 20356 9080 20358
rect 9136 20410 9184 20412
rect 9240 20410 9288 20412
rect 9136 20358 9144 20410
rect 9240 20358 9268 20410
rect 9136 20356 9184 20358
rect 9240 20356 9288 20358
rect 9344 20356 9392 20412
rect 8768 20346 9448 20356
rect 5740 19966 5742 20018
rect 5794 19966 5796 20018
rect 5740 19908 5796 19966
rect 5740 19842 5796 19852
rect 6076 20132 6356 20188
rect 6636 20132 6916 20188
rect 6076 20020 6132 20132
rect 6076 19906 6132 19964
rect 6076 19854 6078 19906
rect 6130 19854 6132 19906
rect 4268 19628 4948 19638
rect 4324 19572 4372 19628
rect 4428 19626 4476 19628
rect 4532 19626 4580 19628
rect 4448 19574 4476 19626
rect 4572 19574 4580 19626
rect 4428 19572 4476 19574
rect 4532 19572 4580 19574
rect 4636 19626 4684 19628
rect 4740 19626 4788 19628
rect 4636 19574 4644 19626
rect 4740 19574 4768 19626
rect 4636 19572 4684 19574
rect 4740 19572 4788 19574
rect 4844 19572 4892 19628
rect 4268 19562 4948 19572
rect 3164 19348 3220 19358
rect 3164 19254 3220 19292
rect 6076 19348 6132 19854
rect 6524 19348 6580 19358
rect 6076 19346 6580 19348
rect 6076 19294 6078 19346
rect 6130 19294 6526 19346
rect 6578 19294 6580 19346
rect 6076 19292 6580 19294
rect 6076 19282 6132 19292
rect 6524 19282 6580 19292
rect 2828 18946 2884 18956
rect 2716 18610 2772 18620
rect 2156 18450 2324 18452
rect 2156 18398 2158 18450
rect 2210 18398 2324 18450
rect 2156 18396 2324 18398
rect 2156 18386 2212 18396
rect 4268 18060 4948 18070
rect 4324 18004 4372 18060
rect 4428 18058 4476 18060
rect 4532 18058 4580 18060
rect 4448 18006 4476 18058
rect 4572 18006 4580 18058
rect 4428 18004 4476 18006
rect 4532 18004 4580 18006
rect 4636 18058 4684 18060
rect 4740 18058 4788 18060
rect 4636 18006 4644 18058
rect 4740 18006 4768 18058
rect 4636 18004 4684 18006
rect 4740 18004 4788 18006
rect 4844 18004 4892 18060
rect 4268 17994 4948 18004
rect 2044 17502 2046 17554
rect 2098 17502 2100 17554
rect 2044 17490 2100 17502
rect 2492 17556 2548 17566
rect 2492 17462 2548 17500
rect 2044 17108 2100 17118
rect 1932 17106 2100 17108
rect 1932 17054 2046 17106
rect 2098 17054 2100 17106
rect 1932 17052 2100 17054
rect 2044 17042 2100 17052
rect 1708 16882 1764 16894
rect 1708 16830 1710 16882
rect 1762 16830 1764 16882
rect 1708 16436 1764 16830
rect 1708 16370 1764 16380
rect 2492 16882 2548 16894
rect 2492 16830 2494 16882
rect 2546 16830 2548 16882
rect 2492 16436 2548 16830
rect 4268 16492 4948 16502
rect 4324 16436 4372 16492
rect 4428 16490 4476 16492
rect 4532 16490 4580 16492
rect 4448 16438 4476 16490
rect 4572 16438 4580 16490
rect 4428 16436 4476 16438
rect 4532 16436 4580 16438
rect 4636 16490 4684 16492
rect 4740 16490 4788 16492
rect 4636 16438 4644 16490
rect 4740 16438 4768 16490
rect 4636 16436 4684 16438
rect 4740 16436 4788 16438
rect 4844 16436 4892 16492
rect 4268 16426 4948 16436
rect 2492 16370 2548 16380
rect 4268 14924 4948 14934
rect 4324 14868 4372 14924
rect 4428 14922 4476 14924
rect 4532 14922 4580 14924
rect 4448 14870 4476 14922
rect 4572 14870 4580 14922
rect 4428 14868 4476 14870
rect 4532 14868 4580 14870
rect 4636 14922 4684 14924
rect 4740 14922 4788 14924
rect 4636 14870 4644 14922
rect 4740 14870 4768 14922
rect 4636 14868 4684 14870
rect 4740 14868 4788 14870
rect 4844 14868 4892 14924
rect 4268 14858 4948 14868
rect 2044 13972 2100 13982
rect 2044 13878 2100 13916
rect 1708 13746 1764 13758
rect 1708 13694 1710 13746
rect 1762 13694 1764 13746
rect 1708 13076 1764 13694
rect 1708 13010 1764 13020
rect 2492 13634 2548 13646
rect 2492 13582 2494 13634
rect 2546 13582 2548 13634
rect 2492 13076 2548 13582
rect 4268 13356 4948 13366
rect 4324 13300 4372 13356
rect 4428 13354 4476 13356
rect 4532 13354 4580 13356
rect 4448 13302 4476 13354
rect 4572 13302 4580 13354
rect 4428 13300 4476 13302
rect 4532 13300 4580 13302
rect 4636 13354 4684 13356
rect 4740 13354 4788 13356
rect 4636 13302 4644 13354
rect 4740 13302 4768 13354
rect 4636 13300 4684 13302
rect 4740 13300 4788 13302
rect 4844 13300 4892 13356
rect 4268 13290 4948 13300
rect 2492 13010 2548 13020
rect 2044 12292 2100 12302
rect 2044 12198 2100 12236
rect 1708 12178 1764 12190
rect 1708 12126 1710 12178
rect 1762 12126 1764 12178
rect 1708 11956 1764 12126
rect 1708 11890 1764 11900
rect 2492 12066 2548 12078
rect 2492 12014 2494 12066
rect 2546 12014 2548 12066
rect 2492 11956 2548 12014
rect 2492 11890 2548 11900
rect 4268 11788 4948 11798
rect 4324 11732 4372 11788
rect 4428 11786 4476 11788
rect 4532 11786 4580 11788
rect 4448 11734 4476 11786
rect 4572 11734 4580 11786
rect 4428 11732 4476 11734
rect 4532 11732 4580 11734
rect 4636 11786 4684 11788
rect 4740 11786 4788 11788
rect 4636 11734 4644 11786
rect 4740 11734 4768 11786
rect 4636 11732 4684 11734
rect 4740 11732 4788 11734
rect 4844 11732 4892 11788
rect 4268 11722 4948 11732
rect 1708 11282 1764 11294
rect 1708 11230 1710 11282
rect 1762 11230 1764 11282
rect 1708 10836 1764 11230
rect 2044 11172 2100 11182
rect 2044 11078 2100 11116
rect 2492 11170 2548 11182
rect 2492 11118 2494 11170
rect 2546 11118 2548 11170
rect 1708 10770 1764 10780
rect 2492 10836 2548 11118
rect 2492 10770 2548 10780
rect 4268 10220 4948 10230
rect 4324 10164 4372 10220
rect 4428 10218 4476 10220
rect 4532 10218 4580 10220
rect 4448 10166 4476 10218
rect 4572 10166 4580 10218
rect 4428 10164 4476 10166
rect 4532 10164 4580 10166
rect 4636 10218 4684 10220
rect 4740 10218 4788 10220
rect 4636 10166 4644 10218
rect 4740 10166 4768 10218
rect 4636 10164 4684 10166
rect 4740 10164 4788 10166
rect 4844 10164 4892 10220
rect 4268 10154 4948 10164
rect 1708 9716 1764 9726
rect 1708 9622 1764 9660
rect 2492 9716 2548 9726
rect 2492 9622 2548 9660
rect 2044 9604 2100 9614
rect 2044 9510 2100 9548
rect 4268 8652 4948 8662
rect 4324 8596 4372 8652
rect 4428 8650 4476 8652
rect 4532 8650 4580 8652
rect 4448 8598 4476 8650
rect 4572 8598 4580 8650
rect 4428 8596 4476 8598
rect 4532 8596 4580 8598
rect 4636 8650 4684 8652
rect 4740 8650 4788 8652
rect 4636 8598 4644 8650
rect 4740 8598 4768 8650
rect 4636 8596 4684 8598
rect 4740 8596 4788 8598
rect 4844 8596 4892 8652
rect 4268 8586 4948 8596
rect 1820 7362 1876 7374
rect 1820 7310 1822 7362
rect 1874 7310 1876 7362
rect 1708 6468 1764 6478
rect 1820 6468 1876 7310
rect 4268 7084 4948 7094
rect 4324 7028 4372 7084
rect 4428 7082 4476 7084
rect 4532 7082 4580 7084
rect 4448 7030 4476 7082
rect 4572 7030 4580 7082
rect 4428 7028 4476 7030
rect 4532 7028 4580 7030
rect 4636 7082 4684 7084
rect 4740 7082 4788 7084
rect 4636 7030 4644 7082
rect 4740 7030 4768 7082
rect 4636 7028 4684 7030
rect 4740 7028 4788 7030
rect 4844 7028 4892 7084
rect 4268 7018 4948 7028
rect 1708 6466 1876 6468
rect 1708 6414 1710 6466
rect 1762 6414 1876 6466
rect 1708 6412 1876 6414
rect 2268 6690 2324 6702
rect 2268 6638 2270 6690
rect 2322 6638 2324 6690
rect 1708 6356 1764 6412
rect 1708 6290 1764 6300
rect 2268 6132 2324 6638
rect 2268 6066 2324 6076
rect 1820 5906 1876 5918
rect 1820 5854 1822 5906
rect 1874 5854 1876 5906
rect 1820 5236 1876 5854
rect 2268 5796 2324 5806
rect 2268 5702 2324 5740
rect 4268 5516 4948 5526
rect 4324 5460 4372 5516
rect 4428 5514 4476 5516
rect 4532 5514 4580 5516
rect 4448 5462 4476 5514
rect 4572 5462 4580 5514
rect 4428 5460 4476 5462
rect 4532 5460 4580 5462
rect 4636 5514 4684 5516
rect 4740 5514 4788 5516
rect 4636 5462 4644 5514
rect 4740 5462 4768 5514
rect 4636 5460 4684 5462
rect 4740 5460 4788 5462
rect 4844 5460 4892 5516
rect 4268 5450 4948 5460
rect 1820 5142 1876 5180
rect 4268 3948 4948 3958
rect 4324 3892 4372 3948
rect 4428 3946 4476 3948
rect 4532 3946 4580 3948
rect 4448 3894 4476 3946
rect 4572 3894 4580 3946
rect 4428 3892 4476 3894
rect 4532 3892 4580 3894
rect 4636 3946 4684 3948
rect 4740 3946 4788 3948
rect 4636 3894 4644 3946
rect 4740 3894 4768 3946
rect 4636 3892 4684 3894
rect 4740 3892 4788 3894
rect 4844 3892 4892 3948
rect 4268 3882 4948 3892
rect 6076 3444 6132 3454
rect 6300 3444 6356 3454
rect 6076 3442 6356 3444
rect 6076 3390 6078 3442
rect 6130 3390 6302 3442
rect 6354 3390 6356 3442
rect 6076 3388 6356 3390
rect 6076 800 6132 3388
rect 6300 3378 6356 3388
rect 6636 3442 6692 20132
rect 7308 19908 7364 19918
rect 7308 19814 7364 19852
rect 8768 18844 9448 18854
rect 8824 18788 8872 18844
rect 8928 18842 8976 18844
rect 9032 18842 9080 18844
rect 8948 18790 8976 18842
rect 9072 18790 9080 18842
rect 8928 18788 8976 18790
rect 9032 18788 9080 18790
rect 9136 18842 9184 18844
rect 9240 18842 9288 18844
rect 9136 18790 9144 18842
rect 9240 18790 9268 18842
rect 9136 18788 9184 18790
rect 9240 18788 9288 18790
rect 9344 18788 9392 18844
rect 8768 18778 9448 18788
rect 8768 17276 9448 17286
rect 8824 17220 8872 17276
rect 8928 17274 8976 17276
rect 9032 17274 9080 17276
rect 8948 17222 8976 17274
rect 9072 17222 9080 17274
rect 8928 17220 8976 17222
rect 9032 17220 9080 17222
rect 9136 17274 9184 17276
rect 9240 17274 9288 17276
rect 9136 17222 9144 17274
rect 9240 17222 9268 17274
rect 9136 17220 9184 17222
rect 9240 17220 9288 17222
rect 9344 17220 9392 17276
rect 8768 17210 9448 17220
rect 8768 15708 9448 15718
rect 8824 15652 8872 15708
rect 8928 15706 8976 15708
rect 9032 15706 9080 15708
rect 8948 15654 8976 15706
rect 9072 15654 9080 15706
rect 8928 15652 8976 15654
rect 9032 15652 9080 15654
rect 9136 15706 9184 15708
rect 9240 15706 9288 15708
rect 9136 15654 9144 15706
rect 9240 15654 9268 15706
rect 9136 15652 9184 15654
rect 9240 15652 9288 15654
rect 9344 15652 9392 15708
rect 8768 15642 9448 15652
rect 8768 14140 9448 14150
rect 8824 14084 8872 14140
rect 8928 14138 8976 14140
rect 9032 14138 9080 14140
rect 8948 14086 8976 14138
rect 9072 14086 9080 14138
rect 8928 14084 8976 14086
rect 9032 14084 9080 14086
rect 9136 14138 9184 14140
rect 9240 14138 9288 14140
rect 9136 14086 9144 14138
rect 9240 14086 9268 14138
rect 9136 14084 9184 14086
rect 9240 14084 9288 14086
rect 9344 14084 9392 14140
rect 8768 14074 9448 14084
rect 9660 13972 9716 23436
rect 10108 23378 10164 33404
rect 10332 24946 10388 42476
rect 12236 42532 12292 42542
rect 12236 42438 12292 42476
rect 12908 42532 12964 42542
rect 12908 42438 12964 42476
rect 13132 41412 13188 43262
rect 13268 43148 13948 43158
rect 13324 43092 13372 43148
rect 13428 43146 13476 43148
rect 13532 43146 13580 43148
rect 13448 43094 13476 43146
rect 13572 43094 13580 43146
rect 13428 43092 13476 43094
rect 13532 43092 13580 43094
rect 13636 43146 13684 43148
rect 13740 43146 13788 43148
rect 13636 43094 13644 43146
rect 13740 43094 13768 43146
rect 13636 43092 13684 43094
rect 13740 43092 13788 43094
rect 13844 43092 13892 43148
rect 13268 43082 13948 43092
rect 13580 42980 13636 42990
rect 13244 42868 13300 42878
rect 13244 41970 13300 42812
rect 13580 42642 13636 42924
rect 14028 42868 14084 43596
rect 14028 42802 14084 42812
rect 13804 42756 13860 42794
rect 13804 42690 13860 42700
rect 14364 42754 14420 42766
rect 14364 42702 14366 42754
rect 14418 42702 14420 42754
rect 13580 42590 13582 42642
rect 13634 42590 13636 42642
rect 13580 42578 13636 42590
rect 13244 41918 13246 41970
rect 13298 41918 13300 41970
rect 13244 41906 13300 41918
rect 13804 42532 13860 42542
rect 13804 41970 13860 42476
rect 14364 42532 14420 42702
rect 15148 42756 15204 45052
rect 15372 45042 15428 45052
rect 15148 42690 15204 42700
rect 14700 42644 14756 42654
rect 14700 42550 14756 42588
rect 15596 42644 15652 49532
rect 17768 48636 18448 48646
rect 17824 48580 17872 48636
rect 17928 48634 17976 48636
rect 18032 48634 18080 48636
rect 17948 48582 17976 48634
rect 18072 48582 18080 48634
rect 17928 48580 17976 48582
rect 18032 48580 18080 48582
rect 18136 48634 18184 48636
rect 18240 48634 18288 48636
rect 18136 48582 18144 48634
rect 18240 48582 18268 48634
rect 18136 48580 18184 48582
rect 18240 48580 18288 48582
rect 18344 48580 18392 48636
rect 17768 48570 18448 48580
rect 19852 48356 19908 48366
rect 19852 48262 19908 48300
rect 20300 48356 20356 48366
rect 15820 48244 15876 48254
rect 15820 48150 15876 48188
rect 20300 48242 20356 48300
rect 20412 48354 20468 50318
rect 20412 48302 20414 48354
rect 20466 48302 20468 48354
rect 20412 48290 20468 48302
rect 20300 48190 20302 48242
rect 20354 48190 20356 48242
rect 20300 48178 20356 48190
rect 16492 48130 16548 48142
rect 20524 48132 20580 50428
rect 20860 50484 20916 50494
rect 20860 50390 20916 50428
rect 26236 49922 26292 51884
rect 26236 49870 26238 49922
rect 26290 49870 26292 49922
rect 26236 49858 26292 49870
rect 25564 49812 25620 49822
rect 25564 49718 25620 49756
rect 26348 49812 26404 52108
rect 26908 52052 26964 52062
rect 26908 51958 26964 51996
rect 27020 51940 27076 51978
rect 27020 51874 27076 51884
rect 27132 51940 27188 53116
rect 27692 53058 27748 53070
rect 27692 53006 27694 53058
rect 27746 53006 27748 53058
rect 27692 52948 27748 53006
rect 27580 52892 27692 52948
rect 27580 52162 27636 52892
rect 27692 52882 27748 52892
rect 27916 52946 27972 52958
rect 27916 52894 27918 52946
rect 27970 52894 27972 52946
rect 27916 52612 27972 52894
rect 28140 52948 28196 52958
rect 28252 52948 28308 53676
rect 28476 53666 28532 53676
rect 29596 53730 29652 53742
rect 29596 53678 29598 53730
rect 29650 53678 29652 53730
rect 29260 53506 29316 53518
rect 29260 53454 29262 53506
rect 29314 53454 29316 53506
rect 29260 53396 29316 53454
rect 29036 53340 29260 53396
rect 29036 53170 29092 53340
rect 29260 53330 29316 53340
rect 29036 53118 29038 53170
rect 29090 53118 29092 53170
rect 29036 53106 29092 53118
rect 29596 53172 29652 53678
rect 30828 53620 30884 53630
rect 30828 53526 30884 53564
rect 32060 53620 32116 55358
rect 32396 55186 32452 56028
rect 32844 56018 32900 56028
rect 43260 56082 43988 56084
rect 43260 56030 43934 56082
rect 43986 56030 43988 56082
rect 43260 56028 43988 56030
rect 40268 55692 40948 55702
rect 40324 55636 40372 55692
rect 40428 55690 40476 55692
rect 40532 55690 40580 55692
rect 40448 55638 40476 55690
rect 40572 55638 40580 55690
rect 40428 55636 40476 55638
rect 40532 55636 40580 55638
rect 40636 55690 40684 55692
rect 40740 55690 40788 55692
rect 40636 55638 40644 55690
rect 40740 55638 40768 55690
rect 40636 55636 40684 55638
rect 40740 55636 40788 55638
rect 40844 55636 40892 55692
rect 40268 55626 40948 55636
rect 36428 55412 36484 55422
rect 36428 55410 36596 55412
rect 36428 55358 36430 55410
rect 36482 55358 36596 55410
rect 36428 55356 36596 55358
rect 36428 55346 36484 55356
rect 33180 55300 33236 55310
rect 33180 55206 33236 55244
rect 33628 55300 33684 55310
rect 33628 55206 33684 55244
rect 32396 55134 32398 55186
rect 32450 55134 32452 55186
rect 32396 55122 32452 55134
rect 32732 55188 32788 55198
rect 34300 55188 34356 55198
rect 32732 55186 33124 55188
rect 32732 55134 32734 55186
rect 32786 55134 33124 55186
rect 32732 55132 33124 55134
rect 32732 55122 32788 55132
rect 32060 53554 32116 53564
rect 29372 53060 29428 53070
rect 28140 52946 28308 52948
rect 28140 52894 28142 52946
rect 28194 52894 28308 52946
rect 28140 52892 28308 52894
rect 28588 52946 28644 52958
rect 28588 52894 28590 52946
rect 28642 52894 28644 52946
rect 28140 52882 28196 52892
rect 28028 52836 28084 52846
rect 28028 52742 28084 52780
rect 28588 52836 28644 52894
rect 28812 52948 28868 52958
rect 28812 52854 28868 52892
rect 29148 52948 29204 52958
rect 29148 52946 29316 52948
rect 29148 52894 29150 52946
rect 29202 52894 29316 52946
rect 29148 52892 29316 52894
rect 29148 52882 29204 52892
rect 28476 52722 28532 52734
rect 28476 52670 28478 52722
rect 28530 52670 28532 52722
rect 28476 52612 28532 52670
rect 27916 52556 28532 52612
rect 27916 52386 27972 52556
rect 28588 52500 28644 52780
rect 28588 52434 28644 52444
rect 27916 52334 27918 52386
rect 27970 52334 27972 52386
rect 27916 52322 27972 52334
rect 28476 52388 28532 52398
rect 28476 52294 28532 52332
rect 28364 52276 28420 52286
rect 28364 52182 28420 52220
rect 29260 52276 29316 52892
rect 29260 52182 29316 52220
rect 27580 52110 27582 52162
rect 27634 52110 27636 52162
rect 27580 52098 27636 52110
rect 28140 52164 28196 52174
rect 28140 52070 28196 52108
rect 28812 52164 28868 52174
rect 27804 52052 27860 52062
rect 27804 51958 27860 51996
rect 27132 51938 27636 51940
rect 27132 51886 27134 51938
rect 27186 51886 27636 51938
rect 27132 51884 27636 51886
rect 27132 51874 27188 51884
rect 26768 51772 27448 51782
rect 26824 51716 26872 51772
rect 26928 51770 26976 51772
rect 27032 51770 27080 51772
rect 26948 51718 26976 51770
rect 27072 51718 27080 51770
rect 26928 51716 26976 51718
rect 27032 51716 27080 51718
rect 27136 51770 27184 51772
rect 27240 51770 27288 51772
rect 27136 51718 27144 51770
rect 27240 51718 27268 51770
rect 27136 51716 27184 51718
rect 27240 51716 27288 51718
rect 27344 51716 27392 51772
rect 26768 51706 27448 51716
rect 27580 50820 27636 51884
rect 28812 51602 28868 52108
rect 28812 51550 28814 51602
rect 28866 51550 28868 51602
rect 28812 51538 28868 51550
rect 27916 50820 27972 50830
rect 27580 50818 27972 50820
rect 27580 50766 27918 50818
rect 27970 50766 27972 50818
rect 27580 50764 27972 50766
rect 27916 50754 27972 50764
rect 29372 50818 29428 53004
rect 29596 53058 29652 53116
rect 29932 53508 29988 53518
rect 29596 53006 29598 53058
rect 29650 53006 29652 53058
rect 29596 52994 29652 53006
rect 29820 53060 29876 53070
rect 29820 52966 29876 53004
rect 29708 52836 29764 52846
rect 29372 50766 29374 50818
rect 29426 50766 29428 50818
rect 29372 50754 29428 50766
rect 29596 52834 29764 52836
rect 29596 52782 29710 52834
rect 29762 52782 29764 52834
rect 29596 52780 29764 52782
rect 28028 50482 28084 50494
rect 28028 50430 28030 50482
rect 28082 50430 28084 50482
rect 28028 50428 28084 50430
rect 29484 50482 29540 50494
rect 29484 50430 29486 50482
rect 29538 50430 29540 50482
rect 28028 50372 28532 50428
rect 28476 50370 28532 50372
rect 28476 50318 28478 50370
rect 28530 50318 28532 50370
rect 26768 50204 27448 50214
rect 26824 50148 26872 50204
rect 26928 50202 26976 50204
rect 27032 50202 27080 50204
rect 26948 50150 26976 50202
rect 27072 50150 27080 50202
rect 26928 50148 26976 50150
rect 27032 50148 27080 50150
rect 27136 50202 27184 50204
rect 27240 50202 27288 50204
rect 27136 50150 27144 50202
rect 27240 50150 27268 50202
rect 27136 50148 27184 50150
rect 27240 50148 27288 50150
rect 27344 50148 27392 50204
rect 26768 50138 27448 50148
rect 26348 49746 26404 49756
rect 28476 49698 28532 50318
rect 29484 50372 29540 50430
rect 29484 50306 29540 50316
rect 29596 49924 29652 52780
rect 29708 52770 29764 52780
rect 29708 52052 29764 52062
rect 29932 52052 29988 53452
rect 30156 53506 30212 53518
rect 30156 53454 30158 53506
rect 30210 53454 30212 53506
rect 30156 53396 30212 53454
rect 30716 53508 30772 53518
rect 30716 53414 30772 53452
rect 31276 53508 31332 53518
rect 31276 53414 31332 53452
rect 30156 53330 30212 53340
rect 31164 53060 31220 53070
rect 31052 53004 31164 53060
rect 30380 52946 30436 52958
rect 30380 52894 30382 52946
rect 30434 52894 30436 52946
rect 30380 52836 30436 52894
rect 30828 52836 30884 52846
rect 30380 52834 30884 52836
rect 30380 52782 30830 52834
rect 30882 52782 30884 52834
rect 30380 52780 30884 52782
rect 30044 52722 30100 52734
rect 30044 52670 30046 52722
rect 30098 52670 30100 52722
rect 30044 52274 30100 52670
rect 30044 52222 30046 52274
rect 30098 52222 30100 52274
rect 30044 52210 30100 52222
rect 30156 52724 30212 52734
rect 30156 52164 30212 52668
rect 30156 52070 30212 52108
rect 30828 52164 30884 52780
rect 30828 52098 30884 52108
rect 31052 52388 31108 53004
rect 31164 52994 31220 53004
rect 31276 52948 31332 52958
rect 31276 52854 31332 52892
rect 31948 52948 32004 52958
rect 32004 52892 32116 52948
rect 31948 52882 32004 52892
rect 31268 52556 31948 52566
rect 31324 52500 31372 52556
rect 31428 52554 31476 52556
rect 31532 52554 31580 52556
rect 31448 52502 31476 52554
rect 31572 52502 31580 52554
rect 31428 52500 31476 52502
rect 31532 52500 31580 52502
rect 31636 52554 31684 52556
rect 31740 52554 31788 52556
rect 31636 52502 31644 52554
rect 31740 52502 31768 52554
rect 31636 52500 31684 52502
rect 31740 52500 31788 52502
rect 31844 52500 31892 52556
rect 31268 52490 31948 52500
rect 32060 52388 32116 52892
rect 29708 52050 29988 52052
rect 29708 51998 29710 52050
rect 29762 51998 29988 52050
rect 29708 51996 29988 51998
rect 31052 52052 31108 52332
rect 31724 52332 32116 52388
rect 32172 52724 32228 52734
rect 32172 52388 32228 52668
rect 33068 52388 33124 55132
rect 34300 55186 34580 55188
rect 34300 55134 34302 55186
rect 34354 55134 34580 55186
rect 34300 55132 34580 55134
rect 34300 55122 34356 55132
rect 33964 53844 34020 53854
rect 33852 53170 33908 53182
rect 33852 53118 33854 53170
rect 33906 53118 33908 53170
rect 33740 53060 33796 53070
rect 33740 52966 33796 53004
rect 33852 52612 33908 53118
rect 31276 52276 31332 52286
rect 31724 52276 31780 52332
rect 31332 52274 31780 52276
rect 31332 52222 31726 52274
rect 31778 52222 31780 52274
rect 31332 52220 31780 52222
rect 31276 52162 31332 52220
rect 31724 52210 31780 52220
rect 32172 52274 32228 52332
rect 32172 52222 32174 52274
rect 32226 52222 32228 52274
rect 32172 52210 32228 52222
rect 32396 52332 33124 52388
rect 31276 52110 31278 52162
rect 31330 52110 31332 52162
rect 31276 52098 31332 52110
rect 31164 52052 31220 52062
rect 31052 52050 31220 52052
rect 31052 51998 31166 52050
rect 31218 51998 31220 52050
rect 31052 51996 31220 51998
rect 29708 51986 29764 51996
rect 31164 51986 31220 51996
rect 31268 50988 31948 50998
rect 31324 50932 31372 50988
rect 31428 50986 31476 50988
rect 31532 50986 31580 50988
rect 31448 50934 31476 50986
rect 31572 50934 31580 50986
rect 31428 50932 31476 50934
rect 31532 50932 31580 50934
rect 31636 50986 31684 50988
rect 31740 50986 31788 50988
rect 31636 50934 31644 50986
rect 31740 50934 31768 50986
rect 31636 50932 31684 50934
rect 31740 50932 31788 50934
rect 31844 50932 31892 50988
rect 31268 50922 31948 50932
rect 32396 50818 32452 52332
rect 32956 52164 33012 52174
rect 33068 52164 33124 52332
rect 33292 52556 33908 52612
rect 33292 52386 33348 52556
rect 33292 52334 33294 52386
rect 33346 52334 33348 52386
rect 33292 52322 33348 52334
rect 33404 52164 33460 52174
rect 33068 52162 33460 52164
rect 33068 52110 33406 52162
rect 33458 52110 33460 52162
rect 33068 52108 33460 52110
rect 32956 52070 33012 52108
rect 33404 52098 33460 52108
rect 33740 52164 33796 52174
rect 33964 52164 34020 53788
rect 34524 53842 34580 55132
rect 35768 54908 36448 54918
rect 35824 54852 35872 54908
rect 35928 54906 35976 54908
rect 36032 54906 36080 54908
rect 35948 54854 35976 54906
rect 36072 54854 36080 54906
rect 35928 54852 35976 54854
rect 36032 54852 36080 54854
rect 36136 54906 36184 54908
rect 36240 54906 36288 54908
rect 36136 54854 36144 54906
rect 36240 54854 36268 54906
rect 36136 54852 36184 54854
rect 36240 54852 36288 54854
rect 36344 54852 36392 54908
rect 35768 54842 36448 54852
rect 35196 54404 35252 54414
rect 34524 53790 34526 53842
rect 34578 53790 34580 53842
rect 34524 53778 34580 53790
rect 34972 54402 35252 54404
rect 34972 54350 35198 54402
rect 35250 54350 35252 54402
rect 34972 54348 35252 54350
rect 34412 53508 34468 53518
rect 34300 52948 34356 52958
rect 34300 52724 34356 52892
rect 34300 52658 34356 52668
rect 34412 52500 34468 53452
rect 34636 53508 34692 53518
rect 34636 53414 34692 53452
rect 34412 52434 34468 52444
rect 34972 52500 35028 54348
rect 35196 54338 35252 54348
rect 36316 54402 36372 54414
rect 36316 54350 36318 54402
rect 36370 54350 36372 54402
rect 36316 54180 36372 54350
rect 36092 54124 36372 54180
rect 35084 53844 35140 53854
rect 35308 53844 35364 53854
rect 35140 53842 35364 53844
rect 35140 53790 35310 53842
rect 35362 53790 35364 53842
rect 35140 53788 35364 53790
rect 35084 53730 35140 53788
rect 35308 53778 35364 53788
rect 35644 53844 35700 53854
rect 35084 53678 35086 53730
rect 35138 53678 35140 53730
rect 35084 53666 35140 53678
rect 35644 53730 35700 53788
rect 35644 53678 35646 53730
rect 35698 53678 35700 53730
rect 35644 53666 35700 53678
rect 35420 53620 35476 53630
rect 35196 53508 35252 53518
rect 35196 53058 35252 53452
rect 35196 53006 35198 53058
rect 35250 53006 35252 53058
rect 35196 52994 35252 53006
rect 35420 53506 35476 53564
rect 35868 53620 35924 53630
rect 36092 53620 36148 54124
rect 36540 54068 36596 55356
rect 42588 55410 42644 55422
rect 42588 55358 42590 55410
rect 42642 55358 42644 55410
rect 37100 55300 37156 55310
rect 37100 55206 37156 55244
rect 39788 55300 39844 55310
rect 39788 55206 39844 55244
rect 40460 55188 40516 55198
rect 40460 55186 41412 55188
rect 40460 55134 40462 55186
rect 40514 55134 41412 55186
rect 40460 55132 41412 55134
rect 40460 55122 40516 55132
rect 40348 54740 40404 54750
rect 41244 54740 41300 54750
rect 40348 54738 41300 54740
rect 40348 54686 40350 54738
rect 40402 54686 41246 54738
rect 41298 54686 41300 54738
rect 40348 54684 41300 54686
rect 40348 54674 40404 54684
rect 38892 54516 38948 54526
rect 36316 54012 36596 54068
rect 36316 53842 36372 54012
rect 36316 53790 36318 53842
rect 36370 53790 36372 53842
rect 36316 53778 36372 53790
rect 36540 53732 36596 54012
rect 36540 53666 36596 53676
rect 36764 54402 36820 54414
rect 36764 54350 36766 54402
rect 36818 54350 36820 54402
rect 36764 53844 36820 54350
rect 35924 53564 36148 53620
rect 35868 53526 35924 53564
rect 35420 53454 35422 53506
rect 35474 53454 35476 53506
rect 34972 52434 35028 52444
rect 35308 52946 35364 52958
rect 35308 52894 35310 52946
rect 35362 52894 35364 52946
rect 35308 52388 35364 52894
rect 35420 52948 35476 53454
rect 36204 53508 36260 53546
rect 36204 53442 36260 53452
rect 36540 53508 36596 53518
rect 35768 53340 36448 53350
rect 35824 53284 35872 53340
rect 35928 53338 35976 53340
rect 36032 53338 36080 53340
rect 35948 53286 35976 53338
rect 36072 53286 36080 53338
rect 35928 53284 35976 53286
rect 36032 53284 36080 53286
rect 36136 53338 36184 53340
rect 36240 53338 36288 53340
rect 36136 53286 36144 53338
rect 36240 53286 36268 53338
rect 36136 53284 36184 53286
rect 36240 53284 36288 53286
rect 36344 53284 36392 53340
rect 35768 53274 36448 53284
rect 35532 53172 35588 53182
rect 35532 53078 35588 53116
rect 35868 53172 35924 53182
rect 35868 53078 35924 53116
rect 35420 52882 35476 52892
rect 35644 53002 35700 53014
rect 35644 52950 35646 53002
rect 35698 52950 35700 53002
rect 35644 52836 35700 52950
rect 36204 52946 36260 52958
rect 36204 52894 36206 52946
rect 36258 52894 36260 52946
rect 36204 52836 36260 52894
rect 36540 52836 36596 53452
rect 36764 53396 36820 53788
rect 37212 53730 37268 53742
rect 37212 53678 37214 53730
rect 37266 53678 37268 53730
rect 36988 53396 37044 53406
rect 36764 53340 36988 53396
rect 36988 53172 37044 53340
rect 36988 53078 37044 53116
rect 37212 52948 37268 53678
rect 38220 53732 38276 53742
rect 38220 53638 38276 53676
rect 37212 52882 37268 52892
rect 37324 53618 37380 53630
rect 37324 53566 37326 53618
rect 37378 53566 37380 53618
rect 36204 52780 36540 52836
rect 35644 52612 35700 52780
rect 36540 52742 36596 52780
rect 35644 52546 35700 52556
rect 35756 52724 35812 52734
rect 33740 52162 34020 52164
rect 33740 52110 33742 52162
rect 33794 52110 34020 52162
rect 33740 52108 34020 52110
rect 34188 52162 34244 52174
rect 34188 52110 34190 52162
rect 34242 52110 34244 52162
rect 33740 52098 33796 52108
rect 34188 52052 34244 52110
rect 35308 52164 35364 52332
rect 35756 52274 35812 52668
rect 37324 52612 37380 53566
rect 38892 53618 38948 54460
rect 40236 54516 40292 54526
rect 40236 54422 40292 54460
rect 39900 54404 39956 54414
rect 39452 54348 39900 54404
rect 38892 53566 38894 53618
rect 38946 53566 38948 53618
rect 38892 53554 38948 53566
rect 39228 53732 39284 53742
rect 38332 53506 38388 53518
rect 38332 53454 38334 53506
rect 38386 53454 38388 53506
rect 38332 53172 38388 53454
rect 38332 53106 38388 53116
rect 39228 53170 39284 53676
rect 39228 53118 39230 53170
rect 39282 53118 39284 53170
rect 39228 53106 39284 53118
rect 39452 53396 39508 54348
rect 39900 54310 39956 54348
rect 40796 54292 40852 54684
rect 41244 54674 41300 54684
rect 41356 54738 41412 55132
rect 41356 54686 41358 54738
rect 41410 54686 41412 54738
rect 41356 54674 41412 54686
rect 41916 54628 41972 54638
rect 40908 54516 40964 54526
rect 40908 54514 41188 54516
rect 40908 54462 40910 54514
rect 40962 54462 41188 54514
rect 40908 54460 41188 54462
rect 40908 54450 40964 54460
rect 40796 54236 41076 54292
rect 40268 54124 40948 54134
rect 40324 54068 40372 54124
rect 40428 54122 40476 54124
rect 40532 54122 40580 54124
rect 40448 54070 40476 54122
rect 40572 54070 40580 54122
rect 40428 54068 40476 54070
rect 40532 54068 40580 54070
rect 40636 54122 40684 54124
rect 40740 54122 40788 54124
rect 40636 54070 40644 54122
rect 40740 54070 40768 54122
rect 40636 54068 40684 54070
rect 40740 54068 40788 54070
rect 40844 54068 40892 54124
rect 40268 54058 40948 54068
rect 39452 53170 39508 53340
rect 40124 53844 40180 53854
rect 39452 53118 39454 53170
rect 39506 53118 39508 53170
rect 39452 53106 39508 53118
rect 39564 53284 39620 53294
rect 37324 52546 37380 52556
rect 38444 52836 38500 52846
rect 35756 52222 35758 52274
rect 35810 52222 35812 52274
rect 35756 52210 35812 52222
rect 35308 52098 35364 52108
rect 36204 52164 36260 52174
rect 34188 51986 34244 51996
rect 32396 50766 32398 50818
rect 32450 50766 32452 50818
rect 32396 50754 32452 50766
rect 32956 51938 33012 51950
rect 32956 51886 32958 51938
rect 33010 51886 33012 51938
rect 29932 50594 29988 50606
rect 29932 50542 29934 50594
rect 29986 50542 29988 50594
rect 29932 50372 29988 50542
rect 32284 50484 32340 50494
rect 32844 50484 32900 50522
rect 32284 50482 32900 50484
rect 32284 50430 32286 50482
rect 32338 50430 32846 50482
rect 32898 50430 32900 50482
rect 32284 50428 32900 50430
rect 32284 50418 32340 50428
rect 29708 49924 29764 49934
rect 29596 49922 29764 49924
rect 29596 49870 29710 49922
rect 29762 49870 29764 49922
rect 29596 49868 29764 49870
rect 29708 49858 29764 49868
rect 28476 49646 28478 49698
rect 28530 49646 28532 49698
rect 22268 49420 22948 49430
rect 22324 49364 22372 49420
rect 22428 49418 22476 49420
rect 22532 49418 22580 49420
rect 22448 49366 22476 49418
rect 22572 49366 22580 49418
rect 22428 49364 22476 49366
rect 22532 49364 22580 49366
rect 22636 49418 22684 49420
rect 22740 49418 22788 49420
rect 22636 49366 22644 49418
rect 22740 49366 22768 49418
rect 22636 49364 22684 49366
rect 22740 49364 22788 49366
rect 22844 49364 22892 49420
rect 22268 49354 22948 49364
rect 20748 48804 20804 48814
rect 20748 48802 20916 48804
rect 20748 48750 20750 48802
rect 20802 48750 20916 48802
rect 20748 48748 20916 48750
rect 20748 48738 20804 48748
rect 16492 48078 16494 48130
rect 16546 48078 16548 48130
rect 16492 48020 16548 48078
rect 16492 47236 16548 47964
rect 20412 48076 20580 48132
rect 16492 47170 16548 47180
rect 17276 47348 17332 47358
rect 17276 47234 17332 47292
rect 17276 47182 17278 47234
rect 17330 47182 17332 47234
rect 17276 47170 17332 47182
rect 17612 47236 17668 47246
rect 17836 47236 17892 47246
rect 17668 47234 17892 47236
rect 17668 47182 17838 47234
rect 17890 47182 17892 47234
rect 17668 47180 17892 47182
rect 17612 46564 17668 47180
rect 17836 47170 17892 47180
rect 18172 47236 18228 47274
rect 20412 47236 20468 48076
rect 20748 48020 20804 48030
rect 20524 47964 20748 48020
rect 20524 47458 20580 47964
rect 20748 47954 20804 47964
rect 20524 47406 20526 47458
rect 20578 47406 20580 47458
rect 20524 47394 20580 47406
rect 20748 47460 20804 47470
rect 20860 47460 20916 48748
rect 26768 48636 27448 48646
rect 26824 48580 26872 48636
rect 26928 48634 26976 48636
rect 27032 48634 27080 48636
rect 26948 48582 26976 48634
rect 27072 48582 27080 48634
rect 26928 48580 26976 48582
rect 27032 48580 27080 48582
rect 27136 48634 27184 48636
rect 27240 48634 27288 48636
rect 27136 48582 27144 48634
rect 27240 48582 27268 48634
rect 27136 48580 27184 48582
rect 27240 48580 27288 48582
rect 27344 48580 27392 48636
rect 26768 48570 27448 48580
rect 21084 48132 21140 48142
rect 21084 48038 21140 48076
rect 22092 48132 22148 48142
rect 21420 48020 21476 48030
rect 21420 47926 21476 47964
rect 21196 47460 21252 47470
rect 20860 47458 21252 47460
rect 20860 47406 21198 47458
rect 21250 47406 21252 47458
rect 20860 47404 21252 47406
rect 20748 47346 20804 47404
rect 21196 47394 21252 47404
rect 21756 47460 21812 47470
rect 21756 47366 21812 47404
rect 20748 47294 20750 47346
rect 20802 47294 20804 47346
rect 20748 47282 20804 47294
rect 20524 47236 20580 47246
rect 20412 47180 20524 47236
rect 18172 47170 18228 47180
rect 20524 47170 20580 47180
rect 22092 47236 22148 48076
rect 22268 47852 22948 47862
rect 22324 47796 22372 47852
rect 22428 47850 22476 47852
rect 22532 47850 22580 47852
rect 22448 47798 22476 47850
rect 22572 47798 22580 47850
rect 22428 47796 22476 47798
rect 22532 47796 22580 47798
rect 22636 47850 22684 47852
rect 22740 47850 22788 47852
rect 22636 47798 22644 47850
rect 22740 47798 22768 47850
rect 22636 47796 22684 47798
rect 22740 47796 22788 47798
rect 22844 47796 22892 47852
rect 22268 47786 22948 47796
rect 22092 47170 22148 47180
rect 24108 47234 24164 47246
rect 24108 47182 24110 47234
rect 24162 47182 24164 47234
rect 20972 47124 21028 47134
rect 17768 47068 18448 47078
rect 17824 47012 17872 47068
rect 17928 47066 17976 47068
rect 18032 47066 18080 47068
rect 17948 47014 17976 47066
rect 18072 47014 18080 47066
rect 17928 47012 17976 47014
rect 18032 47012 18080 47014
rect 18136 47066 18184 47068
rect 18240 47066 18288 47068
rect 18136 47014 18144 47066
rect 18240 47014 18268 47066
rect 18136 47012 18184 47014
rect 18240 47012 18288 47014
rect 18344 47012 18392 47068
rect 17768 47002 18448 47012
rect 20972 46898 21028 47068
rect 20972 46846 20974 46898
rect 21026 46846 21028 46898
rect 20972 46834 21028 46846
rect 21532 47124 21588 47134
rect 17612 46498 17668 46508
rect 21308 45666 21364 45678
rect 21308 45614 21310 45666
rect 21362 45614 21364 45666
rect 17768 45500 18448 45510
rect 17824 45444 17872 45500
rect 17928 45498 17976 45500
rect 18032 45498 18080 45500
rect 17948 45446 17976 45498
rect 18072 45446 18080 45498
rect 17928 45444 17976 45446
rect 18032 45444 18080 45446
rect 18136 45498 18184 45500
rect 18240 45498 18288 45500
rect 18136 45446 18144 45498
rect 18240 45446 18268 45498
rect 18136 45444 18184 45446
rect 18240 45444 18288 45446
rect 18344 45444 18392 45500
rect 17768 45434 18448 45444
rect 20300 45332 20356 45342
rect 20300 45330 21140 45332
rect 20300 45278 20302 45330
rect 20354 45278 21140 45330
rect 20300 45276 21140 45278
rect 20300 45266 20356 45276
rect 17388 45220 17444 45230
rect 16492 45108 16548 45118
rect 16492 45014 16548 45052
rect 16156 44884 16212 44894
rect 16156 44790 16212 44828
rect 17388 44212 17444 45164
rect 19628 45220 19684 45230
rect 19628 45126 19684 45164
rect 20076 45106 20132 45118
rect 20076 45054 20078 45106
rect 20130 45054 20132 45106
rect 17388 44098 17444 44156
rect 17388 44046 17390 44098
rect 17442 44046 17444 44098
rect 17388 44034 17444 44046
rect 17612 44994 17668 45006
rect 17612 44942 17614 44994
rect 17666 44942 17668 44994
rect 17612 44884 17668 44942
rect 17612 44100 17668 44828
rect 20076 44436 20132 45054
rect 20748 45106 20804 45118
rect 20748 45054 20750 45106
rect 20802 45054 20804 45106
rect 20748 44884 20804 45054
rect 21084 45106 21140 45276
rect 21084 45054 21086 45106
rect 21138 45054 21140 45106
rect 21084 45042 21140 45054
rect 21308 44884 21364 45614
rect 20748 44828 21364 44884
rect 20076 44370 20132 44380
rect 21420 44548 21476 44558
rect 21420 44210 21476 44492
rect 21420 44158 21422 44210
rect 21474 44158 21476 44210
rect 21420 44146 21476 44158
rect 17948 44100 18004 44138
rect 17612 44044 17948 44100
rect 17948 44034 18004 44044
rect 20748 44098 20804 44110
rect 20748 44046 20750 44098
rect 20802 44046 20804 44098
rect 17768 43932 18448 43942
rect 17824 43876 17872 43932
rect 17928 43930 17976 43932
rect 18032 43930 18080 43932
rect 17948 43878 17976 43930
rect 18072 43878 18080 43930
rect 17928 43876 17976 43878
rect 18032 43876 18080 43878
rect 18136 43930 18184 43932
rect 18240 43930 18288 43932
rect 18136 43878 18144 43930
rect 18240 43878 18268 43930
rect 18136 43876 18184 43878
rect 18240 43876 18288 43878
rect 18344 43876 18392 43932
rect 17768 43866 18448 43876
rect 20748 43652 20804 44046
rect 20748 42868 20804 43596
rect 20748 42802 20804 42812
rect 18956 42756 19012 42766
rect 18956 42662 19012 42700
rect 19516 42756 19572 42766
rect 19516 42662 19572 42700
rect 20188 42756 20244 42766
rect 20188 42662 20244 42700
rect 15596 42578 15652 42588
rect 19404 42644 19460 42654
rect 19404 42550 19460 42588
rect 14364 42466 14420 42476
rect 15260 42532 15316 42542
rect 15260 42438 15316 42476
rect 16940 42532 16996 42542
rect 20524 42532 20580 42542
rect 21308 42532 21364 42542
rect 13804 41918 13806 41970
rect 13858 41918 13860 41970
rect 13804 41906 13860 41918
rect 16380 42194 16436 42206
rect 16380 42142 16382 42194
rect 16434 42142 16436 42194
rect 16380 41972 16436 42142
rect 16380 41906 16436 41916
rect 16940 41748 16996 42476
rect 20188 42530 20580 42532
rect 20188 42478 20526 42530
rect 20578 42478 20580 42530
rect 20188 42476 20580 42478
rect 17768 42364 18448 42374
rect 17824 42308 17872 42364
rect 17928 42362 17976 42364
rect 18032 42362 18080 42364
rect 17948 42310 17976 42362
rect 18072 42310 18080 42362
rect 17928 42308 17976 42310
rect 18032 42308 18080 42310
rect 18136 42362 18184 42364
rect 18240 42362 18288 42364
rect 18136 42310 18144 42362
rect 18240 42310 18268 42362
rect 18136 42308 18184 42310
rect 18240 42308 18288 42310
rect 18344 42308 18392 42364
rect 17768 42298 18448 42308
rect 17500 41972 17556 41982
rect 17500 41878 17556 41916
rect 19740 41972 19796 41982
rect 19740 41878 19796 41916
rect 20188 41970 20244 42476
rect 20524 42466 20580 42476
rect 20636 42530 21364 42532
rect 20636 42478 21310 42530
rect 21362 42478 21364 42530
rect 20636 42476 21364 42478
rect 20188 41918 20190 41970
rect 20242 41918 20244 41970
rect 20188 41906 20244 41918
rect 20412 42082 20468 42094
rect 20412 42030 20414 42082
rect 20466 42030 20468 42082
rect 17612 41748 17668 41758
rect 16940 41746 17108 41748
rect 16940 41694 16942 41746
rect 16994 41694 17108 41746
rect 16940 41692 17108 41694
rect 16940 41682 16996 41692
rect 13268 41580 13948 41590
rect 13324 41524 13372 41580
rect 13428 41578 13476 41580
rect 13532 41578 13580 41580
rect 13448 41526 13476 41578
rect 13572 41526 13580 41578
rect 13428 41524 13476 41526
rect 13532 41524 13580 41526
rect 13636 41578 13684 41580
rect 13740 41578 13788 41580
rect 13636 41526 13644 41578
rect 13740 41526 13768 41578
rect 13636 41524 13684 41526
rect 13740 41524 13788 41526
rect 13844 41524 13892 41580
rect 13268 41514 13948 41524
rect 13132 41346 13188 41356
rect 12348 40964 12404 40974
rect 12348 40626 12404 40908
rect 12348 40574 12350 40626
rect 12402 40574 12404 40626
rect 12348 40562 12404 40574
rect 16828 40514 16884 40526
rect 16828 40462 16830 40514
rect 16882 40462 16884 40514
rect 13580 40402 13636 40414
rect 13580 40350 13582 40402
rect 13634 40350 13636 40402
rect 13132 40180 13188 40190
rect 11900 40178 13188 40180
rect 11900 40126 13134 40178
rect 13186 40126 13188 40178
rect 11900 40124 13188 40126
rect 11676 39618 11732 39630
rect 11676 39566 11678 39618
rect 11730 39566 11732 39618
rect 11228 39396 11284 39406
rect 11676 39396 11732 39566
rect 11900 39506 11956 40124
rect 13132 40114 13188 40124
rect 13580 40180 13636 40350
rect 16828 40404 16884 40462
rect 16940 40404 16996 40414
rect 16828 40348 16940 40404
rect 13580 40114 13636 40124
rect 16828 40180 16884 40190
rect 13268 40012 13948 40022
rect 12460 39956 12516 39966
rect 13324 39956 13372 40012
rect 13428 40010 13476 40012
rect 13532 40010 13580 40012
rect 13448 39958 13476 40010
rect 13572 39958 13580 40010
rect 13428 39956 13476 39958
rect 13532 39956 13580 39958
rect 13636 40010 13684 40012
rect 13740 40010 13788 40012
rect 13636 39958 13644 40010
rect 13740 39958 13768 40010
rect 13636 39956 13684 39958
rect 13740 39956 13788 39958
rect 13844 39956 13892 40012
rect 13268 39946 13948 39956
rect 12460 39842 12516 39900
rect 12460 39790 12462 39842
rect 12514 39790 12516 39842
rect 12460 39778 12516 39790
rect 15484 39620 15540 39630
rect 11900 39454 11902 39506
rect 11954 39454 11956 39506
rect 11900 39442 11956 39454
rect 12796 39508 12852 39518
rect 12796 39414 12852 39452
rect 13468 39508 13524 39518
rect 13468 39414 13524 39452
rect 11228 39394 11732 39396
rect 11228 39342 11230 39394
rect 11282 39342 11732 39394
rect 11228 39340 11732 39342
rect 11788 39396 11844 39406
rect 10556 37380 10612 37390
rect 10556 37286 10612 37324
rect 11228 37156 11284 39340
rect 11340 37156 11396 37166
rect 11228 37154 11396 37156
rect 11228 37102 11342 37154
rect 11394 37102 11396 37154
rect 11228 37100 11396 37102
rect 11340 36932 11396 37100
rect 11340 36866 11396 36876
rect 11564 36260 11620 36270
rect 11564 36166 11620 36204
rect 11340 34690 11396 34702
rect 11340 34638 11342 34690
rect 11394 34638 11396 34690
rect 11340 34130 11396 34638
rect 11340 34078 11342 34130
rect 11394 34078 11396 34130
rect 11340 34066 11396 34078
rect 11788 34130 11844 39340
rect 13356 39396 13412 39406
rect 13356 38834 13412 39340
rect 13356 38782 13358 38834
rect 13410 38782 13412 38834
rect 13356 38770 13412 38782
rect 13804 39394 13860 39406
rect 13804 39342 13806 39394
rect 13858 39342 13860 39394
rect 13804 38834 13860 39342
rect 14140 39396 14196 39406
rect 14140 39302 14196 39340
rect 13804 38782 13806 38834
rect 13858 38782 13860 38834
rect 13804 38770 13860 38782
rect 13268 38444 13948 38454
rect 13324 38388 13372 38444
rect 13428 38442 13476 38444
rect 13532 38442 13580 38444
rect 13448 38390 13476 38442
rect 13572 38390 13580 38442
rect 13428 38388 13476 38390
rect 13532 38388 13580 38390
rect 13636 38442 13684 38444
rect 13740 38442 13788 38444
rect 13636 38390 13644 38442
rect 13740 38390 13768 38442
rect 13636 38388 13684 38390
rect 13740 38388 13788 38390
rect 13844 38388 13892 38444
rect 13268 38378 13948 38388
rect 15260 37378 15316 37390
rect 15260 37326 15262 37378
rect 15314 37326 15316 37378
rect 11900 37154 11956 37166
rect 11900 37102 11902 37154
rect 11954 37102 11956 37154
rect 11900 37044 11956 37102
rect 11900 36484 11956 36988
rect 13268 36876 13948 36886
rect 13324 36820 13372 36876
rect 13428 36874 13476 36876
rect 13532 36874 13580 36876
rect 13448 36822 13476 36874
rect 13572 36822 13580 36874
rect 13428 36820 13476 36822
rect 13532 36820 13580 36822
rect 13636 36874 13684 36876
rect 13740 36874 13788 36876
rect 13636 36822 13644 36874
rect 13740 36822 13768 36874
rect 13636 36820 13684 36822
rect 13740 36820 13788 36822
rect 13844 36820 13892 36876
rect 13268 36810 13948 36820
rect 12348 36484 12404 36494
rect 14812 36484 14868 36494
rect 11900 36428 12348 36484
rect 12348 36390 12404 36428
rect 14588 36482 14868 36484
rect 14588 36430 14814 36482
rect 14866 36430 14868 36482
rect 14588 36428 14868 36430
rect 15260 36484 15316 37326
rect 15372 36484 15428 36494
rect 15260 36482 15428 36484
rect 15260 36430 15374 36482
rect 15426 36430 15428 36482
rect 15260 36428 15428 36430
rect 14588 36370 14644 36428
rect 14812 36418 14868 36428
rect 15372 36418 15428 36428
rect 14588 36318 14590 36370
rect 14642 36318 14644 36370
rect 14588 36306 14644 36318
rect 15484 35810 15540 39564
rect 16268 39060 16324 39070
rect 16268 38966 16324 39004
rect 16828 38724 16884 40124
rect 16828 38658 16884 38668
rect 16940 38500 16996 40348
rect 17052 38668 17108 41692
rect 20412 41748 20468 42030
rect 20636 41970 20692 42476
rect 21308 42466 21364 42476
rect 21196 41972 21252 41982
rect 20636 41918 20638 41970
rect 20690 41918 20692 41970
rect 20636 41906 20692 41918
rect 20748 41970 21252 41972
rect 20748 41918 21198 41970
rect 21250 41918 21252 41970
rect 20748 41916 21252 41918
rect 20748 41748 20804 41916
rect 21196 41906 21252 41916
rect 21532 41972 21588 47068
rect 24108 47124 24164 47182
rect 24108 47058 24164 47068
rect 24892 47236 24948 47246
rect 24892 46900 24948 47180
rect 26768 47068 27448 47078
rect 26824 47012 26872 47068
rect 26928 47066 26976 47068
rect 27032 47066 27080 47068
rect 26948 47014 26976 47066
rect 27072 47014 27080 47066
rect 26928 47012 26976 47014
rect 27032 47012 27080 47014
rect 27136 47066 27184 47068
rect 27240 47066 27288 47068
rect 27136 47014 27144 47066
rect 27240 47014 27268 47066
rect 27136 47012 27184 47014
rect 27240 47012 27288 47014
rect 27344 47012 27392 47068
rect 26768 47002 27448 47012
rect 24892 46834 24948 46844
rect 25676 46674 25732 46686
rect 25676 46622 25678 46674
rect 25730 46622 25732 46674
rect 22268 46284 22948 46294
rect 22324 46228 22372 46284
rect 22428 46282 22476 46284
rect 22532 46282 22580 46284
rect 22448 46230 22476 46282
rect 22572 46230 22580 46282
rect 22428 46228 22476 46230
rect 22532 46228 22580 46230
rect 22636 46282 22684 46284
rect 22740 46282 22788 46284
rect 22636 46230 22644 46282
rect 22740 46230 22768 46282
rect 22636 46228 22684 46230
rect 22740 46228 22788 46230
rect 22844 46228 22892 46284
rect 22268 46218 22948 46228
rect 25676 45778 25732 46622
rect 26124 46676 26180 46686
rect 26124 46582 26180 46620
rect 26908 46676 26964 46686
rect 25676 45726 25678 45778
rect 25730 45726 25732 45778
rect 25676 45714 25732 45726
rect 26908 45778 26964 46620
rect 27244 46452 27300 46462
rect 27244 45890 27300 46396
rect 27244 45838 27246 45890
rect 27298 45838 27300 45890
rect 27244 45826 27300 45838
rect 26908 45726 26910 45778
rect 26962 45726 26964 45778
rect 26908 45714 26964 45726
rect 28476 45556 28532 49646
rect 29036 49812 29092 49822
rect 29036 49140 29092 49756
rect 29932 49700 29988 50316
rect 29932 49634 29988 49644
rect 31948 49700 32004 49710
rect 32004 49644 32116 49700
rect 31948 49606 32004 49644
rect 31268 49420 31948 49430
rect 31324 49364 31372 49420
rect 31428 49418 31476 49420
rect 31532 49418 31580 49420
rect 31448 49366 31476 49418
rect 31572 49366 31580 49418
rect 31428 49364 31476 49366
rect 31532 49364 31580 49366
rect 31636 49418 31684 49420
rect 31740 49418 31788 49420
rect 31636 49366 31644 49418
rect 31740 49366 31768 49418
rect 31636 49364 31684 49366
rect 31740 49364 31788 49366
rect 31844 49364 31892 49420
rect 31268 49354 31948 49364
rect 29260 49140 29316 49150
rect 29036 49084 29260 49140
rect 29260 49046 29316 49084
rect 31268 47852 31948 47862
rect 31324 47796 31372 47852
rect 31428 47850 31476 47852
rect 31532 47850 31580 47852
rect 31448 47798 31476 47850
rect 31572 47798 31580 47850
rect 31428 47796 31476 47798
rect 31532 47796 31580 47798
rect 31636 47850 31684 47852
rect 31740 47850 31788 47852
rect 31636 47798 31644 47850
rect 31740 47798 31768 47850
rect 31636 47796 31684 47798
rect 31740 47796 31788 47798
rect 31844 47796 31892 47852
rect 31268 47786 31948 47796
rect 30380 47572 30436 47582
rect 26768 45500 27448 45510
rect 26824 45444 26872 45500
rect 26928 45498 26976 45500
rect 27032 45498 27080 45500
rect 26948 45446 26976 45498
rect 27072 45446 27080 45498
rect 26928 45444 26976 45446
rect 27032 45444 27080 45446
rect 27136 45498 27184 45500
rect 27240 45498 27288 45500
rect 27136 45446 27144 45498
rect 27240 45446 27268 45498
rect 27136 45444 27184 45446
rect 27240 45444 27288 45446
rect 27344 45444 27392 45500
rect 26768 45434 27448 45444
rect 28364 45500 28532 45556
rect 28588 46898 28644 46910
rect 28588 46846 28590 46898
rect 28642 46846 28644 46898
rect 28588 45780 28644 46846
rect 30380 46786 30436 47516
rect 31612 47572 31668 47582
rect 31164 47236 31220 47246
rect 30380 46734 30382 46786
rect 30434 46734 30436 46786
rect 30380 46722 30436 46734
rect 31052 47234 31220 47236
rect 31052 47182 31166 47234
rect 31218 47182 31220 47234
rect 31052 47180 31220 47182
rect 30604 46676 30660 46686
rect 31052 46676 31108 47180
rect 31164 47170 31220 47180
rect 31612 46898 31668 47516
rect 31612 46846 31614 46898
rect 31666 46846 31668 46898
rect 31612 46834 31668 46846
rect 30604 46674 30772 46676
rect 30604 46622 30606 46674
rect 30658 46622 30772 46674
rect 30604 46620 30772 46622
rect 30604 46610 30660 46620
rect 29148 46564 29204 46574
rect 29148 46470 29204 46508
rect 29820 46564 29876 46574
rect 29820 46470 29876 46508
rect 29484 46452 29540 46462
rect 29484 46358 29540 46396
rect 23436 45220 23492 45230
rect 23436 45126 23492 45164
rect 24220 44882 24276 44894
rect 24220 44830 24222 44882
rect 24274 44830 24276 44882
rect 22268 44716 22948 44726
rect 22324 44660 22372 44716
rect 22428 44714 22476 44716
rect 22532 44714 22580 44716
rect 22448 44662 22476 44714
rect 22572 44662 22580 44714
rect 22428 44660 22476 44662
rect 22532 44660 22580 44662
rect 22636 44714 22684 44716
rect 22740 44714 22788 44716
rect 22636 44662 22644 44714
rect 22740 44662 22768 44714
rect 22636 44660 22684 44662
rect 22740 44660 22788 44662
rect 22844 44660 22892 44716
rect 22268 44650 22948 44660
rect 22540 44436 22596 44446
rect 22540 44342 22596 44380
rect 21756 44322 21812 44334
rect 21756 44270 21758 44322
rect 21810 44270 21812 44322
rect 21756 43652 21812 44270
rect 22204 44322 22260 44334
rect 22204 44270 22206 44322
rect 22258 44270 22260 44322
rect 22204 44100 22260 44270
rect 22204 44034 22260 44044
rect 23100 44100 23156 44110
rect 23100 44006 23156 44044
rect 24220 44100 24276 44830
rect 24220 44034 24276 44044
rect 26768 43932 27448 43942
rect 26824 43876 26872 43932
rect 26928 43930 26976 43932
rect 27032 43930 27080 43932
rect 26948 43878 26976 43930
rect 27072 43878 27080 43930
rect 26928 43876 26976 43878
rect 27032 43876 27080 43878
rect 27136 43930 27184 43932
rect 27240 43930 27288 43932
rect 27136 43878 27144 43930
rect 27240 43878 27268 43930
rect 27136 43876 27184 43878
rect 27240 43876 27288 43878
rect 27344 43876 27392 43932
rect 26768 43866 27448 43876
rect 21756 43586 21812 43596
rect 25340 43650 25396 43662
rect 25340 43598 25342 43650
rect 25394 43598 25396 43650
rect 25340 43540 25396 43598
rect 25564 43540 25620 43550
rect 25340 43538 25620 43540
rect 25340 43486 25566 43538
rect 25618 43486 25620 43538
rect 25340 43484 25620 43486
rect 25564 43474 25620 43484
rect 26236 43538 26292 43550
rect 26236 43486 26238 43538
rect 26290 43486 26292 43538
rect 22268 43148 22948 43158
rect 22324 43092 22372 43148
rect 22428 43146 22476 43148
rect 22532 43146 22580 43148
rect 22448 43094 22476 43146
rect 22572 43094 22580 43146
rect 22428 43092 22476 43094
rect 22532 43092 22580 43094
rect 22636 43146 22684 43148
rect 22740 43146 22788 43148
rect 22636 43094 22644 43146
rect 22740 43094 22768 43146
rect 22636 43092 22684 43094
rect 22740 43092 22788 43094
rect 22844 43092 22892 43148
rect 22268 43082 22948 43092
rect 21868 42756 21924 42766
rect 21868 42530 21924 42700
rect 26236 42644 26292 43486
rect 27244 43316 27300 43326
rect 27244 42754 27300 43260
rect 27244 42702 27246 42754
rect 27298 42702 27300 42754
rect 27244 42690 27300 42702
rect 28252 42868 28308 42878
rect 26236 42578 26292 42588
rect 26908 42644 26964 42654
rect 26908 42550 26964 42588
rect 21868 42478 21870 42530
rect 21922 42478 21924 42530
rect 21868 42084 21924 42478
rect 26768 42364 27448 42374
rect 26824 42308 26872 42364
rect 26928 42362 26976 42364
rect 27032 42362 27080 42364
rect 26948 42310 26976 42362
rect 27072 42310 27080 42362
rect 26928 42308 26976 42310
rect 27032 42308 27080 42310
rect 27136 42362 27184 42364
rect 27240 42362 27288 42364
rect 27136 42310 27144 42362
rect 27240 42310 27268 42362
rect 27136 42308 27184 42310
rect 27240 42308 27288 42310
rect 27344 42308 27392 42364
rect 26768 42298 27448 42308
rect 21868 42018 21924 42028
rect 23548 42082 23604 42094
rect 23548 42030 23550 42082
rect 23602 42030 23604 42082
rect 21532 41906 21588 41916
rect 21980 41972 22036 41982
rect 20412 41692 20804 41748
rect 17612 40514 17668 41692
rect 18508 41076 18564 41086
rect 17768 40796 18448 40806
rect 17824 40740 17872 40796
rect 17928 40794 17976 40796
rect 18032 40794 18080 40796
rect 17948 40742 17976 40794
rect 18072 40742 18080 40794
rect 17928 40740 17976 40742
rect 18032 40740 18080 40742
rect 18136 40794 18184 40796
rect 18240 40794 18288 40796
rect 18136 40742 18144 40794
rect 18240 40742 18268 40794
rect 18136 40740 18184 40742
rect 18240 40740 18288 40742
rect 18344 40740 18392 40796
rect 17768 40730 18448 40740
rect 18508 40628 18564 41020
rect 19068 41076 19124 41086
rect 19068 40982 19124 41020
rect 17612 40462 17614 40514
rect 17666 40462 17668 40514
rect 17612 40450 17668 40462
rect 18284 40572 18564 40628
rect 21084 40628 21140 40638
rect 17500 40404 17556 40414
rect 17500 40310 17556 40348
rect 18284 40290 18340 40572
rect 18620 40404 18676 40414
rect 18284 40238 18286 40290
rect 18338 40238 18340 40290
rect 18284 40226 18340 40238
rect 18396 40402 18676 40404
rect 18396 40350 18622 40402
rect 18674 40350 18676 40402
rect 18396 40348 18676 40350
rect 18396 39618 18452 40348
rect 18620 40338 18676 40348
rect 19180 40404 19236 40414
rect 19516 40404 19572 40414
rect 19180 40402 19348 40404
rect 19180 40350 19182 40402
rect 19234 40350 19348 40402
rect 19180 40348 19348 40350
rect 19180 40338 19236 40348
rect 18396 39566 18398 39618
rect 18450 39566 18452 39618
rect 18396 39554 18452 39566
rect 19292 39506 19348 40348
rect 19292 39454 19294 39506
rect 19346 39454 19348 39506
rect 19292 39442 19348 39454
rect 19404 40402 19572 40404
rect 19404 40350 19518 40402
rect 19570 40350 19572 40402
rect 19404 40348 19572 40350
rect 18620 39394 18676 39406
rect 18620 39342 18622 39394
rect 18674 39342 18676 39394
rect 18620 39284 18676 39342
rect 19404 39284 19460 40348
rect 19516 40338 19572 40348
rect 17768 39228 18448 39238
rect 18620 39228 19460 39284
rect 17824 39172 17872 39228
rect 17928 39226 17976 39228
rect 18032 39226 18080 39228
rect 17948 39174 17976 39226
rect 18072 39174 18080 39226
rect 17928 39172 17976 39174
rect 18032 39172 18080 39174
rect 18136 39226 18184 39228
rect 18240 39226 18288 39228
rect 18136 39174 18144 39226
rect 18240 39174 18268 39226
rect 18136 39172 18184 39174
rect 18240 39172 18288 39174
rect 18344 39172 18392 39228
rect 17768 39162 18448 39172
rect 17500 39060 17556 39070
rect 17500 38668 17556 39004
rect 21084 39058 21140 40572
rect 21980 40628 22036 41916
rect 23548 41972 23604 42030
rect 24444 42084 24500 42094
rect 24444 41990 24500 42028
rect 23548 41906 23604 41916
rect 22268 41580 22948 41590
rect 22324 41524 22372 41580
rect 22428 41578 22476 41580
rect 22532 41578 22580 41580
rect 22448 41526 22476 41578
rect 22572 41526 22580 41578
rect 22428 41524 22476 41526
rect 22532 41524 22580 41526
rect 22636 41578 22684 41580
rect 22740 41578 22788 41580
rect 22636 41526 22644 41578
rect 22740 41526 22768 41578
rect 22636 41524 22684 41526
rect 22740 41524 22788 41526
rect 22844 41524 22892 41580
rect 22268 41514 22948 41524
rect 21980 40534 22036 40572
rect 22652 41076 22708 41086
rect 22652 40626 22708 41020
rect 25452 40962 25508 40974
rect 25452 40910 25454 40962
rect 25506 40910 25508 40962
rect 22652 40574 22654 40626
rect 22706 40574 22708 40626
rect 22652 40562 22708 40574
rect 22988 40628 23044 40638
rect 22988 40534 23044 40572
rect 25452 40402 25508 40910
rect 26768 40796 27448 40806
rect 26824 40740 26872 40796
rect 26928 40794 26976 40796
rect 27032 40794 27080 40796
rect 26948 40742 26976 40794
rect 27072 40742 27080 40794
rect 26928 40740 26976 40742
rect 27032 40740 27080 40742
rect 27136 40794 27184 40796
rect 27240 40794 27288 40796
rect 27136 40742 27144 40794
rect 27240 40742 27268 40794
rect 27136 40740 27184 40742
rect 27240 40740 27288 40742
rect 27344 40740 27392 40796
rect 26768 40730 27448 40740
rect 28252 40626 28308 42812
rect 28364 41972 28420 45500
rect 28588 43762 28644 45724
rect 29260 45780 29316 45790
rect 29260 45686 29316 45724
rect 30604 45780 30660 45790
rect 30604 45686 30660 45724
rect 30716 45668 30772 46620
rect 30940 46620 31108 46676
rect 30940 45890 30996 46620
rect 31164 46562 31220 46574
rect 31164 46510 31166 46562
rect 31218 46510 31220 46562
rect 31164 46452 31220 46510
rect 30940 45838 30942 45890
rect 30994 45838 30996 45890
rect 30940 45826 30996 45838
rect 31052 46396 31220 46452
rect 31052 45668 31108 46396
rect 31268 46284 31948 46294
rect 31324 46228 31372 46284
rect 31428 46282 31476 46284
rect 31532 46282 31580 46284
rect 31448 46230 31476 46282
rect 31572 46230 31580 46282
rect 31428 46228 31476 46230
rect 31532 46228 31580 46230
rect 31636 46282 31684 46284
rect 31740 46282 31788 46284
rect 31636 46230 31644 46282
rect 31740 46230 31768 46282
rect 31636 46228 31684 46230
rect 31740 46228 31788 46230
rect 31844 46228 31892 46284
rect 31268 46218 31948 46228
rect 31500 46116 31556 46126
rect 31500 45890 31556 46060
rect 31500 45838 31502 45890
rect 31554 45838 31556 45890
rect 31500 45826 31556 45838
rect 32060 45892 32116 49644
rect 32508 49698 32564 49710
rect 32508 49646 32510 49698
rect 32562 49646 32564 49698
rect 32284 49140 32340 49150
rect 32508 49140 32564 49646
rect 32844 49252 32900 50428
rect 32844 49186 32900 49196
rect 32340 49084 32564 49140
rect 32956 49138 33012 51886
rect 36204 51940 36260 52108
rect 37996 52052 38052 52062
rect 36204 51884 36596 51940
rect 35768 51772 36448 51782
rect 35824 51716 35872 51772
rect 35928 51770 35976 51772
rect 36032 51770 36080 51772
rect 35948 51718 35976 51770
rect 36072 51718 36080 51770
rect 35928 51716 35976 51718
rect 36032 51716 36080 51718
rect 36136 51770 36184 51772
rect 36240 51770 36288 51772
rect 36136 51718 36144 51770
rect 36240 51718 36268 51770
rect 36136 51716 36184 51718
rect 36240 51716 36288 51718
rect 36344 51716 36392 51772
rect 35768 51706 36448 51716
rect 36540 51380 36596 51884
rect 37996 51602 38052 51996
rect 37996 51550 37998 51602
rect 38050 51550 38052 51602
rect 37996 51538 38052 51550
rect 38444 51604 38500 52780
rect 38892 52834 38948 52846
rect 38892 52782 38894 52834
rect 38946 52782 38948 52834
rect 38892 52052 38948 52782
rect 39564 52834 39620 53228
rect 39564 52782 39566 52834
rect 39618 52782 39620 52834
rect 39564 52770 39620 52782
rect 39676 52946 39732 52958
rect 39676 52894 39678 52946
rect 39730 52894 39732 52946
rect 38892 51986 38948 51996
rect 39228 52612 39284 52622
rect 38668 51604 38724 51614
rect 38444 51548 38668 51604
rect 38668 51490 38724 51548
rect 38668 51438 38670 51490
rect 38722 51438 38724 51490
rect 36540 51314 36596 51324
rect 38444 51380 38500 51390
rect 38444 51286 38500 51324
rect 38556 50708 38612 50718
rect 38668 50708 38724 51438
rect 38556 50706 38724 50708
rect 38556 50654 38558 50706
rect 38610 50654 38724 50706
rect 38556 50652 38724 50654
rect 39116 51380 39172 51390
rect 39116 50706 39172 51324
rect 39228 51378 39284 52556
rect 39228 51326 39230 51378
rect 39282 51326 39284 51378
rect 39228 51314 39284 51326
rect 39564 52052 39620 52062
rect 39564 51492 39620 51996
rect 39116 50654 39118 50706
rect 39170 50654 39172 50706
rect 38556 50642 38612 50652
rect 39116 50642 39172 50654
rect 39564 50706 39620 51436
rect 39676 51604 39732 52894
rect 40124 52834 40180 53788
rect 40796 53620 40852 53630
rect 41020 53620 41076 54236
rect 40796 53618 41076 53620
rect 40796 53566 40798 53618
rect 40850 53566 41076 53618
rect 40796 53564 41076 53566
rect 40796 53554 40852 53564
rect 41132 53396 41188 54460
rect 41468 54514 41524 54526
rect 41468 54462 41470 54514
rect 41522 54462 41524 54514
rect 41468 54404 41524 54462
rect 41916 54404 41972 54572
rect 42588 54516 42644 55358
rect 42924 55188 42980 55198
rect 42588 54450 42644 54460
rect 42700 55186 42980 55188
rect 42700 55134 42926 55186
rect 42978 55134 42980 55186
rect 42700 55132 42980 55134
rect 41468 54402 41972 54404
rect 41468 54350 41918 54402
rect 41970 54350 41972 54402
rect 41468 54348 41972 54350
rect 41468 53844 41524 54348
rect 41916 54338 41972 54348
rect 41468 53778 41524 53788
rect 41356 53730 41412 53742
rect 41356 53678 41358 53730
rect 41410 53678 41412 53730
rect 40908 53340 41188 53396
rect 41244 53506 41300 53518
rect 41244 53454 41246 53506
rect 41298 53454 41300 53506
rect 40908 53284 40964 53340
rect 40908 53058 40964 53228
rect 40908 53006 40910 53058
rect 40962 53006 40964 53058
rect 40908 52994 40964 53006
rect 41132 52948 41188 52958
rect 41244 52948 41300 53454
rect 41356 53172 41412 53678
rect 41692 53730 41748 53742
rect 41692 53678 41694 53730
rect 41746 53678 41748 53730
rect 41356 53116 41524 53172
rect 41356 52948 41412 52958
rect 41244 52946 41412 52948
rect 41244 52894 41358 52946
rect 41410 52894 41412 52946
rect 41244 52892 41412 52894
rect 41132 52854 41188 52892
rect 41356 52882 41412 52892
rect 40124 52782 40126 52834
rect 40178 52782 40180 52834
rect 40124 52612 40180 52782
rect 41020 52834 41076 52846
rect 41020 52782 41022 52834
rect 41074 52782 41076 52834
rect 40124 52546 40180 52556
rect 40268 52556 40948 52566
rect 40324 52500 40372 52556
rect 40428 52554 40476 52556
rect 40532 52554 40580 52556
rect 40448 52502 40476 52554
rect 40572 52502 40580 52554
rect 40428 52500 40476 52502
rect 40532 52500 40580 52502
rect 40636 52554 40684 52556
rect 40740 52554 40788 52556
rect 40636 52502 40644 52554
rect 40740 52502 40768 52554
rect 40636 52500 40684 52502
rect 40740 52500 40788 52502
rect 40844 52500 40892 52556
rect 40268 52490 40948 52500
rect 41020 51716 41076 52782
rect 41468 52500 41524 53116
rect 41468 52434 41524 52444
rect 41580 52946 41636 52958
rect 41580 52894 41582 52946
rect 41634 52894 41636 52946
rect 41580 52388 41636 52894
rect 41692 52724 41748 53678
rect 42252 53620 42308 53630
rect 41692 52658 41748 52668
rect 41916 53618 42308 53620
rect 41916 53566 42254 53618
rect 42306 53566 42308 53618
rect 41916 53564 42308 53566
rect 41916 53060 41972 53564
rect 42252 53554 42308 53564
rect 41020 51660 41188 51716
rect 39676 51378 39732 51548
rect 39676 51326 39678 51378
rect 39730 51326 39732 51378
rect 39676 51314 39732 51326
rect 40124 51604 40180 51614
rect 39788 51268 39844 51278
rect 39788 51266 40068 51268
rect 39788 51214 39790 51266
rect 39842 51214 40068 51266
rect 39788 51212 40068 51214
rect 39788 51202 39844 51212
rect 39564 50654 39566 50706
rect 39618 50654 39620 50706
rect 39564 50642 39620 50654
rect 39900 50596 39956 50606
rect 32956 49086 32958 49138
rect 33010 49086 33012 49138
rect 32284 49026 32340 49084
rect 32956 49074 33012 49086
rect 33740 50484 33796 50494
rect 32284 48974 32286 49026
rect 32338 48974 32340 49026
rect 32284 48962 32340 48974
rect 32508 47236 32564 47246
rect 32172 46786 32228 46798
rect 32172 46734 32174 46786
rect 32226 46734 32228 46786
rect 32172 46116 32228 46734
rect 32508 46786 32564 47180
rect 33628 47236 33684 47246
rect 33628 47142 33684 47180
rect 32508 46734 32510 46786
rect 32562 46734 32564 46786
rect 32508 46722 32564 46734
rect 33292 46676 33348 46686
rect 33292 46582 33348 46620
rect 32172 46050 32228 46060
rect 32060 45836 32228 45892
rect 30716 45612 31108 45668
rect 30604 44436 30660 44446
rect 28588 43710 28590 43762
rect 28642 43710 28644 43762
rect 28588 42868 28644 43710
rect 30492 44380 30604 44436
rect 30492 43650 30548 44380
rect 30604 44370 30660 44380
rect 30492 43598 30494 43650
rect 30546 43598 30548 43650
rect 30492 43586 30548 43598
rect 29260 43540 29316 43550
rect 29260 43446 29316 43484
rect 29932 43540 29988 43550
rect 29932 43446 29988 43484
rect 30604 43538 30660 43550
rect 30604 43486 30606 43538
rect 30658 43486 30660 43538
rect 30604 43428 30660 43486
rect 30940 43428 30996 45612
rect 31268 44716 31948 44726
rect 31324 44660 31372 44716
rect 31428 44714 31476 44716
rect 31532 44714 31580 44716
rect 31448 44662 31476 44714
rect 31572 44662 31580 44714
rect 31428 44660 31476 44662
rect 31532 44660 31580 44662
rect 31636 44714 31684 44716
rect 31740 44714 31788 44716
rect 31636 44662 31644 44714
rect 31740 44662 31768 44714
rect 31636 44660 31684 44662
rect 31740 44660 31788 44662
rect 31844 44660 31892 44716
rect 31268 44650 31948 44660
rect 31052 44436 31108 44446
rect 31052 44342 31108 44380
rect 31948 43764 32004 43774
rect 31724 43650 31780 43662
rect 31724 43598 31726 43650
rect 31778 43598 31780 43650
rect 31276 43428 31332 43438
rect 30604 43426 31332 43428
rect 30604 43374 31278 43426
rect 31330 43374 31332 43426
rect 30604 43372 31332 43374
rect 29596 43316 29652 43326
rect 29596 43222 29652 43260
rect 28588 42802 28644 42812
rect 29372 42868 29428 42878
rect 29372 42774 29428 42812
rect 28364 41916 28644 41972
rect 28252 40574 28254 40626
rect 28306 40574 28308 40626
rect 25452 40350 25454 40402
rect 25506 40350 25508 40402
rect 25452 40338 25508 40350
rect 25900 40404 25956 40414
rect 25900 40402 26628 40404
rect 25900 40350 25902 40402
rect 25954 40350 26628 40402
rect 25900 40348 26628 40350
rect 25900 40338 25956 40348
rect 22268 40012 22948 40022
rect 22324 39956 22372 40012
rect 22428 40010 22476 40012
rect 22532 40010 22580 40012
rect 22448 39958 22476 40010
rect 22572 39958 22580 40010
rect 22428 39956 22476 39958
rect 22532 39956 22580 39958
rect 22636 40010 22684 40012
rect 22740 40010 22788 40012
rect 22636 39958 22644 40010
rect 22740 39958 22768 40010
rect 22636 39956 22684 39958
rect 22740 39956 22788 39958
rect 22844 39956 22892 40012
rect 22268 39946 22948 39956
rect 26572 39506 26628 40348
rect 28252 40292 28308 40574
rect 28252 40226 28308 40236
rect 26796 40180 26852 40190
rect 26796 39618 26852 40124
rect 26796 39566 26798 39618
rect 26850 39566 26852 39618
rect 26796 39554 26852 39566
rect 26572 39454 26574 39506
rect 26626 39454 26628 39506
rect 26572 39442 26628 39454
rect 26768 39228 27448 39238
rect 26824 39172 26872 39228
rect 26928 39226 26976 39228
rect 27032 39226 27080 39228
rect 26948 39174 26976 39226
rect 27072 39174 27080 39226
rect 26928 39172 26976 39174
rect 27032 39172 27080 39174
rect 27136 39226 27184 39228
rect 27240 39226 27288 39228
rect 27136 39174 27144 39226
rect 27240 39174 27268 39226
rect 27136 39172 27184 39174
rect 27240 39172 27288 39174
rect 27344 39172 27392 39228
rect 26768 39162 27448 39172
rect 21084 39006 21086 39058
rect 21138 39006 21140 39058
rect 17052 38612 17332 38668
rect 17500 38612 17668 38668
rect 16828 38444 16996 38500
rect 15596 37268 15652 37278
rect 15596 37266 16548 37268
rect 15596 37214 15598 37266
rect 15650 37214 16548 37266
rect 15596 37212 16548 37214
rect 15596 37202 15652 37212
rect 15484 35758 15486 35810
rect 15538 35758 15540 35810
rect 15484 35746 15540 35758
rect 16156 36372 16212 36382
rect 15372 35700 15428 35710
rect 14924 35588 14980 35598
rect 15372 35588 15428 35644
rect 16156 35698 16212 36316
rect 16492 35922 16548 37212
rect 16828 36932 16884 38444
rect 17276 38276 17332 38612
rect 17276 38210 17332 38220
rect 16492 35870 16494 35922
rect 16546 35870 16548 35922
rect 16492 35858 16548 35870
rect 16716 36876 16884 36932
rect 16156 35646 16158 35698
rect 16210 35646 16212 35698
rect 16156 35634 16212 35646
rect 16716 35700 16772 36876
rect 17612 36708 17668 38612
rect 20524 38050 20580 38062
rect 20524 37998 20526 38050
rect 20578 37998 20580 38050
rect 20188 37828 20244 37838
rect 17768 37660 18448 37670
rect 17824 37604 17872 37660
rect 17928 37658 17976 37660
rect 18032 37658 18080 37660
rect 17948 37606 17976 37658
rect 18072 37606 18080 37658
rect 17928 37604 17976 37606
rect 18032 37604 18080 37606
rect 18136 37658 18184 37660
rect 18240 37658 18288 37660
rect 18136 37606 18144 37658
rect 18240 37606 18268 37658
rect 18136 37604 18184 37606
rect 18240 37604 18288 37606
rect 18344 37604 18392 37660
rect 17768 37594 18448 37604
rect 18396 37492 18452 37502
rect 18396 37398 18452 37436
rect 19740 37492 19796 37502
rect 19628 37154 19684 37166
rect 19628 37102 19630 37154
rect 19682 37102 19684 37154
rect 19628 36932 19684 37102
rect 17500 36372 17556 36382
rect 17612 36372 17668 36652
rect 18620 36708 18676 36718
rect 17724 36372 17780 36382
rect 17612 36370 17780 36372
rect 17612 36318 17726 36370
rect 17778 36318 17780 36370
rect 17612 36316 17780 36318
rect 17500 35922 17556 36316
rect 17724 36306 17780 36316
rect 18508 36372 18564 36382
rect 18508 36278 18564 36316
rect 17768 36092 18448 36102
rect 17824 36036 17872 36092
rect 17928 36090 17976 36092
rect 18032 36090 18080 36092
rect 17948 36038 17976 36090
rect 18072 36038 18080 36090
rect 17928 36036 17976 36038
rect 18032 36036 18080 36038
rect 18136 36090 18184 36092
rect 18240 36090 18288 36092
rect 18136 36038 18144 36090
rect 18240 36038 18268 36090
rect 18136 36036 18184 36038
rect 18240 36036 18288 36038
rect 18344 36036 18392 36092
rect 17768 36026 18448 36036
rect 17500 35870 17502 35922
rect 17554 35870 17556 35922
rect 17500 35858 17556 35870
rect 18620 35922 18676 36652
rect 18956 36708 19012 36718
rect 18956 36614 19012 36652
rect 18620 35870 18622 35922
rect 18674 35870 18676 35922
rect 18620 35858 18676 35870
rect 19628 35924 19684 36876
rect 19740 36482 19796 37436
rect 20188 37492 20244 37772
rect 20524 37716 20580 37998
rect 20748 38052 20804 38062
rect 20748 37938 20804 37996
rect 20748 37886 20750 37938
rect 20802 37886 20804 37938
rect 20748 37874 20804 37886
rect 20524 37650 20580 37660
rect 20188 37490 20692 37492
rect 20188 37438 20190 37490
rect 20242 37438 20692 37490
rect 20188 37436 20692 37438
rect 20188 37426 20244 37436
rect 20636 37378 20692 37436
rect 20636 37326 20638 37378
rect 20690 37326 20692 37378
rect 20636 37314 20692 37326
rect 20524 37266 20580 37278
rect 20524 37214 20526 37266
rect 20578 37214 20580 37266
rect 20524 36932 20580 37214
rect 20524 36866 20580 36876
rect 20748 37044 20804 37054
rect 19740 36430 19742 36482
rect 19794 36430 19796 36482
rect 19740 36418 19796 36430
rect 20748 36708 20804 36988
rect 21084 37044 21140 39006
rect 21644 38946 21700 38958
rect 21644 38894 21646 38946
rect 21698 38894 21700 38946
rect 21532 38052 21588 38062
rect 21644 38052 21700 38894
rect 28588 38668 28644 41916
rect 30380 40852 30436 40862
rect 30156 40516 30212 40526
rect 28924 40404 28980 40414
rect 28924 40310 28980 40348
rect 29596 40404 29652 40414
rect 29596 40310 29652 40348
rect 30156 40402 30212 40460
rect 30380 40514 30436 40796
rect 30380 40462 30382 40514
rect 30434 40462 30436 40514
rect 30380 40450 30436 40462
rect 30604 40516 30660 43372
rect 31276 43362 31332 43372
rect 31724 43316 31780 43598
rect 31948 43428 32004 43708
rect 31948 43362 32004 43372
rect 32060 43652 32116 43662
rect 31724 43250 31780 43260
rect 31268 43148 31948 43158
rect 31324 43092 31372 43148
rect 31428 43146 31476 43148
rect 31532 43146 31580 43148
rect 31448 43094 31476 43146
rect 31572 43094 31580 43146
rect 31428 43092 31476 43094
rect 31532 43092 31580 43094
rect 31636 43146 31684 43148
rect 31740 43146 31788 43148
rect 31636 43094 31644 43146
rect 31740 43094 31768 43146
rect 31636 43092 31684 43094
rect 31740 43092 31788 43094
rect 31844 43092 31892 43148
rect 31268 43082 31948 43092
rect 31612 42980 31668 42990
rect 30604 40450 30660 40460
rect 30828 42868 30884 42878
rect 30156 40350 30158 40402
rect 30210 40350 30212 40402
rect 29036 40292 29092 40302
rect 29092 40236 29204 40292
rect 29036 40226 29092 40236
rect 29148 39732 29204 40236
rect 29260 40180 29316 40190
rect 29260 40086 29316 40124
rect 29260 39732 29316 39742
rect 29148 39730 29316 39732
rect 29148 39678 29262 39730
rect 29314 39678 29316 39730
rect 29148 39676 29316 39678
rect 28812 38722 28868 38734
rect 28812 38670 28814 38722
rect 28866 38670 28868 38722
rect 28812 38668 28868 38670
rect 28476 38612 28868 38668
rect 22268 38444 22948 38454
rect 22324 38388 22372 38444
rect 22428 38442 22476 38444
rect 22532 38442 22580 38444
rect 22448 38390 22476 38442
rect 22572 38390 22580 38442
rect 22428 38388 22476 38390
rect 22532 38388 22580 38390
rect 22636 38442 22684 38444
rect 22740 38442 22788 38444
rect 22636 38390 22644 38442
rect 22740 38390 22768 38442
rect 22636 38388 22684 38390
rect 22740 38388 22788 38390
rect 22844 38388 22892 38444
rect 22268 38378 22948 38388
rect 21532 38050 21700 38052
rect 21532 37998 21534 38050
rect 21586 37998 21700 38050
rect 21532 37996 21700 37998
rect 21868 38052 21924 38062
rect 21532 37986 21588 37996
rect 21868 37958 21924 37996
rect 27692 38050 27748 38062
rect 27692 37998 27694 38050
rect 27746 37998 27748 38050
rect 24220 37826 24276 37838
rect 24220 37774 24222 37826
rect 24274 37774 24276 37826
rect 21644 37716 21700 37726
rect 21644 37490 21700 37660
rect 21644 37438 21646 37490
rect 21698 37438 21700 37490
rect 21644 37426 21700 37438
rect 21308 37268 21364 37278
rect 21308 37174 21364 37212
rect 21084 36978 21140 36988
rect 24220 37044 24276 37774
rect 25004 37828 25060 37838
rect 25004 37268 25060 37772
rect 26348 37826 26404 37838
rect 26348 37774 26350 37826
rect 26402 37774 26404 37826
rect 25004 37202 25060 37212
rect 26236 37268 26292 37278
rect 26348 37268 26404 37774
rect 27356 37828 27412 37838
rect 27356 37826 27636 37828
rect 27356 37774 27358 37826
rect 27410 37774 27636 37826
rect 27356 37772 27636 37774
rect 27356 37762 27412 37772
rect 26768 37660 27448 37670
rect 26824 37604 26872 37660
rect 26928 37658 26976 37660
rect 27032 37658 27080 37660
rect 26948 37606 26976 37658
rect 27072 37606 27080 37658
rect 26928 37604 26976 37606
rect 27032 37604 27080 37606
rect 27136 37658 27184 37660
rect 27240 37658 27288 37660
rect 27136 37606 27144 37658
rect 27240 37606 27268 37658
rect 27136 37604 27184 37606
rect 27240 37604 27288 37606
rect 27344 37604 27392 37660
rect 26768 37594 27448 37604
rect 26236 37266 26404 37268
rect 26236 37214 26238 37266
rect 26290 37214 26404 37266
rect 26236 37212 26404 37214
rect 26684 37268 26740 37278
rect 26684 37266 27188 37268
rect 26684 37214 26686 37266
rect 26738 37214 27188 37266
rect 26684 37212 27188 37214
rect 26236 37202 26292 37212
rect 26684 37202 26740 37212
rect 22268 36876 22948 36886
rect 22324 36820 22372 36876
rect 22428 36874 22476 36876
rect 22532 36874 22580 36876
rect 22448 36822 22476 36874
rect 22572 36822 22580 36874
rect 22428 36820 22476 36822
rect 22532 36820 22580 36822
rect 22636 36874 22684 36876
rect 22740 36874 22788 36876
rect 22636 36822 22644 36874
rect 22740 36822 22768 36874
rect 22636 36820 22684 36822
rect 22740 36820 22788 36822
rect 22844 36820 22892 36876
rect 22268 36810 22948 36820
rect 19740 35924 19796 35934
rect 19628 35922 20132 35924
rect 19628 35870 19742 35922
rect 19794 35870 20132 35922
rect 19628 35868 20132 35870
rect 16716 35634 16772 35644
rect 14924 35586 15428 35588
rect 14924 35534 14926 35586
rect 14978 35534 15428 35586
rect 14924 35532 15428 35534
rect 14924 35476 14980 35532
rect 14700 35420 14980 35476
rect 13268 35308 13948 35318
rect 13324 35252 13372 35308
rect 13428 35306 13476 35308
rect 13532 35306 13580 35308
rect 13448 35254 13476 35306
rect 13572 35254 13580 35306
rect 13428 35252 13476 35254
rect 13532 35252 13580 35254
rect 13636 35306 13684 35308
rect 13740 35306 13788 35308
rect 13636 35254 13644 35306
rect 13740 35254 13768 35306
rect 13636 35252 13684 35254
rect 13740 35252 13788 35254
rect 13844 35252 13892 35308
rect 13268 35242 13948 35252
rect 11788 34078 11790 34130
rect 11842 34078 11844 34130
rect 11788 34066 11844 34078
rect 12012 34244 12068 34254
rect 12012 33684 12068 34188
rect 14028 34244 14084 34254
rect 14028 34150 14084 34188
rect 13244 34132 13300 34142
rect 12012 29988 12068 33628
rect 13132 34076 13244 34132
rect 13132 32786 13188 34076
rect 13244 34066 13300 34076
rect 13268 33740 13948 33750
rect 13324 33684 13372 33740
rect 13428 33738 13476 33740
rect 13532 33738 13580 33740
rect 13448 33686 13476 33738
rect 13572 33686 13580 33738
rect 13428 33684 13476 33686
rect 13532 33684 13580 33686
rect 13636 33738 13684 33740
rect 13740 33738 13788 33740
rect 13636 33686 13644 33738
rect 13740 33686 13768 33738
rect 13636 33684 13684 33686
rect 13740 33684 13788 33686
rect 13844 33684 13892 33740
rect 13268 33674 13948 33684
rect 14588 33460 14644 33470
rect 14700 33460 14756 35420
rect 17768 34524 18448 34534
rect 17824 34468 17872 34524
rect 17928 34522 17976 34524
rect 18032 34522 18080 34524
rect 17948 34470 17976 34522
rect 18072 34470 18080 34522
rect 17928 34468 17976 34470
rect 18032 34468 18080 34470
rect 18136 34522 18184 34524
rect 18240 34522 18288 34524
rect 18136 34470 18144 34522
rect 18240 34470 18268 34522
rect 18136 34468 18184 34470
rect 18240 34468 18288 34470
rect 18344 34468 18392 34524
rect 17768 34458 18448 34468
rect 19516 34020 19572 34030
rect 14812 33908 14868 33918
rect 14812 33906 15204 33908
rect 14812 33854 14814 33906
rect 14866 33854 15204 33906
rect 14812 33852 15204 33854
rect 14812 33842 14868 33852
rect 14644 33404 15092 33460
rect 14588 33366 14644 33404
rect 15036 33346 15092 33404
rect 15036 33294 15038 33346
rect 15090 33294 15092 33346
rect 15036 33282 15092 33294
rect 15148 33234 15204 33852
rect 19068 33460 19124 33470
rect 19068 33366 19124 33404
rect 15148 33182 15150 33234
rect 15202 33182 15204 33234
rect 15148 33170 15204 33182
rect 15372 33348 15428 33358
rect 13132 32734 13134 32786
rect 13186 32734 13188 32786
rect 13132 32722 13188 32734
rect 12348 32676 12404 32686
rect 12348 32582 12404 32620
rect 14812 32674 14868 32686
rect 14812 32622 14814 32674
rect 14866 32622 14868 32674
rect 14588 32340 14644 32350
rect 13268 32172 13948 32182
rect 13324 32116 13372 32172
rect 13428 32170 13476 32172
rect 13532 32170 13580 32172
rect 13448 32118 13476 32170
rect 13572 32118 13580 32170
rect 13428 32116 13476 32118
rect 13532 32116 13580 32118
rect 13636 32170 13684 32172
rect 13740 32170 13788 32172
rect 13636 32118 13644 32170
rect 13740 32118 13768 32170
rect 13636 32116 13684 32118
rect 13740 32116 13788 32118
rect 13844 32116 13892 32172
rect 13268 32106 13948 32116
rect 14588 31778 14644 32284
rect 14812 31948 14868 32622
rect 15148 32676 15204 32686
rect 15148 32582 15204 32620
rect 14812 31892 14980 31948
rect 14588 31726 14590 31778
rect 14642 31726 14644 31778
rect 14588 31714 14644 31726
rect 14924 31778 14980 31892
rect 14924 31726 14926 31778
rect 14978 31726 14980 31778
rect 14924 31714 14980 31726
rect 14700 30884 14756 30894
rect 14700 30882 14868 30884
rect 14700 30830 14702 30882
rect 14754 30830 14868 30882
rect 14700 30828 14868 30830
rect 14700 30818 14756 30828
rect 13268 30604 13948 30614
rect 13324 30548 13372 30604
rect 13428 30602 13476 30604
rect 13532 30602 13580 30604
rect 13448 30550 13476 30602
rect 13572 30550 13580 30602
rect 13428 30548 13476 30550
rect 13532 30548 13580 30550
rect 13636 30602 13684 30604
rect 13740 30602 13788 30604
rect 13636 30550 13644 30602
rect 13740 30550 13768 30602
rect 13636 30548 13684 30550
rect 13740 30548 13788 30550
rect 13844 30548 13892 30604
rect 13268 30538 13948 30548
rect 14812 30212 14868 30828
rect 15148 30212 15204 30222
rect 14812 30210 15204 30212
rect 14812 30158 15150 30210
rect 15202 30158 15204 30210
rect 14812 30156 15204 30158
rect 14700 30100 14756 30110
rect 14700 30006 14756 30044
rect 12012 29894 12068 29932
rect 12572 29986 12628 29998
rect 13916 29988 13972 29998
rect 14364 29988 14420 29998
rect 12572 29934 12574 29986
rect 12626 29934 12628 29986
rect 12460 27972 12516 27982
rect 12572 27972 12628 29934
rect 13468 29986 13972 29988
rect 13468 29934 13918 29986
rect 13970 29934 13972 29986
rect 13468 29932 13972 29934
rect 13468 29426 13524 29932
rect 13916 29922 13972 29932
rect 14028 29986 14420 29988
rect 14028 29934 14366 29986
rect 14418 29934 14420 29986
rect 14028 29932 14420 29934
rect 13468 29374 13470 29426
rect 13522 29374 13524 29426
rect 13468 29362 13524 29374
rect 13916 29428 13972 29438
rect 14028 29428 14084 29932
rect 14364 29922 14420 29932
rect 13916 29426 14084 29428
rect 13916 29374 13918 29426
rect 13970 29374 14084 29426
rect 13916 29372 14084 29374
rect 13916 29362 13972 29372
rect 13020 29316 13076 29326
rect 13020 29222 13076 29260
rect 13268 29036 13948 29046
rect 13324 28980 13372 29036
rect 13428 29034 13476 29036
rect 13532 29034 13580 29036
rect 13448 28982 13476 29034
rect 13572 28982 13580 29034
rect 13428 28980 13476 28982
rect 13532 28980 13580 28982
rect 13636 29034 13684 29036
rect 13740 29034 13788 29036
rect 13636 28982 13644 29034
rect 13740 28982 13768 29034
rect 13636 28980 13684 28982
rect 13740 28980 13788 28982
rect 13844 28980 13892 29036
rect 13268 28970 13948 28980
rect 13804 28642 13860 28654
rect 13804 28590 13806 28642
rect 13858 28590 13860 28642
rect 12460 27970 12628 27972
rect 12460 27918 12462 27970
rect 12514 27918 12628 27970
rect 12460 27916 12628 27918
rect 13020 28084 13076 28094
rect 12460 27906 12516 27916
rect 12236 27860 12292 27870
rect 11788 27748 11844 27758
rect 12236 27748 12292 27804
rect 13020 27858 13076 28028
rect 13804 28084 13860 28590
rect 13804 28018 13860 28028
rect 14028 28140 14308 28196
rect 13020 27806 13022 27858
rect 13074 27806 13076 27858
rect 13020 27794 13076 27806
rect 13356 27860 13412 27870
rect 13804 27860 13860 27870
rect 13356 27858 13860 27860
rect 13356 27806 13358 27858
rect 13410 27806 13806 27858
rect 13858 27806 13860 27858
rect 13356 27804 13860 27806
rect 13356 27794 13412 27804
rect 13804 27794 13860 27804
rect 11788 27746 12292 27748
rect 11788 27694 11790 27746
rect 11842 27694 12292 27746
rect 11788 27692 12292 27694
rect 11788 27636 11844 27692
rect 11228 27580 11844 27636
rect 10780 26850 10836 26862
rect 10780 26798 10782 26850
rect 10834 26798 10836 26850
rect 10332 24894 10334 24946
rect 10386 24894 10388 24946
rect 10332 24882 10388 24894
rect 10556 25394 10612 25406
rect 10556 25342 10558 25394
rect 10610 25342 10612 25394
rect 10556 24948 10612 25342
rect 10556 24882 10612 24892
rect 10780 24164 10836 26798
rect 10780 24098 10836 24108
rect 10892 26178 10948 26190
rect 10892 26126 10894 26178
rect 10946 26126 10948 26178
rect 10892 24834 10948 26126
rect 11116 25396 11172 25406
rect 11116 25302 11172 25340
rect 10892 24782 10894 24834
rect 10946 24782 10948 24834
rect 10892 23938 10948 24782
rect 11228 24050 11284 27580
rect 13268 27468 13948 27478
rect 13324 27412 13372 27468
rect 13428 27466 13476 27468
rect 13532 27466 13580 27468
rect 13448 27414 13476 27466
rect 13572 27414 13580 27466
rect 13428 27412 13476 27414
rect 13532 27412 13580 27414
rect 13636 27466 13684 27468
rect 13740 27466 13788 27468
rect 13636 27414 13644 27466
rect 13740 27414 13768 27466
rect 13636 27412 13684 27414
rect 13740 27412 13788 27414
rect 13844 27412 13892 27468
rect 13268 27402 13948 27412
rect 13916 27076 13972 27086
rect 14028 27076 14084 28140
rect 14252 28084 14308 28140
rect 14476 28084 14532 28094
rect 14252 28082 14532 28084
rect 14252 28030 14478 28082
rect 14530 28030 14532 28082
rect 14252 28028 14532 28030
rect 14476 28018 14532 28028
rect 13916 27074 14084 27076
rect 13916 27022 13918 27074
rect 13970 27022 14084 27074
rect 13916 27020 14084 27022
rect 14140 27970 14196 27982
rect 14140 27918 14142 27970
rect 14194 27918 14196 27970
rect 14140 27076 14196 27918
rect 15148 27860 15204 30156
rect 15372 30098 15428 33292
rect 15820 33348 15876 33358
rect 16716 33348 16772 33358
rect 15820 33346 16772 33348
rect 15820 33294 15822 33346
rect 15874 33294 16718 33346
rect 16770 33294 16772 33346
rect 15820 33292 16772 33294
rect 15820 33282 15876 33292
rect 16156 33122 16212 33134
rect 16156 33070 16158 33122
rect 16210 33070 16212 33122
rect 15484 32674 15540 32686
rect 15484 32622 15486 32674
rect 15538 32622 15540 32674
rect 15484 32340 15540 32622
rect 16156 32676 16212 33070
rect 16156 32610 16212 32620
rect 15484 32274 15540 32284
rect 16716 31668 16772 33292
rect 19516 33234 19572 33964
rect 19628 33460 19684 35868
rect 19740 35858 19796 35868
rect 20076 35588 20132 35868
rect 20300 35812 20356 35822
rect 20300 35718 20356 35756
rect 20188 35698 20244 35710
rect 20188 35646 20190 35698
rect 20242 35646 20244 35698
rect 20188 35588 20244 35646
rect 20076 35532 20244 35588
rect 20748 35026 20804 36652
rect 21308 36260 21364 36270
rect 21196 36258 21364 36260
rect 21196 36206 21310 36258
rect 21362 36206 21364 36258
rect 21196 36204 21364 36206
rect 20748 34974 20750 35026
rect 20802 34974 20804 35026
rect 20748 34962 20804 34974
rect 20972 35474 21028 35486
rect 20972 35422 20974 35474
rect 21026 35422 21028 35474
rect 20972 34804 21028 35422
rect 21196 34914 21252 36204
rect 21308 36194 21364 36204
rect 22092 35812 22148 35822
rect 21868 35810 22148 35812
rect 21868 35758 22094 35810
rect 22146 35758 22148 35810
rect 21868 35756 22148 35758
rect 21308 35700 21364 35710
rect 21756 35700 21812 35710
rect 21308 35698 21812 35700
rect 21308 35646 21310 35698
rect 21362 35646 21758 35698
rect 21810 35646 21812 35698
rect 21308 35644 21812 35646
rect 21308 35634 21364 35644
rect 21756 35634 21812 35644
rect 21196 34862 21198 34914
rect 21250 34862 21252 34914
rect 21196 34850 21252 34862
rect 21868 34914 21924 35756
rect 22092 35746 22148 35756
rect 22268 35308 22948 35318
rect 22324 35252 22372 35308
rect 22428 35306 22476 35308
rect 22532 35306 22580 35308
rect 22448 35254 22476 35306
rect 22572 35254 22580 35306
rect 22428 35252 22476 35254
rect 22532 35252 22580 35254
rect 22636 35306 22684 35308
rect 22740 35306 22788 35308
rect 22636 35254 22644 35306
rect 22740 35254 22768 35306
rect 22636 35252 22684 35254
rect 22740 35252 22788 35254
rect 22844 35252 22892 35308
rect 22268 35242 22948 35252
rect 21868 34862 21870 34914
rect 21922 34862 21924 34914
rect 21868 34850 21924 34862
rect 20972 34738 21028 34748
rect 24220 34690 24276 36988
rect 27132 36370 27188 37212
rect 27468 36484 27524 36494
rect 27580 36484 27636 37772
rect 27692 37268 27748 37998
rect 28364 38052 28420 38062
rect 28364 37958 28420 37996
rect 28476 37940 28532 38612
rect 28476 37846 28532 37884
rect 29148 37490 29204 39676
rect 29260 39666 29316 39676
rect 29932 38164 29988 38174
rect 29596 37826 29652 37838
rect 29596 37774 29598 37826
rect 29650 37774 29652 37826
rect 29596 37604 29652 37774
rect 29932 37604 29988 38108
rect 30156 38052 30212 40350
rect 30828 39732 30884 42812
rect 31164 42868 31220 42878
rect 31164 42774 31220 42812
rect 31612 42754 31668 42924
rect 31612 42702 31614 42754
rect 31666 42702 31668 42754
rect 31612 42690 31668 42702
rect 32060 42754 32116 43596
rect 32060 42702 32062 42754
rect 32114 42702 32116 42754
rect 32060 42690 32116 42702
rect 31268 41580 31948 41590
rect 31324 41524 31372 41580
rect 31428 41578 31476 41580
rect 31532 41578 31580 41580
rect 31448 41526 31476 41578
rect 31572 41526 31580 41578
rect 31428 41524 31476 41526
rect 31532 41524 31580 41526
rect 31636 41578 31684 41580
rect 31740 41578 31788 41580
rect 31636 41526 31644 41578
rect 31740 41526 31768 41578
rect 31636 41524 31684 41526
rect 31740 41524 31788 41526
rect 31844 41524 31892 41580
rect 31268 41514 31948 41524
rect 31500 40964 31556 40974
rect 31052 40962 31556 40964
rect 31052 40910 31502 40962
rect 31554 40910 31556 40962
rect 31052 40908 31556 40910
rect 30940 40516 30996 40526
rect 30940 40422 30996 40460
rect 30940 39732 30996 39742
rect 30828 39730 30996 39732
rect 30828 39678 30942 39730
rect 30994 39678 30996 39730
rect 30828 39676 30996 39678
rect 30940 39666 30996 39676
rect 31052 39620 31108 40908
rect 31500 40898 31556 40908
rect 31612 40852 31668 40862
rect 31388 40628 31444 40638
rect 31612 40628 31668 40796
rect 32172 40852 32228 45836
rect 33740 45780 33796 50428
rect 35768 50204 36448 50214
rect 35824 50148 35872 50204
rect 35928 50202 35976 50204
rect 36032 50202 36080 50204
rect 35948 50150 35976 50202
rect 36072 50150 36080 50202
rect 35928 50148 35976 50150
rect 36032 50148 36080 50150
rect 36136 50202 36184 50204
rect 36240 50202 36288 50204
rect 36136 50150 36144 50202
rect 36240 50150 36268 50202
rect 36136 50148 36184 50150
rect 36240 50148 36288 50150
rect 36344 50148 36392 50204
rect 35768 50138 36448 50148
rect 37660 49924 37716 49934
rect 37660 49830 37716 49868
rect 38444 49812 38500 49822
rect 38444 49718 38500 49756
rect 35532 49698 35588 49710
rect 35532 49646 35534 49698
rect 35586 49646 35588 49698
rect 35532 49588 35588 49646
rect 39004 49700 39060 49710
rect 39004 49606 39060 49644
rect 35588 49532 35700 49588
rect 35532 49522 35588 49532
rect 35084 49252 35140 49262
rect 35084 49138 35140 49196
rect 35084 49086 35086 49138
rect 35138 49086 35140 49138
rect 34748 47572 34804 47582
rect 33964 47458 34020 47470
rect 33964 47406 33966 47458
rect 34018 47406 34020 47458
rect 33964 46676 34020 47406
rect 34636 47458 34692 47470
rect 34636 47406 34638 47458
rect 34690 47406 34692 47458
rect 34636 47348 34692 47406
rect 34636 47282 34692 47292
rect 34748 47346 34804 47516
rect 34748 47294 34750 47346
rect 34802 47294 34804 47346
rect 34748 47282 34804 47294
rect 33964 46610 34020 46620
rect 34524 46676 34580 46686
rect 34524 46114 34580 46620
rect 34524 46062 34526 46114
rect 34578 46062 34580 46114
rect 34524 46050 34580 46062
rect 34748 46674 34804 46686
rect 34748 46622 34750 46674
rect 34802 46622 34804 46674
rect 33796 45724 34356 45780
rect 33740 45686 33796 45724
rect 34188 44322 34244 44334
rect 34188 44270 34190 44322
rect 34242 44270 34244 44322
rect 33852 44100 33908 44110
rect 33404 44098 33908 44100
rect 33404 44046 33854 44098
rect 33906 44046 33908 44098
rect 33404 44044 33908 44046
rect 33068 43652 33124 43662
rect 33068 43558 33124 43596
rect 33404 43650 33460 44044
rect 33852 44034 33908 44044
rect 33404 43598 33406 43650
rect 33458 43598 33460 43650
rect 33404 43586 33460 43598
rect 33740 43876 33796 43886
rect 32508 43428 32564 43438
rect 32508 43334 32564 43372
rect 33740 41298 33796 43820
rect 34188 42980 34244 44270
rect 34188 42914 34244 42924
rect 33740 41246 33742 41298
rect 33794 41246 33796 41298
rect 32172 40786 32228 40796
rect 33292 40962 33348 40974
rect 33292 40910 33294 40962
rect 33346 40910 33348 40962
rect 33292 40852 33348 40910
rect 33292 40786 33348 40796
rect 33404 40964 33460 40974
rect 31388 40626 31668 40628
rect 31388 40574 31390 40626
rect 31442 40574 31668 40626
rect 31388 40572 31668 40574
rect 31388 40562 31444 40572
rect 33068 40514 33124 40526
rect 33068 40462 33070 40514
rect 33122 40462 33124 40514
rect 31268 40012 31948 40022
rect 31324 39956 31372 40012
rect 31428 40010 31476 40012
rect 31532 40010 31580 40012
rect 31448 39958 31476 40010
rect 31572 39958 31580 40010
rect 31428 39956 31476 39958
rect 31532 39956 31580 39958
rect 31636 40010 31684 40012
rect 31740 40010 31788 40012
rect 31636 39958 31644 40010
rect 31740 39958 31768 40010
rect 31636 39956 31684 39958
rect 31740 39956 31788 39958
rect 31844 39956 31892 40012
rect 31268 39946 31948 39956
rect 31836 39844 31892 39854
rect 31164 39620 31220 39630
rect 31052 39618 31220 39620
rect 31052 39566 31166 39618
rect 31218 39566 31220 39618
rect 31052 39564 31220 39566
rect 31164 39554 31220 39564
rect 31836 39618 31892 39788
rect 33068 39844 33124 40462
rect 33404 40514 33460 40908
rect 33740 40628 33796 41246
rect 34300 42642 34356 45724
rect 34748 43540 34804 46622
rect 34972 46674 35028 46686
rect 34972 46622 34974 46674
rect 35026 46622 35028 46674
rect 34972 46564 35028 46622
rect 34972 46498 35028 46508
rect 35084 45780 35140 49086
rect 35644 47572 35700 49532
rect 35756 49140 35812 49150
rect 35756 49046 35812 49084
rect 38668 49140 38724 49150
rect 35768 48636 36448 48646
rect 35824 48580 35872 48636
rect 35928 48634 35976 48636
rect 36032 48634 36080 48636
rect 35948 48582 35976 48634
rect 36072 48582 36080 48634
rect 35928 48580 35976 48582
rect 36032 48580 36080 48582
rect 36136 48634 36184 48636
rect 36240 48634 36288 48636
rect 36136 48582 36144 48634
rect 36240 48582 36268 48634
rect 36136 48580 36184 48582
rect 36240 48580 36288 48582
rect 36344 48580 36392 48636
rect 35768 48570 36448 48580
rect 36764 48244 36820 48254
rect 36428 48242 36820 48244
rect 36428 48190 36766 48242
rect 36818 48190 36820 48242
rect 36428 48188 36820 48190
rect 35756 47572 35812 47582
rect 35700 47570 35812 47572
rect 35700 47518 35758 47570
rect 35810 47518 35812 47570
rect 35700 47516 35812 47518
rect 35644 47478 35700 47516
rect 35756 47506 35812 47516
rect 35084 44436 35140 45724
rect 34860 44322 34916 44334
rect 34860 44270 34862 44322
rect 34914 44270 34916 44322
rect 34860 44212 34916 44270
rect 34860 44146 34916 44156
rect 34972 44212 35028 44222
rect 35084 44212 35140 44380
rect 34972 44210 35140 44212
rect 34972 44158 34974 44210
rect 35026 44158 35140 44210
rect 34972 44156 35140 44158
rect 35308 47348 35364 47358
rect 35308 47234 35364 47292
rect 36428 47346 36484 48188
rect 36764 48178 36820 48188
rect 37324 48242 37380 48254
rect 37324 48190 37326 48242
rect 37378 48190 37380 48242
rect 36428 47294 36430 47346
rect 36482 47294 36484 47346
rect 36428 47282 36484 47294
rect 37324 47346 37380 48190
rect 38668 47570 38724 49084
rect 39900 49140 39956 50540
rect 40012 50428 40068 51212
rect 40124 50820 40180 51548
rect 40908 51492 40964 51502
rect 40908 51398 40964 51436
rect 41020 51490 41076 51502
rect 41020 51438 41022 51490
rect 41074 51438 41076 51490
rect 40348 51268 40404 51278
rect 41020 51268 41076 51438
rect 40348 51266 41076 51268
rect 40348 51214 40350 51266
rect 40402 51214 41076 51266
rect 40348 51212 41076 51214
rect 40348 51202 40404 51212
rect 40268 50988 40948 50998
rect 40324 50932 40372 50988
rect 40428 50986 40476 50988
rect 40532 50986 40580 50988
rect 40448 50934 40476 50986
rect 40572 50934 40580 50986
rect 40428 50932 40476 50934
rect 40532 50932 40580 50934
rect 40636 50986 40684 50988
rect 40740 50986 40788 50988
rect 40636 50934 40644 50986
rect 40740 50934 40768 50986
rect 40636 50932 40684 50934
rect 40740 50932 40788 50934
rect 40844 50932 40892 50988
rect 40268 50922 40948 50932
rect 41020 50820 41076 51212
rect 40124 50764 40404 50820
rect 40012 50372 40180 50428
rect 39900 49074 39956 49084
rect 39900 48468 39956 48478
rect 39900 48374 39956 48412
rect 38668 47518 38670 47570
rect 38722 47518 38724 47570
rect 38668 47506 38724 47518
rect 40012 48020 40068 48030
rect 37324 47294 37326 47346
rect 37378 47294 37380 47346
rect 37324 47282 37380 47294
rect 37660 47348 37716 47358
rect 37660 47254 37716 47292
rect 39116 47348 39172 47358
rect 35308 47182 35310 47234
rect 35362 47182 35364 47234
rect 35308 44212 35364 47182
rect 35768 47068 36448 47078
rect 35824 47012 35872 47068
rect 35928 47066 35976 47068
rect 36032 47066 36080 47068
rect 35948 47014 35976 47066
rect 36072 47014 36080 47066
rect 35928 47012 35976 47014
rect 36032 47012 36080 47014
rect 36136 47066 36184 47068
rect 36240 47066 36288 47068
rect 36136 47014 36144 47066
rect 36240 47014 36268 47066
rect 36136 47012 36184 47014
rect 36240 47012 36288 47014
rect 36344 47012 36392 47068
rect 35768 47002 36448 47012
rect 38556 47012 38612 47022
rect 38556 46898 38612 46956
rect 38556 46846 38558 46898
rect 38610 46846 38612 46898
rect 38556 46834 38612 46846
rect 39116 46898 39172 47292
rect 39116 46846 39118 46898
rect 39170 46846 39172 46898
rect 39116 46834 39172 46846
rect 36764 46786 36820 46798
rect 36764 46734 36766 46786
rect 36818 46734 36820 46786
rect 35644 46676 35700 46686
rect 35644 46582 35700 46620
rect 36764 46116 36820 46734
rect 37884 46788 37940 46798
rect 38220 46788 38276 46798
rect 37884 46786 38052 46788
rect 37884 46734 37886 46786
rect 37938 46734 38052 46786
rect 37884 46732 38052 46734
rect 37884 46722 37940 46732
rect 36764 46050 36820 46060
rect 35768 45500 36448 45510
rect 35824 45444 35872 45500
rect 35928 45498 35976 45500
rect 36032 45498 36080 45500
rect 35948 45446 35976 45498
rect 36072 45446 36080 45498
rect 35928 45444 35976 45446
rect 36032 45444 36080 45446
rect 36136 45498 36184 45500
rect 36240 45498 36288 45500
rect 36136 45446 36144 45498
rect 36240 45446 36268 45498
rect 36136 45444 36184 45446
rect 36240 45444 36288 45446
rect 36344 45444 36392 45500
rect 35768 45434 36448 45444
rect 37436 45218 37492 45230
rect 37436 45166 37438 45218
rect 37490 45166 37492 45218
rect 35980 44436 36036 44446
rect 35980 44342 36036 44380
rect 37436 44324 37492 45166
rect 37996 45106 38052 46732
rect 38220 46674 38276 46732
rect 40012 46786 40068 47964
rect 40012 46734 40014 46786
rect 40066 46734 40068 46786
rect 40012 46722 40068 46734
rect 38220 46622 38222 46674
rect 38274 46622 38276 46674
rect 38220 46610 38276 46622
rect 39452 46452 39508 46462
rect 39340 46450 39508 46452
rect 39340 46398 39454 46450
rect 39506 46398 39508 46450
rect 39340 46396 39508 46398
rect 39004 46116 39060 46126
rect 38556 45780 38612 45790
rect 38556 45686 38612 45724
rect 37996 45054 37998 45106
rect 38050 45054 38052 45106
rect 37772 44324 37828 44334
rect 37436 44322 37828 44324
rect 37436 44270 37774 44322
rect 37826 44270 37828 44322
rect 37436 44268 37828 44270
rect 37772 44258 37828 44268
rect 35532 44212 35588 44222
rect 35308 44156 35532 44212
rect 34972 44146 35028 44156
rect 35532 44098 35588 44156
rect 35532 44046 35534 44098
rect 35586 44046 35588 44098
rect 35196 43540 35252 43550
rect 34748 43538 35028 43540
rect 34748 43486 34750 43538
rect 34802 43486 35028 43538
rect 34748 43484 35028 43486
rect 34748 43474 34804 43484
rect 34300 42590 34302 42642
rect 34354 42590 34356 42642
rect 34188 40964 34244 40974
rect 34188 40870 34244 40908
rect 33740 40562 33796 40572
rect 33404 40462 33406 40514
rect 33458 40462 33460 40514
rect 33404 40450 33460 40462
rect 33068 39778 33124 39788
rect 31836 39566 31838 39618
rect 31890 39566 31892 39618
rect 31836 39554 31892 39566
rect 34300 39394 34356 42590
rect 34524 41186 34580 41198
rect 34524 41134 34526 41186
rect 34578 41134 34580 41186
rect 34524 40516 34580 41134
rect 34972 40964 35028 43484
rect 35196 43446 35252 43484
rect 35084 42980 35140 42990
rect 35084 42886 35140 42924
rect 35308 41188 35364 41198
rect 35532 41188 35588 44046
rect 35768 43932 36448 43942
rect 35824 43876 35872 43932
rect 35928 43930 35976 43932
rect 36032 43930 36080 43932
rect 35948 43878 35976 43930
rect 36072 43878 36080 43930
rect 35928 43876 35976 43878
rect 36032 43876 36080 43878
rect 36136 43930 36184 43932
rect 36240 43930 36288 43932
rect 36136 43878 36144 43930
rect 36240 43878 36268 43930
rect 36136 43876 36184 43878
rect 36240 43876 36288 43878
rect 36344 43876 36392 43932
rect 35768 43866 36448 43876
rect 37996 43650 38052 45054
rect 38444 45668 38500 45678
rect 38444 44322 38500 45612
rect 39004 45666 39060 46060
rect 39340 45780 39396 46396
rect 39452 46386 39508 46396
rect 40012 46452 40068 46462
rect 39340 45714 39396 45724
rect 39004 45614 39006 45666
rect 39058 45614 39060 45666
rect 38444 44270 38446 44322
rect 38498 44270 38500 44322
rect 38444 44258 38500 44270
rect 38556 45444 38612 45454
rect 38556 43764 38612 45388
rect 38668 43764 38724 43774
rect 38556 43762 38724 43764
rect 38556 43710 38670 43762
rect 38722 43710 38724 43762
rect 38556 43708 38724 43710
rect 38668 43698 38724 43708
rect 37996 43598 37998 43650
rect 38050 43598 38052 43650
rect 35364 41132 35588 41188
rect 35644 43538 35700 43550
rect 35644 43486 35646 43538
rect 35698 43486 35700 43538
rect 34860 40516 34916 40526
rect 34524 40460 34860 40516
rect 34860 39842 34916 40460
rect 34972 40404 35028 40908
rect 35196 41074 35252 41086
rect 35196 41022 35198 41074
rect 35250 41022 35252 41074
rect 35196 40852 35252 41022
rect 34972 40402 35140 40404
rect 34972 40350 34974 40402
rect 35026 40350 35140 40402
rect 34972 40348 35140 40350
rect 34972 40338 35028 40348
rect 34860 39790 34862 39842
rect 34914 39790 34916 39842
rect 34860 39778 34916 39790
rect 34300 39342 34302 39394
rect 34354 39342 34356 39394
rect 34300 39330 34356 39342
rect 35084 38668 35140 40348
rect 35196 39060 35252 40796
rect 35196 38994 35252 39004
rect 34972 38612 35140 38668
rect 31268 38444 31948 38454
rect 31324 38388 31372 38444
rect 31428 38442 31476 38444
rect 31532 38442 31580 38444
rect 31448 38390 31476 38442
rect 31572 38390 31580 38442
rect 31428 38388 31476 38390
rect 31532 38388 31580 38390
rect 31636 38442 31684 38444
rect 31740 38442 31788 38444
rect 31636 38390 31644 38442
rect 31740 38390 31768 38442
rect 31636 38388 31684 38390
rect 31740 38388 31788 38390
rect 31844 38388 31892 38444
rect 31268 38378 31948 38388
rect 33404 38276 33460 38286
rect 33404 38162 33460 38220
rect 33404 38110 33406 38162
rect 33458 38110 33460 38162
rect 33404 38098 33460 38110
rect 30044 37828 30100 37838
rect 30156 37828 30212 37996
rect 34300 38050 34356 38062
rect 34300 37998 34302 38050
rect 34354 37998 34356 38050
rect 32956 37940 33012 37950
rect 32956 37846 33012 37884
rect 33964 37828 34020 37838
rect 30044 37826 30212 37828
rect 30044 37774 30046 37826
rect 30098 37774 30212 37826
rect 30044 37772 30212 37774
rect 30044 37762 30100 37772
rect 29596 37548 29988 37604
rect 29148 37438 29150 37490
rect 29202 37438 29204 37490
rect 29148 37380 29204 37438
rect 29148 37314 29204 37324
rect 29820 37380 29876 37390
rect 27692 37202 27748 37212
rect 29708 37268 29764 37278
rect 29708 37174 29764 37212
rect 27468 36482 27636 36484
rect 27468 36430 27470 36482
rect 27522 36430 27636 36482
rect 27468 36428 27636 36430
rect 29148 37044 29204 37054
rect 27468 36418 27524 36428
rect 27132 36318 27134 36370
rect 27186 36318 27188 36370
rect 27132 36306 27188 36318
rect 26768 36092 27448 36102
rect 26824 36036 26872 36092
rect 26928 36090 26976 36092
rect 27032 36090 27080 36092
rect 26948 36038 26976 36090
rect 27072 36038 27080 36090
rect 26928 36036 26976 36038
rect 27032 36036 27080 36038
rect 27136 36090 27184 36092
rect 27240 36090 27288 36092
rect 27136 36038 27144 36090
rect 27240 36038 27268 36090
rect 27136 36036 27184 36038
rect 27240 36036 27288 36038
rect 27344 36036 27392 36092
rect 26768 36026 27448 36036
rect 24892 34804 24948 34814
rect 24892 34710 24948 34748
rect 24220 34638 24222 34690
rect 24274 34638 24276 34690
rect 24220 34626 24276 34638
rect 26236 34690 26292 34702
rect 26236 34638 26238 34690
rect 26290 34638 26292 34690
rect 20860 34244 20916 34254
rect 19628 33346 19684 33404
rect 20524 34242 20916 34244
rect 20524 34190 20862 34242
rect 20914 34190 20916 34242
rect 20524 34188 20916 34190
rect 19628 33294 19630 33346
rect 19682 33294 19684 33346
rect 19628 33282 19684 33294
rect 20300 33348 20356 33358
rect 20300 33346 20468 33348
rect 20300 33294 20302 33346
rect 20354 33294 20468 33346
rect 20300 33292 20468 33294
rect 20300 33282 20356 33292
rect 19516 33182 19518 33234
rect 19570 33182 19572 33234
rect 19516 33170 19572 33182
rect 17768 32956 18448 32966
rect 17824 32900 17872 32956
rect 17928 32954 17976 32956
rect 18032 32954 18080 32956
rect 17948 32902 17976 32954
rect 18072 32902 18080 32954
rect 17928 32900 17976 32902
rect 18032 32900 18080 32902
rect 18136 32954 18184 32956
rect 18240 32954 18288 32956
rect 18136 32902 18144 32954
rect 18240 32902 18268 32954
rect 18136 32900 18184 32902
rect 18240 32900 18288 32902
rect 18344 32900 18392 32956
rect 17768 32890 18448 32900
rect 20300 32676 20356 32686
rect 20300 31948 20356 32620
rect 20412 32340 20468 33292
rect 20524 32562 20580 34188
rect 20860 34178 20916 34188
rect 22268 33740 22948 33750
rect 22324 33684 22372 33740
rect 22428 33738 22476 33740
rect 22532 33738 22580 33740
rect 22448 33686 22476 33738
rect 22572 33686 22580 33738
rect 22428 33684 22476 33686
rect 22532 33684 22580 33686
rect 22636 33738 22684 33740
rect 22740 33738 22788 33740
rect 22636 33686 22644 33738
rect 22740 33686 22768 33738
rect 22636 33684 22684 33686
rect 22740 33684 22788 33686
rect 22844 33684 22892 33740
rect 22268 33674 22948 33684
rect 20636 33348 20692 33358
rect 21532 33348 21588 33358
rect 20636 33346 21588 33348
rect 20636 33294 20638 33346
rect 20690 33294 21534 33346
rect 21586 33294 21588 33346
rect 20636 33292 21588 33294
rect 20636 33282 20692 33292
rect 21532 33282 21588 33292
rect 21308 33122 21364 33134
rect 21308 33070 21310 33122
rect 21362 33070 21364 33122
rect 20524 32510 20526 32562
rect 20578 32510 20580 32562
rect 20524 32498 20580 32510
rect 21196 32564 21252 32574
rect 21308 32564 21364 33070
rect 23436 32676 23492 32686
rect 23436 32582 23492 32620
rect 21196 32562 21364 32564
rect 21196 32510 21198 32562
rect 21250 32510 21364 32562
rect 21196 32508 21364 32510
rect 26124 32564 26180 32574
rect 26236 32564 26292 34638
rect 27468 34692 27524 34702
rect 27468 34690 27636 34692
rect 27468 34638 27470 34690
rect 27522 34638 27636 34690
rect 27468 34636 27636 34638
rect 27468 34626 27524 34636
rect 26768 34524 27448 34534
rect 26824 34468 26872 34524
rect 26928 34522 26976 34524
rect 27032 34522 27080 34524
rect 26948 34470 26976 34522
rect 27072 34470 27080 34522
rect 26928 34468 26976 34470
rect 27032 34468 27080 34470
rect 27136 34522 27184 34524
rect 27240 34522 27288 34524
rect 27136 34470 27144 34522
rect 27240 34470 27268 34522
rect 27136 34468 27184 34470
rect 27240 34468 27288 34470
rect 27344 34468 27392 34524
rect 26768 34458 27448 34468
rect 27580 34356 27636 34636
rect 27356 34300 27636 34356
rect 27356 34130 27412 34300
rect 27356 34078 27358 34130
rect 27410 34078 27412 34130
rect 27356 34066 27412 34078
rect 27804 34130 27860 34142
rect 27804 34078 27806 34130
rect 27858 34078 27860 34130
rect 27020 34018 27076 34030
rect 27020 33966 27022 34018
rect 27074 33966 27076 34018
rect 27020 33908 27076 33966
rect 27804 33908 27860 34078
rect 27020 33852 27860 33908
rect 26768 32956 27448 32966
rect 26824 32900 26872 32956
rect 26928 32954 26976 32956
rect 27032 32954 27080 32956
rect 26948 32902 26976 32954
rect 27072 32902 27080 32954
rect 26928 32900 26976 32902
rect 27032 32900 27080 32902
rect 27136 32954 27184 32956
rect 27240 32954 27288 32956
rect 27136 32902 27144 32954
rect 27240 32902 27268 32954
rect 27136 32900 27184 32902
rect 27240 32900 27288 32902
rect 27344 32900 27392 32956
rect 26768 32890 27448 32900
rect 26124 32562 26292 32564
rect 26124 32510 26126 32562
rect 26178 32510 26292 32562
rect 26124 32508 26292 32510
rect 26460 32562 26516 32574
rect 26460 32510 26462 32562
rect 26514 32510 26516 32562
rect 21196 32498 21252 32508
rect 26124 32498 26180 32508
rect 25788 32450 25844 32462
rect 25788 32398 25790 32450
rect 25842 32398 25844 32450
rect 20412 32274 20468 32284
rect 24220 32340 24276 32350
rect 24220 32246 24276 32284
rect 25788 32340 25844 32398
rect 26460 32340 26516 32510
rect 25788 32284 26516 32340
rect 22268 32172 22948 32182
rect 22324 32116 22372 32172
rect 22428 32170 22476 32172
rect 22532 32170 22580 32172
rect 22448 32118 22476 32170
rect 22572 32118 22580 32170
rect 22428 32116 22476 32118
rect 22532 32116 22580 32118
rect 22636 32170 22684 32172
rect 22740 32170 22788 32172
rect 22636 32118 22644 32170
rect 22740 32118 22768 32170
rect 22636 32116 22684 32118
rect 22740 32116 22788 32118
rect 22844 32116 22892 32172
rect 22268 32106 22948 32116
rect 20188 31892 20356 31948
rect 19964 31836 20244 31892
rect 16716 31602 16772 31612
rect 18060 31668 18116 31678
rect 18060 31574 18116 31612
rect 17500 31556 17556 31566
rect 18396 31556 18452 31594
rect 17556 31500 17668 31556
rect 17500 31462 17556 31500
rect 15932 30324 15988 30334
rect 15932 30230 15988 30268
rect 16828 30324 16884 30334
rect 15372 30046 15374 30098
rect 15426 30046 15428 30098
rect 15372 30034 15428 30046
rect 16268 30100 16324 30110
rect 16268 30006 16324 30044
rect 16828 29988 16884 30268
rect 16828 29986 16996 29988
rect 16828 29934 16830 29986
rect 16882 29934 16996 29986
rect 16828 29932 16996 29934
rect 16828 29922 16884 29932
rect 16156 29538 16212 29550
rect 16156 29486 16158 29538
rect 16210 29486 16212 29538
rect 16156 29316 16212 29486
rect 16156 29250 16212 29260
rect 16940 29202 16996 29932
rect 16940 29150 16942 29202
rect 16994 29150 16996 29202
rect 16940 28868 16996 29150
rect 16940 28802 16996 28812
rect 15148 27188 15204 27804
rect 17388 28084 17444 28094
rect 17388 27298 17444 28028
rect 17388 27246 17390 27298
rect 17442 27246 17444 27298
rect 17388 27234 17444 27246
rect 15148 27122 15204 27132
rect 17612 27188 17668 31500
rect 18396 31490 18452 31500
rect 19964 31556 20020 31836
rect 17768 31388 18448 31398
rect 17824 31332 17872 31388
rect 17928 31386 17976 31388
rect 18032 31386 18080 31388
rect 17948 31334 17976 31386
rect 18072 31334 18080 31386
rect 17928 31332 17976 31334
rect 18032 31332 18080 31334
rect 18136 31386 18184 31388
rect 18240 31386 18288 31388
rect 18136 31334 18144 31386
rect 18240 31334 18268 31386
rect 18136 31332 18184 31334
rect 18240 31332 18288 31334
rect 18344 31332 18392 31388
rect 17768 31322 18448 31332
rect 19964 31218 20020 31500
rect 19964 31166 19966 31218
rect 20018 31166 20020 31218
rect 19964 30324 20020 31166
rect 20860 31106 20916 31118
rect 20860 31054 20862 31106
rect 20914 31054 20916 31106
rect 20412 30996 20468 31006
rect 20860 30996 20916 31054
rect 23996 31106 24052 31118
rect 23996 31054 23998 31106
rect 24050 31054 24052 31106
rect 21084 30996 21140 31006
rect 20860 30994 21140 30996
rect 20860 30942 21086 30994
rect 21138 30942 21140 30994
rect 20860 30940 21140 30942
rect 20412 30902 20468 30940
rect 21084 30930 21140 30940
rect 21644 30996 21700 31006
rect 21644 30902 21700 30940
rect 22268 30604 22948 30614
rect 22324 30548 22372 30604
rect 22428 30602 22476 30604
rect 22532 30602 22580 30604
rect 22448 30550 22476 30602
rect 22572 30550 22580 30602
rect 22428 30548 22476 30550
rect 22532 30548 22580 30550
rect 22636 30602 22684 30604
rect 22740 30602 22788 30604
rect 22636 30550 22644 30602
rect 22740 30550 22768 30602
rect 22636 30548 22684 30550
rect 22740 30548 22788 30550
rect 22844 30548 22892 30604
rect 22268 30538 22948 30548
rect 19964 30258 20020 30268
rect 21532 30100 21588 30110
rect 17768 29820 18448 29830
rect 17824 29764 17872 29820
rect 17928 29818 17976 29820
rect 18032 29818 18080 29820
rect 17948 29766 17976 29818
rect 18072 29766 18080 29818
rect 17928 29764 17976 29766
rect 18032 29764 18080 29766
rect 18136 29818 18184 29820
rect 18240 29818 18288 29820
rect 18136 29766 18144 29818
rect 18240 29766 18268 29818
rect 18136 29764 18184 29766
rect 18240 29764 18288 29766
rect 18344 29764 18392 29820
rect 17768 29754 18448 29764
rect 21532 29650 21588 30044
rect 21532 29598 21534 29650
rect 21586 29598 21588 29650
rect 21532 29586 21588 29598
rect 22428 30100 22484 30110
rect 22428 29650 22484 30044
rect 23996 30100 24052 31054
rect 24780 30772 24836 30782
rect 24780 30770 25172 30772
rect 24780 30718 24782 30770
rect 24834 30718 25172 30770
rect 24780 30716 25172 30718
rect 24780 30706 24836 30716
rect 23996 30034 24052 30044
rect 22428 29598 22430 29650
rect 22482 29598 22484 29650
rect 22428 29586 22484 29598
rect 18172 29538 18228 29550
rect 18172 29486 18174 29538
rect 18226 29486 18228 29538
rect 17724 29428 17780 29438
rect 18172 29428 18228 29486
rect 18396 29428 18452 29438
rect 18172 29426 18452 29428
rect 18172 29374 18398 29426
rect 18450 29374 18452 29426
rect 18172 29372 18452 29374
rect 17724 29334 17780 29372
rect 18396 29362 18452 29372
rect 18956 29428 19012 29438
rect 18956 29334 19012 29372
rect 22092 29202 22148 29214
rect 22092 29150 22094 29202
rect 22146 29150 22148 29202
rect 21980 28756 22036 28766
rect 17768 28252 18448 28262
rect 17824 28196 17872 28252
rect 17928 28250 17976 28252
rect 18032 28250 18080 28252
rect 17948 28198 17976 28250
rect 18072 28198 18080 28250
rect 17928 28196 17976 28198
rect 18032 28196 18080 28198
rect 18136 28250 18184 28252
rect 18240 28250 18288 28252
rect 18136 28198 18144 28250
rect 18240 28198 18268 28250
rect 18136 28196 18184 28198
rect 18240 28196 18288 28198
rect 18344 28196 18392 28252
rect 17768 28186 18448 28196
rect 17724 27188 17780 27198
rect 17612 27186 17780 27188
rect 17612 27134 17726 27186
rect 17778 27134 17780 27186
rect 17612 27132 17780 27134
rect 14252 27076 14308 27086
rect 14140 27074 14308 27076
rect 14140 27022 14254 27074
rect 14306 27022 14308 27074
rect 14140 27020 14308 27022
rect 13916 27010 13972 27020
rect 14252 27010 14308 27020
rect 16604 26964 16660 26974
rect 16604 26870 16660 26908
rect 17612 26964 17668 27132
rect 17724 27122 17780 27132
rect 20748 27188 20804 27198
rect 20748 27094 20804 27132
rect 21980 27188 22036 28700
rect 21756 27076 21812 27086
rect 21756 26982 21812 27020
rect 12012 26852 12068 26862
rect 11452 26516 11508 26526
rect 12012 26516 12068 26796
rect 11452 26514 12068 26516
rect 11452 26462 11454 26514
rect 11506 26462 12014 26514
rect 12066 26462 12068 26514
rect 11452 26460 12068 26462
rect 11452 26450 11508 26460
rect 12012 26450 12068 26460
rect 17612 26516 17668 26908
rect 21980 26962 22036 27132
rect 21980 26910 21982 26962
rect 22034 26910 22036 26962
rect 21980 26898 22036 26910
rect 22092 26964 22148 29150
rect 22268 29036 22948 29046
rect 22324 28980 22372 29036
rect 22428 29034 22476 29036
rect 22532 29034 22580 29036
rect 22448 28982 22476 29034
rect 22572 28982 22580 29034
rect 22428 28980 22476 28982
rect 22532 28980 22580 28982
rect 22636 29034 22684 29036
rect 22740 29034 22788 29036
rect 22636 28982 22644 29034
rect 22740 28982 22768 29034
rect 22636 28980 22684 28982
rect 22740 28980 22788 28982
rect 22844 28980 22892 29036
rect 22268 28970 22948 28980
rect 24220 28756 24276 28766
rect 24220 28662 24276 28700
rect 24444 28644 24500 28654
rect 24444 27858 24500 28588
rect 25116 28532 25172 30716
rect 25452 30212 25508 30222
rect 25452 28756 25508 30156
rect 25452 28644 25508 28700
rect 25340 28642 25508 28644
rect 25340 28590 25454 28642
rect 25506 28590 25508 28642
rect 25340 28588 25508 28590
rect 25228 28532 25284 28542
rect 25116 28530 25284 28532
rect 25116 28478 25230 28530
rect 25282 28478 25284 28530
rect 25116 28476 25284 28478
rect 25228 28466 25284 28476
rect 24668 28420 24724 28430
rect 24668 28418 24836 28420
rect 24668 28366 24670 28418
rect 24722 28366 24836 28418
rect 24668 28364 24836 28366
rect 24668 28354 24724 28364
rect 24444 27806 24446 27858
rect 24498 27806 24500 27858
rect 24444 27794 24500 27806
rect 24668 27970 24724 27982
rect 24668 27918 24670 27970
rect 24722 27918 24724 27970
rect 24668 27860 24724 27918
rect 24780 27860 24836 28364
rect 25116 27860 25172 27870
rect 24780 27858 25172 27860
rect 24780 27806 25118 27858
rect 25170 27806 25172 27858
rect 24780 27804 25172 27806
rect 24668 27794 24724 27804
rect 25116 27794 25172 27804
rect 22268 27468 22948 27478
rect 22324 27412 22372 27468
rect 22428 27466 22476 27468
rect 22532 27466 22580 27468
rect 22448 27414 22476 27466
rect 22572 27414 22580 27466
rect 22428 27412 22476 27414
rect 22532 27412 22580 27414
rect 22636 27466 22684 27468
rect 22740 27466 22788 27468
rect 22636 27414 22644 27466
rect 22740 27414 22768 27466
rect 22636 27412 22684 27414
rect 22740 27412 22788 27414
rect 22844 27412 22892 27468
rect 22268 27402 22948 27412
rect 23100 27076 23156 27086
rect 22316 26964 22372 26974
rect 22092 26962 22372 26964
rect 22092 26910 22318 26962
rect 22370 26910 22372 26962
rect 22092 26908 22372 26910
rect 22316 26898 22372 26908
rect 19740 26850 19796 26862
rect 21420 26852 21476 26862
rect 19740 26798 19742 26850
rect 19794 26798 19796 26850
rect 17768 26684 18448 26694
rect 17824 26628 17872 26684
rect 17928 26682 17976 26684
rect 18032 26682 18080 26684
rect 17948 26630 17976 26682
rect 18072 26630 18080 26682
rect 17928 26628 17976 26630
rect 18032 26628 18080 26630
rect 18136 26682 18184 26684
rect 18240 26682 18288 26684
rect 18136 26630 18144 26682
rect 18240 26630 18268 26682
rect 18136 26628 18184 26630
rect 18240 26628 18288 26630
rect 18344 26628 18392 26684
rect 17768 26618 18448 26628
rect 17612 26450 17668 26460
rect 19180 26516 19236 26526
rect 19628 26516 19684 26526
rect 19180 26422 19236 26460
rect 19516 26460 19628 26516
rect 13268 25900 13948 25910
rect 13324 25844 13372 25900
rect 13428 25898 13476 25900
rect 13532 25898 13580 25900
rect 13448 25846 13476 25898
rect 13572 25846 13580 25898
rect 13428 25844 13476 25846
rect 13532 25844 13580 25846
rect 13636 25898 13684 25900
rect 13740 25898 13788 25900
rect 13636 25846 13644 25898
rect 13740 25846 13768 25898
rect 13636 25844 13684 25846
rect 13740 25844 13788 25846
rect 13844 25844 13892 25900
rect 13268 25834 13948 25844
rect 16156 25732 16212 25742
rect 11340 25506 11396 25518
rect 11340 25454 11342 25506
rect 11394 25454 11396 25506
rect 11340 25284 11396 25454
rect 11340 25218 11396 25228
rect 11564 25396 11620 25406
rect 11228 23998 11230 24050
rect 11282 23998 11284 24050
rect 11228 23986 11284 23998
rect 10892 23886 10894 23938
rect 10946 23886 10948 23938
rect 10108 23326 10110 23378
rect 10162 23326 10164 23378
rect 10108 23314 10164 23326
rect 10444 23826 10500 23838
rect 10444 23774 10446 23826
rect 10498 23774 10500 23826
rect 10220 23268 10276 23278
rect 10220 23174 10276 23212
rect 9884 22260 9940 22270
rect 9772 22204 9884 22260
rect 9772 21028 9828 22204
rect 9884 22194 9940 22204
rect 9884 21698 9940 21710
rect 9884 21646 9886 21698
rect 9938 21646 9940 21698
rect 9884 21588 9940 21646
rect 10108 21588 10164 21598
rect 9884 21586 10164 21588
rect 9884 21534 10110 21586
rect 10162 21534 10164 21586
rect 9884 21532 10164 21534
rect 10108 21522 10164 21532
rect 9884 21028 9940 21038
rect 9772 21026 9940 21028
rect 9772 20974 9886 21026
rect 9938 20974 9940 21026
rect 9772 20972 9940 20974
rect 9884 20962 9940 20972
rect 10444 20132 10500 23774
rect 10892 23154 10948 23886
rect 10892 23102 10894 23154
rect 10946 23102 10948 23154
rect 10892 22370 10948 23102
rect 10892 22318 10894 22370
rect 10946 22318 10948 22370
rect 10892 22306 10948 22318
rect 10780 22260 10836 22270
rect 10780 22166 10836 22204
rect 11564 22148 11620 25340
rect 12348 25396 12404 25406
rect 12348 25302 12404 25340
rect 11676 25282 11732 25294
rect 11676 25230 11678 25282
rect 11730 25230 11732 25282
rect 11676 24722 11732 25230
rect 12684 25284 12740 25294
rect 12684 25190 12740 25228
rect 15148 25284 15204 25294
rect 11900 24948 11956 24958
rect 11900 24854 11956 24892
rect 13244 24948 13300 24958
rect 11676 24670 11678 24722
rect 11730 24670 11732 24722
rect 11676 24658 11732 24670
rect 12460 24834 12516 24846
rect 12460 24782 12462 24834
rect 12514 24782 12516 24834
rect 12460 24724 12516 24782
rect 12684 24724 12740 24734
rect 12460 24722 12740 24724
rect 12460 24670 12686 24722
rect 12738 24670 12740 24722
rect 12460 24668 12740 24670
rect 12684 24658 12740 24668
rect 13244 24722 13300 24892
rect 13244 24670 13246 24722
rect 13298 24670 13300 24722
rect 13244 24658 13300 24670
rect 13268 24332 13948 24342
rect 13324 24276 13372 24332
rect 13428 24330 13476 24332
rect 13532 24330 13580 24332
rect 13448 24278 13476 24330
rect 13572 24278 13580 24330
rect 13428 24276 13476 24278
rect 13532 24276 13580 24278
rect 13636 24330 13684 24332
rect 13740 24330 13788 24332
rect 13636 24278 13644 24330
rect 13740 24278 13768 24330
rect 13636 24276 13684 24278
rect 13740 24276 13788 24278
rect 13844 24276 13892 24332
rect 13268 24266 13948 24276
rect 15148 24052 15204 25228
rect 15148 23986 15204 23996
rect 15596 24834 15652 24846
rect 15596 24782 15598 24834
rect 15650 24782 15652 24834
rect 12460 23716 12516 23726
rect 11676 22148 11732 22158
rect 11564 22092 11676 22148
rect 11676 22054 11732 22092
rect 12460 21812 12516 23660
rect 15596 23716 15652 24782
rect 15820 23938 15876 23950
rect 15820 23886 15822 23938
rect 15874 23886 15876 23938
rect 15820 23716 15876 23886
rect 16156 23938 16212 25676
rect 17768 25116 18448 25126
rect 17824 25060 17872 25116
rect 17928 25114 17976 25116
rect 18032 25114 18080 25116
rect 17948 25062 17976 25114
rect 18072 25062 18080 25114
rect 17928 25060 17976 25062
rect 18032 25060 18080 25062
rect 18136 25114 18184 25116
rect 18240 25114 18288 25116
rect 18136 25062 18144 25114
rect 18240 25062 18268 25114
rect 18136 25060 18184 25062
rect 18240 25060 18288 25062
rect 18344 25060 18392 25116
rect 17768 25050 18448 25060
rect 16604 24834 16660 24846
rect 16604 24782 16606 24834
rect 16658 24782 16660 24834
rect 16380 24498 16436 24510
rect 16380 24446 16382 24498
rect 16434 24446 16436 24498
rect 16380 24052 16436 24446
rect 16380 23986 16436 23996
rect 16156 23886 16158 23938
rect 16210 23886 16212 23938
rect 16156 23874 16212 23886
rect 16604 23828 16660 24782
rect 19516 24052 19572 26460
rect 19628 26450 19684 26460
rect 19628 26292 19684 26302
rect 19740 26292 19796 26798
rect 20860 26850 21476 26852
rect 20860 26798 21422 26850
rect 21474 26798 21476 26850
rect 20860 26796 21476 26798
rect 19628 26290 19796 26292
rect 19628 26238 19630 26290
rect 19682 26238 19796 26290
rect 19628 26236 19796 26238
rect 20076 26292 20132 26302
rect 20076 26290 20356 26292
rect 20076 26238 20078 26290
rect 20130 26238 20356 26290
rect 20076 26236 20356 26238
rect 19628 26226 19684 26236
rect 20076 26226 20132 26236
rect 20076 25340 20244 25396
rect 19628 24052 19684 24062
rect 16268 23772 16660 23828
rect 18732 24050 19684 24052
rect 18732 23998 19630 24050
rect 19682 23998 19684 24050
rect 18732 23996 19684 23998
rect 16268 23716 16324 23772
rect 15820 23660 16324 23716
rect 18732 23714 18788 23996
rect 18732 23662 18734 23714
rect 18786 23662 18788 23714
rect 15596 23650 15652 23660
rect 17768 23548 18448 23558
rect 17824 23492 17872 23548
rect 17928 23546 17976 23548
rect 18032 23546 18080 23548
rect 17948 23494 17976 23546
rect 18072 23494 18080 23546
rect 17928 23492 17976 23494
rect 18032 23492 18080 23494
rect 18136 23546 18184 23548
rect 18240 23546 18288 23548
rect 18136 23494 18144 23546
rect 18240 23494 18268 23546
rect 18136 23492 18184 23494
rect 18240 23492 18288 23494
rect 18344 23492 18392 23548
rect 17768 23482 18448 23492
rect 13268 22764 13948 22774
rect 13324 22708 13372 22764
rect 13428 22762 13476 22764
rect 13532 22762 13580 22764
rect 13448 22710 13476 22762
rect 13572 22710 13580 22762
rect 13428 22708 13476 22710
rect 13532 22708 13580 22710
rect 13636 22762 13684 22764
rect 13740 22762 13788 22764
rect 13636 22710 13644 22762
rect 13740 22710 13768 22762
rect 13636 22708 13684 22710
rect 13740 22708 13788 22710
rect 13844 22708 13892 22764
rect 13268 22698 13948 22708
rect 14588 22148 14644 22158
rect 14644 22092 14756 22148
rect 14588 22054 14644 22092
rect 12460 21746 12516 21756
rect 13020 21812 13076 21822
rect 14700 21812 14756 22092
rect 14924 22146 14980 22158
rect 14924 22094 14926 22146
rect 14978 22094 14980 22146
rect 14812 21812 14868 21822
rect 14700 21756 14812 21812
rect 13020 21718 13076 21756
rect 14812 21746 14868 21756
rect 13804 21700 13860 21710
rect 13804 21606 13860 21644
rect 14588 21698 14644 21710
rect 14588 21646 14590 21698
rect 14642 21646 14644 21698
rect 10668 21588 10724 21598
rect 10668 21494 10724 21532
rect 14364 21588 14420 21598
rect 14364 21494 14420 21532
rect 13268 21196 13948 21206
rect 13324 21140 13372 21196
rect 13428 21194 13476 21196
rect 13532 21194 13580 21196
rect 13448 21142 13476 21194
rect 13572 21142 13580 21194
rect 13428 21140 13476 21142
rect 13532 21140 13580 21142
rect 13636 21194 13684 21196
rect 13740 21194 13788 21196
rect 13636 21142 13644 21194
rect 13740 21142 13768 21194
rect 13636 21140 13684 21142
rect 13740 21140 13788 21142
rect 13844 21140 13892 21196
rect 13268 21130 13948 21140
rect 14588 20804 14644 21646
rect 14588 20738 14644 20748
rect 14924 20802 14980 22094
rect 17768 21980 18448 21990
rect 17824 21924 17872 21980
rect 17928 21978 17976 21980
rect 18032 21978 18080 21980
rect 17948 21926 17976 21978
rect 18072 21926 18080 21978
rect 17928 21924 17976 21926
rect 18032 21924 18080 21926
rect 18136 21978 18184 21980
rect 18240 21978 18288 21980
rect 18136 21926 18144 21978
rect 18240 21926 18268 21978
rect 18136 21924 18184 21926
rect 18240 21924 18288 21926
rect 18344 21924 18392 21980
rect 17768 21914 18448 21924
rect 15596 21812 15652 21822
rect 15148 21700 15204 21710
rect 15148 21606 15204 21644
rect 15596 21698 15652 21756
rect 15596 21646 15598 21698
rect 15650 21646 15652 21698
rect 15596 21634 15652 21646
rect 16156 21588 16212 21598
rect 16156 21494 16212 21532
rect 17836 21586 17892 21598
rect 17836 21534 17838 21586
rect 17890 21534 17892 21586
rect 16828 21474 16884 21486
rect 16828 21422 16830 21474
rect 16882 21422 16884 21474
rect 15820 21362 15876 21374
rect 15820 21310 15822 21362
rect 15874 21310 15876 21362
rect 15820 20916 15876 21310
rect 15820 20850 15876 20860
rect 16828 20916 16884 21422
rect 16828 20850 16884 20860
rect 17500 21476 17556 21486
rect 17836 21476 17892 21534
rect 17500 21474 17892 21476
rect 17500 21422 17502 21474
rect 17554 21422 17892 21474
rect 17500 21420 17892 21422
rect 18732 21474 18788 23662
rect 19292 23716 19348 23726
rect 19292 23622 19348 23660
rect 19628 23268 19684 23996
rect 19628 23202 19684 23212
rect 20076 21812 20132 25340
rect 20188 24052 20244 25340
rect 20300 25394 20356 26236
rect 20860 26068 20916 26796
rect 21420 26786 21476 26796
rect 23100 26850 23156 27020
rect 23100 26798 23102 26850
rect 23154 26798 23156 26850
rect 22316 26516 22372 26526
rect 22316 26422 22372 26460
rect 23100 26516 23156 26798
rect 23100 26422 23156 26460
rect 20636 26012 20916 26068
rect 20636 25506 20692 26012
rect 22268 25900 22948 25910
rect 22324 25844 22372 25900
rect 22428 25898 22476 25900
rect 22532 25898 22580 25900
rect 22448 25846 22476 25898
rect 22572 25846 22580 25898
rect 22428 25844 22476 25846
rect 22532 25844 22580 25846
rect 22636 25898 22684 25900
rect 22740 25898 22788 25900
rect 22636 25846 22644 25898
rect 22740 25846 22768 25898
rect 22636 25844 22684 25846
rect 22740 25844 22788 25846
rect 22844 25844 22892 25900
rect 22268 25834 22948 25844
rect 25228 25620 25284 25630
rect 25340 25620 25396 28588
rect 25452 28578 25508 28588
rect 25676 27860 25732 27870
rect 25676 27766 25732 27804
rect 25228 25618 25396 25620
rect 25228 25566 25230 25618
rect 25282 25566 25396 25618
rect 25228 25564 25396 25566
rect 25228 25554 25284 25564
rect 20636 25454 20638 25506
rect 20690 25454 20692 25506
rect 20636 25442 20692 25454
rect 25340 25508 25396 25564
rect 25676 25620 25732 25630
rect 25676 25526 25732 25564
rect 25340 25442 25396 25452
rect 20300 25342 20302 25394
rect 20354 25342 20356 25394
rect 20300 25330 20356 25342
rect 22268 24332 22948 24342
rect 22324 24276 22372 24332
rect 22428 24330 22476 24332
rect 22532 24330 22580 24332
rect 22448 24278 22476 24330
rect 22572 24278 22580 24330
rect 22428 24276 22476 24278
rect 22532 24276 22580 24278
rect 22636 24330 22684 24332
rect 22740 24330 22788 24332
rect 22636 24278 22644 24330
rect 22740 24278 22768 24330
rect 22636 24276 22684 24278
rect 22740 24276 22788 24278
rect 22844 24276 22892 24332
rect 22268 24266 22948 24276
rect 20300 24052 20356 24062
rect 20188 24050 21588 24052
rect 20188 23998 20302 24050
rect 20354 23998 21588 24050
rect 20188 23996 21588 23998
rect 20300 23986 20356 23996
rect 21532 23938 21588 23996
rect 21532 23886 21534 23938
rect 21586 23886 21588 23938
rect 21532 23874 21588 23886
rect 22204 23938 22260 23950
rect 22204 23886 22206 23938
rect 22258 23886 22260 23938
rect 21420 23826 21476 23838
rect 21420 23774 21422 23826
rect 21474 23774 21476 23826
rect 20636 23714 20692 23726
rect 20636 23662 20638 23714
rect 20690 23662 20692 23714
rect 20300 23268 20356 23278
rect 20300 23174 20356 23212
rect 20636 23154 20692 23662
rect 21420 23716 21476 23774
rect 21420 23650 21476 23660
rect 21644 23716 21700 23726
rect 20636 23102 20638 23154
rect 20690 23102 20692 23154
rect 20636 23090 20692 23102
rect 21196 23156 21252 23166
rect 21196 23154 21364 23156
rect 21196 23102 21198 23154
rect 21250 23102 21364 23154
rect 21196 23100 21364 23102
rect 21196 23090 21252 23100
rect 21308 22258 21364 23100
rect 21644 22370 21700 23660
rect 21644 22318 21646 22370
rect 21698 22318 21700 22370
rect 21644 22306 21700 22318
rect 21756 23268 21812 23278
rect 21308 22206 21310 22258
rect 21362 22206 21364 22258
rect 21308 22194 21364 22206
rect 20076 21746 20132 21756
rect 18732 21422 18734 21474
rect 18786 21422 18788 21474
rect 14924 20750 14926 20802
rect 14978 20750 14980 20802
rect 14924 20738 14980 20750
rect 15260 20804 15316 20814
rect 15260 20710 15316 20748
rect 10444 20066 10500 20076
rect 17500 19908 17556 21420
rect 18396 20916 18452 20926
rect 18396 20822 18452 20860
rect 18732 20914 18788 21422
rect 18732 20862 18734 20914
rect 18786 20862 18788 20914
rect 17836 20692 17892 20702
rect 18732 20692 18788 20862
rect 17836 20578 17892 20636
rect 17836 20526 17838 20578
rect 17890 20526 17892 20578
rect 17836 20514 17892 20526
rect 18508 20636 18732 20692
rect 17768 20412 18448 20422
rect 17824 20356 17872 20412
rect 17928 20410 17976 20412
rect 18032 20410 18080 20412
rect 17948 20358 17976 20410
rect 18072 20358 18080 20410
rect 17928 20356 17976 20358
rect 18032 20356 18080 20358
rect 18136 20410 18184 20412
rect 18240 20410 18288 20412
rect 18136 20358 18144 20410
rect 18240 20358 18268 20410
rect 18136 20356 18184 20358
rect 18240 20356 18288 20358
rect 18344 20356 18392 20412
rect 17768 20346 18448 20356
rect 18172 20244 18228 20254
rect 18508 20244 18564 20636
rect 18732 20626 18788 20636
rect 18172 20242 18564 20244
rect 18172 20190 18174 20242
rect 18226 20190 18564 20242
rect 18172 20188 18564 20190
rect 19068 20578 19124 20590
rect 19068 20526 19070 20578
rect 19122 20526 19124 20578
rect 18172 20178 18228 20188
rect 18956 20020 19012 20030
rect 19068 20020 19124 20526
rect 21756 20242 21812 23212
rect 22204 23156 22260 23886
rect 22540 23716 22596 23726
rect 22540 23622 22596 23660
rect 23100 23714 23156 23726
rect 23100 23662 23102 23714
rect 23154 23662 23156 23714
rect 22204 23090 22260 23100
rect 23100 23156 23156 23662
rect 23436 23268 23492 23278
rect 23436 23174 23492 23212
rect 23100 23090 23156 23100
rect 24220 23156 24276 23166
rect 24220 23062 24276 23100
rect 22268 22764 22948 22774
rect 22324 22708 22372 22764
rect 22428 22762 22476 22764
rect 22532 22762 22580 22764
rect 22448 22710 22476 22762
rect 22572 22710 22580 22762
rect 22428 22708 22476 22710
rect 22532 22708 22580 22710
rect 22636 22762 22684 22764
rect 22740 22762 22788 22764
rect 22636 22710 22644 22762
rect 22740 22710 22768 22762
rect 22636 22708 22684 22710
rect 22740 22708 22788 22710
rect 22844 22708 22892 22764
rect 22268 22698 22948 22708
rect 23100 21812 23156 21822
rect 22268 21196 22948 21206
rect 22324 21140 22372 21196
rect 22428 21194 22476 21196
rect 22532 21194 22580 21196
rect 22448 21142 22476 21194
rect 22572 21142 22580 21194
rect 22428 21140 22476 21142
rect 22532 21140 22580 21142
rect 22636 21194 22684 21196
rect 22740 21194 22788 21196
rect 22636 21142 22644 21194
rect 22740 21142 22768 21194
rect 22636 21140 22684 21142
rect 22740 21140 22788 21142
rect 22844 21140 22892 21196
rect 22268 21130 22948 21140
rect 22988 20804 23044 20814
rect 23100 20804 23156 21756
rect 25228 21698 25284 21710
rect 25228 21646 25230 21698
rect 25282 21646 25284 21698
rect 23044 20748 23156 20804
rect 24220 20804 24276 20814
rect 22988 20710 23044 20748
rect 24220 20710 24276 20748
rect 25116 20804 25172 20814
rect 25228 20804 25284 21646
rect 25116 20802 25284 20804
rect 25116 20750 25118 20802
rect 25170 20750 25284 20802
rect 25116 20748 25284 20750
rect 25564 20802 25620 20814
rect 25564 20750 25566 20802
rect 25618 20750 25620 20802
rect 25116 20738 25172 20748
rect 21756 20190 21758 20242
rect 21810 20190 21812 20242
rect 21756 20178 21812 20190
rect 22428 20692 22484 20702
rect 22428 20130 22484 20636
rect 23436 20692 23492 20702
rect 23436 20598 23492 20636
rect 23996 20692 24052 20702
rect 23996 20598 24052 20636
rect 24556 20580 24612 20590
rect 24556 20486 24612 20524
rect 25340 20580 25396 20590
rect 22428 20078 22430 20130
rect 22482 20078 22484 20130
rect 22428 20066 22484 20078
rect 18956 20018 19124 20020
rect 18956 19966 18958 20018
rect 19010 19966 19124 20018
rect 18956 19964 19124 19966
rect 19292 20018 19348 20030
rect 19292 19966 19294 20018
rect 19346 19966 19348 20018
rect 18956 19954 19012 19964
rect 17500 19842 17556 19852
rect 18508 19906 18564 19918
rect 18508 19854 18510 19906
rect 18562 19854 18564 19906
rect 13268 19628 13948 19638
rect 13324 19572 13372 19628
rect 13428 19626 13476 19628
rect 13532 19626 13580 19628
rect 13448 19574 13476 19626
rect 13572 19574 13580 19626
rect 13428 19572 13476 19574
rect 13532 19572 13580 19574
rect 13636 19626 13684 19628
rect 13740 19626 13788 19628
rect 13636 19574 13644 19626
rect 13740 19574 13768 19626
rect 13636 19572 13684 19574
rect 13740 19572 13788 19574
rect 13844 19572 13892 19628
rect 13268 19562 13948 19572
rect 18508 19460 18564 19854
rect 18508 19394 18564 19404
rect 19292 19460 19348 19966
rect 25340 20018 25396 20524
rect 25564 20242 25620 20750
rect 25564 20190 25566 20242
rect 25618 20190 25620 20242
rect 25564 20178 25620 20190
rect 25340 19966 25342 20018
rect 25394 19966 25396 20018
rect 25340 19954 25396 19966
rect 22268 19628 22948 19638
rect 22324 19572 22372 19628
rect 22428 19626 22476 19628
rect 22532 19626 22580 19628
rect 22448 19574 22476 19626
rect 22572 19574 22580 19626
rect 22428 19572 22476 19574
rect 22532 19572 22580 19574
rect 22636 19626 22684 19628
rect 22740 19626 22788 19628
rect 22636 19574 22644 19626
rect 22740 19574 22768 19626
rect 22636 19572 22684 19574
rect 22740 19572 22788 19574
rect 22844 19572 22892 19628
rect 22268 19562 22948 19572
rect 19292 19394 19348 19404
rect 17768 18844 18448 18854
rect 17824 18788 17872 18844
rect 17928 18842 17976 18844
rect 18032 18842 18080 18844
rect 17948 18790 17976 18842
rect 18072 18790 18080 18842
rect 17928 18788 17976 18790
rect 18032 18788 18080 18790
rect 18136 18842 18184 18844
rect 18240 18842 18288 18844
rect 18136 18790 18144 18842
rect 18240 18790 18268 18842
rect 18136 18788 18184 18790
rect 18240 18788 18288 18790
rect 18344 18788 18392 18844
rect 17768 18778 18448 18788
rect 13268 18060 13948 18070
rect 13324 18004 13372 18060
rect 13428 18058 13476 18060
rect 13532 18058 13580 18060
rect 13448 18006 13476 18058
rect 13572 18006 13580 18058
rect 13428 18004 13476 18006
rect 13532 18004 13580 18006
rect 13636 18058 13684 18060
rect 13740 18058 13788 18060
rect 13636 18006 13644 18058
rect 13740 18006 13768 18058
rect 13636 18004 13684 18006
rect 13740 18004 13788 18006
rect 13844 18004 13892 18060
rect 13268 17994 13948 18004
rect 22268 18060 22948 18070
rect 22324 18004 22372 18060
rect 22428 18058 22476 18060
rect 22532 18058 22580 18060
rect 22448 18006 22476 18058
rect 22572 18006 22580 18058
rect 22428 18004 22476 18006
rect 22532 18004 22580 18006
rect 22636 18058 22684 18060
rect 22740 18058 22788 18060
rect 22636 18006 22644 18058
rect 22740 18006 22768 18058
rect 22636 18004 22684 18006
rect 22740 18004 22788 18006
rect 22844 18004 22892 18060
rect 22268 17994 22948 18004
rect 17768 17276 18448 17286
rect 17824 17220 17872 17276
rect 17928 17274 17976 17276
rect 18032 17274 18080 17276
rect 17948 17222 17976 17274
rect 18072 17222 18080 17274
rect 17928 17220 17976 17222
rect 18032 17220 18080 17222
rect 18136 17274 18184 17276
rect 18240 17274 18288 17276
rect 18136 17222 18144 17274
rect 18240 17222 18268 17274
rect 18136 17220 18184 17222
rect 18240 17220 18288 17222
rect 18344 17220 18392 17276
rect 17768 17210 18448 17220
rect 13268 16492 13948 16502
rect 13324 16436 13372 16492
rect 13428 16490 13476 16492
rect 13532 16490 13580 16492
rect 13448 16438 13476 16490
rect 13572 16438 13580 16490
rect 13428 16436 13476 16438
rect 13532 16436 13580 16438
rect 13636 16490 13684 16492
rect 13740 16490 13788 16492
rect 13636 16438 13644 16490
rect 13740 16438 13768 16490
rect 13636 16436 13684 16438
rect 13740 16436 13788 16438
rect 13844 16436 13892 16492
rect 13268 16426 13948 16436
rect 22268 16492 22948 16502
rect 22324 16436 22372 16492
rect 22428 16490 22476 16492
rect 22532 16490 22580 16492
rect 22448 16438 22476 16490
rect 22572 16438 22580 16490
rect 22428 16436 22476 16438
rect 22532 16436 22580 16438
rect 22636 16490 22684 16492
rect 22740 16490 22788 16492
rect 22636 16438 22644 16490
rect 22740 16438 22768 16490
rect 22636 16436 22684 16438
rect 22740 16436 22788 16438
rect 22844 16436 22892 16492
rect 22268 16426 22948 16436
rect 17768 15708 18448 15718
rect 17824 15652 17872 15708
rect 17928 15706 17976 15708
rect 18032 15706 18080 15708
rect 17948 15654 17976 15706
rect 18072 15654 18080 15706
rect 17928 15652 17976 15654
rect 18032 15652 18080 15654
rect 18136 15706 18184 15708
rect 18240 15706 18288 15708
rect 18136 15654 18144 15706
rect 18240 15654 18268 15706
rect 18136 15652 18184 15654
rect 18240 15652 18288 15654
rect 18344 15652 18392 15708
rect 17768 15642 18448 15652
rect 13268 14924 13948 14934
rect 13324 14868 13372 14924
rect 13428 14922 13476 14924
rect 13532 14922 13580 14924
rect 13448 14870 13476 14922
rect 13572 14870 13580 14922
rect 13428 14868 13476 14870
rect 13532 14868 13580 14870
rect 13636 14922 13684 14924
rect 13740 14922 13788 14924
rect 13636 14870 13644 14922
rect 13740 14870 13768 14922
rect 13636 14868 13684 14870
rect 13740 14868 13788 14870
rect 13844 14868 13892 14924
rect 13268 14858 13948 14868
rect 22268 14924 22948 14934
rect 22324 14868 22372 14924
rect 22428 14922 22476 14924
rect 22532 14922 22580 14924
rect 22448 14870 22476 14922
rect 22572 14870 22580 14922
rect 22428 14868 22476 14870
rect 22532 14868 22580 14870
rect 22636 14922 22684 14924
rect 22740 14922 22788 14924
rect 22636 14870 22644 14922
rect 22740 14870 22768 14922
rect 22636 14868 22684 14870
rect 22740 14868 22788 14870
rect 22844 14868 22892 14924
rect 22268 14858 22948 14868
rect 20748 14532 20804 14542
rect 20748 14306 20804 14476
rect 21420 14532 21476 14542
rect 21420 14438 21476 14476
rect 20748 14254 20750 14306
rect 20802 14254 20804 14306
rect 17768 14140 18448 14150
rect 17824 14084 17872 14140
rect 17928 14138 17976 14140
rect 18032 14138 18080 14140
rect 17948 14086 17976 14138
rect 18072 14086 18080 14138
rect 17928 14084 17976 14086
rect 18032 14084 18080 14086
rect 18136 14138 18184 14140
rect 18240 14138 18288 14140
rect 18136 14086 18144 14138
rect 18240 14086 18268 14138
rect 18136 14084 18184 14086
rect 18240 14084 18288 14086
rect 18344 14084 18392 14140
rect 17768 14074 18448 14084
rect 9660 13906 9716 13916
rect 13268 13356 13948 13366
rect 13324 13300 13372 13356
rect 13428 13354 13476 13356
rect 13532 13354 13580 13356
rect 13448 13302 13476 13354
rect 13572 13302 13580 13354
rect 13428 13300 13476 13302
rect 13532 13300 13580 13302
rect 13636 13354 13684 13356
rect 13740 13354 13788 13356
rect 13636 13302 13644 13354
rect 13740 13302 13768 13354
rect 13636 13300 13684 13302
rect 13740 13300 13788 13302
rect 13844 13300 13892 13356
rect 13268 13290 13948 13300
rect 8768 12572 9448 12582
rect 8824 12516 8872 12572
rect 8928 12570 8976 12572
rect 9032 12570 9080 12572
rect 8948 12518 8976 12570
rect 9072 12518 9080 12570
rect 8928 12516 8976 12518
rect 9032 12516 9080 12518
rect 9136 12570 9184 12572
rect 9240 12570 9288 12572
rect 9136 12518 9144 12570
rect 9240 12518 9268 12570
rect 9136 12516 9184 12518
rect 9240 12516 9288 12518
rect 9344 12516 9392 12572
rect 8768 12506 9448 12516
rect 17768 12572 18448 12582
rect 17824 12516 17872 12572
rect 17928 12570 17976 12572
rect 18032 12570 18080 12572
rect 17948 12518 17976 12570
rect 18072 12518 18080 12570
rect 17928 12516 17976 12518
rect 18032 12516 18080 12518
rect 18136 12570 18184 12572
rect 18240 12570 18288 12572
rect 18136 12518 18144 12570
rect 18240 12518 18268 12570
rect 18136 12516 18184 12518
rect 18240 12516 18288 12518
rect 18344 12516 18392 12572
rect 17768 12506 18448 12516
rect 13268 11788 13948 11798
rect 13324 11732 13372 11788
rect 13428 11786 13476 11788
rect 13532 11786 13580 11788
rect 13448 11734 13476 11786
rect 13572 11734 13580 11786
rect 13428 11732 13476 11734
rect 13532 11732 13580 11734
rect 13636 11786 13684 11788
rect 13740 11786 13788 11788
rect 13636 11734 13644 11786
rect 13740 11734 13768 11786
rect 13636 11732 13684 11734
rect 13740 11732 13788 11734
rect 13844 11732 13892 11788
rect 13268 11722 13948 11732
rect 8768 11004 9448 11014
rect 8824 10948 8872 11004
rect 8928 11002 8976 11004
rect 9032 11002 9080 11004
rect 8948 10950 8976 11002
rect 9072 10950 9080 11002
rect 8928 10948 8976 10950
rect 9032 10948 9080 10950
rect 9136 11002 9184 11004
rect 9240 11002 9288 11004
rect 9136 10950 9144 11002
rect 9240 10950 9268 11002
rect 9136 10948 9184 10950
rect 9240 10948 9288 10950
rect 9344 10948 9392 11004
rect 8768 10938 9448 10948
rect 17768 11004 18448 11014
rect 17824 10948 17872 11004
rect 17928 11002 17976 11004
rect 18032 11002 18080 11004
rect 17948 10950 17976 11002
rect 18072 10950 18080 11002
rect 17928 10948 17976 10950
rect 18032 10948 18080 10950
rect 18136 11002 18184 11004
rect 18240 11002 18288 11004
rect 18136 10950 18144 11002
rect 18240 10950 18268 11002
rect 18136 10948 18184 10950
rect 18240 10948 18288 10950
rect 18344 10948 18392 11004
rect 17768 10938 18448 10948
rect 13268 10220 13948 10230
rect 13324 10164 13372 10220
rect 13428 10218 13476 10220
rect 13532 10218 13580 10220
rect 13448 10166 13476 10218
rect 13572 10166 13580 10218
rect 13428 10164 13476 10166
rect 13532 10164 13580 10166
rect 13636 10218 13684 10220
rect 13740 10218 13788 10220
rect 13636 10166 13644 10218
rect 13740 10166 13768 10218
rect 13636 10164 13684 10166
rect 13740 10164 13788 10166
rect 13844 10164 13892 10220
rect 13268 10154 13948 10164
rect 8768 9436 9448 9446
rect 8824 9380 8872 9436
rect 8928 9434 8976 9436
rect 9032 9434 9080 9436
rect 8948 9382 8976 9434
rect 9072 9382 9080 9434
rect 8928 9380 8976 9382
rect 9032 9380 9080 9382
rect 9136 9434 9184 9436
rect 9240 9434 9288 9436
rect 9136 9382 9144 9434
rect 9240 9382 9268 9434
rect 9136 9380 9184 9382
rect 9240 9380 9288 9382
rect 9344 9380 9392 9436
rect 8768 9370 9448 9380
rect 17768 9436 18448 9446
rect 17824 9380 17872 9436
rect 17928 9434 17976 9436
rect 18032 9434 18080 9436
rect 17948 9382 17976 9434
rect 18072 9382 18080 9434
rect 17928 9380 17976 9382
rect 18032 9380 18080 9382
rect 18136 9434 18184 9436
rect 18240 9434 18288 9436
rect 18136 9382 18144 9434
rect 18240 9382 18268 9434
rect 18136 9380 18184 9382
rect 18240 9380 18288 9382
rect 18344 9380 18392 9436
rect 17768 9370 18448 9380
rect 13268 8652 13948 8662
rect 13324 8596 13372 8652
rect 13428 8650 13476 8652
rect 13532 8650 13580 8652
rect 13448 8598 13476 8650
rect 13572 8598 13580 8650
rect 13428 8596 13476 8598
rect 13532 8596 13580 8598
rect 13636 8650 13684 8652
rect 13740 8650 13788 8652
rect 13636 8598 13644 8650
rect 13740 8598 13768 8650
rect 13636 8596 13684 8598
rect 13740 8596 13788 8598
rect 13844 8596 13892 8652
rect 13268 8586 13948 8596
rect 8768 7868 9448 7878
rect 8824 7812 8872 7868
rect 8928 7866 8976 7868
rect 9032 7866 9080 7868
rect 8948 7814 8976 7866
rect 9072 7814 9080 7866
rect 8928 7812 8976 7814
rect 9032 7812 9080 7814
rect 9136 7866 9184 7868
rect 9240 7866 9288 7868
rect 9136 7814 9144 7866
rect 9240 7814 9268 7866
rect 9136 7812 9184 7814
rect 9240 7812 9288 7814
rect 9344 7812 9392 7868
rect 8768 7802 9448 7812
rect 17768 7868 18448 7878
rect 17824 7812 17872 7868
rect 17928 7866 17976 7868
rect 18032 7866 18080 7868
rect 17948 7814 17976 7866
rect 18072 7814 18080 7866
rect 17928 7812 17976 7814
rect 18032 7812 18080 7814
rect 18136 7866 18184 7868
rect 18240 7866 18288 7868
rect 18136 7814 18144 7866
rect 18240 7814 18268 7866
rect 18136 7812 18184 7814
rect 18240 7812 18288 7814
rect 18344 7812 18392 7868
rect 17768 7802 18448 7812
rect 13268 7084 13948 7094
rect 13324 7028 13372 7084
rect 13428 7082 13476 7084
rect 13532 7082 13580 7084
rect 13448 7030 13476 7082
rect 13572 7030 13580 7082
rect 13428 7028 13476 7030
rect 13532 7028 13580 7030
rect 13636 7082 13684 7084
rect 13740 7082 13788 7084
rect 13636 7030 13644 7082
rect 13740 7030 13768 7082
rect 13636 7028 13684 7030
rect 13740 7028 13788 7030
rect 13844 7028 13892 7084
rect 13268 7018 13948 7028
rect 8768 6300 9448 6310
rect 8824 6244 8872 6300
rect 8928 6298 8976 6300
rect 9032 6298 9080 6300
rect 8948 6246 8976 6298
rect 9072 6246 9080 6298
rect 8928 6244 8976 6246
rect 9032 6244 9080 6246
rect 9136 6298 9184 6300
rect 9240 6298 9288 6300
rect 9136 6246 9144 6298
rect 9240 6246 9268 6298
rect 9136 6244 9184 6246
rect 9240 6244 9288 6246
rect 9344 6244 9392 6300
rect 8768 6234 9448 6244
rect 17768 6300 18448 6310
rect 17824 6244 17872 6300
rect 17928 6298 17976 6300
rect 18032 6298 18080 6300
rect 17948 6246 17976 6298
rect 18072 6246 18080 6298
rect 17928 6244 17976 6246
rect 18032 6244 18080 6246
rect 18136 6298 18184 6300
rect 18240 6298 18288 6300
rect 18136 6246 18144 6298
rect 18240 6246 18268 6298
rect 18136 6244 18184 6246
rect 18240 6244 18288 6246
rect 18344 6244 18392 6300
rect 17768 6234 18448 6244
rect 13268 5516 13948 5526
rect 13324 5460 13372 5516
rect 13428 5514 13476 5516
rect 13532 5514 13580 5516
rect 13448 5462 13476 5514
rect 13572 5462 13580 5514
rect 13428 5460 13476 5462
rect 13532 5460 13580 5462
rect 13636 5514 13684 5516
rect 13740 5514 13788 5516
rect 13636 5462 13644 5514
rect 13740 5462 13768 5514
rect 13636 5460 13684 5462
rect 13740 5460 13788 5462
rect 13844 5460 13892 5516
rect 13268 5450 13948 5460
rect 8768 4732 9448 4742
rect 8824 4676 8872 4732
rect 8928 4730 8976 4732
rect 9032 4730 9080 4732
rect 8948 4678 8976 4730
rect 9072 4678 9080 4730
rect 8928 4676 8976 4678
rect 9032 4676 9080 4678
rect 9136 4730 9184 4732
rect 9240 4730 9288 4732
rect 9136 4678 9144 4730
rect 9240 4678 9268 4730
rect 9136 4676 9184 4678
rect 9240 4676 9288 4678
rect 9344 4676 9392 4732
rect 8768 4666 9448 4676
rect 17768 4732 18448 4742
rect 17824 4676 17872 4732
rect 17928 4730 17976 4732
rect 18032 4730 18080 4732
rect 17948 4678 17976 4730
rect 18072 4678 18080 4730
rect 17928 4676 17976 4678
rect 18032 4676 18080 4678
rect 18136 4730 18184 4732
rect 18240 4730 18288 4732
rect 18136 4678 18144 4730
rect 18240 4678 18268 4730
rect 18136 4676 18184 4678
rect 18240 4676 18288 4678
rect 18344 4676 18392 4732
rect 17768 4666 18448 4676
rect 20748 4116 20804 14254
rect 22268 13356 22948 13366
rect 22324 13300 22372 13356
rect 22428 13354 22476 13356
rect 22532 13354 22580 13356
rect 22448 13302 22476 13354
rect 22572 13302 22580 13354
rect 22428 13300 22476 13302
rect 22532 13300 22580 13302
rect 22636 13354 22684 13356
rect 22740 13354 22788 13356
rect 22636 13302 22644 13354
rect 22740 13302 22768 13354
rect 22636 13300 22684 13302
rect 22740 13300 22788 13302
rect 22844 13300 22892 13356
rect 22268 13290 22948 13300
rect 22268 11788 22948 11798
rect 22324 11732 22372 11788
rect 22428 11786 22476 11788
rect 22532 11786 22580 11788
rect 22448 11734 22476 11786
rect 22572 11734 22580 11786
rect 22428 11732 22476 11734
rect 22532 11732 22580 11734
rect 22636 11786 22684 11788
rect 22740 11786 22788 11788
rect 22636 11734 22644 11786
rect 22740 11734 22768 11786
rect 22636 11732 22684 11734
rect 22740 11732 22788 11734
rect 22844 11732 22892 11788
rect 22268 11722 22948 11732
rect 25788 11172 25844 32284
rect 27132 31780 27188 31790
rect 27132 31686 27188 31724
rect 26460 31556 26516 31566
rect 26796 31556 26852 31566
rect 26460 30994 26516 31500
rect 26460 30942 26462 30994
rect 26514 30942 26516 30994
rect 26460 30930 26516 30942
rect 26572 31554 26852 31556
rect 26572 31502 26798 31554
rect 26850 31502 26852 31554
rect 26572 31500 26852 31502
rect 26572 30996 26628 31500
rect 26796 31490 26852 31500
rect 27468 31556 27524 31594
rect 27468 31490 27524 31500
rect 26768 31388 27448 31398
rect 26824 31332 26872 31388
rect 26928 31386 26976 31388
rect 27032 31386 27080 31388
rect 26948 31334 26976 31386
rect 27072 31334 27080 31386
rect 26928 31332 26976 31334
rect 27032 31332 27080 31334
rect 27136 31386 27184 31388
rect 27240 31386 27288 31388
rect 27136 31334 27144 31386
rect 27240 31334 27268 31386
rect 27136 31332 27184 31334
rect 27240 31332 27288 31334
rect 27344 31332 27392 31388
rect 26768 31322 27448 31332
rect 26796 30996 26852 31006
rect 26572 30994 26852 30996
rect 26572 30942 26798 30994
rect 26850 30942 26852 30994
rect 26572 30940 26852 30942
rect 26796 30930 26852 30940
rect 26236 30212 26292 30222
rect 26236 30118 26292 30156
rect 27244 30212 27300 30222
rect 27244 30118 27300 30156
rect 27132 30098 27188 30110
rect 27132 30046 27134 30098
rect 27186 30046 27188 30098
rect 26684 29988 26740 29998
rect 27132 29988 27188 30046
rect 26572 29986 27188 29988
rect 26572 29934 26686 29986
rect 26738 29934 27188 29986
rect 26572 29932 27188 29934
rect 26572 29652 26628 29932
rect 26684 29922 26740 29932
rect 26768 29820 27448 29830
rect 26824 29764 26872 29820
rect 26928 29818 26976 29820
rect 27032 29818 27080 29820
rect 26948 29766 26976 29818
rect 27072 29766 27080 29818
rect 26928 29764 26976 29766
rect 27032 29764 27080 29766
rect 27136 29818 27184 29820
rect 27240 29818 27288 29820
rect 27136 29766 27144 29818
rect 27240 29766 27268 29818
rect 27136 29764 27184 29766
rect 27240 29764 27288 29766
rect 27344 29764 27392 29820
rect 26768 29754 27448 29764
rect 26572 29586 26628 29596
rect 25900 28756 25956 28766
rect 25900 28662 25956 28700
rect 26236 28644 26292 28654
rect 26236 28550 26292 28588
rect 26796 28644 26852 28654
rect 26796 28550 26852 28588
rect 26768 28252 27448 28262
rect 26824 28196 26872 28252
rect 26928 28250 26976 28252
rect 27032 28250 27080 28252
rect 26948 28198 26976 28250
rect 27072 28198 27080 28250
rect 26928 28196 26976 28198
rect 27032 28196 27080 28198
rect 27136 28250 27184 28252
rect 27240 28250 27288 28252
rect 27136 28198 27144 28250
rect 27240 28198 27268 28250
rect 27136 28196 27184 28198
rect 27240 28196 27288 28198
rect 27344 28196 27392 28252
rect 26768 28186 27448 28196
rect 26768 26684 27448 26694
rect 26824 26628 26872 26684
rect 26928 26682 26976 26684
rect 27032 26682 27080 26684
rect 26948 26630 26976 26682
rect 27072 26630 27080 26682
rect 26928 26628 26976 26630
rect 27032 26628 27080 26630
rect 27136 26682 27184 26684
rect 27240 26682 27288 26684
rect 27136 26630 27144 26682
rect 27240 26630 27268 26682
rect 27136 26628 27184 26630
rect 27240 26628 27288 26630
rect 27344 26628 27392 26684
rect 26768 26618 27448 26628
rect 26684 26404 26740 26414
rect 26572 26402 26740 26404
rect 26572 26350 26686 26402
rect 26738 26350 26740 26402
rect 26572 26348 26740 26350
rect 26460 26292 26516 26302
rect 26460 26198 26516 26236
rect 26124 25620 26180 25630
rect 26124 25394 26180 25564
rect 26236 25508 26292 25518
rect 26236 25414 26292 25452
rect 26124 25342 26126 25394
rect 26178 25342 26180 25394
rect 26124 25330 26180 25342
rect 26460 25284 26516 25294
rect 26460 24722 26516 25228
rect 26572 24948 26628 26348
rect 26684 26338 26740 26348
rect 27244 26292 27300 26302
rect 27244 25730 27300 26236
rect 27804 26068 27860 33852
rect 29036 32786 29092 32798
rect 29036 32734 29038 32786
rect 29090 32734 29092 32786
rect 29036 32452 29092 32734
rect 29036 32386 29092 32396
rect 29148 32228 29204 36988
rect 29820 36260 29876 37324
rect 29932 37266 29988 37548
rect 29932 37214 29934 37266
rect 29986 37214 29988 37266
rect 29932 37044 29988 37214
rect 29932 36978 29988 36988
rect 30044 36260 30100 36270
rect 29820 36258 30044 36260
rect 29820 36206 29822 36258
rect 29874 36206 30044 36258
rect 29820 36204 30044 36206
rect 29820 36194 29876 36204
rect 30044 36194 30100 36204
rect 30156 36036 30212 37772
rect 33516 37826 34020 37828
rect 33516 37774 33966 37826
rect 34018 37774 34020 37826
rect 33516 37772 34020 37774
rect 31724 37378 31780 37390
rect 33068 37380 33124 37390
rect 31724 37326 31726 37378
rect 31778 37326 31780 37378
rect 30940 37042 30996 37054
rect 30940 36990 30942 37042
rect 30994 36990 30996 37042
rect 30940 36260 30996 36990
rect 31724 37044 31780 37326
rect 31724 36978 31780 36988
rect 32060 37378 33124 37380
rect 32060 37326 33070 37378
rect 33122 37326 33124 37378
rect 32060 37324 33124 37326
rect 31268 36876 31948 36886
rect 31324 36820 31372 36876
rect 31428 36874 31476 36876
rect 31532 36874 31580 36876
rect 31448 36822 31476 36874
rect 31572 36822 31580 36874
rect 31428 36820 31476 36822
rect 31532 36820 31580 36822
rect 31636 36874 31684 36876
rect 31740 36874 31788 36876
rect 31636 36822 31644 36874
rect 31740 36822 31768 36874
rect 31636 36820 31684 36822
rect 31740 36820 31788 36822
rect 31844 36820 31892 36876
rect 31268 36810 31948 36820
rect 31612 36708 31668 36718
rect 31612 36482 31668 36652
rect 31612 36430 31614 36482
rect 31666 36430 31668 36482
rect 31612 36418 31668 36430
rect 32060 36482 32116 37324
rect 33068 37314 33124 37324
rect 33404 37380 33460 37390
rect 33516 37380 33572 37772
rect 33964 37762 34020 37772
rect 33404 37378 33572 37380
rect 33404 37326 33406 37378
rect 33458 37326 33572 37378
rect 33404 37324 33572 37326
rect 33404 37314 33460 37324
rect 34300 37044 34356 37998
rect 34860 37940 34916 37950
rect 34860 37492 34916 37884
rect 34860 37426 34916 37436
rect 34860 37268 34916 37278
rect 34972 37268 35028 38612
rect 35084 38050 35140 38062
rect 35084 37998 35086 38050
rect 35138 37998 35140 38050
rect 35084 37828 35140 37998
rect 35308 37828 35364 41132
rect 35420 40404 35476 40414
rect 35644 40404 35700 43486
rect 35868 43538 35924 43550
rect 35868 43486 35870 43538
rect 35922 43486 35924 43538
rect 35868 42980 35924 43486
rect 35868 42914 35924 42924
rect 35768 42364 36448 42374
rect 35824 42308 35872 42364
rect 35928 42362 35976 42364
rect 36032 42362 36080 42364
rect 35948 42310 35976 42362
rect 36072 42310 36080 42362
rect 35928 42308 35976 42310
rect 36032 42308 36080 42310
rect 36136 42362 36184 42364
rect 36240 42362 36288 42364
rect 36136 42310 36144 42362
rect 36240 42310 36268 42362
rect 36136 42308 36184 42310
rect 36240 42308 36288 42310
rect 36344 42308 36392 42364
rect 35768 42298 36448 42308
rect 35868 41188 35924 41198
rect 35868 41094 35924 41132
rect 37100 41076 37156 41086
rect 35768 40796 36448 40806
rect 35824 40740 35872 40796
rect 35928 40794 35976 40796
rect 36032 40794 36080 40796
rect 35948 40742 35976 40794
rect 36072 40742 36080 40794
rect 35928 40740 35976 40742
rect 36032 40740 36080 40742
rect 36136 40794 36184 40796
rect 36240 40794 36288 40796
rect 36136 40742 36144 40794
rect 36240 40742 36268 40794
rect 36136 40740 36184 40742
rect 36240 40740 36288 40742
rect 36344 40740 36392 40796
rect 35768 40730 36448 40740
rect 36092 40516 36148 40526
rect 35756 40404 35812 40414
rect 35644 40402 36036 40404
rect 35644 40350 35758 40402
rect 35810 40350 36036 40402
rect 35644 40348 36036 40350
rect 35420 40310 35476 40348
rect 35756 40338 35812 40348
rect 35980 40180 36036 40348
rect 36092 40402 36148 40460
rect 36092 40350 36094 40402
rect 36146 40350 36148 40402
rect 36092 40338 36148 40350
rect 35980 40124 36932 40180
rect 36540 39620 36596 39630
rect 36540 39526 36596 39564
rect 36204 39508 36260 39518
rect 35868 39396 35924 39434
rect 36204 39414 36260 39452
rect 35644 39340 35868 39396
rect 35644 38724 35700 39340
rect 35868 39330 35924 39340
rect 36316 39396 36372 39434
rect 36316 39330 36372 39340
rect 35768 39228 36448 39238
rect 35824 39172 35872 39228
rect 35928 39226 35976 39228
rect 36032 39226 36080 39228
rect 35948 39174 35976 39226
rect 36072 39174 36080 39226
rect 35928 39172 35976 39174
rect 36032 39172 36080 39174
rect 36136 39226 36184 39228
rect 36240 39226 36288 39228
rect 36136 39174 36144 39226
rect 36240 39174 36268 39226
rect 36136 39172 36184 39174
rect 36240 39172 36288 39174
rect 36344 39172 36392 39228
rect 35768 39162 36448 39172
rect 35644 38658 35700 38668
rect 35644 37828 35700 37838
rect 35084 37826 35700 37828
rect 35084 37774 35646 37826
rect 35698 37774 35700 37826
rect 35084 37772 35700 37774
rect 34860 37266 35028 37268
rect 34860 37214 34862 37266
rect 34914 37214 35028 37266
rect 34860 37212 35028 37214
rect 35084 37268 35140 37278
rect 34860 37202 34916 37212
rect 35084 37174 35140 37212
rect 35644 37156 35700 37772
rect 35768 37660 36448 37670
rect 35824 37604 35872 37660
rect 35928 37658 35976 37660
rect 36032 37658 36080 37660
rect 35948 37606 35976 37658
rect 36072 37606 36080 37658
rect 35928 37604 35976 37606
rect 36032 37604 36080 37606
rect 36136 37658 36184 37660
rect 36240 37658 36288 37660
rect 36136 37606 36144 37658
rect 36240 37606 36268 37658
rect 36136 37604 36184 37606
rect 36240 37604 36288 37606
rect 36344 37604 36392 37660
rect 35768 37594 36448 37604
rect 36876 37378 36932 40124
rect 37100 39844 37156 41020
rect 37996 40514 38052 43598
rect 38444 43538 38500 43550
rect 38444 43486 38446 43538
rect 38498 43486 38500 43538
rect 38444 43428 38500 43486
rect 39004 43428 39060 45614
rect 39452 45668 39508 45678
rect 39900 45668 39956 45678
rect 39452 45666 39732 45668
rect 39452 45614 39454 45666
rect 39506 45614 39732 45666
rect 39452 45612 39732 45614
rect 39452 45602 39508 45612
rect 39676 43652 39732 45612
rect 39900 45574 39956 45612
rect 40012 44994 40068 46396
rect 40012 44942 40014 44994
rect 40066 44942 40068 44994
rect 39676 43650 39956 43652
rect 39676 43598 39678 43650
rect 39730 43598 39956 43650
rect 39676 43596 39956 43598
rect 39676 43586 39732 43596
rect 39228 43428 39284 43438
rect 39004 43426 39396 43428
rect 39004 43374 39230 43426
rect 39282 43374 39396 43426
rect 39004 43372 39396 43374
rect 38444 43362 38500 43372
rect 39228 43362 39284 43372
rect 38556 42082 38612 42094
rect 38556 42030 38558 42082
rect 38610 42030 38612 42082
rect 38556 41186 38612 42030
rect 38556 41134 38558 41186
rect 38610 41134 38612 41186
rect 38556 41122 38612 41134
rect 38780 42084 38836 42094
rect 37996 40462 37998 40514
rect 38050 40462 38052 40514
rect 37100 39788 37716 39844
rect 36876 37326 36878 37378
rect 36930 37326 36932 37378
rect 35644 37090 35700 37100
rect 35756 37266 35812 37278
rect 35756 37214 35758 37266
rect 35810 37214 35812 37266
rect 34300 36978 34356 36988
rect 35084 37044 35140 37054
rect 35084 36706 35140 36988
rect 35756 37044 35812 37214
rect 36876 37156 36932 37326
rect 36876 37090 36932 37100
rect 36988 39508 37044 39518
rect 36988 37938 37044 39452
rect 37100 39506 37156 39788
rect 37660 39730 37716 39788
rect 37660 39678 37662 39730
rect 37714 39678 37716 39730
rect 37660 39666 37716 39678
rect 37324 39620 37380 39630
rect 37324 39526 37380 39564
rect 37100 39454 37102 39506
rect 37154 39454 37156 39506
rect 37100 39442 37156 39454
rect 36988 37886 36990 37938
rect 37042 37886 37044 37938
rect 35756 36978 35812 36988
rect 35084 36654 35086 36706
rect 35138 36654 35140 36706
rect 35084 36642 35140 36654
rect 36876 36708 36932 36718
rect 32060 36430 32062 36482
rect 32114 36430 32116 36482
rect 32060 36418 32116 36430
rect 36764 36372 36820 36382
rect 31164 36260 31220 36270
rect 30940 36204 31164 36260
rect 31164 36166 31220 36204
rect 34300 36260 34356 36270
rect 34300 36166 34356 36204
rect 30044 35980 30212 36036
rect 35768 36092 36448 36102
rect 35824 36036 35872 36092
rect 35928 36090 35976 36092
rect 36032 36090 36080 36092
rect 35948 36038 35976 36090
rect 36072 36038 36080 36090
rect 35928 36036 35976 36038
rect 36032 36036 36080 36038
rect 36136 36090 36184 36092
rect 36240 36090 36288 36092
rect 36136 36038 36144 36090
rect 36240 36038 36268 36090
rect 36136 36036 36184 36038
rect 36240 36036 36288 36038
rect 36344 36036 36392 36092
rect 35768 36026 36448 36036
rect 29708 33908 29764 33918
rect 29708 32674 29764 33852
rect 29708 32622 29710 32674
rect 29762 32622 29764 32674
rect 29708 32610 29764 32622
rect 30044 32564 30100 35980
rect 36764 35924 36820 36316
rect 36764 35830 36820 35868
rect 35868 35700 35924 35710
rect 31268 35308 31948 35318
rect 31324 35252 31372 35308
rect 31428 35306 31476 35308
rect 31532 35306 31580 35308
rect 31448 35254 31476 35306
rect 31572 35254 31580 35306
rect 31428 35252 31476 35254
rect 31532 35252 31580 35254
rect 31636 35306 31684 35308
rect 31740 35306 31788 35308
rect 31636 35254 31644 35306
rect 31740 35254 31768 35306
rect 31636 35252 31684 35254
rect 31740 35252 31788 35254
rect 31844 35252 31892 35308
rect 31268 35242 31948 35252
rect 35308 35028 35364 35038
rect 35868 35028 35924 35644
rect 36652 35700 36708 35710
rect 36652 35606 36708 35644
rect 30940 34692 30996 34702
rect 30044 32498 30100 32508
rect 30156 34354 30212 34366
rect 30156 34302 30158 34354
rect 30210 34302 30212 34354
rect 30156 34020 30212 34302
rect 30940 34242 30996 34636
rect 30940 34190 30942 34242
rect 30994 34190 30996 34242
rect 30940 34178 30996 34190
rect 32508 34242 32564 34254
rect 32508 34190 32510 34242
rect 32562 34190 32564 34242
rect 32508 34132 32564 34190
rect 32956 34132 33012 34142
rect 33516 34132 33572 34142
rect 32508 34130 33012 34132
rect 32508 34078 32958 34130
rect 33010 34078 33012 34130
rect 32508 34076 33012 34078
rect 32956 34066 33012 34076
rect 33404 34130 33572 34132
rect 33404 34078 33518 34130
rect 33570 34078 33572 34130
rect 33404 34076 33572 34078
rect 29036 32172 29204 32228
rect 30156 32452 30212 33964
rect 31388 34020 31444 34030
rect 31388 33926 31444 33964
rect 32172 34020 32228 34030
rect 32172 33926 32228 33964
rect 33404 34020 33460 34076
rect 33516 34066 33572 34076
rect 31268 33740 31948 33750
rect 31324 33684 31372 33740
rect 31428 33738 31476 33740
rect 31532 33738 31580 33740
rect 31448 33686 31476 33738
rect 31572 33686 31580 33738
rect 31428 33684 31476 33686
rect 31532 33684 31580 33686
rect 31636 33738 31684 33740
rect 31740 33738 31788 33740
rect 31636 33686 31644 33738
rect 31740 33686 31768 33738
rect 31636 33684 31684 33686
rect 31740 33684 31788 33686
rect 31844 33684 31892 33740
rect 31268 33674 31948 33684
rect 28140 31780 28196 31790
rect 28196 31724 28308 31780
rect 28140 31714 28196 31724
rect 27916 30772 27972 30782
rect 27916 30434 27972 30716
rect 27916 30382 27918 30434
rect 27970 30382 27972 30434
rect 27916 30370 27972 30382
rect 28252 30434 28308 31724
rect 28252 30382 28254 30434
rect 28306 30382 28308 30434
rect 28252 30370 28308 30382
rect 28812 28644 28868 28654
rect 28252 28532 28308 28542
rect 28252 28082 28308 28476
rect 28252 28030 28254 28082
rect 28306 28030 28308 28082
rect 28252 26908 28308 28030
rect 28812 27636 28868 28588
rect 28812 27542 28868 27580
rect 28140 26852 28308 26908
rect 27804 26012 28084 26068
rect 27244 25678 27246 25730
rect 27298 25678 27300 25730
rect 27244 25666 27300 25678
rect 26908 25508 26964 25518
rect 26908 25414 26964 25452
rect 27692 25284 27748 25294
rect 27692 25190 27748 25228
rect 26768 25116 27448 25126
rect 26824 25060 26872 25116
rect 26928 25114 26976 25116
rect 27032 25114 27080 25116
rect 26948 25062 26976 25114
rect 27072 25062 27080 25114
rect 26928 25060 26976 25062
rect 27032 25060 27080 25062
rect 27136 25114 27184 25116
rect 27240 25114 27288 25116
rect 27136 25062 27144 25114
rect 27240 25062 27268 25114
rect 27136 25060 27184 25062
rect 27240 25060 27288 25062
rect 27344 25060 27392 25116
rect 26768 25050 27448 25060
rect 26572 24892 26964 24948
rect 26460 24670 26462 24722
rect 26514 24670 26516 24722
rect 26460 24658 26516 24670
rect 26908 24724 26964 24892
rect 27020 24724 27076 24734
rect 26908 24722 27076 24724
rect 26908 24670 27022 24722
rect 27074 24670 27076 24722
rect 26908 24668 27076 24670
rect 27020 24658 27076 24668
rect 26908 23716 26964 23726
rect 26572 23714 26964 23716
rect 26572 23662 26910 23714
rect 26962 23662 26964 23714
rect 26572 23660 26964 23662
rect 26348 23380 26404 23390
rect 26348 23286 26404 23324
rect 26572 23154 26628 23660
rect 26908 23650 26964 23660
rect 26768 23548 27448 23558
rect 26824 23492 26872 23548
rect 26928 23546 26976 23548
rect 27032 23546 27080 23548
rect 26948 23494 26976 23546
rect 27072 23494 27080 23546
rect 26928 23492 26976 23494
rect 27032 23492 27080 23494
rect 27136 23546 27184 23548
rect 27240 23546 27288 23548
rect 27136 23494 27144 23546
rect 27240 23494 27268 23546
rect 27136 23492 27184 23494
rect 27240 23492 27288 23494
rect 27344 23492 27392 23548
rect 26768 23482 27448 23492
rect 26572 23102 26574 23154
rect 26626 23102 26628 23154
rect 26572 23090 26628 23102
rect 27132 23380 27188 23390
rect 27132 23154 27188 23324
rect 27132 23102 27134 23154
rect 27186 23102 27188 23154
rect 27132 23090 27188 23102
rect 27804 22258 27860 22270
rect 27804 22206 27806 22258
rect 27858 22206 27860 22258
rect 26768 21980 27448 21990
rect 26824 21924 26872 21980
rect 26928 21978 26976 21980
rect 27032 21978 27080 21980
rect 26948 21926 26976 21978
rect 27072 21926 27080 21978
rect 26928 21924 26976 21926
rect 27032 21924 27080 21926
rect 27136 21978 27184 21980
rect 27240 21978 27288 21980
rect 27136 21926 27144 21978
rect 27240 21926 27268 21978
rect 27136 21924 27184 21926
rect 27240 21924 27288 21926
rect 27344 21924 27392 21980
rect 26768 21914 27448 21924
rect 27356 21586 27412 21598
rect 27356 21534 27358 21586
rect 27410 21534 27412 21586
rect 26572 21474 26628 21486
rect 26572 21422 26574 21474
rect 26626 21422 26628 21474
rect 26572 21028 26628 21422
rect 27020 21476 27076 21486
rect 27020 21382 27076 21420
rect 26572 20962 26628 20972
rect 27356 21028 27412 21534
rect 27356 20962 27412 20972
rect 27804 20690 27860 22206
rect 27804 20638 27806 20690
rect 27858 20638 27860 20690
rect 26768 20412 27448 20422
rect 26824 20356 26872 20412
rect 26928 20410 26976 20412
rect 27032 20410 27080 20412
rect 26948 20358 26976 20410
rect 27072 20358 27080 20410
rect 26928 20356 26976 20358
rect 27032 20356 27080 20358
rect 27136 20410 27184 20412
rect 27240 20410 27288 20412
rect 27136 20358 27144 20410
rect 27240 20358 27268 20410
rect 27136 20356 27184 20358
rect 27240 20356 27288 20358
rect 27344 20356 27392 20412
rect 26768 20346 27448 20356
rect 27804 20132 27860 20638
rect 27804 20066 27860 20076
rect 26768 18844 27448 18854
rect 26824 18788 26872 18844
rect 26928 18842 26976 18844
rect 27032 18842 27080 18844
rect 26948 18790 26976 18842
rect 27072 18790 27080 18842
rect 26928 18788 26976 18790
rect 27032 18788 27080 18790
rect 27136 18842 27184 18844
rect 27240 18842 27288 18844
rect 27136 18790 27144 18842
rect 27240 18790 27268 18842
rect 27136 18788 27184 18790
rect 27240 18788 27288 18790
rect 27344 18788 27392 18844
rect 26768 18778 27448 18788
rect 26768 17276 27448 17286
rect 26824 17220 26872 17276
rect 26928 17274 26976 17276
rect 27032 17274 27080 17276
rect 26948 17222 26976 17274
rect 27072 17222 27080 17274
rect 26928 17220 26976 17222
rect 27032 17220 27080 17222
rect 27136 17274 27184 17276
rect 27240 17274 27288 17276
rect 27136 17222 27144 17274
rect 27240 17222 27268 17274
rect 27136 17220 27184 17222
rect 27240 17220 27288 17222
rect 27344 17220 27392 17276
rect 26768 17210 27448 17220
rect 26768 15708 27448 15718
rect 26824 15652 26872 15708
rect 26928 15706 26976 15708
rect 27032 15706 27080 15708
rect 26948 15654 26976 15706
rect 27072 15654 27080 15706
rect 26928 15652 26976 15654
rect 27032 15652 27080 15654
rect 27136 15706 27184 15708
rect 27240 15706 27288 15708
rect 27136 15654 27144 15706
rect 27240 15654 27268 15706
rect 27136 15652 27184 15654
rect 27240 15652 27288 15654
rect 27344 15652 27392 15708
rect 26768 15642 27448 15652
rect 27692 14308 27748 14318
rect 27692 14214 27748 14252
rect 26768 14140 27448 14150
rect 26824 14084 26872 14140
rect 26928 14138 26976 14140
rect 27032 14138 27080 14140
rect 26948 14086 26976 14138
rect 27072 14086 27080 14138
rect 26928 14084 26976 14086
rect 27032 14084 27080 14086
rect 27136 14138 27184 14140
rect 27240 14138 27288 14140
rect 27136 14086 27144 14138
rect 27240 14086 27268 14138
rect 27136 14084 27184 14086
rect 27240 14084 27288 14086
rect 27344 14084 27392 14140
rect 26768 14074 27448 14084
rect 26768 12572 27448 12582
rect 26824 12516 26872 12572
rect 26928 12570 26976 12572
rect 27032 12570 27080 12572
rect 26948 12518 26976 12570
rect 27072 12518 27080 12570
rect 26928 12516 26976 12518
rect 27032 12516 27080 12518
rect 27136 12570 27184 12572
rect 27240 12570 27288 12572
rect 27136 12518 27144 12570
rect 27240 12518 27268 12570
rect 27136 12516 27184 12518
rect 27240 12516 27288 12518
rect 27344 12516 27392 12572
rect 26768 12506 27448 12516
rect 25788 11106 25844 11116
rect 26768 11004 27448 11014
rect 26824 10948 26872 11004
rect 26928 11002 26976 11004
rect 27032 11002 27080 11004
rect 26948 10950 26976 11002
rect 27072 10950 27080 11002
rect 26928 10948 26976 10950
rect 27032 10948 27080 10950
rect 27136 11002 27184 11004
rect 27240 11002 27288 11004
rect 27136 10950 27144 11002
rect 27240 10950 27268 11002
rect 27136 10948 27184 10950
rect 27240 10948 27288 10950
rect 27344 10948 27392 11004
rect 26768 10938 27448 10948
rect 22268 10220 22948 10230
rect 22324 10164 22372 10220
rect 22428 10218 22476 10220
rect 22532 10218 22580 10220
rect 22448 10166 22476 10218
rect 22572 10166 22580 10218
rect 22428 10164 22476 10166
rect 22532 10164 22580 10166
rect 22636 10218 22684 10220
rect 22740 10218 22788 10220
rect 22636 10166 22644 10218
rect 22740 10166 22768 10218
rect 22636 10164 22684 10166
rect 22740 10164 22788 10166
rect 22844 10164 22892 10220
rect 22268 10154 22948 10164
rect 28028 9604 28084 26012
rect 28140 22260 28196 26852
rect 28252 25508 28308 25518
rect 28252 25284 28308 25452
rect 28252 25282 28644 25284
rect 28252 25230 28254 25282
rect 28306 25230 28644 25282
rect 28252 25228 28644 25230
rect 28252 25218 28308 25228
rect 28588 24948 28644 25228
rect 28588 24882 28644 24892
rect 28588 22260 28644 22270
rect 28140 22204 28588 22260
rect 28588 22166 28644 22204
rect 28364 21812 28420 21822
rect 28364 21474 28420 21756
rect 29036 21812 29092 32172
rect 30044 31554 30100 31566
rect 30044 31502 30046 31554
rect 30098 31502 30100 31554
rect 29372 31220 29428 31230
rect 30044 31220 30100 31502
rect 29372 31218 30100 31220
rect 29372 31166 29374 31218
rect 29426 31166 30100 31218
rect 29372 31164 30100 31166
rect 29372 31154 29428 31164
rect 29932 30772 29988 30782
rect 29932 30678 29988 30716
rect 29596 28756 29652 28766
rect 29260 28642 29316 28654
rect 29260 28590 29262 28642
rect 29314 28590 29316 28642
rect 29260 28532 29316 28590
rect 29260 28466 29316 28476
rect 29148 28420 29204 28430
rect 29148 27858 29204 28364
rect 29148 27806 29150 27858
rect 29202 27806 29204 27858
rect 29148 27794 29204 27806
rect 29596 27858 29652 28700
rect 30044 28644 30100 31164
rect 30044 28578 30100 28588
rect 29596 27806 29598 27858
rect 29650 27806 29652 27858
rect 29596 27794 29652 27806
rect 29932 27300 29988 27310
rect 29484 27188 29540 27198
rect 29484 27094 29540 27132
rect 29932 27186 29988 27244
rect 29932 27134 29934 27186
rect 29986 27134 29988 27186
rect 29932 27122 29988 27134
rect 29708 26964 29764 26974
rect 29372 26852 29764 26908
rect 30156 26964 30212 32396
rect 32508 33124 32564 33134
rect 32508 32452 32564 33068
rect 32508 32386 32564 32396
rect 31268 32172 31948 32182
rect 31324 32116 31372 32172
rect 31428 32170 31476 32172
rect 31532 32170 31580 32172
rect 31448 32118 31476 32170
rect 31572 32118 31580 32170
rect 31428 32116 31476 32118
rect 31532 32116 31580 32118
rect 31636 32170 31684 32172
rect 31740 32170 31788 32172
rect 31636 32118 31644 32170
rect 31740 32118 31768 32170
rect 31636 32116 31684 32118
rect 31740 32116 31788 32118
rect 31844 32116 31892 32172
rect 31268 32106 31948 32116
rect 30604 31892 30660 31902
rect 30604 31220 30660 31836
rect 32732 31554 32788 31566
rect 32732 31502 32734 31554
rect 32786 31502 32788 31554
rect 30604 31218 31108 31220
rect 30604 31166 30606 31218
rect 30658 31166 31108 31218
rect 30604 31164 31108 31166
rect 30604 31154 30660 31164
rect 31052 31106 31108 31164
rect 31052 31054 31054 31106
rect 31106 31054 31108 31106
rect 31052 31042 31108 31054
rect 30940 30994 30996 31006
rect 30940 30942 30942 30994
rect 30994 30942 30996 30994
rect 30268 30212 30324 30222
rect 30940 30212 30996 30942
rect 32172 30996 32228 31006
rect 32732 30996 32788 31502
rect 32956 30996 33012 31006
rect 32732 30994 33012 30996
rect 32732 30942 32958 30994
rect 33010 30942 33012 30994
rect 32732 30940 33012 30942
rect 31724 30884 31780 30894
rect 31724 30790 31780 30828
rect 32060 30770 32116 30782
rect 32060 30718 32062 30770
rect 32114 30718 32116 30770
rect 31268 30604 31948 30614
rect 31324 30548 31372 30604
rect 31428 30602 31476 30604
rect 31532 30602 31580 30604
rect 31448 30550 31476 30602
rect 31572 30550 31580 30602
rect 31428 30548 31476 30550
rect 31532 30548 31580 30550
rect 31636 30602 31684 30604
rect 31740 30602 31788 30604
rect 31636 30550 31644 30602
rect 31740 30550 31768 30602
rect 31636 30548 31684 30550
rect 31740 30548 31788 30550
rect 31844 30548 31892 30604
rect 31268 30538 31948 30548
rect 32060 30436 32116 30718
rect 30324 30156 30436 30212
rect 30268 30118 30324 30156
rect 30268 28756 30324 28766
rect 30268 28530 30324 28700
rect 30268 28478 30270 28530
rect 30322 28478 30324 28530
rect 30268 28466 30324 28478
rect 30380 27188 30436 30156
rect 30940 30146 30996 30156
rect 31836 30380 32116 30436
rect 31836 30210 31892 30380
rect 32172 30324 32228 30940
rect 32956 30930 33012 30940
rect 31836 30158 31838 30210
rect 31890 30158 31892 30210
rect 31836 30146 31892 30158
rect 32060 30268 32228 30324
rect 33180 30884 33236 30894
rect 32060 30098 32116 30268
rect 32732 30212 32788 30222
rect 32732 30118 32788 30156
rect 33068 30212 33124 30222
rect 32060 30046 32062 30098
rect 32114 30046 32116 30098
rect 32060 30034 32116 30046
rect 31268 29036 31948 29046
rect 31324 28980 31372 29036
rect 31428 29034 31476 29036
rect 31532 29034 31580 29036
rect 31448 28982 31476 29034
rect 31572 28982 31580 29034
rect 31428 28980 31476 28982
rect 31532 28980 31580 28982
rect 31636 29034 31684 29036
rect 31740 29034 31788 29036
rect 31636 28982 31644 29034
rect 31740 28982 31768 29034
rect 31636 28980 31684 28982
rect 31740 28980 31788 28982
rect 31844 28980 31892 29036
rect 31268 28970 31948 28980
rect 30604 28532 30660 28542
rect 32060 28532 32116 28542
rect 30604 28530 30884 28532
rect 30604 28478 30606 28530
rect 30658 28478 30884 28530
rect 30604 28476 30884 28478
rect 30604 28466 30660 28476
rect 30828 27412 30884 28476
rect 30940 28420 30996 28430
rect 30940 28326 30996 28364
rect 32060 28196 32116 28476
rect 32060 28082 32116 28140
rect 32060 28030 32062 28082
rect 32114 28030 32116 28082
rect 32060 28018 32116 28030
rect 33068 28196 33124 30156
rect 33180 29986 33236 30828
rect 33180 29934 33182 29986
rect 33234 29934 33236 29986
rect 33180 29652 33236 29934
rect 33180 29586 33236 29596
rect 33068 28084 33124 28140
rect 33180 28084 33236 28094
rect 33068 28082 33236 28084
rect 33068 28030 33182 28082
rect 33234 28030 33236 28082
rect 33068 28028 33236 28030
rect 33180 28018 33236 28028
rect 32620 27634 32676 27646
rect 32620 27582 32622 27634
rect 32674 27582 32676 27634
rect 31268 27468 31948 27478
rect 31324 27412 31372 27468
rect 31428 27466 31476 27468
rect 31532 27466 31580 27468
rect 31448 27414 31476 27466
rect 31572 27414 31580 27466
rect 31428 27412 31476 27414
rect 31532 27412 31580 27414
rect 31636 27466 31684 27468
rect 31740 27466 31788 27468
rect 31636 27414 31644 27466
rect 31740 27414 31768 27466
rect 31636 27412 31684 27414
rect 31740 27412 31788 27414
rect 31844 27412 31892 27468
rect 30828 27356 31108 27412
rect 31268 27402 31948 27412
rect 30380 27074 30436 27132
rect 30380 27022 30382 27074
rect 30434 27022 30436 27074
rect 30380 27010 30436 27022
rect 30492 27300 30548 27310
rect 31052 27300 31108 27356
rect 31500 27300 31556 27310
rect 31052 27298 31556 27300
rect 31052 27246 31502 27298
rect 31554 27246 31556 27298
rect 31052 27244 31556 27246
rect 30156 26898 30212 26908
rect 30492 26962 30548 27244
rect 31500 27234 31556 27244
rect 32060 27300 32116 27310
rect 32060 27186 32116 27244
rect 32620 27300 32676 27582
rect 32620 27234 32676 27244
rect 32060 27134 32062 27186
rect 32114 27134 32116 27186
rect 31164 27076 31220 27086
rect 31164 26982 31220 27020
rect 32060 27076 32116 27134
rect 32060 27010 32116 27020
rect 30492 26910 30494 26962
rect 30546 26910 30548 26962
rect 30492 26898 30548 26910
rect 33404 26908 33460 33964
rect 35308 33908 35364 34972
rect 35644 34972 35924 35028
rect 35532 34690 35588 34702
rect 35532 34638 35534 34690
rect 35586 34638 35588 34690
rect 35532 34356 35588 34638
rect 35532 34290 35588 34300
rect 35308 33842 35364 33852
rect 35644 32564 35700 34972
rect 35868 34914 35924 34972
rect 35868 34862 35870 34914
rect 35922 34862 35924 34914
rect 35868 34850 35924 34862
rect 36204 35586 36260 35598
rect 36204 35534 36206 35586
rect 36258 35534 36260 35586
rect 35756 34804 35812 34814
rect 35756 34710 35812 34748
rect 36204 34692 36260 35534
rect 36764 35476 36820 35486
rect 36876 35476 36932 36652
rect 36988 36370 37044 37886
rect 37100 37828 37156 37838
rect 37100 37734 37156 37772
rect 37324 37826 37380 37838
rect 37324 37774 37326 37826
rect 37378 37774 37380 37826
rect 37324 37492 37380 37774
rect 37324 37426 37380 37436
rect 37996 37380 38052 40462
rect 38556 40628 38612 40638
rect 38556 40404 38612 40572
rect 38668 40404 38724 40414
rect 38556 40402 38724 40404
rect 38556 40350 38670 40402
rect 38722 40350 38724 40402
rect 38556 40348 38724 40350
rect 38668 40338 38724 40348
rect 38556 38946 38612 38958
rect 38556 38894 38558 38946
rect 38610 38894 38612 38946
rect 37996 37286 38052 37324
rect 38332 38276 38388 38286
rect 38332 37266 38388 38220
rect 38444 38052 38500 38062
rect 38444 37492 38500 37996
rect 38556 38050 38612 38894
rect 38780 38668 38836 42028
rect 39228 42082 39284 42094
rect 39228 42030 39230 42082
rect 39282 42030 39284 42082
rect 39228 41636 39284 42030
rect 39004 41580 39284 41636
rect 39004 41186 39060 41580
rect 39004 41134 39006 41186
rect 39058 41134 39060 41186
rect 39004 41122 39060 41134
rect 39004 40628 39060 40638
rect 39004 40534 39060 40572
rect 39340 40404 39396 43372
rect 39564 41972 39620 41982
rect 39564 41878 39620 41916
rect 39900 40964 39956 43596
rect 39900 40626 39956 40908
rect 39900 40574 39902 40626
rect 39954 40574 39956 40626
rect 39452 40404 39508 40414
rect 39340 40402 39620 40404
rect 39340 40350 39454 40402
rect 39506 40350 39620 40402
rect 39340 40348 39620 40350
rect 39452 40338 39508 40348
rect 38556 37998 38558 38050
rect 38610 37998 38612 38050
rect 38556 37986 38612 37998
rect 38668 38612 38836 38668
rect 38556 37492 38612 37502
rect 38444 37490 38612 37492
rect 38444 37438 38558 37490
rect 38610 37438 38612 37490
rect 38444 37436 38612 37438
rect 38556 37426 38612 37436
rect 38332 37214 38334 37266
rect 38386 37214 38388 37266
rect 38332 37202 38388 37214
rect 36988 36318 36990 36370
rect 37042 36318 37044 36370
rect 36988 35700 37044 36318
rect 37100 36484 37156 36494
rect 37100 36370 37156 36428
rect 37324 36484 37380 36494
rect 37324 36390 37380 36428
rect 38668 36484 38724 38612
rect 39004 38052 39060 38062
rect 39004 38050 39508 38052
rect 39004 37998 39006 38050
rect 39058 37998 39508 38050
rect 39004 37996 39508 37998
rect 39004 37986 39060 37996
rect 39452 37490 39508 37996
rect 39452 37438 39454 37490
rect 39506 37438 39508 37490
rect 39452 37426 39508 37438
rect 39228 37380 39284 37390
rect 39116 37156 39172 37166
rect 39116 37062 39172 37100
rect 38668 36428 39172 36484
rect 37100 36318 37102 36370
rect 37154 36318 37156 36370
rect 37100 36306 37156 36318
rect 37660 36372 37716 36382
rect 37660 36278 37716 36316
rect 37324 35924 37380 35934
rect 37324 35830 37380 35868
rect 38668 35922 38724 36428
rect 38668 35870 38670 35922
rect 38722 35870 38724 35922
rect 36988 35634 37044 35644
rect 36764 35474 36932 35476
rect 36764 35422 36766 35474
rect 36818 35422 36932 35474
rect 36764 35420 36932 35422
rect 36764 35410 36820 35420
rect 38668 35140 38724 35870
rect 38892 36258 38948 36270
rect 38892 36206 38894 36258
rect 38946 36206 38948 36258
rect 38892 35140 38948 36206
rect 39116 35922 39172 36428
rect 39116 35870 39118 35922
rect 39170 35870 39172 35922
rect 39116 35858 39172 35870
rect 38668 35084 38836 35140
rect 37212 34916 37268 34926
rect 36988 34802 37044 34814
rect 36988 34750 36990 34802
rect 37042 34750 37044 34802
rect 36204 34626 36260 34636
rect 36428 34692 36484 34702
rect 36988 34692 37044 34750
rect 36428 34690 37044 34692
rect 36428 34638 36430 34690
rect 36482 34638 37044 34690
rect 36428 34636 37044 34638
rect 36428 34626 36484 34636
rect 35768 34524 36448 34534
rect 35824 34468 35872 34524
rect 35928 34522 35976 34524
rect 36032 34522 36080 34524
rect 35948 34470 35976 34522
rect 36072 34470 36080 34522
rect 35928 34468 35976 34470
rect 36032 34468 36080 34470
rect 36136 34522 36184 34524
rect 36240 34522 36288 34524
rect 36136 34470 36144 34522
rect 36240 34470 36268 34522
rect 36136 34468 36184 34470
rect 36240 34468 36288 34470
rect 36344 34468 36392 34524
rect 35768 34458 36448 34468
rect 35868 34242 35924 34254
rect 35868 34190 35870 34242
rect 35922 34190 35924 34242
rect 35868 33124 35924 34190
rect 36428 34132 36484 34142
rect 36540 34132 36596 34636
rect 36988 34580 37044 34636
rect 36988 34514 37044 34524
rect 37100 34356 37156 34366
rect 37212 34356 37268 34860
rect 38668 34916 38724 34926
rect 38668 34822 38724 34860
rect 37100 34354 37268 34356
rect 37100 34302 37102 34354
rect 37154 34302 37268 34354
rect 37100 34300 37268 34302
rect 38668 34356 38724 34366
rect 38780 34356 38836 35084
rect 38892 35074 38948 35084
rect 39004 35700 39060 35710
rect 39228 35700 39284 37324
rect 39564 37156 39620 40348
rect 39788 37268 39844 37278
rect 39788 37174 39844 37212
rect 39564 37090 39620 37100
rect 39564 35812 39620 35822
rect 39452 35810 39620 35812
rect 39452 35758 39566 35810
rect 39618 35758 39620 35810
rect 39452 35756 39620 35758
rect 39004 35698 39284 35700
rect 39004 35646 39006 35698
rect 39058 35646 39284 35698
rect 39004 35644 39284 35646
rect 39340 35700 39396 35710
rect 39004 35026 39060 35644
rect 39340 35606 39396 35644
rect 39004 34974 39006 35026
rect 39058 34974 39060 35026
rect 39004 34962 39060 34974
rect 39116 34914 39172 34926
rect 39116 34862 39118 34914
rect 39170 34862 39172 34914
rect 39116 34804 39172 34862
rect 39116 34738 39172 34748
rect 39452 34580 39508 35756
rect 39564 35746 39620 35756
rect 39900 35140 39956 40574
rect 39900 35074 39956 35084
rect 39116 34524 39508 34580
rect 38668 34354 39060 34356
rect 38668 34302 38670 34354
rect 38722 34302 39060 34354
rect 38668 34300 39060 34302
rect 37100 34290 37156 34300
rect 38668 34290 38724 34300
rect 36484 34076 36596 34132
rect 36428 34066 36484 34076
rect 38220 34018 38276 34030
rect 38220 33966 38222 34018
rect 38274 33966 38276 34018
rect 38220 33572 38276 33966
rect 38444 33572 38500 33582
rect 38220 33516 38444 33572
rect 35868 33058 35924 33068
rect 35768 32956 36448 32966
rect 35824 32900 35872 32956
rect 35928 32954 35976 32956
rect 36032 32954 36080 32956
rect 35948 32902 35976 32954
rect 36072 32902 36080 32954
rect 35928 32900 35976 32902
rect 36032 32900 36080 32902
rect 36136 32954 36184 32956
rect 36240 32954 36288 32956
rect 36136 32902 36144 32954
rect 36240 32902 36268 32954
rect 36136 32900 36184 32902
rect 36240 32900 36288 32902
rect 36344 32900 36392 32956
rect 35768 32890 36448 32900
rect 35980 32676 36036 32686
rect 35980 32582 36036 32620
rect 35868 32564 35924 32574
rect 35644 32562 35924 32564
rect 35644 32510 35870 32562
rect 35922 32510 35924 32562
rect 35644 32508 35924 32510
rect 35868 31892 35924 32508
rect 36204 32564 36260 32574
rect 36204 32562 36932 32564
rect 36204 32510 36206 32562
rect 36258 32510 36932 32562
rect 36204 32508 36932 32510
rect 36204 32498 36260 32508
rect 35868 31836 36820 31892
rect 36204 31778 36260 31836
rect 36204 31726 36206 31778
rect 36258 31726 36260 31778
rect 36204 31714 36260 31726
rect 35868 31668 35924 31678
rect 35868 31574 35924 31612
rect 36316 31668 36372 31678
rect 36316 31574 36372 31612
rect 36540 31668 36596 31678
rect 36540 31574 36596 31612
rect 35768 31388 36448 31398
rect 35824 31332 35872 31388
rect 35928 31386 35976 31388
rect 36032 31386 36080 31388
rect 35948 31334 35976 31386
rect 36072 31334 36080 31386
rect 35928 31332 35976 31334
rect 36032 31332 36080 31334
rect 36136 31386 36184 31388
rect 36240 31386 36288 31388
rect 36136 31334 36144 31386
rect 36240 31334 36268 31386
rect 36136 31332 36184 31334
rect 36240 31332 36288 31334
rect 36344 31332 36392 31388
rect 35768 31322 36448 31332
rect 35868 31106 35924 31118
rect 35868 31054 35870 31106
rect 35922 31054 35924 31106
rect 33516 30996 33572 31006
rect 33516 30902 33572 30940
rect 35868 30212 35924 31054
rect 35868 30146 35924 30156
rect 36652 30770 36708 30782
rect 36652 30718 36654 30770
rect 36706 30718 36708 30770
rect 35768 29820 36448 29830
rect 35824 29764 35872 29820
rect 35928 29818 35976 29820
rect 36032 29818 36080 29820
rect 35948 29766 35976 29818
rect 36072 29766 36080 29818
rect 35928 29764 35976 29766
rect 36032 29764 36080 29766
rect 36136 29818 36184 29820
rect 36240 29818 36288 29820
rect 36136 29766 36144 29818
rect 36240 29766 36268 29818
rect 36136 29764 36184 29766
rect 36240 29764 36288 29766
rect 36344 29764 36392 29820
rect 35768 29754 36448 29764
rect 36652 29652 36708 30718
rect 36764 30212 36820 31836
rect 36876 31220 36932 32508
rect 38444 32450 38500 33516
rect 38444 32398 38446 32450
rect 38498 32398 38500 32450
rect 38444 31556 38500 32398
rect 38556 33122 38612 33134
rect 38556 33070 38558 33122
rect 38610 33070 38612 33122
rect 38556 32340 38612 33070
rect 38780 32788 38836 34300
rect 39004 34130 39060 34300
rect 39004 34078 39006 34130
rect 39058 34078 39060 34130
rect 39004 34066 39060 34078
rect 39116 33908 39172 34524
rect 39564 34468 39620 34478
rect 39564 34354 39620 34412
rect 40012 34356 40068 44942
rect 40124 34468 40180 50372
rect 40348 50034 40404 50764
rect 40908 50764 41076 50820
rect 40796 50596 40852 50606
rect 40796 50502 40852 50540
rect 40460 50484 40516 50494
rect 40460 50390 40516 50428
rect 40348 49982 40350 50034
rect 40402 49982 40404 50034
rect 40348 49970 40404 49982
rect 40908 49588 40964 50764
rect 41132 49924 41188 51660
rect 41580 51492 41636 52332
rect 41580 51426 41636 51436
rect 41692 52500 41748 52510
rect 41692 51490 41748 52444
rect 41916 52386 41972 53004
rect 42700 52948 42756 55132
rect 42924 55122 42980 55132
rect 43260 55186 43316 56028
rect 43932 56018 43988 56028
rect 44380 55970 44436 56590
rect 56028 56642 56084 59200
rect 56028 56590 56030 56642
rect 56082 56590 56084 56642
rect 56028 56578 56084 56590
rect 57036 56642 57092 56654
rect 57036 56590 57038 56642
rect 57090 56590 57092 56642
rect 44768 56476 45448 56486
rect 44824 56420 44872 56476
rect 44928 56474 44976 56476
rect 45032 56474 45080 56476
rect 44948 56422 44976 56474
rect 45072 56422 45080 56474
rect 44928 56420 44976 56422
rect 45032 56420 45080 56422
rect 45136 56474 45184 56476
rect 45240 56474 45288 56476
rect 45136 56422 45144 56474
rect 45240 56422 45268 56474
rect 45136 56420 45184 56422
rect 45240 56420 45288 56422
rect 45344 56420 45392 56476
rect 44768 56410 45448 56420
rect 53768 56476 54448 56486
rect 53824 56420 53872 56476
rect 53928 56474 53976 56476
rect 54032 56474 54080 56476
rect 53948 56422 53976 56474
rect 54072 56422 54080 56474
rect 53928 56420 53976 56422
rect 54032 56420 54080 56422
rect 54136 56474 54184 56476
rect 54240 56474 54288 56476
rect 54136 56422 54144 56474
rect 54240 56422 54268 56474
rect 54136 56420 54184 56422
rect 54240 56420 54288 56422
rect 54344 56420 54392 56476
rect 53768 56410 54448 56420
rect 57036 56306 57092 56590
rect 62768 56476 63448 56486
rect 62824 56420 62872 56476
rect 62928 56474 62976 56476
rect 63032 56474 63080 56476
rect 62948 56422 62976 56474
rect 63072 56422 63080 56474
rect 62928 56420 62976 56422
rect 63032 56420 63080 56422
rect 63136 56474 63184 56476
rect 63240 56474 63288 56476
rect 63136 56422 63144 56474
rect 63240 56422 63268 56474
rect 63136 56420 63184 56422
rect 63240 56420 63288 56422
rect 63344 56420 63392 56476
rect 62768 56410 63448 56420
rect 57036 56254 57038 56306
rect 57090 56254 57092 56306
rect 57036 56242 57092 56254
rect 68348 56308 68404 59200
rect 80668 56642 80724 59200
rect 80668 56590 80670 56642
rect 80722 56590 80724 56642
rect 80668 56578 80724 56590
rect 82236 56642 82292 56654
rect 82236 56590 82238 56642
rect 82290 56590 82292 56642
rect 71768 56476 72448 56486
rect 71824 56420 71872 56476
rect 71928 56474 71976 56476
rect 72032 56474 72080 56476
rect 71948 56422 71976 56474
rect 72072 56422 72080 56474
rect 71928 56420 71976 56422
rect 72032 56420 72080 56422
rect 72136 56474 72184 56476
rect 72240 56474 72288 56476
rect 72136 56422 72144 56474
rect 72240 56422 72268 56474
rect 72136 56420 72184 56422
rect 72240 56420 72288 56422
rect 72344 56420 72392 56476
rect 71768 56410 72448 56420
rect 80768 56476 81448 56486
rect 80824 56420 80872 56476
rect 80928 56474 80976 56476
rect 81032 56474 81080 56476
rect 80948 56422 80976 56474
rect 81072 56422 81080 56474
rect 80928 56420 80976 56422
rect 81032 56420 81080 56422
rect 81136 56474 81184 56476
rect 81240 56474 81288 56476
rect 81136 56422 81144 56474
rect 81240 56422 81268 56474
rect 81136 56420 81184 56422
rect 81240 56420 81288 56422
rect 81344 56420 81392 56476
rect 80768 56410 81448 56420
rect 68348 56242 68404 56252
rect 69020 56308 69076 56318
rect 44380 55918 44382 55970
rect 44434 55918 44436 55970
rect 44380 55906 44436 55918
rect 56252 56082 56308 56094
rect 56252 56030 56254 56082
rect 56306 56030 56308 56082
rect 49268 55692 49948 55702
rect 49324 55636 49372 55692
rect 49428 55690 49476 55692
rect 49532 55690 49580 55692
rect 49448 55638 49476 55690
rect 49572 55638 49580 55690
rect 49428 55636 49476 55638
rect 49532 55636 49580 55638
rect 49636 55690 49684 55692
rect 49740 55690 49788 55692
rect 49636 55638 49644 55690
rect 49740 55638 49768 55690
rect 49636 55636 49684 55638
rect 49740 55636 49788 55638
rect 49844 55636 49892 55692
rect 49268 55626 49948 55636
rect 56252 55468 56308 56030
rect 67116 56084 67172 56094
rect 58268 55692 58948 55702
rect 58324 55636 58372 55692
rect 58428 55690 58476 55692
rect 58532 55690 58580 55692
rect 58448 55638 58476 55690
rect 58572 55638 58580 55690
rect 58428 55636 58476 55638
rect 58532 55636 58580 55638
rect 58636 55690 58684 55692
rect 58740 55690 58788 55692
rect 58636 55638 58644 55690
rect 58740 55638 58768 55690
rect 58636 55636 58684 55638
rect 58740 55636 58788 55638
rect 58844 55636 58892 55692
rect 58268 55626 58948 55636
rect 48076 55410 48132 55422
rect 48076 55358 48078 55410
rect 48130 55358 48132 55410
rect 43260 55134 43262 55186
rect 43314 55134 43316 55186
rect 43260 55122 43316 55134
rect 43596 55300 43652 55310
rect 43260 54514 43316 54526
rect 43260 54462 43262 54514
rect 43314 54462 43316 54514
rect 43260 54404 43316 54462
rect 43260 54180 43316 54348
rect 43260 54114 43316 54124
rect 41916 52334 41918 52386
rect 41970 52334 41972 52386
rect 41916 52322 41972 52334
rect 42028 52724 42084 52734
rect 41692 51438 41694 51490
rect 41746 51438 41748 51490
rect 41244 51380 41300 51390
rect 41468 51380 41524 51390
rect 41244 51378 41524 51380
rect 41244 51326 41246 51378
rect 41298 51326 41470 51378
rect 41522 51326 41524 51378
rect 41244 51324 41524 51326
rect 41244 51314 41300 51324
rect 41468 51314 41524 51324
rect 41692 51380 41748 51438
rect 41692 51314 41748 51324
rect 42028 52164 42084 52668
rect 42028 51378 42084 52108
rect 42700 51602 42756 52892
rect 42700 51550 42702 51602
rect 42754 51550 42756 51602
rect 42700 51538 42756 51550
rect 43260 52164 43316 52174
rect 43260 51602 43316 52108
rect 43260 51550 43262 51602
rect 43314 51550 43316 51602
rect 43260 51538 43316 51550
rect 42028 51326 42030 51378
rect 42082 51326 42084 51378
rect 42028 51314 42084 51326
rect 42252 51380 42308 51390
rect 42252 51286 42308 51324
rect 42812 51266 42868 51278
rect 42812 51214 42814 51266
rect 42866 51214 42868 51266
rect 41580 51156 41636 51166
rect 41244 51154 41636 51156
rect 41244 51102 41582 51154
rect 41634 51102 41636 51154
rect 41244 51100 41636 51102
rect 41244 50594 41300 51100
rect 41580 51090 41636 51100
rect 41244 50542 41246 50594
rect 41298 50542 41300 50594
rect 41244 50530 41300 50542
rect 41132 49858 41188 49868
rect 42364 49812 42420 49822
rect 42812 49812 42868 51214
rect 43596 50820 43652 55244
rect 43708 55300 43764 55310
rect 43708 55206 43764 55244
rect 44268 55300 44324 55310
rect 44268 55206 44324 55244
rect 45164 55300 45220 55310
rect 45164 55206 45220 55244
rect 45948 55188 46004 55198
rect 45948 55094 46004 55132
rect 44768 54908 45448 54918
rect 44824 54852 44872 54908
rect 44928 54906 44976 54908
rect 45032 54906 45080 54908
rect 44948 54854 44976 54906
rect 45072 54854 45080 54906
rect 44928 54852 44976 54854
rect 45032 54852 45080 54854
rect 45136 54906 45184 54908
rect 45240 54906 45288 54908
rect 45136 54854 45144 54906
rect 45240 54854 45268 54906
rect 45136 54852 45184 54854
rect 45240 54852 45288 54854
rect 45344 54852 45392 54908
rect 44768 54842 45448 54852
rect 47740 54740 47796 54750
rect 44156 54628 44212 54638
rect 44156 54404 44212 54572
rect 44604 54628 44660 54638
rect 44604 54534 44660 54572
rect 47740 54626 47796 54684
rect 47740 54574 47742 54626
rect 47794 54574 47796 54626
rect 47740 54562 47796 54574
rect 47964 54628 48020 54638
rect 48076 54628 48132 55358
rect 56028 55412 56308 55468
rect 55804 55298 55860 55310
rect 55804 55246 55806 55298
rect 55858 55246 55860 55298
rect 48860 55188 48916 55198
rect 48020 54572 48132 54628
rect 48636 55074 48692 55086
rect 48636 55022 48638 55074
rect 48690 55022 48692 55074
rect 47964 54534 48020 54572
rect 44156 54310 44212 54348
rect 44828 54514 44884 54526
rect 44828 54462 44830 54514
rect 44882 54462 44884 54514
rect 44828 54180 44884 54462
rect 45164 54514 45220 54526
rect 45164 54462 45166 54514
rect 45218 54462 45220 54514
rect 45164 54404 45220 54462
rect 47292 54514 47348 54526
rect 47292 54462 47294 54514
rect 47346 54462 47348 54514
rect 45500 54404 45556 54414
rect 45164 54402 45556 54404
rect 45164 54350 45502 54402
rect 45554 54350 45556 54402
rect 45164 54348 45556 54350
rect 44940 54292 44996 54302
rect 44940 54198 44996 54236
rect 44828 53732 44884 54124
rect 44940 53732 44996 53742
rect 44828 53676 44940 53732
rect 44940 53638 44996 53676
rect 43820 53508 43876 53518
rect 43708 53506 43876 53508
rect 43708 53454 43822 53506
rect 43874 53454 43876 53506
rect 43708 53452 43876 53454
rect 43708 52164 43764 53452
rect 43820 53442 43876 53452
rect 44268 53506 44324 53518
rect 44268 53454 44270 53506
rect 44322 53454 44324 53506
rect 43708 52098 43764 52108
rect 43820 53060 43876 53070
rect 43820 52162 43876 53004
rect 43820 52110 43822 52162
rect 43874 52110 43876 52162
rect 43820 52098 43876 52110
rect 43932 52500 43988 52510
rect 44268 52500 44324 53454
rect 45500 53508 45556 54348
rect 45948 54402 46004 54414
rect 45948 54350 45950 54402
rect 46002 54350 46004 54402
rect 45948 53732 46004 54350
rect 47068 54290 47124 54302
rect 47068 54238 47070 54290
rect 47122 54238 47124 54290
rect 46732 53956 46788 53966
rect 45948 53666 46004 53676
rect 46060 53730 46116 53742
rect 46060 53678 46062 53730
rect 46114 53678 46116 53730
rect 45500 53452 45780 53508
rect 44768 53340 45448 53350
rect 44824 53284 44872 53340
rect 44928 53338 44976 53340
rect 45032 53338 45080 53340
rect 44948 53286 44976 53338
rect 45072 53286 45080 53338
rect 44928 53284 44976 53286
rect 45032 53284 45080 53286
rect 45136 53338 45184 53340
rect 45240 53338 45288 53340
rect 45136 53286 45144 53338
rect 45240 53286 45268 53338
rect 45136 53284 45184 53286
rect 45240 53284 45288 53286
rect 45344 53284 45392 53340
rect 44768 53274 45448 53284
rect 45500 53060 45556 53070
rect 45500 52966 45556 53004
rect 44716 52612 44772 52622
rect 43988 52444 44324 52500
rect 44604 52556 44716 52612
rect 43708 51604 43764 51614
rect 43932 51604 43988 52444
rect 43708 51602 43988 51604
rect 43708 51550 43710 51602
rect 43762 51550 43988 51602
rect 43708 51548 43988 51550
rect 44604 51604 44660 52556
rect 44716 52546 44772 52556
rect 45612 52612 45668 52622
rect 45724 52612 45780 53452
rect 46060 53060 46116 53678
rect 46060 52994 46116 53004
rect 45668 52556 45780 52612
rect 46620 52946 46676 52958
rect 46620 52894 46622 52946
rect 46674 52894 46676 52946
rect 45612 52274 45668 52556
rect 45612 52222 45614 52274
rect 45666 52222 45668 52274
rect 45612 52210 45668 52222
rect 46172 52500 46228 52510
rect 45948 52164 46004 52174
rect 45948 52070 46004 52108
rect 46172 52162 46228 52444
rect 46172 52110 46174 52162
rect 46226 52110 46228 52162
rect 46172 52098 46228 52110
rect 46620 52164 46676 52894
rect 46396 52052 46452 52062
rect 46172 51940 46228 51950
rect 44768 51772 45448 51782
rect 44824 51716 44872 51772
rect 44928 51770 44976 51772
rect 45032 51770 45080 51772
rect 44948 51718 44976 51770
rect 45072 51718 45080 51770
rect 44928 51716 44976 51718
rect 45032 51716 45080 51718
rect 45136 51770 45184 51772
rect 45240 51770 45288 51772
rect 45136 51718 45144 51770
rect 45240 51718 45268 51770
rect 45136 51716 45184 51718
rect 45240 51716 45288 51718
rect 45344 51716 45392 51772
rect 44768 51706 45448 51716
rect 44716 51604 44772 51614
rect 44660 51602 44772 51604
rect 44660 51550 44718 51602
rect 44770 51550 44772 51602
rect 44660 51548 44772 51550
rect 43708 51538 43764 51548
rect 44604 51510 44660 51548
rect 44716 51538 44772 51548
rect 43596 50754 43652 50764
rect 44268 51378 44324 51390
rect 44268 51326 44270 51378
rect 44322 51326 44324 51378
rect 44268 50818 44324 51326
rect 46172 51378 46228 51884
rect 46172 51326 46174 51378
rect 46226 51326 46228 51378
rect 46172 51314 46228 51326
rect 46396 51380 46452 51996
rect 46396 51286 46452 51324
rect 44268 50766 44270 50818
rect 44322 50766 44324 50818
rect 44268 50754 44324 50766
rect 45500 50596 45556 50606
rect 45500 50502 45556 50540
rect 46172 50596 46228 50606
rect 46172 50502 46228 50540
rect 43596 50484 43652 50494
rect 43596 50370 43652 50428
rect 46060 50484 46116 50494
rect 46060 50390 46116 50428
rect 43596 50318 43598 50370
rect 43650 50318 43652 50370
rect 43596 50306 43652 50318
rect 44768 50204 45448 50214
rect 44824 50148 44872 50204
rect 44928 50202 44976 50204
rect 45032 50202 45080 50204
rect 44948 50150 44976 50202
rect 45072 50150 45080 50202
rect 44928 50148 44976 50150
rect 45032 50148 45080 50150
rect 45136 50202 45184 50204
rect 45240 50202 45288 50204
rect 45136 50150 45144 50202
rect 45240 50150 45268 50202
rect 45136 50148 45184 50150
rect 45240 50148 45288 50150
rect 45344 50148 45392 50204
rect 44768 50138 45448 50148
rect 42364 49810 42868 49812
rect 42364 49758 42366 49810
rect 42418 49758 42868 49810
rect 42364 49756 42868 49758
rect 42364 49746 42420 49756
rect 42252 49700 42308 49710
rect 40908 49532 41188 49588
rect 40268 49420 40948 49430
rect 40324 49364 40372 49420
rect 40428 49418 40476 49420
rect 40532 49418 40580 49420
rect 40448 49366 40476 49418
rect 40572 49366 40580 49418
rect 40428 49364 40476 49366
rect 40532 49364 40580 49366
rect 40636 49418 40684 49420
rect 40740 49418 40788 49420
rect 40636 49366 40644 49418
rect 40740 49366 40768 49418
rect 40636 49364 40684 49366
rect 40740 49364 40788 49366
rect 40844 49364 40892 49420
rect 40268 49354 40948 49364
rect 41020 48468 41076 48478
rect 40460 48020 40516 48058
rect 40460 47954 40516 47964
rect 40268 47852 40948 47862
rect 40324 47796 40372 47852
rect 40428 47850 40476 47852
rect 40532 47850 40580 47852
rect 40448 47798 40476 47850
rect 40572 47798 40580 47850
rect 40428 47796 40476 47798
rect 40532 47796 40580 47798
rect 40636 47850 40684 47852
rect 40740 47850 40788 47852
rect 40636 47798 40644 47850
rect 40740 47798 40768 47850
rect 40636 47796 40684 47798
rect 40740 47796 40788 47798
rect 40844 47796 40892 47852
rect 40268 47786 40948 47796
rect 41020 47124 41076 48412
rect 41020 47058 41076 47068
rect 40236 46674 40292 46686
rect 40236 46622 40238 46674
rect 40290 46622 40292 46674
rect 40236 46564 40292 46622
rect 40236 46498 40292 46508
rect 41020 46564 41076 46574
rect 41020 46470 41076 46508
rect 40268 46284 40948 46294
rect 40324 46228 40372 46284
rect 40428 46282 40476 46284
rect 40532 46282 40580 46284
rect 40448 46230 40476 46282
rect 40572 46230 40580 46282
rect 40428 46228 40476 46230
rect 40532 46228 40580 46230
rect 40636 46282 40684 46284
rect 40740 46282 40788 46284
rect 40636 46230 40644 46282
rect 40740 46230 40768 46282
rect 40636 46228 40684 46230
rect 40740 46228 40788 46230
rect 40844 46228 40892 46284
rect 40268 46218 40948 46228
rect 40684 45892 40740 45902
rect 40684 45798 40740 45836
rect 40236 45780 40292 45790
rect 40236 45686 40292 45724
rect 41020 45780 41076 45790
rect 41020 45330 41076 45724
rect 41020 45278 41022 45330
rect 41074 45278 41076 45330
rect 41020 45266 41076 45278
rect 40268 44716 40948 44726
rect 40324 44660 40372 44716
rect 40428 44714 40476 44716
rect 40532 44714 40580 44716
rect 40448 44662 40476 44714
rect 40572 44662 40580 44714
rect 40428 44660 40476 44662
rect 40532 44660 40580 44662
rect 40636 44714 40684 44716
rect 40740 44714 40788 44716
rect 40636 44662 40644 44714
rect 40740 44662 40768 44714
rect 40636 44660 40684 44662
rect 40740 44660 40788 44662
rect 40844 44660 40892 44716
rect 40268 44650 40948 44660
rect 40908 44212 40964 44222
rect 40908 44098 40964 44156
rect 40908 44046 40910 44098
rect 40962 44046 40964 44098
rect 40908 44034 40964 44046
rect 40268 43148 40948 43158
rect 40324 43092 40372 43148
rect 40428 43146 40476 43148
rect 40532 43146 40580 43148
rect 40448 43094 40476 43146
rect 40572 43094 40580 43146
rect 40428 43092 40476 43094
rect 40532 43092 40580 43094
rect 40636 43146 40684 43148
rect 40740 43146 40788 43148
rect 40636 43094 40644 43146
rect 40740 43094 40768 43146
rect 40636 43092 40684 43094
rect 40740 43092 40788 43094
rect 40844 43092 40892 43148
rect 40268 43082 40948 43092
rect 41020 41972 41076 41982
rect 40268 41580 40948 41590
rect 40324 41524 40372 41580
rect 40428 41578 40476 41580
rect 40532 41578 40580 41580
rect 40448 41526 40476 41578
rect 40572 41526 40580 41578
rect 40428 41524 40476 41526
rect 40532 41524 40580 41526
rect 40636 41578 40684 41580
rect 40740 41578 40788 41580
rect 40636 41526 40644 41578
rect 40740 41526 40768 41578
rect 40636 41524 40684 41526
rect 40740 41524 40788 41526
rect 40844 41524 40892 41580
rect 40268 41514 40948 41524
rect 41020 40626 41076 41916
rect 41020 40574 41022 40626
rect 41074 40574 41076 40626
rect 41020 40562 41076 40574
rect 40348 40292 40404 40302
rect 40348 40198 40404 40236
rect 40268 40012 40948 40022
rect 40324 39956 40372 40012
rect 40428 40010 40476 40012
rect 40532 40010 40580 40012
rect 40448 39958 40476 40010
rect 40572 39958 40580 40010
rect 40428 39956 40476 39958
rect 40532 39956 40580 39958
rect 40636 40010 40684 40012
rect 40740 40010 40788 40012
rect 40636 39958 40644 40010
rect 40740 39958 40768 40010
rect 40636 39956 40684 39958
rect 40740 39956 40788 39958
rect 40844 39956 40892 40012
rect 40268 39946 40948 39956
rect 40268 38444 40948 38454
rect 40324 38388 40372 38444
rect 40428 38442 40476 38444
rect 40532 38442 40580 38444
rect 40448 38390 40476 38442
rect 40572 38390 40580 38442
rect 40428 38388 40476 38390
rect 40532 38388 40580 38390
rect 40636 38442 40684 38444
rect 40740 38442 40788 38444
rect 40636 38390 40644 38442
rect 40740 38390 40768 38442
rect 40636 38388 40684 38390
rect 40740 38388 40788 38390
rect 40844 38388 40892 38444
rect 40268 38378 40948 38388
rect 40460 37604 40516 37614
rect 40460 37490 40516 37548
rect 40460 37438 40462 37490
rect 40514 37438 40516 37490
rect 40460 37426 40516 37438
rect 41020 37268 41076 37278
rect 41020 37174 41076 37212
rect 40268 36876 40948 36886
rect 40324 36820 40372 36876
rect 40428 36874 40476 36876
rect 40532 36874 40580 36876
rect 40448 36822 40476 36874
rect 40572 36822 40580 36874
rect 40428 36820 40476 36822
rect 40532 36820 40580 36822
rect 40636 36874 40684 36876
rect 40740 36874 40788 36876
rect 40636 36822 40644 36874
rect 40740 36822 40768 36874
rect 40636 36820 40684 36822
rect 40740 36820 40788 36822
rect 40844 36820 40892 36876
rect 40268 36810 40948 36820
rect 40268 35308 40948 35318
rect 40324 35252 40372 35308
rect 40428 35306 40476 35308
rect 40532 35306 40580 35308
rect 40448 35254 40476 35306
rect 40572 35254 40580 35306
rect 40428 35252 40476 35254
rect 40532 35252 40580 35254
rect 40636 35306 40684 35308
rect 40740 35306 40788 35308
rect 40636 35254 40644 35306
rect 40740 35254 40768 35306
rect 40636 35252 40684 35254
rect 40740 35252 40788 35254
rect 40844 35252 40892 35308
rect 40268 35242 40948 35252
rect 40796 35028 40852 35038
rect 40796 34802 40852 34972
rect 40796 34750 40798 34802
rect 40850 34750 40852 34802
rect 40796 34738 40852 34750
rect 40124 34402 40180 34412
rect 41020 34356 41076 34366
rect 41132 34356 41188 49532
rect 41804 47124 41860 47134
rect 41580 46564 41636 46574
rect 41356 45108 41412 45118
rect 41412 45052 41524 45108
rect 41356 45014 41412 45052
rect 41468 44546 41524 45052
rect 41468 44494 41470 44546
rect 41522 44494 41524 44546
rect 41468 44482 41524 44494
rect 41468 41300 41524 41310
rect 41468 40962 41524 41244
rect 41468 40910 41470 40962
rect 41522 40910 41524 40962
rect 41468 40898 41524 40910
rect 41580 40516 41636 46508
rect 41804 44434 41860 47068
rect 41916 45892 41972 45902
rect 41916 45332 41972 45836
rect 41916 45220 41972 45276
rect 42028 45220 42084 45230
rect 41916 45218 42084 45220
rect 41916 45166 42030 45218
rect 42082 45166 42084 45218
rect 41916 45164 42084 45166
rect 42028 45154 42084 45164
rect 42140 45106 42196 45118
rect 42140 45054 42142 45106
rect 42194 45054 42196 45106
rect 42140 44996 42196 45054
rect 42140 44930 42196 44940
rect 41804 44382 41806 44434
rect 41858 44382 41860 44434
rect 41804 44212 41860 44382
rect 41804 44146 41860 44156
rect 42140 41300 42196 41310
rect 41580 40422 41636 40460
rect 42028 41076 42084 41086
rect 42028 40514 42084 41020
rect 42028 40462 42030 40514
rect 42082 40462 42084 40514
rect 42028 40450 42084 40462
rect 41244 40292 41300 40302
rect 41300 40236 41412 40292
rect 41244 38612 41300 40236
rect 41356 40178 41412 40236
rect 41356 40126 41358 40178
rect 41410 40126 41412 40178
rect 41356 40114 41412 40126
rect 42140 39058 42196 41244
rect 42140 39006 42142 39058
rect 42194 39006 42196 39058
rect 42140 38668 42196 39006
rect 41244 37604 41300 38556
rect 41916 38612 42196 38668
rect 41244 37538 41300 37548
rect 41356 38276 41412 38286
rect 41356 37266 41412 38220
rect 41468 37828 41524 37838
rect 41468 37734 41524 37772
rect 41916 37828 41972 38612
rect 42028 38276 42084 38286
rect 42252 38276 42308 49644
rect 42812 49588 42868 49756
rect 42812 49522 42868 49532
rect 44768 48636 45448 48646
rect 44824 48580 44872 48636
rect 44928 48634 44976 48636
rect 45032 48634 45080 48636
rect 44948 48582 44976 48634
rect 45072 48582 45080 48634
rect 44928 48580 44976 48582
rect 45032 48580 45080 48582
rect 45136 48634 45184 48636
rect 45240 48634 45288 48636
rect 45136 48582 45144 48634
rect 45240 48582 45268 48634
rect 45136 48580 45184 48582
rect 45240 48580 45288 48582
rect 45344 48580 45392 48636
rect 44768 48570 45448 48580
rect 43484 48354 43540 48366
rect 43484 48302 43486 48354
rect 43538 48302 43540 48354
rect 43260 47460 43316 47470
rect 43260 47366 43316 47404
rect 42812 47012 42868 47022
rect 42868 46956 43092 47012
rect 42812 46946 42868 46956
rect 43036 46898 43092 46956
rect 43036 46846 43038 46898
rect 43090 46846 43092 46898
rect 43036 46834 43092 46846
rect 43484 46674 43540 48302
rect 43932 48354 43988 48366
rect 43932 48302 43934 48354
rect 43986 48302 43988 48354
rect 43484 46622 43486 46674
rect 43538 46622 43540 46674
rect 43484 46610 43540 46622
rect 43708 47460 43764 47470
rect 43708 47234 43764 47404
rect 43708 47182 43710 47234
rect 43762 47182 43764 47234
rect 43596 45220 43652 45230
rect 42700 44996 42756 45006
rect 42756 44940 42868 44996
rect 42700 44902 42756 44940
rect 42364 44212 42420 44222
rect 42364 41972 42420 44156
rect 42364 41300 42420 41916
rect 42364 41206 42420 41244
rect 42700 40516 42756 40526
rect 42588 39396 42644 39406
rect 42588 38946 42644 39340
rect 42588 38894 42590 38946
rect 42642 38894 42644 38946
rect 42588 38668 42644 38894
rect 42028 38182 42084 38220
rect 42140 38220 42308 38276
rect 42364 38612 42644 38668
rect 41916 37762 41972 37772
rect 41916 37604 41972 37614
rect 41356 37214 41358 37266
rect 41410 37214 41412 37266
rect 41356 37202 41412 37214
rect 41692 37380 41748 37390
rect 41692 37044 41748 37324
rect 41916 37378 41972 37548
rect 41916 37326 41918 37378
rect 41970 37326 41972 37378
rect 41916 37314 41972 37326
rect 42028 37268 42084 37278
rect 42028 37174 42084 37212
rect 41692 36978 41748 36988
rect 39564 34302 39566 34354
rect 39618 34302 39620 34354
rect 39564 34290 39620 34302
rect 39676 34300 40068 34356
rect 40236 34354 41188 34356
rect 40236 34302 41022 34354
rect 41074 34302 41188 34354
rect 40236 34300 41188 34302
rect 41244 34916 41300 34926
rect 41244 34690 41300 34860
rect 41244 34638 41246 34690
rect 41298 34638 41300 34690
rect 39340 34132 39396 34142
rect 38892 33852 39172 33908
rect 39228 34130 39396 34132
rect 39228 34078 39342 34130
rect 39394 34078 39396 34130
rect 39228 34076 39396 34078
rect 38892 33346 38948 33852
rect 38892 33294 38894 33346
rect 38946 33294 38948 33346
rect 38892 33282 38948 33294
rect 39228 33572 39284 34076
rect 39340 34066 39396 34076
rect 38892 32788 38948 32798
rect 38780 32786 38948 32788
rect 38780 32734 38894 32786
rect 38946 32734 38948 32786
rect 38780 32732 38948 32734
rect 38556 32274 38612 32284
rect 38892 32452 38948 32732
rect 39228 32674 39284 33516
rect 39452 34018 39508 34030
rect 39452 33966 39454 34018
rect 39506 33966 39508 34018
rect 39340 33348 39396 33358
rect 39452 33348 39508 33966
rect 39340 33346 39508 33348
rect 39340 33294 39342 33346
rect 39394 33294 39508 33346
rect 39340 33292 39508 33294
rect 39340 33282 39396 33292
rect 39676 32788 39732 34300
rect 40236 34242 40292 34300
rect 40236 34190 40238 34242
rect 40290 34190 40292 34242
rect 40236 34178 40292 34190
rect 39788 34132 39844 34142
rect 40124 34132 40180 34142
rect 39788 34130 40180 34132
rect 39788 34078 39790 34130
rect 39842 34078 40126 34130
rect 40178 34078 40180 34130
rect 39788 34076 40180 34078
rect 39788 34066 39844 34076
rect 40124 34066 40180 34076
rect 40268 33740 40948 33750
rect 40324 33684 40372 33740
rect 40428 33738 40476 33740
rect 40532 33738 40580 33740
rect 40448 33686 40476 33738
rect 40572 33686 40580 33738
rect 40428 33684 40476 33686
rect 40532 33684 40580 33686
rect 40636 33738 40684 33740
rect 40740 33738 40788 33740
rect 40636 33686 40644 33738
rect 40740 33686 40768 33738
rect 40636 33684 40684 33686
rect 40740 33684 40788 33686
rect 40844 33684 40892 33740
rect 40268 33674 40948 33684
rect 39228 32622 39230 32674
rect 39282 32622 39284 32674
rect 39228 32610 39284 32622
rect 39564 32732 39732 32788
rect 39900 32788 39956 32798
rect 39340 32562 39396 32574
rect 39340 32510 39342 32562
rect 39394 32510 39396 32562
rect 39340 32452 39396 32510
rect 38892 32396 39396 32452
rect 38892 31890 38948 32396
rect 38892 31838 38894 31890
rect 38946 31838 38948 31890
rect 38892 31826 38948 31838
rect 39228 31778 39284 32396
rect 39228 31726 39230 31778
rect 39282 31726 39284 31778
rect 38892 31556 38948 31566
rect 38444 31554 38612 31556
rect 38444 31502 38446 31554
rect 38498 31502 38612 31554
rect 38444 31500 38612 31502
rect 38444 31490 38500 31500
rect 36876 31154 36932 31164
rect 37100 30772 37156 30782
rect 36988 30212 37044 30222
rect 36764 30156 36988 30212
rect 36652 29586 36708 29596
rect 36988 30098 37044 30156
rect 36988 30046 36990 30098
rect 37042 30046 37044 30098
rect 35420 28420 35476 28430
rect 35308 28418 35476 28420
rect 35308 28366 35422 28418
rect 35474 28366 35476 28418
rect 35308 28364 35476 28366
rect 34860 27972 34916 27982
rect 34860 27878 34916 27916
rect 35196 27972 35252 27982
rect 33292 26852 33460 26908
rect 35196 26964 35252 27916
rect 35308 27858 35364 28364
rect 35420 28354 35476 28364
rect 35768 28252 36448 28262
rect 35824 28196 35872 28252
rect 35928 28250 35976 28252
rect 36032 28250 36080 28252
rect 35948 28198 35976 28250
rect 36072 28198 36080 28250
rect 35928 28196 35976 28198
rect 36032 28196 36080 28198
rect 36136 28250 36184 28252
rect 36240 28250 36288 28252
rect 36136 28198 36144 28250
rect 36240 28198 36268 28250
rect 36136 28196 36184 28198
rect 36240 28196 36288 28198
rect 36344 28196 36392 28252
rect 35768 28186 36448 28196
rect 35308 27806 35310 27858
rect 35362 27806 35364 27858
rect 35308 27794 35364 27806
rect 35644 27858 35700 27870
rect 35644 27806 35646 27858
rect 35698 27806 35700 27858
rect 29372 24946 29428 26852
rect 31268 25900 31948 25910
rect 31324 25844 31372 25900
rect 31428 25898 31476 25900
rect 31532 25898 31580 25900
rect 31448 25846 31476 25898
rect 31572 25846 31580 25898
rect 31428 25844 31476 25846
rect 31532 25844 31580 25846
rect 31636 25898 31684 25900
rect 31740 25898 31788 25900
rect 31636 25846 31644 25898
rect 31740 25846 31768 25898
rect 31636 25844 31684 25846
rect 31740 25844 31788 25846
rect 31844 25844 31892 25900
rect 31268 25834 31948 25844
rect 33068 25396 33124 25406
rect 33068 25302 33124 25340
rect 30492 25060 30548 25070
rect 29372 24894 29374 24946
rect 29426 24894 29428 24946
rect 29372 24836 29428 24894
rect 30156 24948 30212 24958
rect 30156 24854 30212 24892
rect 29372 23380 29428 24780
rect 30492 24836 30548 25004
rect 32060 25060 32116 25070
rect 32060 24946 32116 25004
rect 32060 24894 32062 24946
rect 32114 24894 32116 24946
rect 32060 24882 32116 24894
rect 30548 24780 30660 24836
rect 30492 24742 30548 24780
rect 29484 23380 29540 23390
rect 29372 23378 29540 23380
rect 29372 23326 29486 23378
rect 29538 23326 29540 23378
rect 29372 23324 29540 23326
rect 29484 23314 29540 23324
rect 30604 23378 30660 24780
rect 32508 24834 32564 24846
rect 32508 24782 32510 24834
rect 32562 24782 32564 24834
rect 32508 24724 32564 24782
rect 32956 24724 33012 24734
rect 32508 24722 33012 24724
rect 32508 24670 32958 24722
rect 33010 24670 33012 24722
rect 32508 24668 33012 24670
rect 32956 24658 33012 24668
rect 31268 24332 31948 24342
rect 31324 24276 31372 24332
rect 31428 24330 31476 24332
rect 31532 24330 31580 24332
rect 31448 24278 31476 24330
rect 31572 24278 31580 24330
rect 31428 24276 31476 24278
rect 31532 24276 31580 24278
rect 31636 24330 31684 24332
rect 31740 24330 31788 24332
rect 31636 24278 31644 24330
rect 31740 24278 31768 24330
rect 31636 24276 31684 24278
rect 31740 24276 31788 24278
rect 31844 24276 31892 24332
rect 31268 24266 31948 24276
rect 32620 23828 32676 23838
rect 32620 23734 32676 23772
rect 33068 23828 33124 23838
rect 33068 23734 33124 23772
rect 30604 23326 30606 23378
rect 30658 23326 30660 23378
rect 30268 22932 30324 22942
rect 30268 22838 30324 22876
rect 29708 22260 29764 22270
rect 29036 21746 29092 21756
rect 29148 22146 29204 22158
rect 29148 22094 29150 22146
rect 29202 22094 29204 22146
rect 29036 21588 29092 21598
rect 29148 21588 29204 22094
rect 29708 22146 29764 22204
rect 29708 22094 29710 22146
rect 29762 22094 29764 22146
rect 29036 21586 29204 21588
rect 29036 21534 29038 21586
rect 29090 21534 29204 21586
rect 29036 21532 29204 21534
rect 29372 21586 29428 21598
rect 29372 21534 29374 21586
rect 29426 21534 29428 21586
rect 29036 21522 29092 21532
rect 28364 21422 28366 21474
rect 28418 21422 28420 21474
rect 28364 21410 28420 21422
rect 29372 21476 29428 21534
rect 29372 21410 29428 21420
rect 29148 21028 29204 21038
rect 29708 21028 29764 22094
rect 30604 21812 30660 23326
rect 32172 23714 32228 23726
rect 32172 23662 32174 23714
rect 32226 23662 32228 23714
rect 32172 23380 32228 23662
rect 32284 23380 32340 23390
rect 32172 23324 32284 23380
rect 32284 23314 32340 23324
rect 32620 23380 32676 23390
rect 31268 22764 31948 22774
rect 31324 22708 31372 22764
rect 31428 22762 31476 22764
rect 31532 22762 31580 22764
rect 31448 22710 31476 22762
rect 31572 22710 31580 22762
rect 31428 22708 31476 22710
rect 31532 22708 31580 22710
rect 31636 22762 31684 22764
rect 31740 22762 31788 22764
rect 31636 22710 31644 22762
rect 31740 22710 31768 22762
rect 31636 22708 31684 22710
rect 31740 22708 31788 22710
rect 31844 22708 31892 22764
rect 31268 22698 31948 22708
rect 30156 21028 30212 21038
rect 29708 20972 30156 21028
rect 28588 20804 28644 20814
rect 29148 20804 29204 20972
rect 30156 20934 30212 20972
rect 28588 20244 28644 20748
rect 28588 20178 28644 20188
rect 28924 20802 29204 20804
rect 28924 20750 29150 20802
rect 29202 20750 29204 20802
rect 28924 20748 29204 20750
rect 28924 20242 28980 20748
rect 29148 20738 29204 20748
rect 28924 20190 28926 20242
rect 28978 20190 28980 20242
rect 28924 20178 28980 20190
rect 28476 20132 28532 20142
rect 28476 20038 28532 20076
rect 29372 20132 29428 20142
rect 29372 20038 29428 20076
rect 30604 20132 30660 21756
rect 31948 21812 32004 21822
rect 31948 21718 32004 21756
rect 32508 21364 32564 21374
rect 32508 21270 32564 21308
rect 31268 21196 31948 21206
rect 31324 21140 31372 21196
rect 31428 21194 31476 21196
rect 31532 21194 31580 21196
rect 31448 21142 31476 21194
rect 31572 21142 31580 21194
rect 31428 21140 31476 21142
rect 31532 21140 31580 21142
rect 31636 21194 31684 21196
rect 31740 21194 31788 21196
rect 31636 21142 31644 21194
rect 31740 21142 31768 21194
rect 31636 21140 31684 21142
rect 31740 21140 31788 21142
rect 31844 21140 31892 21196
rect 31268 21130 31948 21140
rect 32620 20914 32676 23324
rect 32620 20862 32622 20914
rect 32674 20862 32676 20914
rect 32620 20804 32676 20862
rect 33068 21700 33124 21710
rect 33068 20914 33124 21644
rect 33068 20862 33070 20914
rect 33122 20862 33124 20914
rect 33068 20850 33124 20862
rect 32620 20738 32676 20748
rect 30604 20066 30660 20076
rect 31268 19628 31948 19638
rect 31324 19572 31372 19628
rect 31428 19626 31476 19628
rect 31532 19626 31580 19628
rect 31448 19574 31476 19626
rect 31572 19574 31580 19626
rect 31428 19572 31476 19574
rect 31532 19572 31580 19574
rect 31636 19626 31684 19628
rect 31740 19626 31788 19628
rect 31636 19574 31644 19626
rect 31740 19574 31768 19626
rect 31636 19572 31684 19574
rect 31740 19572 31788 19574
rect 31844 19572 31892 19628
rect 31268 19562 31948 19572
rect 31268 18060 31948 18070
rect 31324 18004 31372 18060
rect 31428 18058 31476 18060
rect 31532 18058 31580 18060
rect 31448 18006 31476 18058
rect 31572 18006 31580 18058
rect 31428 18004 31476 18006
rect 31532 18004 31580 18006
rect 31636 18058 31684 18060
rect 31740 18058 31788 18060
rect 31636 18006 31644 18058
rect 31740 18006 31768 18058
rect 31636 18004 31684 18006
rect 31740 18004 31788 18006
rect 31844 18004 31892 18060
rect 31268 17994 31948 18004
rect 31268 16492 31948 16502
rect 31324 16436 31372 16492
rect 31428 16490 31476 16492
rect 31532 16490 31580 16492
rect 31448 16438 31476 16490
rect 31572 16438 31580 16490
rect 31428 16436 31476 16438
rect 31532 16436 31580 16438
rect 31636 16490 31684 16492
rect 31740 16490 31788 16492
rect 31636 16438 31644 16490
rect 31740 16438 31768 16490
rect 31636 16436 31684 16438
rect 31740 16436 31788 16438
rect 31844 16436 31892 16492
rect 31268 16426 31948 16436
rect 31268 14924 31948 14934
rect 31324 14868 31372 14924
rect 31428 14922 31476 14924
rect 31532 14922 31580 14924
rect 31448 14870 31476 14922
rect 31572 14870 31580 14922
rect 31428 14868 31476 14870
rect 31532 14868 31580 14870
rect 31636 14922 31684 14924
rect 31740 14922 31788 14924
rect 31636 14870 31644 14922
rect 31740 14870 31768 14922
rect 31636 14868 31684 14870
rect 31740 14868 31788 14870
rect 31844 14868 31892 14924
rect 31268 14858 31948 14868
rect 31268 13356 31948 13366
rect 31324 13300 31372 13356
rect 31428 13354 31476 13356
rect 31532 13354 31580 13356
rect 31448 13302 31476 13354
rect 31572 13302 31580 13354
rect 31428 13300 31476 13302
rect 31532 13300 31580 13302
rect 31636 13354 31684 13356
rect 31740 13354 31788 13356
rect 31636 13302 31644 13354
rect 31740 13302 31768 13354
rect 31636 13300 31684 13302
rect 31740 13300 31788 13302
rect 31844 13300 31892 13356
rect 31268 13290 31948 13300
rect 33292 12292 33348 26852
rect 34860 25506 34916 25518
rect 35084 25508 35140 25518
rect 34860 25454 34862 25506
rect 34914 25454 34916 25506
rect 34188 25396 34244 25406
rect 33404 25284 33460 25294
rect 34076 25284 34132 25294
rect 33404 25282 33684 25284
rect 33404 25230 33406 25282
rect 33458 25230 33684 25282
rect 33404 25228 33684 25230
rect 33404 25218 33460 25228
rect 33628 24722 33684 25228
rect 34076 25190 34132 25228
rect 33628 24670 33630 24722
rect 33682 24670 33684 24722
rect 33628 24658 33684 24670
rect 33852 24724 33908 24734
rect 33852 24162 33908 24668
rect 33852 24110 33854 24162
rect 33906 24110 33908 24162
rect 33852 24098 33908 24110
rect 34188 24162 34244 25340
rect 34860 25396 34916 25454
rect 34188 24110 34190 24162
rect 34242 24110 34244 24162
rect 34188 24098 34244 24110
rect 34524 25284 34580 25294
rect 34860 25284 34916 25340
rect 34524 25282 34916 25284
rect 34524 25230 34526 25282
rect 34578 25230 34916 25282
rect 34524 25228 34916 25230
rect 34972 25506 35140 25508
rect 34972 25454 35086 25506
rect 35138 25454 35140 25506
rect 34972 25452 35140 25454
rect 34972 25284 35028 25452
rect 35084 25442 35140 25452
rect 33516 23826 33572 23838
rect 33516 23774 33518 23826
rect 33570 23774 33572 23826
rect 33516 23380 33572 23774
rect 33628 23380 33684 23390
rect 33516 23324 33628 23380
rect 33628 23314 33684 23324
rect 33628 22372 33684 22382
rect 33628 22278 33684 22316
rect 33404 22148 33460 22158
rect 33404 21586 33460 22092
rect 33404 21534 33406 21586
rect 33458 21534 33460 21586
rect 33404 21522 33460 21534
rect 33852 22146 33908 22158
rect 33852 22094 33854 22146
rect 33906 22094 33908 22146
rect 33852 21586 33908 22094
rect 34188 22148 34244 22158
rect 34188 22054 34244 22092
rect 33852 21534 33854 21586
rect 33906 21534 33908 21586
rect 33852 21522 33908 21534
rect 33628 21364 33684 21374
rect 33628 20690 33684 21308
rect 33740 20804 33796 20814
rect 33740 20710 33796 20748
rect 34412 20802 34468 20814
rect 34412 20750 34414 20802
rect 34466 20750 34468 20802
rect 33628 20638 33630 20690
rect 33682 20638 33684 20690
rect 33628 20626 33684 20638
rect 34412 20692 34468 20750
rect 34412 20626 34468 20636
rect 34524 20188 34580 25228
rect 34748 24724 34804 24734
rect 34748 24050 34804 24668
rect 34748 23998 34750 24050
rect 34802 23998 34804 24050
rect 34748 23986 34804 23998
rect 34636 22372 34692 22382
rect 34692 22316 34804 22372
rect 34636 22306 34692 22316
rect 34748 21026 34804 22316
rect 34748 20974 34750 21026
rect 34802 20974 34804 21026
rect 34748 20962 34804 20974
rect 33628 20132 34580 20188
rect 33628 15148 33684 20132
rect 33628 15092 33908 15148
rect 33292 12226 33348 12236
rect 30940 12068 30996 12078
rect 28028 9538 28084 9548
rect 28476 9716 28532 9726
rect 26768 9436 27448 9446
rect 26824 9380 26872 9436
rect 26928 9434 26976 9436
rect 27032 9434 27080 9436
rect 26948 9382 26976 9434
rect 27072 9382 27080 9434
rect 26928 9380 26976 9382
rect 27032 9380 27080 9382
rect 27136 9434 27184 9436
rect 27240 9434 27288 9436
rect 27136 9382 27144 9434
rect 27240 9382 27268 9434
rect 27136 9380 27184 9382
rect 27240 9380 27288 9382
rect 27344 9380 27392 9436
rect 26768 9370 27448 9380
rect 22268 8652 22948 8662
rect 22324 8596 22372 8652
rect 22428 8650 22476 8652
rect 22532 8650 22580 8652
rect 22448 8598 22476 8650
rect 22572 8598 22580 8650
rect 22428 8596 22476 8598
rect 22532 8596 22580 8598
rect 22636 8650 22684 8652
rect 22740 8650 22788 8652
rect 22636 8598 22644 8650
rect 22740 8598 22768 8650
rect 22636 8596 22684 8598
rect 22740 8596 22788 8598
rect 22844 8596 22892 8652
rect 22268 8586 22948 8596
rect 26768 7868 27448 7878
rect 26824 7812 26872 7868
rect 26928 7866 26976 7868
rect 27032 7866 27080 7868
rect 26948 7814 26976 7866
rect 27072 7814 27080 7866
rect 26928 7812 26976 7814
rect 27032 7812 27080 7814
rect 27136 7866 27184 7868
rect 27240 7866 27288 7868
rect 27136 7814 27144 7866
rect 27240 7814 27268 7866
rect 27136 7812 27184 7814
rect 27240 7812 27288 7814
rect 27344 7812 27392 7868
rect 26768 7802 27448 7812
rect 22268 7084 22948 7094
rect 22324 7028 22372 7084
rect 22428 7082 22476 7084
rect 22532 7082 22580 7084
rect 22448 7030 22476 7082
rect 22572 7030 22580 7082
rect 22428 7028 22476 7030
rect 22532 7028 22580 7030
rect 22636 7082 22684 7084
rect 22740 7082 22788 7084
rect 22636 7030 22644 7082
rect 22740 7030 22768 7082
rect 22636 7028 22684 7030
rect 22740 7028 22788 7030
rect 22844 7028 22892 7084
rect 22268 7018 22948 7028
rect 25116 6692 25172 6702
rect 25116 6598 25172 6636
rect 25900 6692 25956 6702
rect 22268 5516 22948 5526
rect 22324 5460 22372 5516
rect 22428 5514 22476 5516
rect 22532 5514 22580 5516
rect 22448 5462 22476 5514
rect 22572 5462 22580 5514
rect 22428 5460 22476 5462
rect 22532 5460 22580 5462
rect 22636 5514 22684 5516
rect 22740 5514 22788 5516
rect 22636 5462 22644 5514
rect 22740 5462 22768 5514
rect 22636 5460 22684 5462
rect 22740 5460 22788 5462
rect 22844 5460 22892 5516
rect 22268 5450 22948 5460
rect 20748 4050 20804 4060
rect 13268 3948 13948 3958
rect 13324 3892 13372 3948
rect 13428 3946 13476 3948
rect 13532 3946 13580 3948
rect 13448 3894 13476 3946
rect 13572 3894 13580 3946
rect 13428 3892 13476 3894
rect 13532 3892 13580 3894
rect 13636 3946 13684 3948
rect 13740 3946 13788 3948
rect 13636 3894 13644 3946
rect 13740 3894 13768 3946
rect 13636 3892 13684 3894
rect 13740 3892 13788 3894
rect 13844 3892 13892 3948
rect 13268 3882 13948 3892
rect 22268 3948 22948 3958
rect 22324 3892 22372 3948
rect 22428 3946 22476 3948
rect 22532 3946 22580 3948
rect 22448 3894 22476 3946
rect 22572 3894 22580 3946
rect 22428 3892 22476 3894
rect 22532 3892 22580 3894
rect 22636 3946 22684 3948
rect 22740 3946 22788 3948
rect 22636 3894 22644 3946
rect 22740 3894 22768 3946
rect 22636 3892 22684 3894
rect 22740 3892 22788 3894
rect 22844 3892 22892 3948
rect 22268 3882 22948 3892
rect 25900 3780 25956 6636
rect 26796 6690 26852 6702
rect 26796 6638 26798 6690
rect 26850 6638 26852 6690
rect 26796 6468 26852 6638
rect 28364 6692 28420 6702
rect 28364 6598 28420 6636
rect 27916 6578 27972 6590
rect 27916 6526 27918 6578
rect 27970 6526 27972 6578
rect 26796 6402 26852 6412
rect 27580 6466 27636 6478
rect 27580 6414 27582 6466
rect 27634 6414 27636 6466
rect 26768 6300 27448 6310
rect 26824 6244 26872 6300
rect 26928 6298 26976 6300
rect 27032 6298 27080 6300
rect 26948 6246 26976 6298
rect 27072 6246 27080 6298
rect 26928 6244 26976 6246
rect 27032 6244 27080 6246
rect 27136 6298 27184 6300
rect 27240 6298 27288 6300
rect 27136 6246 27144 6298
rect 27240 6246 27268 6298
rect 27136 6244 27184 6246
rect 27240 6244 27288 6246
rect 27344 6244 27392 6300
rect 26768 6234 27448 6244
rect 27580 5906 27636 6414
rect 27580 5854 27582 5906
rect 27634 5854 27636 5906
rect 27580 5842 27636 5854
rect 26572 5236 26628 5246
rect 26572 5142 26628 5180
rect 27916 5124 27972 6526
rect 27916 5058 27972 5068
rect 28476 5122 28532 9660
rect 30044 9044 30100 9054
rect 30044 7586 30100 8988
rect 30044 7534 30046 7586
rect 30098 7534 30100 7586
rect 30044 7522 30100 7534
rect 30156 8930 30212 8942
rect 30156 8878 30158 8930
rect 30210 8878 30212 8930
rect 29372 6468 29428 6478
rect 29372 6374 29428 6412
rect 28476 5070 28478 5122
rect 28530 5070 28532 5122
rect 28476 5058 28532 5070
rect 30156 5012 30212 8878
rect 30716 6692 30772 6702
rect 30716 5346 30772 6636
rect 30716 5294 30718 5346
rect 30770 5294 30772 5346
rect 30716 5282 30772 5294
rect 30156 4946 30212 4956
rect 26768 4732 27448 4742
rect 26824 4676 26872 4732
rect 26928 4730 26976 4732
rect 27032 4730 27080 4732
rect 26948 4678 26976 4730
rect 27072 4678 27080 4730
rect 26928 4676 26976 4678
rect 27032 4676 27080 4678
rect 27136 4730 27184 4732
rect 27240 4730 27288 4732
rect 27136 4678 27144 4730
rect 27240 4678 27268 4730
rect 27136 4676 27184 4678
rect 27240 4676 27288 4678
rect 27344 4676 27392 4732
rect 26768 4666 27448 4676
rect 30156 4452 30212 4462
rect 30156 4358 30212 4396
rect 30940 4340 30996 12012
rect 31268 11788 31948 11798
rect 31324 11732 31372 11788
rect 31428 11786 31476 11788
rect 31532 11786 31580 11788
rect 31448 11734 31476 11786
rect 31572 11734 31580 11786
rect 31428 11732 31476 11734
rect 31532 11732 31580 11734
rect 31636 11786 31684 11788
rect 31740 11786 31788 11788
rect 31636 11734 31644 11786
rect 31740 11734 31768 11786
rect 31636 11732 31684 11734
rect 31740 11732 31788 11734
rect 31844 11732 31892 11788
rect 31268 11722 31948 11732
rect 31164 11396 31220 11406
rect 31052 11340 31164 11396
rect 31052 6018 31108 11340
rect 31164 11302 31220 11340
rect 31268 10220 31948 10230
rect 31324 10164 31372 10220
rect 31428 10218 31476 10220
rect 31532 10218 31580 10220
rect 31448 10166 31476 10218
rect 31572 10166 31580 10218
rect 31428 10164 31476 10166
rect 31532 10164 31580 10166
rect 31636 10218 31684 10220
rect 31740 10218 31788 10220
rect 31636 10166 31644 10218
rect 31740 10166 31768 10218
rect 31636 10164 31684 10166
rect 31740 10164 31788 10166
rect 31844 10164 31892 10220
rect 31268 10154 31948 10164
rect 31948 9716 32004 9726
rect 31948 9622 32004 9660
rect 31836 9044 31892 9054
rect 31836 8950 31892 8988
rect 31268 8652 31948 8662
rect 31324 8596 31372 8652
rect 31428 8650 31476 8652
rect 31532 8650 31580 8652
rect 31448 8598 31476 8650
rect 31572 8598 31580 8650
rect 31428 8596 31476 8598
rect 31532 8596 31580 8598
rect 31636 8650 31684 8652
rect 31740 8650 31788 8652
rect 31636 8598 31644 8650
rect 31740 8598 31768 8650
rect 31636 8596 31684 8598
rect 31740 8596 31788 8598
rect 31844 8596 31892 8652
rect 31268 8586 31948 8596
rect 33516 7586 33572 7598
rect 33516 7534 33518 7586
rect 33570 7534 33572 7586
rect 32508 7476 32564 7486
rect 32508 7382 32564 7420
rect 31268 7084 31948 7094
rect 31324 7028 31372 7084
rect 31428 7082 31476 7084
rect 31532 7082 31580 7084
rect 31448 7030 31476 7082
rect 31572 7030 31580 7082
rect 31428 7028 31476 7030
rect 31532 7028 31580 7030
rect 31636 7082 31684 7084
rect 31740 7082 31788 7084
rect 31636 7030 31644 7082
rect 31740 7030 31768 7082
rect 31636 7028 31684 7030
rect 31740 7028 31788 7030
rect 31844 7028 31892 7084
rect 31268 7018 31948 7028
rect 33516 6804 33572 7534
rect 33516 6738 33572 6748
rect 33740 6244 33796 6254
rect 31052 5966 31054 6018
rect 31106 5966 31108 6018
rect 31052 5954 31108 5966
rect 33516 6020 33572 6030
rect 33516 6018 33684 6020
rect 33516 5966 33518 6018
rect 33570 5966 33684 6018
rect 33516 5964 33684 5966
rect 33516 5954 33572 5964
rect 33404 5908 33460 5918
rect 31268 5516 31948 5526
rect 31324 5460 31372 5516
rect 31428 5514 31476 5516
rect 31532 5514 31580 5516
rect 31448 5462 31476 5514
rect 31572 5462 31580 5514
rect 31428 5460 31476 5462
rect 31532 5460 31580 5462
rect 31636 5514 31684 5516
rect 31740 5514 31788 5516
rect 31636 5462 31644 5514
rect 31740 5462 31768 5514
rect 31636 5460 31684 5462
rect 31740 5460 31788 5462
rect 31844 5460 31892 5516
rect 31268 5450 31948 5460
rect 33292 5348 33348 5358
rect 31052 4340 31108 4350
rect 30940 4338 31108 4340
rect 30940 4286 31054 4338
rect 31106 4286 31108 4338
rect 30940 4284 31108 4286
rect 25900 3714 25956 3724
rect 28812 3780 28868 3790
rect 31052 3780 31108 4284
rect 32508 4340 32564 4350
rect 31268 3948 31948 3958
rect 31324 3892 31372 3948
rect 31428 3946 31476 3948
rect 31532 3946 31580 3948
rect 31448 3894 31476 3946
rect 31572 3894 31580 3946
rect 31428 3892 31476 3894
rect 31532 3892 31580 3894
rect 31636 3946 31684 3948
rect 31740 3946 31788 3948
rect 31636 3894 31644 3946
rect 31740 3894 31768 3946
rect 31636 3892 31684 3894
rect 31740 3892 31788 3894
rect 31844 3892 31892 3948
rect 31268 3882 31948 3892
rect 31052 3724 31332 3780
rect 17836 3668 17892 3678
rect 17836 3574 17892 3612
rect 28812 3666 28868 3724
rect 28812 3614 28814 3666
rect 28866 3614 28868 3666
rect 28812 3602 28868 3614
rect 31276 3666 31332 3724
rect 31276 3614 31278 3666
rect 31330 3614 31332 3666
rect 31276 3602 31332 3614
rect 32508 3666 32564 4284
rect 32508 3614 32510 3666
rect 32562 3614 32564 3666
rect 31724 3556 31780 3566
rect 31724 3462 31780 3500
rect 32508 3556 32564 3614
rect 33068 4228 33124 4238
rect 33068 3666 33124 4172
rect 33292 4004 33348 5292
rect 33404 4226 33460 5852
rect 33628 4340 33684 5964
rect 33740 4452 33796 6188
rect 33852 6132 33908 15092
rect 34860 13746 34916 13758
rect 34860 13694 34862 13746
rect 34914 13694 34916 13746
rect 33964 11282 34020 11294
rect 33964 11230 33966 11282
rect 34018 11230 34020 11282
rect 33964 7028 34020 11230
rect 34524 8932 34580 8942
rect 34412 8930 34580 8932
rect 34412 8878 34526 8930
rect 34578 8878 34580 8930
rect 34412 8876 34580 8878
rect 34300 8148 34356 8158
rect 34300 8054 34356 8092
rect 34300 7588 34356 7598
rect 34412 7588 34468 8876
rect 34524 8866 34580 8876
rect 34300 7586 34468 7588
rect 34300 7534 34302 7586
rect 34354 7534 34468 7586
rect 34300 7532 34468 7534
rect 34636 7588 34692 7598
rect 34188 7250 34244 7262
rect 34188 7198 34190 7250
rect 34242 7198 34244 7250
rect 33964 6972 34132 7028
rect 33852 6066 33908 6076
rect 33964 6804 34020 6814
rect 33852 5908 33908 5918
rect 33852 5814 33908 5852
rect 33964 5460 34020 6748
rect 34076 5684 34132 6972
rect 34188 5906 34244 7198
rect 34300 6244 34356 7532
rect 34636 7494 34692 7532
rect 34748 7250 34804 7262
rect 34748 7198 34750 7250
rect 34802 7198 34804 7250
rect 34748 6916 34804 7198
rect 34748 6850 34804 6860
rect 34412 6580 34468 6590
rect 34412 6486 34468 6524
rect 34300 6178 34356 6188
rect 34860 6130 34916 13694
rect 34972 6356 35028 25228
rect 35196 24836 35252 26908
rect 35420 27074 35476 27086
rect 35420 27022 35422 27074
rect 35474 27022 35476 27074
rect 35420 25730 35476 27022
rect 35644 26962 35700 27806
rect 36988 27300 37044 30046
rect 37100 30098 37156 30716
rect 37100 30046 37102 30098
rect 37154 30046 37156 30098
rect 37100 30034 37156 30046
rect 38556 30436 38612 31500
rect 38892 31220 38948 31500
rect 38780 31218 38948 31220
rect 38780 31166 38894 31218
rect 38946 31166 38948 31218
rect 38780 31164 38948 31166
rect 38780 30436 38836 31164
rect 38892 31154 38948 31164
rect 39228 30770 39284 31726
rect 39564 31332 39620 32732
rect 39788 32676 39844 32686
rect 39676 32620 39788 32676
rect 39676 32562 39732 32620
rect 39788 32610 39844 32620
rect 39676 32510 39678 32562
rect 39730 32510 39732 32562
rect 39676 32498 39732 32510
rect 39900 32562 39956 32732
rect 41020 32788 41076 34300
rect 41244 33908 41300 34638
rect 41244 33842 41300 33852
rect 41468 34468 41524 34478
rect 41468 34354 41524 34412
rect 41468 34302 41470 34354
rect 41522 34302 41524 34354
rect 41020 32694 41076 32732
rect 41468 32786 41524 34302
rect 41804 33122 41860 33134
rect 41804 33070 41806 33122
rect 41858 33070 41860 33122
rect 41468 32734 41470 32786
rect 41522 32734 41524 32786
rect 41468 32676 41524 32734
rect 39900 32510 39902 32562
rect 39954 32510 39956 32562
rect 39900 32498 39956 32510
rect 40236 32564 40292 32574
rect 40236 32470 40292 32508
rect 39900 32340 39956 32350
rect 39228 30718 39230 30770
rect 39282 30718 39284 30770
rect 39228 30706 39284 30718
rect 39340 31276 39620 31332
rect 39788 31556 39844 31566
rect 38556 30380 38836 30436
rect 37324 29986 37380 29998
rect 37324 29934 37326 29986
rect 37378 29934 37380 29986
rect 37324 28756 37380 29934
rect 37324 28690 37380 28700
rect 37996 27972 38052 27982
rect 37996 27878 38052 27916
rect 37324 27300 37380 27310
rect 36988 27298 37380 27300
rect 36988 27246 37326 27298
rect 37378 27246 37380 27298
rect 36988 27244 37380 27246
rect 37324 27234 37380 27244
rect 37548 27188 37604 27198
rect 37548 27094 37604 27132
rect 38108 27188 38164 27198
rect 38108 27094 38164 27132
rect 35644 26910 35646 26962
rect 35698 26910 35700 26962
rect 35644 26898 35700 26910
rect 36988 26852 37044 26862
rect 36988 26758 37044 26796
rect 35768 26684 36448 26694
rect 35824 26628 35872 26684
rect 35928 26682 35976 26684
rect 36032 26682 36080 26684
rect 35948 26630 35976 26682
rect 36072 26630 36080 26682
rect 35928 26628 35976 26630
rect 36032 26628 36080 26630
rect 36136 26682 36184 26684
rect 36240 26682 36288 26684
rect 36136 26630 36144 26682
rect 36240 26630 36268 26682
rect 36136 26628 36184 26630
rect 36240 26628 36288 26630
rect 36344 26628 36392 26684
rect 35768 26618 36448 26628
rect 35420 25678 35422 25730
rect 35474 25678 35476 25730
rect 35420 25666 35476 25678
rect 35768 25116 36448 25126
rect 35824 25060 35872 25116
rect 35928 25114 35976 25116
rect 36032 25114 36080 25116
rect 35948 25062 35976 25114
rect 36072 25062 36080 25114
rect 35928 25060 35976 25062
rect 36032 25060 36080 25062
rect 36136 25114 36184 25116
rect 36240 25114 36288 25116
rect 36136 25062 36144 25114
rect 36240 25062 36268 25114
rect 36136 25060 36184 25062
rect 36240 25060 36288 25062
rect 36344 25060 36392 25116
rect 35768 25050 36448 25060
rect 38556 25060 38612 30380
rect 38780 30212 38836 30222
rect 38780 29538 38836 30156
rect 39340 29652 39396 31276
rect 39788 31218 39844 31500
rect 39788 31166 39790 31218
rect 39842 31166 39844 31218
rect 39788 31154 39844 31166
rect 39676 30994 39732 31006
rect 39676 30942 39678 30994
rect 39730 30942 39732 30994
rect 39452 30884 39508 30894
rect 39676 30884 39732 30942
rect 39452 30882 39732 30884
rect 39452 30830 39454 30882
rect 39506 30830 39732 30882
rect 39452 30828 39732 30830
rect 39452 30770 39508 30828
rect 39452 30718 39454 30770
rect 39506 30718 39508 30770
rect 39452 30706 39508 30718
rect 39788 29652 39844 29662
rect 39340 29650 39844 29652
rect 39340 29598 39342 29650
rect 39394 29598 39790 29650
rect 39842 29598 39844 29650
rect 39340 29596 39844 29598
rect 39340 29586 39396 29596
rect 38780 29486 38782 29538
rect 38834 29486 38836 29538
rect 38780 29474 38836 29486
rect 38780 27634 38836 27646
rect 38780 27582 38782 27634
rect 38834 27582 38836 27634
rect 38780 27188 38836 27582
rect 38780 27122 38836 27132
rect 38892 25508 38948 25518
rect 38892 25506 39620 25508
rect 38892 25454 38894 25506
rect 38946 25454 39620 25506
rect 38892 25452 39620 25454
rect 38892 25442 38948 25452
rect 39116 25282 39172 25294
rect 39452 25284 39508 25294
rect 39116 25230 39118 25282
rect 39170 25230 39172 25282
rect 38556 25004 38724 25060
rect 35196 24770 35252 24780
rect 35868 24836 35924 24846
rect 35868 24742 35924 24780
rect 37548 24836 37604 24846
rect 37548 24834 38276 24836
rect 37548 24782 37550 24834
rect 37602 24782 38276 24834
rect 37548 24780 38276 24782
rect 37548 24770 37604 24780
rect 36652 24724 36708 24734
rect 36652 24630 36708 24668
rect 35768 23548 36448 23558
rect 35824 23492 35872 23548
rect 35928 23546 35976 23548
rect 36032 23546 36080 23548
rect 35948 23494 35976 23546
rect 36072 23494 36080 23546
rect 35928 23492 35976 23494
rect 36032 23492 36080 23494
rect 36136 23546 36184 23548
rect 36240 23546 36288 23548
rect 36136 23494 36144 23546
rect 36240 23494 36268 23546
rect 36136 23492 36184 23494
rect 36240 23492 36288 23494
rect 36344 23492 36392 23548
rect 35768 23482 36448 23492
rect 37996 23380 38052 24780
rect 38220 24724 38276 24780
rect 38556 24834 38612 24846
rect 38556 24782 38558 24834
rect 38610 24782 38612 24834
rect 38444 24724 38500 24734
rect 38220 24722 38500 24724
rect 38220 24670 38446 24722
rect 38498 24670 38500 24722
rect 38220 24668 38500 24670
rect 38444 24658 38500 24668
rect 38108 24610 38164 24622
rect 38108 24558 38110 24610
rect 38162 24558 38164 24610
rect 38108 24500 38164 24558
rect 38556 24500 38612 24782
rect 38108 24444 38612 24500
rect 38108 24164 38164 24444
rect 38668 24388 38724 25004
rect 38556 24332 38724 24388
rect 38556 24276 38612 24332
rect 38108 24098 38164 24108
rect 38332 24220 38612 24276
rect 37996 22484 38052 23324
rect 38108 22484 38164 22494
rect 37996 22428 38108 22484
rect 38108 22390 38164 22428
rect 35768 21980 36448 21990
rect 35824 21924 35872 21980
rect 35928 21978 35976 21980
rect 36032 21978 36080 21980
rect 35948 21926 35976 21978
rect 36072 21926 36080 21978
rect 35928 21924 35976 21926
rect 36032 21924 36080 21926
rect 36136 21978 36184 21980
rect 36240 21978 36288 21980
rect 36136 21926 36144 21978
rect 36240 21926 36268 21978
rect 36136 21924 36184 21926
rect 36240 21924 36288 21926
rect 36344 21924 36392 21980
rect 35768 21914 36448 21924
rect 36204 21700 36260 21710
rect 36204 21606 36260 21644
rect 36988 21362 37044 21374
rect 36988 21310 36990 21362
rect 37042 21310 37044 21362
rect 36988 20692 37044 21310
rect 36988 20626 37044 20636
rect 35768 20412 36448 20422
rect 35824 20356 35872 20412
rect 35928 20410 35976 20412
rect 36032 20410 36080 20412
rect 35948 20358 35976 20410
rect 36072 20358 36080 20410
rect 35928 20356 35976 20358
rect 36032 20356 36080 20358
rect 36136 20410 36184 20412
rect 36240 20410 36288 20412
rect 36136 20358 36144 20410
rect 36240 20358 36268 20410
rect 36136 20356 36184 20358
rect 36240 20356 36288 20358
rect 36344 20356 36392 20412
rect 35768 20346 36448 20356
rect 35768 18844 36448 18854
rect 35824 18788 35872 18844
rect 35928 18842 35976 18844
rect 36032 18842 36080 18844
rect 35948 18790 35976 18842
rect 36072 18790 36080 18842
rect 35928 18788 35976 18790
rect 36032 18788 36080 18790
rect 36136 18842 36184 18844
rect 36240 18842 36288 18844
rect 36136 18790 36144 18842
rect 36240 18790 36268 18842
rect 36136 18788 36184 18790
rect 36240 18788 36288 18790
rect 36344 18788 36392 18844
rect 35768 18778 36448 18788
rect 35768 17276 36448 17286
rect 35824 17220 35872 17276
rect 35928 17274 35976 17276
rect 36032 17274 36080 17276
rect 35948 17222 35976 17274
rect 36072 17222 36080 17274
rect 35928 17220 35976 17222
rect 36032 17220 36080 17222
rect 36136 17274 36184 17276
rect 36240 17274 36288 17276
rect 36136 17222 36144 17274
rect 36240 17222 36268 17274
rect 36136 17220 36184 17222
rect 36240 17220 36288 17222
rect 36344 17220 36392 17276
rect 35768 17210 36448 17220
rect 35768 15708 36448 15718
rect 35824 15652 35872 15708
rect 35928 15706 35976 15708
rect 36032 15706 36080 15708
rect 35948 15654 35976 15706
rect 36072 15654 36080 15706
rect 35928 15652 35976 15654
rect 36032 15652 36080 15654
rect 36136 15706 36184 15708
rect 36240 15706 36288 15708
rect 36136 15654 36144 15706
rect 36240 15654 36268 15706
rect 36136 15652 36184 15654
rect 36240 15652 36288 15654
rect 36344 15652 36392 15708
rect 35768 15642 36448 15652
rect 38332 15148 38388 24220
rect 38892 23938 38948 23950
rect 38892 23886 38894 23938
rect 38946 23886 38948 23938
rect 38444 23714 38500 23726
rect 38444 23662 38446 23714
rect 38498 23662 38500 23714
rect 38444 23604 38500 23662
rect 38892 23716 38948 23886
rect 39116 23940 39172 25230
rect 39340 25282 39508 25284
rect 39340 25230 39454 25282
rect 39506 25230 39508 25282
rect 39340 25228 39508 25230
rect 39228 24500 39284 24510
rect 39228 24406 39284 24444
rect 39228 23940 39284 23950
rect 39116 23938 39284 23940
rect 39116 23886 39230 23938
rect 39282 23886 39284 23938
rect 39116 23884 39284 23886
rect 39228 23874 39284 23884
rect 39340 23716 39396 25228
rect 39452 25218 39508 25228
rect 39564 24946 39620 25452
rect 39564 24894 39566 24946
rect 39618 24894 39620 24946
rect 39564 24882 39620 24894
rect 39788 24500 39844 29596
rect 39900 28082 39956 32284
rect 40268 32172 40948 32182
rect 40324 32116 40372 32172
rect 40428 32170 40476 32172
rect 40532 32170 40580 32172
rect 40448 32118 40476 32170
rect 40572 32118 40580 32170
rect 40428 32116 40476 32118
rect 40532 32116 40580 32118
rect 40636 32170 40684 32172
rect 40740 32170 40788 32172
rect 40636 32118 40644 32170
rect 40740 32118 40768 32170
rect 40636 32116 40684 32118
rect 40740 32116 40788 32118
rect 40844 32116 40892 32172
rect 40268 32106 40948 32116
rect 41468 31780 41524 32620
rect 41468 31686 41524 31724
rect 41580 32788 41636 32798
rect 40684 31666 40740 31678
rect 40684 31614 40686 31666
rect 40738 31614 40740 31666
rect 40684 31556 40740 31614
rect 41580 31666 41636 32732
rect 41804 32340 41860 33070
rect 42140 32788 42196 38220
rect 42364 38164 42420 38612
rect 42700 38500 42756 40460
rect 42812 38668 42868 44940
rect 43260 44212 43316 44222
rect 43260 43652 43316 44156
rect 43260 43558 43316 43596
rect 43596 43538 43652 45164
rect 43596 43486 43598 43538
rect 43650 43486 43652 43538
rect 43596 43474 43652 43486
rect 43596 38948 43652 38958
rect 42812 38612 43092 38668
rect 42700 38444 42980 38500
rect 42364 38050 42420 38108
rect 42364 37998 42366 38050
rect 42418 37998 42420 38050
rect 42364 37986 42420 37998
rect 42700 37156 42756 37166
rect 42700 37062 42756 37100
rect 42924 36260 42980 38444
rect 43036 37156 43092 38612
rect 43372 37938 43428 37950
rect 43372 37886 43374 37938
rect 43426 37886 43428 37938
rect 43372 37828 43428 37886
rect 43372 37380 43428 37772
rect 43372 37286 43428 37324
rect 43596 37266 43652 38892
rect 43596 37214 43598 37266
rect 43650 37214 43652 37266
rect 43596 37202 43652 37214
rect 43036 37090 43092 37100
rect 42924 36194 42980 36204
rect 43036 34802 43092 34814
rect 43036 34750 43038 34802
rect 43090 34750 43092 34802
rect 41804 32274 41860 32284
rect 42028 32732 42196 32788
rect 42364 33122 42420 33134
rect 42364 33070 42366 33122
rect 42418 33070 42420 33122
rect 42364 32788 42420 33070
rect 41580 31614 41582 31666
rect 41634 31614 41636 31666
rect 41580 31602 41636 31614
rect 41692 32004 41748 32014
rect 40684 31490 40740 31500
rect 40012 30994 40068 31006
rect 40012 30942 40014 30994
rect 40066 30942 40068 30994
rect 40012 29764 40068 30942
rect 40268 30604 40948 30614
rect 40324 30548 40372 30604
rect 40428 30602 40476 30604
rect 40532 30602 40580 30604
rect 40448 30550 40476 30602
rect 40572 30550 40580 30602
rect 40428 30548 40476 30550
rect 40532 30548 40580 30550
rect 40636 30602 40684 30604
rect 40740 30602 40788 30604
rect 40636 30550 40644 30602
rect 40740 30550 40768 30602
rect 40636 30548 40684 30550
rect 40740 30548 40788 30550
rect 40844 30548 40892 30604
rect 40268 30538 40948 30548
rect 41580 30100 41636 30110
rect 41692 30100 41748 31948
rect 41580 30098 41748 30100
rect 41580 30046 41582 30098
rect 41634 30046 41748 30098
rect 41580 30044 41748 30046
rect 41580 30034 41636 30044
rect 40012 29698 40068 29708
rect 41692 29204 41748 29214
rect 40268 29036 40948 29046
rect 40324 28980 40372 29036
rect 40428 29034 40476 29036
rect 40532 29034 40580 29036
rect 40448 28982 40476 29034
rect 40572 28982 40580 29034
rect 40428 28980 40476 28982
rect 40532 28980 40580 28982
rect 40636 29034 40684 29036
rect 40740 29034 40788 29036
rect 40636 28982 40644 29034
rect 40740 28982 40768 29034
rect 40636 28980 40684 28982
rect 40740 28980 40788 28982
rect 40844 28980 40892 29036
rect 40268 28970 40948 28980
rect 41692 28642 41748 29148
rect 41692 28590 41694 28642
rect 41746 28590 41748 28642
rect 41692 28578 41748 28590
rect 39900 28030 39902 28082
rect 39954 28030 39956 28082
rect 39900 26908 39956 28030
rect 41356 28418 41412 28430
rect 41356 28366 41358 28418
rect 41410 28366 41412 28418
rect 40348 27970 40404 27982
rect 40348 27918 40350 27970
rect 40402 27918 40404 27970
rect 40348 27860 40404 27918
rect 40796 27860 40852 27870
rect 40348 27858 40852 27860
rect 40348 27806 40798 27858
rect 40850 27806 40852 27858
rect 40348 27804 40852 27806
rect 40796 27794 40852 27804
rect 41356 27858 41412 28366
rect 41356 27806 41358 27858
rect 41410 27806 41412 27858
rect 41356 27794 41412 27806
rect 40268 27468 40948 27478
rect 40324 27412 40372 27468
rect 40428 27466 40476 27468
rect 40532 27466 40580 27468
rect 40448 27414 40476 27466
rect 40572 27414 40580 27466
rect 40428 27412 40476 27414
rect 40532 27412 40580 27414
rect 40636 27466 40684 27468
rect 40740 27466 40788 27468
rect 40636 27414 40644 27466
rect 40740 27414 40768 27466
rect 40636 27412 40684 27414
rect 40740 27412 40788 27414
rect 40844 27412 40892 27468
rect 40268 27402 40948 27412
rect 39900 26852 40068 26908
rect 39788 24444 39956 24500
rect 38892 23660 39396 23716
rect 38780 23604 38836 23614
rect 38444 23548 38780 23604
rect 38668 22932 38724 22942
rect 38556 22484 38612 22494
rect 38556 22370 38612 22428
rect 38556 22318 38558 22370
rect 38610 22318 38612 22370
rect 38556 22306 38612 22318
rect 38668 22258 38724 22876
rect 38668 22206 38670 22258
rect 38722 22206 38724 22258
rect 38668 22194 38724 22206
rect 38780 21028 38836 23548
rect 39340 22372 39396 22382
rect 39004 22370 39396 22372
rect 39004 22318 39342 22370
rect 39394 22318 39396 22370
rect 39004 22316 39396 22318
rect 39004 21588 39060 22316
rect 39340 22306 39396 22316
rect 39676 22148 39732 22158
rect 39004 21522 39060 21532
rect 39116 22146 39732 22148
rect 39116 22094 39678 22146
rect 39730 22094 39732 22146
rect 39116 22092 39732 22094
rect 39116 21586 39172 22092
rect 39676 22082 39732 22092
rect 39900 21812 39956 24444
rect 40012 23604 40068 26852
rect 40268 25900 40948 25910
rect 40324 25844 40372 25900
rect 40428 25898 40476 25900
rect 40532 25898 40580 25900
rect 40448 25846 40476 25898
rect 40572 25846 40580 25898
rect 40428 25844 40476 25846
rect 40532 25844 40580 25846
rect 40636 25898 40684 25900
rect 40740 25898 40788 25900
rect 40636 25846 40644 25898
rect 40740 25846 40768 25898
rect 40636 25844 40684 25846
rect 40740 25844 40788 25846
rect 40844 25844 40892 25900
rect 40268 25834 40948 25844
rect 41580 24836 41636 24846
rect 40236 24612 40292 24622
rect 40124 24610 40292 24612
rect 40124 24558 40238 24610
rect 40290 24558 40292 24610
rect 40124 24556 40292 24558
rect 40124 24500 40180 24556
rect 40236 24546 40292 24556
rect 40124 23716 40180 24444
rect 40268 24332 40948 24342
rect 40324 24276 40372 24332
rect 40428 24330 40476 24332
rect 40532 24330 40580 24332
rect 40448 24278 40476 24330
rect 40572 24278 40580 24330
rect 40428 24276 40476 24278
rect 40532 24276 40580 24278
rect 40636 24330 40684 24332
rect 40740 24330 40788 24332
rect 40636 24278 40644 24330
rect 40740 24278 40768 24330
rect 40636 24276 40684 24278
rect 40740 24276 40788 24278
rect 40844 24276 40892 24332
rect 40268 24266 40948 24276
rect 40236 23716 40292 23726
rect 40124 23660 40236 23716
rect 40236 23650 40292 23660
rect 41580 23714 41636 24780
rect 41580 23662 41582 23714
rect 41634 23662 41636 23714
rect 40012 23538 40068 23548
rect 41580 23604 41636 23662
rect 41580 23538 41636 23548
rect 40268 22764 40948 22774
rect 40324 22708 40372 22764
rect 40428 22762 40476 22764
rect 40532 22762 40580 22764
rect 40448 22710 40476 22762
rect 40572 22710 40580 22762
rect 40428 22708 40476 22710
rect 40532 22708 40580 22710
rect 40636 22762 40684 22764
rect 40740 22762 40788 22764
rect 40636 22710 40644 22762
rect 40740 22710 40768 22762
rect 40636 22708 40684 22710
rect 40740 22708 40788 22710
rect 40844 22708 40892 22764
rect 40268 22698 40948 22708
rect 39116 21534 39118 21586
rect 39170 21534 39172 21586
rect 39116 21522 39172 21534
rect 39340 21698 39396 21710
rect 39340 21646 39342 21698
rect 39394 21646 39396 21698
rect 39004 21028 39060 21038
rect 38780 20972 39004 21028
rect 39004 20914 39060 20972
rect 39004 20862 39006 20914
rect 39058 20862 39060 20914
rect 39004 20850 39060 20862
rect 39228 20804 39284 20814
rect 39340 20804 39396 21646
rect 39788 20804 39844 20814
rect 39340 20802 39844 20804
rect 39340 20750 39790 20802
rect 39842 20750 39844 20802
rect 39340 20748 39844 20750
rect 39228 20710 39284 20748
rect 39788 20738 39844 20748
rect 39900 20132 39956 21756
rect 40124 22146 40180 22158
rect 40124 22094 40126 22146
rect 40178 22094 40180 22146
rect 40124 20804 40180 22094
rect 40268 21196 40948 21206
rect 40324 21140 40372 21196
rect 40428 21194 40476 21196
rect 40532 21194 40580 21196
rect 40448 21142 40476 21194
rect 40572 21142 40580 21194
rect 40428 21140 40476 21142
rect 40532 21140 40580 21142
rect 40636 21194 40684 21196
rect 40740 21194 40788 21196
rect 40636 21142 40644 21194
rect 40740 21142 40768 21194
rect 40636 21140 40684 21142
rect 40740 21140 40788 21142
rect 40844 21140 40892 21196
rect 40268 21130 40948 21140
rect 40124 20738 40180 20748
rect 40236 20244 40292 20254
rect 40124 20132 40180 20142
rect 39900 20130 40180 20132
rect 39900 20078 39902 20130
rect 39954 20078 40126 20130
rect 40178 20078 40180 20130
rect 39900 20076 40180 20078
rect 39900 20066 39956 20076
rect 40124 20066 40180 20076
rect 40236 20130 40292 20188
rect 40236 20078 40238 20130
rect 40290 20078 40292 20130
rect 40236 20066 40292 20078
rect 40460 20020 40516 20030
rect 40460 19926 40516 19964
rect 40268 19628 40948 19638
rect 40324 19572 40372 19628
rect 40428 19626 40476 19628
rect 40532 19626 40580 19628
rect 40448 19574 40476 19626
rect 40572 19574 40580 19626
rect 40428 19572 40476 19574
rect 40532 19572 40580 19574
rect 40636 19626 40684 19628
rect 40740 19626 40788 19628
rect 40636 19574 40644 19626
rect 40740 19574 40768 19626
rect 40636 19572 40684 19574
rect 40740 19572 40788 19574
rect 40844 19572 40892 19628
rect 40268 19562 40948 19572
rect 40012 19236 40068 19246
rect 40012 19142 40068 19180
rect 42028 19122 42084 32732
rect 42364 32722 42420 32732
rect 42924 32788 42980 32798
rect 42364 32004 42420 32014
rect 42364 31910 42420 31948
rect 42924 31890 42980 32732
rect 42924 31838 42926 31890
rect 42978 31838 42980 31890
rect 42924 31826 42980 31838
rect 42700 31780 42756 31790
rect 42700 31218 42756 31724
rect 42700 31166 42702 31218
rect 42754 31166 42756 31218
rect 42700 31154 42756 31166
rect 43036 30322 43092 34750
rect 43372 32002 43428 32014
rect 43372 31950 43374 32002
rect 43426 31950 43428 32002
rect 43372 31780 43428 31950
rect 43036 30270 43038 30322
rect 43090 30270 43092 30322
rect 43036 30258 43092 30270
rect 43148 31724 43372 31780
rect 42140 30212 42196 30222
rect 42140 30118 42196 30156
rect 42476 30100 42532 30110
rect 42476 29426 42532 30044
rect 43148 29538 43204 31724
rect 43372 31714 43428 31724
rect 43596 31778 43652 31790
rect 43596 31726 43598 31778
rect 43650 31726 43652 31778
rect 43596 30100 43652 31726
rect 43596 30006 43652 30044
rect 43148 29486 43150 29538
rect 43202 29486 43204 29538
rect 43148 29474 43204 29486
rect 43708 29988 43764 47182
rect 43932 46674 43988 48302
rect 44268 48244 44324 48254
rect 44268 48242 44996 48244
rect 44268 48190 44270 48242
rect 44322 48190 44996 48242
rect 44268 48188 44996 48190
rect 44268 48178 44324 48188
rect 44940 47682 44996 48188
rect 46396 48132 46452 48142
rect 44940 47630 44942 47682
rect 44994 47630 44996 47682
rect 44940 47618 44996 47630
rect 45948 48130 46564 48132
rect 45948 48078 46398 48130
rect 46450 48078 46564 48130
rect 45948 48076 46564 48078
rect 45276 47458 45332 47470
rect 45276 47406 45278 47458
rect 45330 47406 45332 47458
rect 43932 46622 43934 46674
rect 43986 46622 43988 46674
rect 43932 46610 43988 46622
rect 44268 47236 44324 47246
rect 45276 47236 45332 47406
rect 45948 47458 46004 48076
rect 46396 48066 46452 48076
rect 45948 47406 45950 47458
rect 46002 47406 46004 47458
rect 45948 47394 46004 47406
rect 46060 47348 46116 47358
rect 46060 47254 46116 47292
rect 44268 47234 45332 47236
rect 44268 47182 44270 47234
rect 44322 47182 45332 47234
rect 44268 47180 45332 47182
rect 44268 45332 44324 47180
rect 44768 47068 45448 47078
rect 44824 47012 44872 47068
rect 44928 47066 44976 47068
rect 45032 47066 45080 47068
rect 44948 47014 44976 47066
rect 45072 47014 45080 47066
rect 44928 47012 44976 47014
rect 45032 47012 45080 47014
rect 45136 47066 45184 47068
rect 45240 47066 45288 47068
rect 45136 47014 45144 47066
rect 45240 47014 45268 47066
rect 45136 47012 45184 47014
rect 45240 47012 45288 47014
rect 45344 47012 45392 47068
rect 44768 47002 45448 47012
rect 46172 46786 46228 46798
rect 46172 46734 46174 46786
rect 46226 46734 46228 46786
rect 44768 45500 45448 45510
rect 44824 45444 44872 45500
rect 44928 45498 44976 45500
rect 45032 45498 45080 45500
rect 44948 45446 44976 45498
rect 45072 45446 45080 45498
rect 44928 45444 44976 45446
rect 45032 45444 45080 45446
rect 45136 45498 45184 45500
rect 45240 45498 45288 45500
rect 45136 45446 45144 45498
rect 45240 45446 45268 45498
rect 45136 45444 45184 45446
rect 45240 45444 45288 45446
rect 45344 45444 45392 45500
rect 44768 45434 45448 45444
rect 44492 45332 44548 45342
rect 44268 45276 44492 45332
rect 44492 45238 44548 45276
rect 45276 45332 45332 45342
rect 43820 45220 43876 45230
rect 43820 45126 43876 45164
rect 45276 44546 45332 45276
rect 46172 44660 46228 46734
rect 45276 44494 45278 44546
rect 45330 44494 45332 44546
rect 45276 44482 45332 44494
rect 45836 44604 46228 44660
rect 44268 44212 44324 44222
rect 44940 44212 44996 44222
rect 44268 44210 44996 44212
rect 44268 44158 44270 44210
rect 44322 44158 44942 44210
rect 44994 44158 44996 44210
rect 44268 44156 44996 44158
rect 44268 44146 44324 44156
rect 44940 44146 44996 44156
rect 43932 44098 43988 44110
rect 43932 44046 43934 44098
rect 43986 44046 43988 44098
rect 43932 43540 43988 44046
rect 44768 43932 45448 43942
rect 44824 43876 44872 43932
rect 44928 43930 44976 43932
rect 45032 43930 45080 43932
rect 44948 43878 44976 43930
rect 45072 43878 45080 43930
rect 44928 43876 44976 43878
rect 45032 43876 45080 43878
rect 45136 43930 45184 43932
rect 45240 43930 45288 43932
rect 45136 43878 45144 43930
rect 45240 43878 45268 43930
rect 45136 43876 45184 43878
rect 45240 43876 45288 43878
rect 45344 43876 45392 43932
rect 44768 43866 45448 43876
rect 45836 43652 45892 44604
rect 46396 44548 46452 44558
rect 45948 44546 46452 44548
rect 45948 44494 46398 44546
rect 46450 44494 46452 44546
rect 45948 44492 46452 44494
rect 45948 44322 46004 44492
rect 46396 44482 46452 44492
rect 45948 44270 45950 44322
rect 46002 44270 46004 44322
rect 45948 44258 46004 44270
rect 46060 44324 46116 44334
rect 46060 44210 46116 44268
rect 46060 44158 46062 44210
rect 46114 44158 46116 44210
rect 46060 44146 46116 44158
rect 45836 43586 45892 43596
rect 46396 43652 46452 43662
rect 46396 43558 46452 43596
rect 44044 43540 44100 43550
rect 43932 43538 44100 43540
rect 43932 43486 44046 43538
rect 44098 43486 44100 43538
rect 43932 43484 44100 43486
rect 44044 43474 44100 43484
rect 44768 42364 45448 42374
rect 44824 42308 44872 42364
rect 44928 42362 44976 42364
rect 45032 42362 45080 42364
rect 44948 42310 44976 42362
rect 45072 42310 45080 42362
rect 44928 42308 44976 42310
rect 45032 42308 45080 42310
rect 45136 42362 45184 42364
rect 45240 42362 45288 42364
rect 45136 42310 45144 42362
rect 45240 42310 45268 42362
rect 45136 42308 45184 42310
rect 45240 42308 45288 42310
rect 45344 42308 45392 42364
rect 44768 42298 45448 42308
rect 44044 42082 44100 42094
rect 44044 42030 44046 42082
rect 44098 42030 44100 42082
rect 44044 41636 44100 42030
rect 44492 41972 44548 41982
rect 44492 41878 44548 41916
rect 44044 41580 44436 41636
rect 44044 41188 44100 41198
rect 44268 41188 44324 41198
rect 44044 41186 44212 41188
rect 44044 41134 44046 41186
rect 44098 41134 44212 41186
rect 44044 41132 44212 41134
rect 44044 41122 44100 41132
rect 44156 40740 44212 41132
rect 44380 41188 44436 41580
rect 44716 41188 44772 41198
rect 44380 41186 44772 41188
rect 44380 41134 44718 41186
rect 44770 41134 44772 41186
rect 44380 41132 44772 41134
rect 44268 41074 44324 41132
rect 44716 41122 44772 41132
rect 45276 41188 45332 41198
rect 45276 41094 45332 41132
rect 44268 41022 44270 41074
rect 44322 41022 44324 41074
rect 44268 41010 44324 41022
rect 44768 40796 45448 40806
rect 44824 40740 44872 40796
rect 44928 40794 44976 40796
rect 45032 40794 45080 40796
rect 44948 40742 44976 40794
rect 45072 40742 45080 40794
rect 44928 40740 44976 40742
rect 45032 40740 45080 40742
rect 45136 40794 45184 40796
rect 45240 40794 45288 40796
rect 45136 40742 45144 40794
rect 45240 40742 45268 40794
rect 45136 40740 45184 40742
rect 45240 40740 45288 40742
rect 45344 40740 45392 40796
rect 46508 40740 46564 48076
rect 44156 40684 44660 40740
rect 44768 40730 45448 40740
rect 44604 40628 44660 40684
rect 45836 40684 46564 40740
rect 44828 40628 44884 40638
rect 44604 40626 44884 40628
rect 44604 40574 44830 40626
rect 44882 40574 44884 40626
rect 44604 40572 44884 40574
rect 44828 40562 44884 40572
rect 45836 40402 45892 40684
rect 46508 40626 46564 40684
rect 46508 40574 46510 40626
rect 46562 40574 46564 40626
rect 46508 40562 46564 40574
rect 45948 40516 46004 40526
rect 45948 40422 46004 40460
rect 45836 40350 45838 40402
rect 45890 40350 45892 40402
rect 44380 40292 44436 40302
rect 45164 40292 45220 40302
rect 44380 40290 45220 40292
rect 44380 40238 44382 40290
rect 44434 40238 45166 40290
rect 45218 40238 45220 40290
rect 44380 40236 45220 40238
rect 44380 40226 44436 40236
rect 44492 39058 44548 40236
rect 45164 40226 45220 40236
rect 44768 39228 45448 39238
rect 44824 39172 44872 39228
rect 44928 39226 44976 39228
rect 45032 39226 45080 39228
rect 44948 39174 44976 39226
rect 45072 39174 45080 39226
rect 44928 39172 44976 39174
rect 45032 39172 45080 39174
rect 45136 39226 45184 39228
rect 45240 39226 45288 39228
rect 45136 39174 45144 39226
rect 45240 39174 45268 39226
rect 45136 39172 45184 39174
rect 45240 39172 45288 39174
rect 45344 39172 45392 39228
rect 44768 39162 45448 39172
rect 44492 39006 44494 39058
rect 44546 39006 44548 39058
rect 43820 38948 43876 38958
rect 43820 38854 43876 38892
rect 44492 38612 44548 39006
rect 44492 38546 44548 38556
rect 45276 38612 45332 38622
rect 45276 38274 45332 38556
rect 45276 38222 45278 38274
rect 45330 38222 45332 38274
rect 45276 38210 45332 38222
rect 44268 37940 44324 37950
rect 44940 37940 44996 37950
rect 44268 37938 44996 37940
rect 44268 37886 44270 37938
rect 44322 37886 44942 37938
rect 44994 37886 44996 37938
rect 44268 37884 44996 37886
rect 44268 37874 44324 37884
rect 44940 37874 44996 37884
rect 43932 37826 43988 37838
rect 43932 37774 43934 37826
rect 43986 37774 43988 37826
rect 43932 37268 43988 37774
rect 44768 37660 45448 37670
rect 44824 37604 44872 37660
rect 44928 37658 44976 37660
rect 45032 37658 45080 37660
rect 44948 37606 44976 37658
rect 45072 37606 45080 37658
rect 44928 37604 44976 37606
rect 45032 37604 45080 37606
rect 45136 37658 45184 37660
rect 45240 37658 45288 37660
rect 45136 37606 45144 37658
rect 45240 37606 45268 37658
rect 45136 37604 45184 37606
rect 45240 37604 45288 37606
rect 45344 37604 45392 37660
rect 44768 37594 45448 37604
rect 44044 37268 44100 37278
rect 43932 37266 44100 37268
rect 43932 37214 44046 37266
rect 44098 37214 44100 37266
rect 43932 37212 44100 37214
rect 44044 37202 44100 37212
rect 45612 37268 45668 37278
rect 45668 37212 45780 37268
rect 45612 37202 45668 37212
rect 44156 37156 44212 37166
rect 44044 36260 44100 36270
rect 44044 35138 44100 36204
rect 44044 35086 44046 35138
rect 44098 35086 44100 35138
rect 44044 35074 44100 35086
rect 44156 33572 44212 37100
rect 44768 36092 45448 36102
rect 44824 36036 44872 36092
rect 44928 36090 44976 36092
rect 45032 36090 45080 36092
rect 44948 36038 44976 36090
rect 45072 36038 45080 36090
rect 44928 36036 44976 36038
rect 45032 36036 45080 36038
rect 45136 36090 45184 36092
rect 45240 36090 45288 36092
rect 45136 36038 45144 36090
rect 45240 36038 45268 36090
rect 45136 36036 45184 36038
rect 45240 36036 45288 36038
rect 45344 36036 45392 36092
rect 44768 36026 45448 36036
rect 45052 35588 45108 35598
rect 44604 34804 44660 34814
rect 44604 34244 44660 34748
rect 44940 34804 44996 34814
rect 45052 34804 45108 35532
rect 44996 34748 45108 34804
rect 45388 35588 45444 35598
rect 45500 35588 45556 35598
rect 45388 35586 45556 35588
rect 45388 35534 45390 35586
rect 45442 35534 45502 35586
rect 45554 35534 45556 35586
rect 45388 35532 45556 35534
rect 44940 34710 44996 34748
rect 45388 34692 45444 35532
rect 45500 35522 45556 35532
rect 45500 34916 45556 34926
rect 45500 34914 45668 34916
rect 45500 34862 45502 34914
rect 45554 34862 45668 34914
rect 45500 34860 45668 34862
rect 45500 34850 45556 34860
rect 45388 34626 45444 34636
rect 44768 34524 45448 34534
rect 44824 34468 44872 34524
rect 44928 34522 44976 34524
rect 45032 34522 45080 34524
rect 44948 34470 44976 34522
rect 45072 34470 45080 34522
rect 44928 34468 44976 34470
rect 45032 34468 45080 34470
rect 45136 34522 45184 34524
rect 45240 34522 45288 34524
rect 45136 34470 45144 34522
rect 45240 34470 45268 34522
rect 45136 34468 45184 34470
rect 45240 34468 45288 34470
rect 45344 34468 45392 34524
rect 44768 34458 45448 34468
rect 44604 34188 44772 34244
rect 44604 34020 44660 34030
rect 44156 33506 44212 33516
rect 44268 34018 44660 34020
rect 44268 33966 44606 34018
rect 44658 33966 44660 34018
rect 44268 33964 44660 33966
rect 44268 33346 44324 33964
rect 44604 33954 44660 33964
rect 44268 33294 44270 33346
rect 44322 33294 44324 33346
rect 43932 33234 43988 33246
rect 43932 33182 43934 33234
rect 43986 33182 43988 33234
rect 43820 32564 43876 32574
rect 43820 31556 43876 32508
rect 43820 31106 43876 31500
rect 43820 31054 43822 31106
rect 43874 31054 43876 31106
rect 43820 31042 43876 31054
rect 43932 30996 43988 33182
rect 44044 33122 44100 33134
rect 44044 33070 44046 33122
rect 44098 33070 44100 33122
rect 44044 32674 44100 33070
rect 44044 32622 44046 32674
rect 44098 32622 44100 32674
rect 44044 32610 44100 32622
rect 44044 31892 44100 31902
rect 44044 31780 44100 31836
rect 44044 31778 44212 31780
rect 44044 31726 44046 31778
rect 44098 31726 44212 31778
rect 44044 31724 44212 31726
rect 44044 31714 44100 31724
rect 44044 30996 44100 31006
rect 43932 30994 44100 30996
rect 43932 30942 44046 30994
rect 44098 30942 44100 30994
rect 43932 30940 44100 30942
rect 42476 29374 42478 29426
rect 42530 29374 42532 29426
rect 42476 29362 42532 29374
rect 43260 29426 43316 29438
rect 43260 29374 43262 29426
rect 43314 29374 43316 29426
rect 43260 29316 43316 29374
rect 43260 29250 43316 29260
rect 42140 29204 42196 29214
rect 42140 29110 42196 29148
rect 43708 28644 43764 29932
rect 44044 30212 44100 30940
rect 44044 29650 44100 30156
rect 44156 30324 44212 31724
rect 44156 30210 44212 30268
rect 44156 30158 44158 30210
rect 44210 30158 44212 30210
rect 44156 30146 44212 30158
rect 44044 29598 44046 29650
rect 44098 29598 44100 29650
rect 44044 29586 44100 29598
rect 44156 29764 44212 29774
rect 44156 29540 44212 29708
rect 44156 29446 44212 29484
rect 44268 29428 44324 33294
rect 44604 33572 44660 33582
rect 44492 32452 44548 32462
rect 44492 30882 44548 32396
rect 44604 32450 44660 33516
rect 44716 33460 44772 34188
rect 45276 34018 45332 34030
rect 45276 33966 45278 34018
rect 45330 33966 45332 34018
rect 44716 33394 44772 33404
rect 44940 33908 44996 33918
rect 45276 33908 45332 33966
rect 44996 33852 45332 33908
rect 44940 33124 44996 33852
rect 45500 33572 45556 33582
rect 45612 33572 45668 34860
rect 45500 33570 45668 33572
rect 45500 33518 45502 33570
rect 45554 33518 45668 33570
rect 45500 33516 45668 33518
rect 45724 33572 45780 37212
rect 45836 34916 45892 40350
rect 46620 38668 46676 52108
rect 46732 52274 46788 53900
rect 47068 52388 47124 54238
rect 47292 53172 47348 54462
rect 48636 54516 48692 55022
rect 48860 54738 48916 55132
rect 51772 55076 51828 55086
rect 49644 54740 49700 54750
rect 48860 54686 48862 54738
rect 48914 54686 48916 54738
rect 48860 54674 48916 54686
rect 49308 54738 49700 54740
rect 49308 54686 49646 54738
rect 49698 54686 49700 54738
rect 49308 54684 49700 54686
rect 48748 54516 48804 54526
rect 48972 54516 49028 54526
rect 49308 54516 49364 54684
rect 49644 54674 49700 54684
rect 49756 54628 49812 54638
rect 49756 54534 49812 54572
rect 51772 54626 51828 55020
rect 52220 55076 52276 55086
rect 52668 55076 52724 55086
rect 52220 55074 52724 55076
rect 52220 55022 52222 55074
rect 52274 55022 52670 55074
rect 52722 55022 52724 55074
rect 52220 55020 52724 55022
rect 52220 55010 52276 55020
rect 51772 54574 51774 54626
rect 51826 54574 51828 54626
rect 51772 54562 51828 54574
rect 48636 54460 48748 54516
rect 48748 54422 48804 54460
rect 48860 54514 49364 54516
rect 48860 54462 48974 54514
rect 49026 54462 49364 54514
rect 48860 54460 49364 54462
rect 49420 54514 49476 54526
rect 49420 54462 49422 54514
rect 49474 54462 49476 54514
rect 48076 54404 48132 54414
rect 48076 54310 48132 54348
rect 48748 53842 48804 53854
rect 48748 53790 48750 53842
rect 48802 53790 48804 53842
rect 47292 53106 47348 53116
rect 47740 53508 47796 53518
rect 46732 52222 46734 52274
rect 46786 52222 46788 52274
rect 46732 51940 46788 52222
rect 46956 52332 47124 52388
rect 47740 52612 47796 53452
rect 46956 52052 47012 52332
rect 47180 52276 47236 52286
rect 47180 52182 47236 52220
rect 47740 52162 47796 52556
rect 47740 52110 47742 52162
rect 47794 52110 47796 52162
rect 47740 52098 47796 52110
rect 48188 52948 48244 52958
rect 48748 52948 48804 53790
rect 48860 53170 48916 54460
rect 48972 54450 49028 54460
rect 49420 54292 49476 54462
rect 50988 54514 51044 54526
rect 50988 54462 50990 54514
rect 51042 54462 51044 54514
rect 50652 54404 50708 54414
rect 50988 54404 51044 54462
rect 52668 54516 52724 55020
rect 52780 55076 52836 55086
rect 52780 54982 52836 55020
rect 52892 55074 52948 55086
rect 52892 55022 52894 55074
rect 52946 55022 52948 55074
rect 52668 54450 52724 54460
rect 50652 54402 51044 54404
rect 50652 54350 50654 54402
rect 50706 54350 51044 54402
rect 50652 54348 51044 54350
rect 52892 54404 52948 55022
rect 53116 55076 53172 55086
rect 53116 54982 53172 55020
rect 53768 54908 54448 54918
rect 53824 54852 53872 54908
rect 53928 54906 53976 54908
rect 54032 54906 54080 54908
rect 53948 54854 53976 54906
rect 54072 54854 54080 54906
rect 53928 54852 53976 54854
rect 54032 54852 54080 54854
rect 54136 54906 54184 54908
rect 54240 54906 54288 54908
rect 54136 54854 54144 54906
rect 54240 54854 54268 54906
rect 54136 54852 54184 54854
rect 54240 54852 54288 54854
rect 54344 54852 54392 54908
rect 53768 54842 54448 54852
rect 54348 54516 54404 54526
rect 54124 54514 54404 54516
rect 54124 54462 54350 54514
rect 54402 54462 54404 54514
rect 54124 54460 54404 54462
rect 49420 54236 50260 54292
rect 49268 54124 49948 54134
rect 49324 54068 49372 54124
rect 49428 54122 49476 54124
rect 49532 54122 49580 54124
rect 49448 54070 49476 54122
rect 49572 54070 49580 54122
rect 49428 54068 49476 54070
rect 49532 54068 49580 54070
rect 49636 54122 49684 54124
rect 49740 54122 49788 54124
rect 49636 54070 49644 54122
rect 49740 54070 49768 54122
rect 49636 54068 49684 54070
rect 49740 54068 49788 54070
rect 49844 54068 49892 54124
rect 49268 54058 49948 54068
rect 50092 53732 50148 53742
rect 48860 53118 48862 53170
rect 48914 53118 48916 53170
rect 48860 53106 48916 53118
rect 48972 53172 49028 53182
rect 48972 53170 49700 53172
rect 48972 53118 48974 53170
rect 49026 53118 49700 53170
rect 48972 53116 49700 53118
rect 48972 53106 49028 53116
rect 49644 53060 49700 53116
rect 49756 53060 49812 53070
rect 49644 53058 49812 53060
rect 49644 53006 49758 53058
rect 49810 53006 49812 53058
rect 49644 53004 49812 53006
rect 49756 52994 49812 53004
rect 49084 52948 49140 52958
rect 48748 52946 49140 52948
rect 48748 52894 49086 52946
rect 49138 52894 49140 52946
rect 48748 52892 49140 52894
rect 48188 52834 48244 52892
rect 48188 52782 48190 52834
rect 48242 52782 48244 52834
rect 46956 51986 47012 51996
rect 46732 51874 46788 51884
rect 47852 51940 47908 51950
rect 48188 51940 48244 52782
rect 49084 52836 49140 52892
rect 49420 52948 49476 52958
rect 49420 52854 49476 52892
rect 49084 52770 49140 52780
rect 49980 52724 50036 52762
rect 49980 52658 50036 52668
rect 49084 52612 49140 52622
rect 48748 52500 48804 52510
rect 48748 52386 48804 52444
rect 48748 52334 48750 52386
rect 48802 52334 48804 52386
rect 48300 52276 48356 52286
rect 48300 52182 48356 52220
rect 48748 52274 48804 52334
rect 48748 52222 48750 52274
rect 48802 52222 48804 52274
rect 48748 52210 48804 52222
rect 49084 52276 49140 52556
rect 49268 52556 49948 52566
rect 49324 52500 49372 52556
rect 49428 52554 49476 52556
rect 49532 52554 49580 52556
rect 49448 52502 49476 52554
rect 49572 52502 49580 52554
rect 49428 52500 49476 52502
rect 49532 52500 49580 52502
rect 49636 52554 49684 52556
rect 49740 52554 49788 52556
rect 49636 52502 49644 52554
rect 49740 52502 49768 52554
rect 49636 52500 49684 52502
rect 49740 52500 49788 52502
rect 49844 52500 49892 52556
rect 49268 52490 49948 52500
rect 50092 52500 50148 53676
rect 50204 53172 50260 54236
rect 50204 52946 50260 53116
rect 50428 53620 50484 53630
rect 50428 53058 50484 53564
rect 50428 53006 50430 53058
rect 50482 53006 50484 53058
rect 50428 52994 50484 53006
rect 50204 52894 50206 52946
rect 50258 52894 50260 52946
rect 50204 52882 50260 52894
rect 50316 52834 50372 52846
rect 50316 52782 50318 52834
rect 50370 52782 50372 52834
rect 50204 52500 50260 52510
rect 50092 52444 50204 52500
rect 49756 52388 49812 52398
rect 49756 52294 49812 52332
rect 49196 52276 49252 52286
rect 49084 52274 49252 52276
rect 49084 52222 49198 52274
rect 49250 52222 49252 52274
rect 49084 52220 49252 52222
rect 49196 52210 49252 52220
rect 50204 52274 50260 52444
rect 50204 52222 50206 52274
rect 50258 52222 50260 52274
rect 50204 52210 50260 52222
rect 49644 52164 49700 52174
rect 49644 52070 49700 52108
rect 47908 51884 48244 51940
rect 49980 52050 50036 52062
rect 49980 51998 49982 52050
rect 50034 51998 50036 52050
rect 47852 51602 47908 51884
rect 47852 51550 47854 51602
rect 47906 51550 47908 51602
rect 47852 51538 47908 51550
rect 47068 51492 47124 51502
rect 46844 51490 47124 51492
rect 46844 51438 47070 51490
rect 47122 51438 47124 51490
rect 46844 51436 47124 51438
rect 46732 51380 46788 51390
rect 46732 51286 46788 51324
rect 46844 50594 46900 51436
rect 47068 51426 47124 51436
rect 47404 51380 47460 51390
rect 47404 51286 47460 51324
rect 49980 51380 50036 51998
rect 49980 51378 50148 51380
rect 49980 51326 49982 51378
rect 50034 51326 50148 51378
rect 49980 51324 50148 51326
rect 49980 51314 50036 51324
rect 49268 50988 49948 50998
rect 49324 50932 49372 50988
rect 49428 50986 49476 50988
rect 49532 50986 49580 50988
rect 49448 50934 49476 50986
rect 49572 50934 49580 50986
rect 49428 50932 49476 50934
rect 49532 50932 49580 50934
rect 49636 50986 49684 50988
rect 49740 50986 49788 50988
rect 49636 50934 49644 50986
rect 49740 50934 49768 50986
rect 49636 50932 49684 50934
rect 49740 50932 49788 50934
rect 49844 50932 49892 50988
rect 49268 50922 49948 50932
rect 49868 50820 49924 50830
rect 50092 50820 50148 51324
rect 49868 50818 50148 50820
rect 49868 50766 49870 50818
rect 49922 50766 50148 50818
rect 49868 50764 50148 50766
rect 49868 50754 49924 50764
rect 46844 50542 46846 50594
rect 46898 50542 46900 50594
rect 46844 50530 46900 50542
rect 49084 50484 49140 50494
rect 49084 50390 49140 50428
rect 50316 49924 50372 52782
rect 50428 52388 50484 52398
rect 50428 51602 50484 52332
rect 50428 51550 50430 51602
rect 50482 51550 50484 51602
rect 50428 51538 50484 51550
rect 50316 49858 50372 49868
rect 50428 50596 50484 50606
rect 50428 49812 50484 50540
rect 50652 49812 50708 54348
rect 52892 54180 52948 54348
rect 51212 53732 51268 53742
rect 50764 53508 50820 53518
rect 50764 53058 50820 53452
rect 51100 53508 51156 53518
rect 50764 53006 50766 53058
rect 50818 53006 50820 53058
rect 50764 52994 50820 53006
rect 50876 53172 50932 53182
rect 50876 52834 50932 53116
rect 50876 52782 50878 52834
rect 50930 52782 50932 52834
rect 50876 52770 50932 52782
rect 50988 52946 51044 52958
rect 50988 52894 50990 52946
rect 51042 52894 51044 52946
rect 50764 52500 50820 52510
rect 50988 52500 51044 52894
rect 50820 52444 51044 52500
rect 50764 52274 50820 52444
rect 50764 52222 50766 52274
rect 50818 52222 50820 52274
rect 50764 52210 50820 52222
rect 51100 52276 51156 53452
rect 51212 53170 51268 53676
rect 52780 53730 52836 53742
rect 52780 53678 52782 53730
rect 52834 53678 52836 53730
rect 51212 53118 51214 53170
rect 51266 53118 51268 53170
rect 51212 53106 51268 53118
rect 51660 53620 51716 53630
rect 51660 53170 51716 53564
rect 51660 53118 51662 53170
rect 51714 53118 51716 53170
rect 51660 53106 51716 53118
rect 52108 53506 52164 53518
rect 52108 53454 52110 53506
rect 52162 53454 52164 53506
rect 51212 52276 51268 52286
rect 51100 52274 51268 52276
rect 51100 52222 51214 52274
rect 51266 52222 51268 52274
rect 51100 52220 51268 52222
rect 51212 52210 51268 52220
rect 52108 52276 52164 53454
rect 52444 52836 52500 52846
rect 52780 52836 52836 53678
rect 52892 53618 52948 54124
rect 53900 54404 53956 54414
rect 54124 54404 54180 54460
rect 54348 54450 54404 54460
rect 55580 54516 55636 54526
rect 55580 54422 55636 54460
rect 53900 54402 54180 54404
rect 53900 54350 53902 54402
rect 53954 54350 54180 54402
rect 53900 54348 54180 54350
rect 53900 53732 53956 54348
rect 54236 54290 54292 54302
rect 54236 54238 54238 54290
rect 54290 54238 54292 54290
rect 54236 54180 54292 54238
rect 54236 54114 54292 54124
rect 53900 53666 53956 53676
rect 52892 53566 52894 53618
rect 52946 53566 52948 53618
rect 52892 53554 52948 53566
rect 53768 53340 54448 53350
rect 53824 53284 53872 53340
rect 53928 53338 53976 53340
rect 54032 53338 54080 53340
rect 53948 53286 53976 53338
rect 54072 53286 54080 53338
rect 53928 53284 53976 53286
rect 54032 53284 54080 53286
rect 54136 53338 54184 53340
rect 54240 53338 54288 53340
rect 54136 53286 54144 53338
rect 54240 53286 54268 53338
rect 54136 53284 54184 53286
rect 54240 53284 54288 53286
rect 54344 53284 54392 53340
rect 53768 53274 54448 53284
rect 55580 52948 55636 52958
rect 52444 52834 52836 52836
rect 52444 52782 52446 52834
rect 52498 52782 52836 52834
rect 52444 52780 52836 52782
rect 54460 52836 54516 52846
rect 52444 52388 52500 52780
rect 52444 52322 52500 52332
rect 53340 52388 53396 52398
rect 52108 52210 52164 52220
rect 53340 52274 53396 52332
rect 53340 52222 53342 52274
rect 53394 52222 53396 52274
rect 53340 52210 53396 52222
rect 53788 52276 53844 52286
rect 53788 52182 53844 52220
rect 54348 52276 54404 52286
rect 54348 52162 54404 52220
rect 54348 52110 54350 52162
rect 54402 52110 54404 52162
rect 54348 52098 54404 52110
rect 54460 52050 54516 52780
rect 55132 52836 55188 52846
rect 55020 52722 55076 52734
rect 55020 52670 55022 52722
rect 55074 52670 55076 52722
rect 55020 52276 55076 52670
rect 55132 52388 55188 52780
rect 55580 52722 55636 52892
rect 55580 52670 55582 52722
rect 55634 52670 55636 52722
rect 55580 52658 55636 52670
rect 55188 52332 55412 52388
rect 55132 52322 55188 52332
rect 55020 52210 55076 52220
rect 55356 52162 55412 52332
rect 55356 52110 55358 52162
rect 55410 52110 55412 52162
rect 55356 52098 55412 52110
rect 55692 52274 55748 52286
rect 55692 52222 55694 52274
rect 55746 52222 55748 52274
rect 55692 52164 55748 52222
rect 55692 52098 55748 52108
rect 54460 51998 54462 52050
rect 54514 51998 54516 52050
rect 54460 51986 54516 51998
rect 55804 52052 55860 55246
rect 56028 55186 56084 55412
rect 66892 55298 66948 55310
rect 66892 55246 66894 55298
rect 66946 55246 66948 55298
rect 56028 55134 56030 55186
rect 56082 55134 56084 55186
rect 56028 55122 56084 55134
rect 58492 55186 58548 55198
rect 58492 55134 58494 55186
rect 58546 55134 58548 55186
rect 57260 55076 57316 55086
rect 57484 55076 57540 55086
rect 57260 55074 57540 55076
rect 57260 55022 57262 55074
rect 57314 55022 57486 55074
rect 57538 55022 57540 55074
rect 57260 55020 57540 55022
rect 56812 54628 56868 54638
rect 57260 54628 57316 55020
rect 57484 55010 57540 55020
rect 57596 55076 57652 55086
rect 57596 54982 57652 55020
rect 57708 55074 57764 55086
rect 57708 55022 57710 55074
rect 57762 55022 57764 55074
rect 56812 54626 57428 54628
rect 56812 54574 56814 54626
rect 56866 54574 57428 54626
rect 56812 54572 57428 54574
rect 56028 54516 56084 54526
rect 56588 54516 56644 54526
rect 56028 54514 56644 54516
rect 56028 54462 56030 54514
rect 56082 54462 56590 54514
rect 56642 54462 56644 54514
rect 56028 54460 56644 54462
rect 56028 53508 56084 54460
rect 56588 54450 56644 54460
rect 56812 54516 56868 54572
rect 56812 54450 56868 54460
rect 56028 53442 56084 53452
rect 56140 54292 56196 54302
rect 56028 52834 56084 52846
rect 56028 52782 56030 52834
rect 56082 52782 56084 52834
rect 56028 52724 56084 52782
rect 56028 52658 56084 52668
rect 56140 52164 56196 54236
rect 56812 54292 56868 54302
rect 56588 53730 56644 53742
rect 56588 53678 56590 53730
rect 56642 53678 56644 53730
rect 56476 53618 56532 53630
rect 56476 53566 56478 53618
rect 56530 53566 56532 53618
rect 56364 53508 56420 53518
rect 56364 53414 56420 53452
rect 56476 53284 56532 53566
rect 56476 53218 56532 53228
rect 56588 52948 56644 53678
rect 56812 53730 56868 54236
rect 56812 53678 56814 53730
rect 56866 53678 56868 53730
rect 56812 53666 56868 53678
rect 57372 53844 57428 54572
rect 57484 54626 57540 54638
rect 57484 54574 57486 54626
rect 57538 54574 57540 54626
rect 57484 54292 57540 54574
rect 57708 54628 57764 55022
rect 57932 55074 57988 55086
rect 57932 55022 57934 55074
rect 57986 55022 57988 55074
rect 57708 54562 57764 54572
rect 57820 54852 57876 54862
rect 57820 54404 57876 54796
rect 57820 54310 57876 54348
rect 57484 54226 57540 54236
rect 57372 53732 57428 53788
rect 57484 53732 57540 53742
rect 57932 53732 57988 55022
rect 58380 55074 58436 55086
rect 58380 55022 58382 55074
rect 58434 55022 58436 55074
rect 58380 54628 58436 55022
rect 58380 54562 58436 54572
rect 58380 54404 58436 54414
rect 58492 54404 58548 55134
rect 60508 55076 60564 55086
rect 58380 54402 58548 54404
rect 58380 54350 58382 54402
rect 58434 54350 58548 54402
rect 58380 54348 58548 54350
rect 59164 54740 59220 54750
rect 58380 54292 58436 54348
rect 58380 54226 58436 54236
rect 58268 54124 58948 54134
rect 58324 54068 58372 54124
rect 58428 54122 58476 54124
rect 58532 54122 58580 54124
rect 58448 54070 58476 54122
rect 58572 54070 58580 54122
rect 58428 54068 58476 54070
rect 58532 54068 58580 54070
rect 58636 54122 58684 54124
rect 58740 54122 58788 54124
rect 58636 54070 58644 54122
rect 58740 54070 58768 54122
rect 58636 54068 58684 54070
rect 58740 54068 58788 54070
rect 58844 54068 58892 54124
rect 58268 54058 58948 54068
rect 57372 53730 57540 53732
rect 57372 53678 57486 53730
rect 57538 53678 57540 53730
rect 57372 53676 57540 53678
rect 57484 53666 57540 53676
rect 57820 53676 57988 53732
rect 58044 53844 58100 53854
rect 57820 53620 57876 53676
rect 57260 53506 57316 53518
rect 57260 53454 57262 53506
rect 57314 53454 57316 53506
rect 57148 53060 57204 53070
rect 56924 52948 56980 52958
rect 57148 52948 57204 53004
rect 56644 52946 56980 52948
rect 56644 52894 56926 52946
rect 56978 52894 56980 52946
rect 56644 52892 56980 52894
rect 56588 52854 56644 52892
rect 56924 52882 56980 52892
rect 57036 52892 57204 52948
rect 56924 52724 56980 52734
rect 57036 52724 57092 52892
rect 56980 52668 57092 52724
rect 56812 52388 56868 52398
rect 56700 52332 56812 52388
rect 56140 52108 56420 52164
rect 53768 51772 54448 51782
rect 53824 51716 53872 51772
rect 53928 51770 53976 51772
rect 54032 51770 54080 51772
rect 53948 51718 53976 51770
rect 54072 51718 54080 51770
rect 53928 51716 53976 51718
rect 54032 51716 54080 51718
rect 54136 51770 54184 51772
rect 54240 51770 54288 51772
rect 54136 51718 54144 51770
rect 54240 51718 54268 51770
rect 54136 51716 54184 51718
rect 54240 51716 54288 51718
rect 54344 51716 54392 51772
rect 53768 51706 54448 51716
rect 55804 51602 55860 51996
rect 56028 52050 56084 52062
rect 56028 51998 56030 52050
rect 56082 51998 56084 52050
rect 56028 51828 56084 51998
rect 56364 52050 56420 52108
rect 56588 52162 56644 52174
rect 56588 52110 56590 52162
rect 56642 52110 56644 52162
rect 56364 51998 56366 52050
rect 56418 51998 56420 52050
rect 56364 51986 56420 51998
rect 56476 52052 56532 52062
rect 56588 52052 56644 52110
rect 56532 51996 56644 52052
rect 56476 51986 56532 51996
rect 56700 51828 56756 52332
rect 56812 52322 56868 52332
rect 56812 52164 56868 52174
rect 56812 52070 56868 52108
rect 56924 52162 56980 52668
rect 57260 52388 57316 53454
rect 57372 53506 57428 53518
rect 57372 53454 57374 53506
rect 57426 53454 57428 53506
rect 57372 52724 57428 53454
rect 57372 52658 57428 52668
rect 57484 53396 57540 53406
rect 57260 52322 57316 52332
rect 56924 52110 56926 52162
rect 56978 52110 56980 52162
rect 56924 52098 56980 52110
rect 57484 52164 57540 53340
rect 57708 53172 57764 53182
rect 57596 52164 57652 52174
rect 57484 52162 57652 52164
rect 57484 52110 57598 52162
rect 57650 52110 57652 52162
rect 57484 52108 57652 52110
rect 57148 51940 57204 51950
rect 57148 51938 57428 51940
rect 57148 51886 57150 51938
rect 57202 51886 57428 51938
rect 57148 51884 57428 51886
rect 57148 51874 57204 51884
rect 56028 51772 56756 51828
rect 55804 51550 55806 51602
rect 55858 51550 55860 51602
rect 55804 51538 55860 51550
rect 54796 51268 54852 51278
rect 53768 50204 54448 50214
rect 53824 50148 53872 50204
rect 53928 50202 53976 50204
rect 54032 50202 54080 50204
rect 53948 50150 53976 50202
rect 54072 50150 54080 50202
rect 53928 50148 53976 50150
rect 54032 50148 54080 50150
rect 54136 50202 54184 50204
rect 54240 50202 54288 50204
rect 54136 50150 54144 50202
rect 54240 50150 54268 50202
rect 54136 50148 54184 50150
rect 54240 50148 54288 50150
rect 54344 50148 54392 50204
rect 53768 50138 54448 50148
rect 51548 49924 51604 49934
rect 51548 49830 51604 49868
rect 50764 49812 50820 49822
rect 50428 49810 50820 49812
rect 50428 49758 50430 49810
rect 50482 49758 50766 49810
rect 50818 49758 50820 49810
rect 50428 49756 50820 49758
rect 50428 49746 50484 49756
rect 50764 49746 50820 49756
rect 53788 49700 53844 49710
rect 54796 49700 54852 51212
rect 55468 51268 55524 51278
rect 55692 51268 55748 51278
rect 55468 51266 55748 51268
rect 55468 51214 55470 51266
rect 55522 51214 55694 51266
rect 55746 51214 55748 51266
rect 55468 51212 55748 51214
rect 55244 50708 55300 50718
rect 55468 50708 55524 51212
rect 55692 51202 55748 51212
rect 57148 51266 57204 51278
rect 57148 51214 57150 51266
rect 57202 51214 57204 51266
rect 57148 51154 57204 51214
rect 57148 51102 57150 51154
rect 57202 51102 57204 51154
rect 57148 51090 57204 51102
rect 55244 50706 55524 50708
rect 55244 50654 55246 50706
rect 55298 50654 55524 50706
rect 55244 50652 55524 50654
rect 57372 50706 57428 51884
rect 57484 51154 57540 52108
rect 57596 52098 57652 52108
rect 57708 51828 57764 53116
rect 57820 52386 57876 53564
rect 57932 53508 57988 53518
rect 58044 53508 58100 53788
rect 59164 53842 59220 54684
rect 59500 54628 59556 54638
rect 59276 54292 59332 54302
rect 59276 53954 59332 54236
rect 59276 53902 59278 53954
rect 59330 53902 59332 53954
rect 59276 53890 59332 53902
rect 59164 53790 59166 53842
rect 59218 53790 59220 53842
rect 59164 53778 59220 53790
rect 57932 53506 58100 53508
rect 57932 53454 57934 53506
rect 57986 53454 58100 53506
rect 57932 53452 58100 53454
rect 59052 53506 59108 53518
rect 59052 53454 59054 53506
rect 59106 53454 59108 53506
rect 57932 53442 57988 53452
rect 58044 53284 58100 53294
rect 58044 53058 58100 53228
rect 58044 53006 58046 53058
rect 58098 53006 58100 53058
rect 58044 52994 58100 53006
rect 58940 52948 58996 52958
rect 58940 52854 58996 52892
rect 58268 52556 58948 52566
rect 57820 52334 57822 52386
rect 57874 52334 57876 52386
rect 57820 52322 57876 52334
rect 57932 52500 57988 52510
rect 58324 52500 58372 52556
rect 58428 52554 58476 52556
rect 58532 52554 58580 52556
rect 58448 52502 58476 52554
rect 58572 52502 58580 52554
rect 58428 52500 58476 52502
rect 58532 52500 58580 52502
rect 58636 52554 58684 52556
rect 58740 52554 58788 52556
rect 58636 52502 58644 52554
rect 58740 52502 58768 52554
rect 58636 52500 58684 52502
rect 58740 52500 58788 52502
rect 58844 52500 58892 52556
rect 58268 52490 58948 52500
rect 57932 52052 57988 52444
rect 58492 52388 58548 52398
rect 58492 52294 58548 52332
rect 58156 52276 58212 52286
rect 57484 51102 57486 51154
rect 57538 51102 57540 51154
rect 57484 51090 57540 51102
rect 57596 51772 57764 51828
rect 57820 52050 57988 52052
rect 57820 51998 57934 52050
rect 57986 51998 57988 52050
rect 57820 51996 57988 51998
rect 57372 50654 57374 50706
rect 57426 50654 57428 50706
rect 55244 50428 55300 50652
rect 57372 50642 57428 50654
rect 53788 49698 54852 49700
rect 53788 49646 53790 49698
rect 53842 49646 54852 49698
rect 53788 49644 54852 49646
rect 53788 49634 53844 49644
rect 49268 49420 49948 49430
rect 49324 49364 49372 49420
rect 49428 49418 49476 49420
rect 49532 49418 49580 49420
rect 49448 49366 49476 49418
rect 49572 49366 49580 49418
rect 49428 49364 49476 49366
rect 49532 49364 49580 49366
rect 49636 49418 49684 49420
rect 49740 49418 49788 49420
rect 49636 49366 49644 49418
rect 49740 49366 49768 49418
rect 49636 49364 49684 49366
rect 49740 49364 49788 49366
rect 49844 49364 49892 49420
rect 49268 49354 49948 49364
rect 53768 48636 54448 48646
rect 53824 48580 53872 48636
rect 53928 48634 53976 48636
rect 54032 48634 54080 48636
rect 53948 48582 53976 48634
rect 54072 48582 54080 48634
rect 53928 48580 53976 48582
rect 54032 48580 54080 48582
rect 54136 48634 54184 48636
rect 54240 48634 54288 48636
rect 54136 48582 54144 48634
rect 54240 48582 54268 48634
rect 54136 48580 54184 48582
rect 54240 48580 54288 48582
rect 54344 48580 54392 48636
rect 53768 48570 54448 48580
rect 52332 48468 52388 48478
rect 52332 48374 52388 48412
rect 52668 48468 52724 48478
rect 48972 48354 49028 48366
rect 48972 48302 48974 48354
rect 49026 48302 49028 48354
rect 48972 48244 49028 48302
rect 49196 48244 49252 48254
rect 48972 48242 49252 48244
rect 48972 48190 49198 48242
rect 49250 48190 49252 48242
rect 48972 48188 49252 48190
rect 49196 48178 49252 48188
rect 49868 48244 49924 48254
rect 49868 48242 50596 48244
rect 49868 48190 49870 48242
rect 49922 48190 50596 48242
rect 49868 48188 50596 48190
rect 49868 48178 49924 48188
rect 47740 48020 47796 48030
rect 47404 47460 47460 47470
rect 47404 47366 47460 47404
rect 47740 47458 47796 47964
rect 49268 47852 49948 47862
rect 49324 47796 49372 47852
rect 49428 47850 49476 47852
rect 49532 47850 49580 47852
rect 49448 47798 49476 47850
rect 49572 47798 49580 47850
rect 49428 47796 49476 47798
rect 49532 47796 49580 47798
rect 49636 47850 49684 47852
rect 49740 47850 49788 47852
rect 49636 47798 49644 47850
rect 49740 47798 49768 47850
rect 49636 47796 49684 47798
rect 49740 47796 49788 47798
rect 49844 47796 49892 47852
rect 49268 47786 49948 47796
rect 47740 47406 47742 47458
rect 47794 47406 47796 47458
rect 47740 47394 47796 47406
rect 48188 47572 48244 47582
rect 46956 47348 47012 47358
rect 46956 46898 47012 47292
rect 46956 46846 46958 46898
rect 47010 46846 47012 46898
rect 46956 46834 47012 46846
rect 47964 47234 48020 47246
rect 47964 47182 47966 47234
rect 48018 47182 48020 47234
rect 47404 45892 47460 45902
rect 47292 45836 47404 45892
rect 47292 45330 47348 45836
rect 47404 45826 47460 45836
rect 47516 45890 47572 45902
rect 47516 45838 47518 45890
rect 47570 45838 47572 45890
rect 47516 45668 47572 45838
rect 47964 45780 48020 47182
rect 48188 47234 48244 47516
rect 48748 47572 48804 47582
rect 48748 47478 48804 47516
rect 50092 47572 50148 47582
rect 48188 47182 48190 47234
rect 48242 47182 48244 47234
rect 48188 47170 48244 47182
rect 48860 47460 48916 47470
rect 48076 45780 48132 45790
rect 47964 45778 48132 45780
rect 47964 45726 48078 45778
rect 48130 45726 48132 45778
rect 47964 45724 48132 45726
rect 48076 45714 48132 45724
rect 47516 45602 47572 45612
rect 47292 45278 47294 45330
rect 47346 45278 47348 45330
rect 47292 45266 47348 45278
rect 47516 45218 47572 45230
rect 47516 45166 47518 45218
rect 47570 45166 47572 45218
rect 47516 45108 47572 45166
rect 47516 45042 47572 45052
rect 47628 45108 47684 45118
rect 48076 45108 48132 45118
rect 47628 45106 48356 45108
rect 47628 45054 47630 45106
rect 47682 45054 48078 45106
rect 48130 45054 48356 45106
rect 47628 45052 48356 45054
rect 47628 45042 47684 45052
rect 48076 45042 48132 45052
rect 46508 38612 46676 38668
rect 46732 44546 46788 44558
rect 46732 44494 46734 44546
rect 46786 44494 46788 44546
rect 46732 44098 46788 44494
rect 46732 44046 46734 44098
rect 46786 44046 46788 44098
rect 46396 38276 46452 38286
rect 45948 38274 46452 38276
rect 45948 38222 46398 38274
rect 46450 38222 46452 38274
rect 45948 38220 46452 38222
rect 45948 38050 46004 38220
rect 46396 38210 46452 38220
rect 45948 37998 45950 38050
rect 46002 37998 46004 38050
rect 45948 37986 46004 37998
rect 46060 37938 46116 37950
rect 46060 37886 46062 37938
rect 46114 37886 46116 37938
rect 46060 37828 46116 37886
rect 46060 37762 46116 37772
rect 46396 37380 46452 37390
rect 46396 37286 46452 37324
rect 46508 36596 46564 38612
rect 46732 38274 46788 44046
rect 47180 44324 47236 44334
rect 47180 43650 47236 44268
rect 48076 44324 48132 44334
rect 48076 44230 48132 44268
rect 47740 44212 47796 44222
rect 47740 44118 47796 44156
rect 47180 43598 47182 43650
rect 47234 43598 47236 43650
rect 47180 43586 47236 43598
rect 47628 43652 47684 43662
rect 47628 41074 47684 43596
rect 47628 41022 47630 41074
rect 47682 41022 47684 41074
rect 47628 41010 47684 41022
rect 48300 39732 48356 45052
rect 48636 44212 48692 44222
rect 48636 44118 48692 44156
rect 48860 41186 48916 47404
rect 49196 47460 49252 47470
rect 49196 47366 49252 47404
rect 49268 46284 49948 46294
rect 49324 46228 49372 46284
rect 49428 46282 49476 46284
rect 49532 46282 49580 46284
rect 49448 46230 49476 46282
rect 49572 46230 49580 46282
rect 49428 46228 49476 46230
rect 49532 46228 49580 46230
rect 49636 46282 49684 46284
rect 49740 46282 49788 46284
rect 49636 46230 49644 46282
rect 49740 46230 49768 46282
rect 49636 46228 49684 46230
rect 49740 46228 49788 46230
rect 49844 46228 49892 46284
rect 49268 46218 49948 46228
rect 49196 45892 49252 45902
rect 49196 45798 49252 45836
rect 49084 45778 49140 45790
rect 49084 45726 49086 45778
rect 49138 45726 49140 45778
rect 49084 44434 49140 45726
rect 49268 44716 49948 44726
rect 49324 44660 49372 44716
rect 49428 44714 49476 44716
rect 49532 44714 49580 44716
rect 49448 44662 49476 44714
rect 49572 44662 49580 44714
rect 49428 44660 49476 44662
rect 49532 44660 49580 44662
rect 49636 44714 49684 44716
rect 49740 44714 49788 44716
rect 49636 44662 49644 44714
rect 49740 44662 49768 44714
rect 49636 44660 49684 44662
rect 49740 44660 49788 44662
rect 49844 44660 49892 44716
rect 49268 44650 49948 44660
rect 50092 44548 50148 47516
rect 50540 47346 50596 48188
rect 50540 47294 50542 47346
rect 50594 47294 50596 47346
rect 50540 47282 50596 47294
rect 50876 47348 50932 47358
rect 50876 47346 51940 47348
rect 50876 47294 50878 47346
rect 50930 47294 51940 47346
rect 50876 47292 51940 47294
rect 50876 47282 50932 47292
rect 51436 46900 51492 46910
rect 51436 46806 51492 46844
rect 51884 46898 51940 47292
rect 51884 46846 51886 46898
rect 51938 46846 51940 46898
rect 51884 46834 51940 46846
rect 52444 46900 52500 46910
rect 52444 46786 52500 46844
rect 52444 46734 52446 46786
rect 52498 46734 52500 46786
rect 52220 46452 52276 46462
rect 52220 46358 52276 46396
rect 50316 46002 50372 46014
rect 50316 45950 50318 46002
rect 50370 45950 50372 46002
rect 50316 45332 50372 45950
rect 52444 45444 52500 46734
rect 52444 45378 52500 45388
rect 50316 45266 50372 45276
rect 49084 44382 49086 44434
rect 49138 44382 49140 44434
rect 49084 44370 49140 44382
rect 49980 44492 50148 44548
rect 50204 45218 50260 45230
rect 50204 45166 50206 45218
rect 50258 45166 50260 45218
rect 48972 44212 49028 44222
rect 49028 44156 49140 44212
rect 48972 44146 49028 44156
rect 48860 41134 48862 41186
rect 48914 41134 48916 41186
rect 48748 41074 48804 41086
rect 48748 41022 48750 41074
rect 48802 41022 48804 41074
rect 48412 40964 48468 40974
rect 48748 40964 48804 41022
rect 48412 40962 48804 40964
rect 48412 40910 48414 40962
rect 48466 40910 48804 40962
rect 48412 40908 48804 40910
rect 48412 40516 48468 40908
rect 48412 40450 48468 40460
rect 48860 40626 48916 41134
rect 48860 40574 48862 40626
rect 48914 40574 48916 40626
rect 48412 39732 48468 39742
rect 47964 39730 48468 39732
rect 47964 39678 48414 39730
rect 48466 39678 48468 39730
rect 47964 39676 48468 39678
rect 47740 38948 47796 38958
rect 47740 38854 47796 38892
rect 47964 38946 48020 39676
rect 48412 39666 48468 39676
rect 47964 38894 47966 38946
rect 48018 38894 48020 38946
rect 46732 38222 46734 38274
rect 46786 38222 46788 38274
rect 46172 36540 46564 36596
rect 46620 37828 46676 37838
rect 46732 37828 46788 38222
rect 46620 37826 46788 37828
rect 46620 37774 46622 37826
rect 46674 37774 46788 37826
rect 46620 37772 46788 37774
rect 47180 37828 47236 37838
rect 46620 36596 46676 37772
rect 47180 37490 47236 37772
rect 47180 37438 47182 37490
rect 47234 37438 47236 37490
rect 47180 37426 47236 37438
rect 46620 36540 46900 36596
rect 45948 36258 46004 36270
rect 45948 36206 45950 36258
rect 46002 36206 46004 36258
rect 45948 36148 46004 36206
rect 45948 36082 46004 36092
rect 45948 35586 46004 35598
rect 45948 35534 45950 35586
rect 46002 35534 46004 35586
rect 45948 35474 46004 35534
rect 45948 35422 45950 35474
rect 46002 35422 46004 35474
rect 45948 35410 46004 35422
rect 46172 35308 46228 36540
rect 46732 36370 46788 36382
rect 46732 36318 46734 36370
rect 46786 36318 46788 36370
rect 46396 36260 46452 36270
rect 46732 36260 46788 36318
rect 46396 36258 46788 36260
rect 46396 36206 46398 36258
rect 46450 36206 46788 36258
rect 46396 36204 46788 36206
rect 46396 36148 46452 36204
rect 46844 36148 46900 36540
rect 46060 35252 46228 35308
rect 46284 35476 46340 35486
rect 46396 35476 46452 36092
rect 46732 36092 46900 36148
rect 46956 36594 47012 36606
rect 46956 36542 46958 36594
rect 47010 36542 47012 36594
rect 46508 35810 46564 35822
rect 46508 35758 46510 35810
rect 46562 35758 46564 35810
rect 46508 35588 46564 35758
rect 46508 35522 46564 35532
rect 46284 35474 46452 35476
rect 46284 35422 46286 35474
rect 46338 35422 46452 35474
rect 46284 35420 46452 35422
rect 46620 35476 46676 35486
rect 46284 35364 46340 35420
rect 46620 35382 46676 35420
rect 46284 35298 46340 35308
rect 46620 35252 46676 35262
rect 46060 35140 46116 35252
rect 46060 35084 46452 35140
rect 46060 34916 46116 34926
rect 45836 34860 46060 34916
rect 46060 34822 46116 34860
rect 46284 34354 46340 34366
rect 46284 34302 46286 34354
rect 46338 34302 46340 34354
rect 46284 34244 46340 34302
rect 46284 34178 46340 34188
rect 45724 33516 45892 33572
rect 45500 33506 45556 33516
rect 45052 33346 45108 33358
rect 45052 33294 45054 33346
rect 45106 33294 45108 33346
rect 45052 33124 45108 33294
rect 45164 33348 45220 33358
rect 45164 33254 45220 33292
rect 45388 33348 45444 33358
rect 45388 33346 45780 33348
rect 45388 33294 45390 33346
rect 45442 33294 45780 33346
rect 45388 33292 45780 33294
rect 45388 33282 45444 33292
rect 45052 33068 45668 33124
rect 44940 33058 44996 33068
rect 44768 32956 45448 32966
rect 44824 32900 44872 32956
rect 44928 32954 44976 32956
rect 45032 32954 45080 32956
rect 44948 32902 44976 32954
rect 45072 32902 45080 32954
rect 44928 32900 44976 32902
rect 45032 32900 45080 32902
rect 45136 32954 45184 32956
rect 45240 32954 45288 32956
rect 45136 32902 45144 32954
rect 45240 32902 45268 32954
rect 45136 32900 45184 32902
rect 45240 32900 45288 32902
rect 45344 32900 45392 32956
rect 44768 32890 45448 32900
rect 44604 32398 44606 32450
rect 44658 32398 44660 32450
rect 44604 32386 44660 32398
rect 45612 32004 45668 33068
rect 44828 31780 44884 31790
rect 44828 31686 44884 31724
rect 45388 31666 45444 31678
rect 45388 31614 45390 31666
rect 45442 31614 45444 31666
rect 45388 31556 45444 31614
rect 45388 31490 45444 31500
rect 44768 31388 45448 31398
rect 44824 31332 44872 31388
rect 44928 31386 44976 31388
rect 45032 31386 45080 31388
rect 44948 31334 44976 31386
rect 45072 31334 45080 31386
rect 44928 31332 44976 31334
rect 45032 31332 45080 31334
rect 45136 31386 45184 31388
rect 45240 31386 45288 31388
rect 45136 31334 45144 31386
rect 45240 31334 45268 31386
rect 45136 31332 45184 31334
rect 45240 31332 45288 31334
rect 45344 31332 45392 31388
rect 44768 31322 45448 31332
rect 45052 31106 45108 31118
rect 45052 31054 45054 31106
rect 45106 31054 45108 31106
rect 45052 30996 45108 31054
rect 44492 30830 44494 30882
rect 44546 30830 44548 30882
rect 44492 30818 44548 30830
rect 44940 30940 45052 30996
rect 44492 30324 44548 30334
rect 44492 29650 44548 30268
rect 44492 29598 44494 29650
rect 44546 29598 44548 29650
rect 44492 29586 44548 29598
rect 44604 30100 44660 30110
rect 44604 29652 44660 30044
rect 44940 30100 44996 30940
rect 45052 30930 45108 30940
rect 45052 30212 45108 30222
rect 45052 30118 45108 30156
rect 44940 30034 44996 30044
rect 45612 30098 45668 31948
rect 45724 32562 45780 33292
rect 45724 32510 45726 32562
rect 45778 32510 45780 32562
rect 45724 30996 45780 32510
rect 45836 32004 45892 33516
rect 45948 33460 46004 33470
rect 45948 33366 46004 33404
rect 45836 31890 45892 31948
rect 46172 33348 46228 33358
rect 46396 33348 46452 35084
rect 46620 35028 46676 35196
rect 46620 34962 46676 34972
rect 46620 34244 46676 34254
rect 46732 34244 46788 36092
rect 46956 34916 47012 36542
rect 47964 36596 48020 38894
rect 48076 38946 48132 38958
rect 48076 38894 48078 38946
rect 48130 38894 48132 38946
rect 48076 38276 48132 38894
rect 48300 38834 48356 38846
rect 48300 38782 48302 38834
rect 48354 38782 48356 38834
rect 48300 38668 48356 38782
rect 48748 38834 48804 38846
rect 48748 38782 48750 38834
rect 48802 38782 48804 38834
rect 48300 38612 48468 38668
rect 48076 38210 48132 38220
rect 48188 38052 48244 38062
rect 48188 37958 48244 37996
rect 48412 38052 48468 38612
rect 48412 37986 48468 37996
rect 48748 37828 48804 38782
rect 48748 37762 48804 37772
rect 47964 36540 48132 36596
rect 47740 36484 47796 36494
rect 47740 36482 48020 36484
rect 47740 36430 47742 36482
rect 47794 36430 48020 36482
rect 47740 36428 48020 36430
rect 47740 36418 47796 36428
rect 47740 35812 47796 35822
rect 47740 35718 47796 35756
rect 47180 35698 47236 35710
rect 47180 35646 47182 35698
rect 47234 35646 47236 35698
rect 47068 35588 47124 35598
rect 47068 35028 47124 35532
rect 47180 35476 47236 35646
rect 47180 35140 47236 35420
rect 47180 35084 47572 35140
rect 47068 34972 47348 35028
rect 46956 34860 47124 34916
rect 46844 34802 46900 34814
rect 46844 34750 46846 34802
rect 46898 34750 46900 34802
rect 46844 34692 46900 34750
rect 47068 34804 47124 34860
rect 47292 34914 47348 34972
rect 47292 34862 47294 34914
rect 47346 34862 47348 34914
rect 47292 34850 47348 34862
rect 47068 34738 47124 34748
rect 46844 34626 46900 34636
rect 46956 34690 47012 34702
rect 46956 34638 46958 34690
rect 47010 34638 47012 34690
rect 46676 34188 46788 34244
rect 46620 34178 46676 34188
rect 46844 34130 46900 34142
rect 46844 34078 46846 34130
rect 46898 34078 46900 34130
rect 46396 33292 46676 33348
rect 46172 32786 46228 33292
rect 46396 33124 46452 33134
rect 46396 33030 46452 33068
rect 46172 32734 46174 32786
rect 46226 32734 46228 32786
rect 46172 32004 46228 32734
rect 46172 31938 46228 31948
rect 46396 32674 46452 32686
rect 46396 32622 46398 32674
rect 46450 32622 46452 32674
rect 45836 31838 45838 31890
rect 45890 31838 45892 31890
rect 45836 31826 45892 31838
rect 46396 31892 46452 32622
rect 45724 30930 45780 30940
rect 46396 30994 46452 31836
rect 46396 30942 46398 30994
rect 46450 30942 46452 30994
rect 46396 30930 46452 30942
rect 46508 32562 46564 32574
rect 46508 32510 46510 32562
rect 46562 32510 46564 32562
rect 46508 31778 46564 32510
rect 46508 31726 46510 31778
rect 46562 31726 46564 31778
rect 46284 30884 46340 30894
rect 45612 30046 45614 30098
rect 45666 30046 45668 30098
rect 45612 30034 45668 30046
rect 45724 30212 45780 30222
rect 44768 29820 45448 29830
rect 44824 29764 44872 29820
rect 44928 29818 44976 29820
rect 45032 29818 45080 29820
rect 44948 29766 44976 29818
rect 45072 29766 45080 29818
rect 44928 29764 44976 29766
rect 45032 29764 45080 29766
rect 45136 29818 45184 29820
rect 45240 29818 45288 29820
rect 45136 29766 45144 29818
rect 45240 29766 45268 29818
rect 45136 29764 45184 29766
rect 45240 29764 45288 29766
rect 45344 29764 45392 29820
rect 44768 29754 45448 29764
rect 44604 29596 45108 29652
rect 44716 29428 44772 29438
rect 44268 29372 44716 29428
rect 44716 29334 44772 29372
rect 44044 29316 44100 29326
rect 44044 29202 44100 29260
rect 44044 29150 44046 29202
rect 44098 29150 44100 29202
rect 44044 29138 44100 29150
rect 45052 28866 45108 29596
rect 45500 29428 45556 29438
rect 45500 29334 45556 29372
rect 45052 28814 45054 28866
rect 45106 28814 45108 28866
rect 45052 28802 45108 28814
rect 44380 28644 44436 28654
rect 43708 28588 44100 28644
rect 43932 28082 43988 28094
rect 43932 28030 43934 28082
rect 43986 28030 43988 28082
rect 43148 25508 43204 25518
rect 43148 25414 43204 25452
rect 43372 25506 43428 25518
rect 43372 25454 43374 25506
rect 43426 25454 43428 25506
rect 43036 25394 43092 25406
rect 43036 25342 43038 25394
rect 43090 25342 43092 25394
rect 42700 25284 42756 25294
rect 43036 25284 43092 25342
rect 42756 25228 43092 25284
rect 43260 25396 43316 25406
rect 42700 25190 42756 25228
rect 43036 24948 43092 24958
rect 43260 24948 43316 25340
rect 43036 24946 43316 24948
rect 43036 24894 43038 24946
rect 43090 24894 43316 24946
rect 43036 24892 43316 24894
rect 43036 24882 43092 24892
rect 43260 24724 43316 24892
rect 43372 24946 43428 25454
rect 43820 25396 43876 25406
rect 43820 25284 43876 25340
rect 43372 24894 43374 24946
rect 43426 24894 43428 24946
rect 43372 24882 43428 24894
rect 43484 25228 43876 25284
rect 43484 24724 43540 25228
rect 43932 25172 43988 28030
rect 43932 24836 43988 25116
rect 43932 24770 43988 24780
rect 43260 24722 43540 24724
rect 43260 24670 43486 24722
rect 43538 24670 43540 24722
rect 43260 24668 43540 24670
rect 43484 24658 43540 24668
rect 42364 23716 42420 23726
rect 42364 23622 42420 23660
rect 43372 21812 43428 21822
rect 43820 21812 43876 21822
rect 43428 21756 43540 21812
rect 43372 21718 43428 21756
rect 42924 21588 42980 21598
rect 42140 21028 42196 21038
rect 42140 20690 42196 20972
rect 42924 21026 42980 21532
rect 42924 20974 42926 21026
rect 42978 20974 42980 21026
rect 42924 20962 42980 20974
rect 43484 21476 43540 21756
rect 43820 21718 43876 21756
rect 43708 21586 43764 21598
rect 43708 21534 43710 21586
rect 43762 21534 43764 21586
rect 43596 21476 43652 21486
rect 43708 21476 43764 21534
rect 43484 21420 43596 21476
rect 43652 21420 43764 21476
rect 43484 20914 43540 21420
rect 43596 21382 43652 21420
rect 43484 20862 43486 20914
rect 43538 20862 43540 20914
rect 43484 20850 43540 20862
rect 43708 20804 43764 21420
rect 43820 21364 43876 21374
rect 43820 21270 43876 21308
rect 43820 20804 43876 20814
rect 43708 20802 43876 20804
rect 43708 20750 43822 20802
rect 43874 20750 43876 20802
rect 43708 20748 43876 20750
rect 43820 20738 43876 20748
rect 42140 20638 42142 20690
rect 42194 20638 42196 20690
rect 42140 20626 42196 20638
rect 43932 20692 43988 20702
rect 43932 20598 43988 20636
rect 44044 20188 44100 28588
rect 44380 28084 44436 28588
rect 44768 28252 45448 28262
rect 44824 28196 44872 28252
rect 44928 28250 44976 28252
rect 45032 28250 45080 28252
rect 44948 28198 44976 28250
rect 45072 28198 45080 28250
rect 44928 28196 44976 28198
rect 45032 28196 45080 28198
rect 45136 28250 45184 28252
rect 45240 28250 45288 28252
rect 45136 28198 45144 28250
rect 45240 28198 45268 28250
rect 45136 28196 45184 28198
rect 45240 28196 45288 28198
rect 45344 28196 45392 28252
rect 44768 28186 45448 28196
rect 44492 28084 44548 28094
rect 44380 28082 44548 28084
rect 44380 28030 44494 28082
rect 44546 28030 44548 28082
rect 44380 28028 44548 28030
rect 44492 26180 44548 28028
rect 45724 27746 45780 30156
rect 46172 30100 46228 30110
rect 46172 29650 46228 30044
rect 46172 29598 46174 29650
rect 46226 29598 46228 29650
rect 46172 29586 46228 29598
rect 46284 29650 46340 30828
rect 46508 30212 46564 31726
rect 46508 30146 46564 30156
rect 46284 29598 46286 29650
rect 46338 29598 46340 29650
rect 46284 29586 46340 29598
rect 46396 29540 46452 29550
rect 45836 29426 45892 29438
rect 45836 29374 45838 29426
rect 45890 29374 45892 29426
rect 45836 29316 45892 29374
rect 46060 29428 46116 29438
rect 46060 29334 46116 29372
rect 46396 29426 46452 29484
rect 46396 29374 46398 29426
rect 46450 29374 46452 29426
rect 45836 29250 45892 29260
rect 46396 28756 46452 29374
rect 46508 28756 46564 28766
rect 46396 28754 46564 28756
rect 46396 28702 46510 28754
rect 46562 28702 46564 28754
rect 46396 28700 46564 28702
rect 46508 28690 46564 28700
rect 45836 28644 45892 28654
rect 45836 28550 45892 28588
rect 45724 27694 45726 27746
rect 45778 27694 45780 27746
rect 45724 27682 45780 27694
rect 46396 27858 46452 27870
rect 46396 27806 46398 27858
rect 46450 27806 46452 27858
rect 46396 27748 46452 27806
rect 46396 27682 46452 27692
rect 44768 26684 45448 26694
rect 44824 26628 44872 26684
rect 44928 26682 44976 26684
rect 45032 26682 45080 26684
rect 44948 26630 44976 26682
rect 45072 26630 45080 26682
rect 44928 26628 44976 26630
rect 45032 26628 45080 26630
rect 45136 26682 45184 26684
rect 45240 26682 45288 26684
rect 45136 26630 45144 26682
rect 45240 26630 45268 26682
rect 45136 26628 45184 26630
rect 45240 26628 45288 26630
rect 45344 26628 45392 26684
rect 44768 26618 45448 26628
rect 44156 26124 44548 26180
rect 44156 24724 44212 26124
rect 44268 25564 44548 25620
rect 44268 25394 44324 25564
rect 44492 25508 44548 25564
rect 44716 25508 44772 25518
rect 44492 25506 44772 25508
rect 44492 25454 44718 25506
rect 44770 25454 44772 25506
rect 44492 25452 44772 25454
rect 44716 25442 44772 25452
rect 45276 25506 45332 25518
rect 45276 25454 45278 25506
rect 45330 25454 45332 25506
rect 44268 25342 44270 25394
rect 44322 25342 44324 25394
rect 44268 25330 44324 25342
rect 45276 25396 45332 25454
rect 45276 25330 45332 25340
rect 44268 25172 44324 25182
rect 44268 24946 44324 25116
rect 44768 25116 45448 25126
rect 44824 25060 44872 25116
rect 44928 25114 44976 25116
rect 45032 25114 45080 25116
rect 44948 25062 44976 25114
rect 45072 25062 45080 25114
rect 44928 25060 44976 25062
rect 45032 25060 45080 25062
rect 45136 25114 45184 25116
rect 45240 25114 45288 25116
rect 45136 25062 45144 25114
rect 45240 25062 45268 25114
rect 45136 25060 45184 25062
rect 45240 25060 45288 25062
rect 45344 25060 45392 25116
rect 44768 25050 45448 25060
rect 44268 24894 44270 24946
rect 44322 24894 44324 24946
rect 44268 24882 44324 24894
rect 44156 24668 44436 24724
rect 44156 20580 44212 20590
rect 44156 20486 44212 20524
rect 44044 20132 44324 20188
rect 44268 19236 44324 20132
rect 44268 19142 44324 19180
rect 42028 19070 42030 19122
rect 42082 19070 42084 19122
rect 40268 18060 40948 18070
rect 40324 18004 40372 18060
rect 40428 18058 40476 18060
rect 40532 18058 40580 18060
rect 40448 18006 40476 18058
rect 40572 18006 40580 18058
rect 40428 18004 40476 18006
rect 40532 18004 40580 18006
rect 40636 18058 40684 18060
rect 40740 18058 40788 18060
rect 40636 18006 40644 18058
rect 40740 18006 40768 18058
rect 40636 18004 40684 18006
rect 40740 18004 40788 18006
rect 40844 18004 40892 18060
rect 40268 17994 40948 18004
rect 40268 16492 40948 16502
rect 40324 16436 40372 16492
rect 40428 16490 40476 16492
rect 40532 16490 40580 16492
rect 40448 16438 40476 16490
rect 40572 16438 40580 16490
rect 40428 16436 40476 16438
rect 40532 16436 40580 16438
rect 40636 16490 40684 16492
rect 40740 16490 40788 16492
rect 40636 16438 40644 16490
rect 40740 16438 40768 16490
rect 40636 16436 40684 16438
rect 40740 16436 40788 16438
rect 40844 16436 40892 16492
rect 40268 16426 40948 16436
rect 41692 15316 41748 15326
rect 41692 15314 41860 15316
rect 41692 15262 41694 15314
rect 41746 15262 41860 15314
rect 41692 15260 41860 15262
rect 41692 15250 41748 15260
rect 38220 15092 38388 15148
rect 41132 15204 41188 15214
rect 41244 15204 41300 15214
rect 41132 15202 41244 15204
rect 41132 15150 41134 15202
rect 41186 15150 41244 15202
rect 41132 15148 41244 15150
rect 41132 15092 41300 15148
rect 35768 14140 36448 14150
rect 35824 14084 35872 14140
rect 35928 14138 35976 14140
rect 36032 14138 36080 14140
rect 35948 14086 35976 14138
rect 36072 14086 36080 14138
rect 35928 14084 35976 14086
rect 36032 14084 36080 14086
rect 36136 14138 36184 14140
rect 36240 14138 36288 14140
rect 36136 14086 36144 14138
rect 36240 14086 36268 14138
rect 36136 14084 36184 14086
rect 36240 14084 36288 14086
rect 36344 14084 36392 14140
rect 35768 14074 36448 14084
rect 37212 13634 37268 13646
rect 37212 13582 37214 13634
rect 37266 13582 37268 13634
rect 37212 12962 37268 13582
rect 37212 12910 37214 12962
rect 37266 12910 37268 12962
rect 35768 12572 36448 12582
rect 35824 12516 35872 12572
rect 35928 12570 35976 12572
rect 36032 12570 36080 12572
rect 35948 12518 35976 12570
rect 36072 12518 36080 12570
rect 35928 12516 35976 12518
rect 36032 12516 36080 12518
rect 36136 12570 36184 12572
rect 36240 12570 36288 12572
rect 36136 12518 36144 12570
rect 36240 12518 36268 12570
rect 36136 12516 36184 12518
rect 36240 12516 36288 12518
rect 36344 12516 36392 12572
rect 35768 12506 36448 12516
rect 36876 12066 36932 12078
rect 36876 12014 36878 12066
rect 36930 12014 36932 12066
rect 35768 11004 36448 11014
rect 35824 10948 35872 11004
rect 35928 11002 35976 11004
rect 36032 11002 36080 11004
rect 35948 10950 35976 11002
rect 36072 10950 36080 11002
rect 35928 10948 35976 10950
rect 36032 10948 36080 10950
rect 36136 11002 36184 11004
rect 36240 11002 36288 11004
rect 36136 10950 36144 11002
rect 36240 10950 36268 11002
rect 36136 10948 36184 10950
rect 36240 10948 36288 10950
rect 36344 10948 36392 11004
rect 35768 10938 36448 10948
rect 35308 10610 35364 10622
rect 35308 10558 35310 10610
rect 35362 10558 35364 10610
rect 35308 9044 35364 10558
rect 35308 8978 35364 8988
rect 35420 9826 35476 9838
rect 35420 9774 35422 9826
rect 35474 9774 35476 9826
rect 34972 6290 35028 6300
rect 35084 7476 35140 7486
rect 34860 6078 34862 6130
rect 34914 6078 34916 6130
rect 34860 6066 34916 6078
rect 34748 5908 34804 5918
rect 34188 5854 34190 5906
rect 34242 5854 34244 5906
rect 34188 5842 34244 5854
rect 34524 5906 34804 5908
rect 34524 5854 34750 5906
rect 34802 5854 34804 5906
rect 34524 5852 34804 5854
rect 34524 5794 34580 5852
rect 34524 5742 34526 5794
rect 34578 5742 34580 5794
rect 34524 5730 34580 5742
rect 34300 5684 34356 5694
rect 34076 5682 34356 5684
rect 34076 5630 34302 5682
rect 34354 5630 34356 5682
rect 34076 5628 34356 5630
rect 34300 5618 34356 5628
rect 34748 5460 34804 5852
rect 34972 5460 35028 5470
rect 33964 5404 34356 5460
rect 34076 5236 34132 5246
rect 33852 5012 33908 5022
rect 33908 4956 34020 5012
rect 33852 4946 33908 4956
rect 33740 4396 33908 4452
rect 33852 4340 33908 4396
rect 33628 4284 33796 4340
rect 33404 4174 33406 4226
rect 33458 4174 33460 4226
rect 33404 4162 33460 4174
rect 33740 4114 33796 4284
rect 33852 4246 33908 4284
rect 33740 4062 33742 4114
rect 33794 4062 33796 4114
rect 33740 4050 33796 4062
rect 33292 3948 33460 4004
rect 33068 3614 33070 3666
rect 33122 3614 33124 3666
rect 33068 3602 33124 3614
rect 33292 3780 33348 3790
rect 32508 3490 32564 3500
rect 33292 3554 33348 3724
rect 33404 3666 33460 3948
rect 33404 3614 33406 3666
rect 33458 3614 33460 3666
rect 33404 3602 33460 3614
rect 33292 3502 33294 3554
rect 33346 3502 33348 3554
rect 6636 3390 6638 3442
rect 6690 3390 6692 3442
rect 6636 3378 6692 3390
rect 16492 3444 16548 3454
rect 16492 3442 16884 3444
rect 16492 3390 16494 3442
rect 16546 3390 16884 3442
rect 16492 3388 16884 3390
rect 16492 3378 16548 3388
rect 16828 3332 16884 3388
rect 17276 3442 17332 3454
rect 17276 3390 17278 3442
rect 17330 3390 17332 3442
rect 17276 3332 17332 3390
rect 27916 3444 27972 3454
rect 28364 3444 28420 3454
rect 27916 3442 28420 3444
rect 27916 3390 27918 3442
rect 27970 3390 28366 3442
rect 28418 3390 28420 3442
rect 27916 3388 28420 3390
rect 27916 3378 27972 3388
rect 16828 3276 17332 3332
rect 8768 3164 9448 3174
rect 8824 3108 8872 3164
rect 8928 3162 8976 3164
rect 9032 3162 9080 3164
rect 8948 3110 8976 3162
rect 9072 3110 9080 3162
rect 8928 3108 8976 3110
rect 9032 3108 9080 3110
rect 9136 3162 9184 3164
rect 9240 3162 9288 3164
rect 9136 3110 9144 3162
rect 9240 3110 9268 3162
rect 9136 3108 9184 3110
rect 9240 3108 9288 3110
rect 9344 3108 9392 3164
rect 8768 3098 9448 3108
rect 17052 800 17108 3276
rect 17768 3164 18448 3174
rect 17824 3108 17872 3164
rect 17928 3162 17976 3164
rect 18032 3162 18080 3164
rect 17948 3110 17976 3162
rect 18072 3110 18080 3162
rect 17928 3108 17976 3110
rect 18032 3108 18080 3110
rect 18136 3162 18184 3164
rect 18240 3162 18288 3164
rect 18136 3110 18144 3162
rect 18240 3110 18268 3162
rect 18136 3108 18184 3110
rect 18240 3108 18288 3110
rect 18344 3108 18392 3164
rect 17768 3098 18448 3108
rect 26768 3164 27448 3174
rect 26824 3108 26872 3164
rect 26928 3162 26976 3164
rect 27032 3162 27080 3164
rect 26948 3110 26976 3162
rect 27072 3110 27080 3162
rect 26928 3108 26976 3110
rect 27032 3108 27080 3110
rect 27136 3162 27184 3164
rect 27240 3162 27288 3164
rect 27136 3110 27144 3162
rect 27240 3110 27268 3162
rect 27136 3108 27184 3110
rect 27240 3108 27288 3110
rect 27344 3108 27392 3164
rect 26768 3098 27448 3108
rect 28028 800 28084 3388
rect 28364 3378 28420 3388
rect 33292 3388 33348 3502
rect 33628 3442 33684 3454
rect 33628 3390 33630 3442
rect 33682 3390 33684 3442
rect 33628 3388 33684 3390
rect 33292 3332 33684 3388
rect 33964 3442 34020 4956
rect 34076 4450 34132 5180
rect 34076 4398 34078 4450
rect 34130 4398 34132 4450
rect 34076 4386 34132 4398
rect 34188 4340 34244 4350
rect 34188 3778 34244 4284
rect 34188 3726 34190 3778
rect 34242 3726 34244 3778
rect 34188 3556 34244 3726
rect 34300 3778 34356 5404
rect 34524 5404 34972 5460
rect 34412 5236 34468 5246
rect 34412 5142 34468 5180
rect 34524 4788 34580 5404
rect 34972 5394 35028 5404
rect 34412 4732 34580 4788
rect 34636 5292 34916 5348
rect 34412 4450 34468 4732
rect 34524 4564 34580 4574
rect 34636 4564 34692 5292
rect 34860 5236 34916 5292
rect 35084 5236 35140 7420
rect 35420 5348 35476 9774
rect 35532 9716 35588 9726
rect 35532 9042 35588 9660
rect 35768 9436 36448 9446
rect 35824 9380 35872 9436
rect 35928 9434 35976 9436
rect 36032 9434 36080 9436
rect 35948 9382 35976 9434
rect 36072 9382 36080 9434
rect 35928 9380 35976 9382
rect 36032 9380 36080 9382
rect 36136 9434 36184 9436
rect 36240 9434 36288 9436
rect 36136 9382 36144 9434
rect 36240 9382 36268 9434
rect 36136 9380 36184 9382
rect 36240 9380 36288 9382
rect 36344 9380 36392 9436
rect 35768 9370 36448 9380
rect 36876 9380 36932 12014
rect 36876 9324 37156 9380
rect 35532 8990 35534 9042
rect 35586 8990 35588 9042
rect 35532 8978 35588 8990
rect 36428 9268 36484 9278
rect 36428 8258 36484 9212
rect 36428 8206 36430 8258
rect 36482 8206 36484 8258
rect 36428 8194 36484 8206
rect 35768 7868 36448 7878
rect 35824 7812 35872 7868
rect 35928 7866 35976 7868
rect 36032 7866 36080 7868
rect 35948 7814 35976 7866
rect 36072 7814 36080 7866
rect 35928 7812 35976 7814
rect 36032 7812 36080 7814
rect 36136 7866 36184 7868
rect 36240 7866 36288 7868
rect 36136 7814 36144 7866
rect 36240 7814 36268 7866
rect 36136 7812 36184 7814
rect 36240 7812 36288 7814
rect 36344 7812 36392 7868
rect 35768 7802 36448 7812
rect 37100 6914 37156 9324
rect 37212 9268 37268 12910
rect 37660 11284 37716 11294
rect 37548 11228 37660 11284
rect 37436 9828 37492 9838
rect 37212 9202 37268 9212
rect 37324 9772 37436 9828
rect 37212 8930 37268 8942
rect 37212 8878 37214 8930
rect 37266 8878 37268 8930
rect 37212 7588 37268 8878
rect 37212 7522 37268 7532
rect 37324 7364 37380 9772
rect 37436 9762 37492 9772
rect 37100 6862 37102 6914
rect 37154 6862 37156 6914
rect 37100 6850 37156 6862
rect 37212 7308 37380 7364
rect 37436 8148 37492 8158
rect 35644 6690 35700 6702
rect 37212 6692 37268 7308
rect 37324 6916 37380 6926
rect 37324 6822 37380 6860
rect 37436 6914 37492 8092
rect 37436 6862 37438 6914
rect 37490 6862 37492 6914
rect 37436 6850 37492 6862
rect 35644 6638 35646 6690
rect 35698 6638 35700 6690
rect 35644 6020 35700 6638
rect 37100 6636 37268 6692
rect 36988 6578 37044 6590
rect 36988 6526 36990 6578
rect 37042 6526 37044 6578
rect 35768 6300 36448 6310
rect 35824 6244 35872 6300
rect 35928 6298 35976 6300
rect 36032 6298 36080 6300
rect 35948 6246 35976 6298
rect 36072 6246 36080 6298
rect 35928 6244 35976 6246
rect 36032 6244 36080 6246
rect 36136 6298 36184 6300
rect 36240 6298 36288 6300
rect 36136 6246 36144 6298
rect 36240 6246 36268 6298
rect 36136 6244 36184 6246
rect 36240 6244 36288 6246
rect 36344 6244 36392 6300
rect 35768 6234 36448 6244
rect 35644 5926 35700 5964
rect 36540 5460 36596 5470
rect 35420 5282 35476 5292
rect 36428 5348 36484 5358
rect 34860 5180 35140 5236
rect 34524 4562 34692 4564
rect 34524 4510 34526 4562
rect 34578 4510 34692 4562
rect 34524 4508 34692 4510
rect 34748 5124 34804 5134
rect 34524 4498 34580 4508
rect 34412 4398 34414 4450
rect 34466 4398 34468 4450
rect 34412 4340 34468 4398
rect 34636 4340 34692 4350
rect 34412 4284 34636 4340
rect 34636 4246 34692 4284
rect 34300 3726 34302 3778
rect 34354 3726 34356 3778
rect 34300 3714 34356 3726
rect 34636 3780 34692 3790
rect 34748 3780 34804 5068
rect 36428 5122 36484 5292
rect 36428 5070 36430 5122
rect 36482 5070 36484 5122
rect 36428 5058 36484 5070
rect 35768 4732 36448 4742
rect 35824 4676 35872 4732
rect 35928 4730 35976 4732
rect 36032 4730 36080 4732
rect 35948 4678 35976 4730
rect 36072 4678 36080 4730
rect 35928 4676 35976 4678
rect 36032 4676 36080 4678
rect 36136 4730 36184 4732
rect 36240 4730 36288 4732
rect 36136 4678 36144 4730
rect 36240 4678 36268 4730
rect 36136 4676 36184 4678
rect 36240 4676 36288 4678
rect 36344 4676 36392 4732
rect 35768 4666 36448 4676
rect 34636 3778 34804 3780
rect 34636 3726 34638 3778
rect 34690 3726 34804 3778
rect 34636 3724 34804 3726
rect 35196 4340 35252 4350
rect 34636 3714 34692 3724
rect 35196 3666 35252 4284
rect 35196 3614 35198 3666
rect 35250 3614 35252 3666
rect 35196 3602 35252 3614
rect 36540 3666 36596 5404
rect 36988 5122 37044 6526
rect 36988 5070 36990 5122
rect 37042 5070 37044 5122
rect 36988 5058 37044 5070
rect 37100 4898 37156 6636
rect 37212 5348 37268 5358
rect 37548 5348 37604 11228
rect 37660 11218 37716 11228
rect 38108 10498 38164 10510
rect 38108 10446 38110 10498
rect 38162 10446 38164 10498
rect 37996 6466 38052 6478
rect 37996 6414 37998 6466
rect 38050 6414 38052 6466
rect 37996 5460 38052 6414
rect 37996 5394 38052 5404
rect 37212 5346 37604 5348
rect 37212 5294 37214 5346
rect 37266 5294 37604 5346
rect 37212 5292 37604 5294
rect 37212 5282 37268 5292
rect 37436 5124 37492 5134
rect 37884 5124 37940 5134
rect 37436 5122 37940 5124
rect 37436 5070 37438 5122
rect 37490 5070 37886 5122
rect 37938 5070 37940 5122
rect 37436 5068 37940 5070
rect 37436 5058 37492 5068
rect 37884 5058 37940 5068
rect 37996 5124 38052 5134
rect 38108 5124 38164 10446
rect 37996 5122 38164 5124
rect 37996 5070 37998 5122
rect 38050 5070 38164 5122
rect 37996 5068 38164 5070
rect 37996 5058 38052 5068
rect 37100 4846 37102 4898
rect 37154 4846 37156 4898
rect 37100 4834 37156 4846
rect 38220 3892 38276 15092
rect 40268 14924 40948 14934
rect 40324 14868 40372 14924
rect 40428 14922 40476 14924
rect 40532 14922 40580 14924
rect 40448 14870 40476 14922
rect 40572 14870 40580 14922
rect 40428 14868 40476 14870
rect 40532 14868 40580 14870
rect 40636 14922 40684 14924
rect 40740 14922 40788 14924
rect 40636 14870 40644 14922
rect 40740 14870 40768 14922
rect 40636 14868 40684 14870
rect 40740 14868 40788 14870
rect 40844 14868 40892 14924
rect 40268 14858 40948 14868
rect 40268 13356 40948 13366
rect 40324 13300 40372 13356
rect 40428 13354 40476 13356
rect 40532 13354 40580 13356
rect 40448 13302 40476 13354
rect 40572 13302 40580 13354
rect 40428 13300 40476 13302
rect 40532 13300 40580 13302
rect 40636 13354 40684 13356
rect 40740 13354 40788 13356
rect 40636 13302 40644 13354
rect 40740 13302 40768 13354
rect 40636 13300 40684 13302
rect 40740 13300 40788 13302
rect 40844 13300 40892 13356
rect 40268 13290 40948 13300
rect 40012 12178 40068 12190
rect 40012 12126 40014 12178
rect 40066 12126 40068 12178
rect 39004 11396 39060 11406
rect 39004 11302 39060 11340
rect 39004 9828 39060 9838
rect 39004 9734 39060 9772
rect 40012 9716 40068 12126
rect 40268 11788 40948 11798
rect 40324 11732 40372 11788
rect 40428 11786 40476 11788
rect 40532 11786 40580 11788
rect 40448 11734 40476 11786
rect 40572 11734 40580 11786
rect 40428 11732 40476 11734
rect 40532 11732 40580 11734
rect 40636 11786 40684 11788
rect 40740 11786 40788 11788
rect 40636 11734 40644 11786
rect 40740 11734 40768 11786
rect 40636 11732 40684 11734
rect 40740 11732 40788 11734
rect 40844 11732 40892 11788
rect 40268 11722 40948 11732
rect 41020 11284 41076 11294
rect 41020 11190 41076 11228
rect 40268 10220 40948 10230
rect 40324 10164 40372 10220
rect 40428 10218 40476 10220
rect 40532 10218 40580 10220
rect 40448 10166 40476 10218
rect 40572 10166 40580 10218
rect 40428 10164 40476 10166
rect 40532 10164 40580 10166
rect 40636 10218 40684 10220
rect 40740 10218 40788 10220
rect 40636 10166 40644 10218
rect 40740 10166 40768 10218
rect 40636 10164 40684 10166
rect 40740 10164 40788 10166
rect 40844 10164 40892 10220
rect 40268 10154 40948 10164
rect 40012 8258 40068 9660
rect 41020 9716 41076 9726
rect 41020 9622 41076 9660
rect 40268 8652 40948 8662
rect 40324 8596 40372 8652
rect 40428 8650 40476 8652
rect 40532 8650 40580 8652
rect 40448 8598 40476 8650
rect 40572 8598 40580 8650
rect 40428 8596 40476 8598
rect 40532 8596 40580 8598
rect 40636 8650 40684 8652
rect 40740 8650 40788 8652
rect 40636 8598 40644 8650
rect 40740 8598 40768 8650
rect 40636 8596 40684 8598
rect 40740 8596 40788 8598
rect 40844 8596 40892 8652
rect 40268 8586 40948 8596
rect 40012 8206 40014 8258
rect 40066 8206 40068 8258
rect 40012 8194 40068 8206
rect 40124 7474 40180 7486
rect 40124 7422 40126 7474
rect 40178 7422 40180 7474
rect 38332 7364 38388 7374
rect 38332 7270 38388 7308
rect 40124 6804 40180 7422
rect 41020 7252 41076 7262
rect 40268 7084 40948 7094
rect 40324 7028 40372 7084
rect 40428 7082 40476 7084
rect 40532 7082 40580 7084
rect 40448 7030 40476 7082
rect 40572 7030 40580 7082
rect 40428 7028 40476 7030
rect 40532 7028 40580 7030
rect 40636 7082 40684 7084
rect 40740 7082 40788 7084
rect 40636 7030 40644 7082
rect 40740 7030 40768 7082
rect 40636 7028 40684 7030
rect 40740 7028 40788 7030
rect 40844 7028 40892 7084
rect 40268 7018 40948 7028
rect 40124 6738 40180 6748
rect 40908 6692 40964 6702
rect 40908 6018 40964 6636
rect 41020 6130 41076 7196
rect 41020 6078 41022 6130
rect 41074 6078 41076 6130
rect 41020 6066 41076 6078
rect 40908 5966 40910 6018
rect 40962 5966 40964 6018
rect 40908 5954 40964 5966
rect 40124 5906 40180 5918
rect 40124 5854 40126 5906
rect 40178 5854 40180 5906
rect 38780 5460 38836 5470
rect 38668 4898 38724 4910
rect 38668 4846 38670 4898
rect 38722 4846 38724 4898
rect 38332 4452 38388 4462
rect 38332 4358 38388 4396
rect 38220 3826 38276 3836
rect 36540 3614 36542 3666
rect 36594 3614 36596 3666
rect 36540 3602 36596 3614
rect 37100 3778 37156 3790
rect 37100 3726 37102 3778
rect 37154 3726 37156 3778
rect 34748 3556 34804 3566
rect 34188 3500 34748 3556
rect 34748 3462 34804 3500
rect 36092 3556 36148 3566
rect 36092 3462 36148 3500
rect 33964 3390 33966 3442
rect 34018 3390 34020 3442
rect 33964 3378 34020 3390
rect 37100 3442 37156 3726
rect 38556 3778 38612 3790
rect 38556 3726 38558 3778
rect 38610 3726 38612 3778
rect 37436 3556 37492 3566
rect 37436 3462 37492 3500
rect 37884 3556 37940 3566
rect 38332 3556 38388 3566
rect 37940 3500 38332 3556
rect 37884 3462 37940 3500
rect 38332 3462 38388 3500
rect 37100 3390 37102 3442
rect 37154 3390 37156 3442
rect 37100 3378 37156 3390
rect 38556 3444 38612 3726
rect 38668 3668 38724 4846
rect 38668 3602 38724 3612
rect 38780 4116 38836 5404
rect 38780 3666 38836 4060
rect 39228 5012 39284 5022
rect 38780 3614 38782 3666
rect 38834 3614 38836 3666
rect 38780 3602 38836 3614
rect 39116 3780 39172 3790
rect 39116 3554 39172 3724
rect 39228 3778 39284 4956
rect 40124 4564 40180 5854
rect 40268 5516 40948 5526
rect 40324 5460 40372 5516
rect 40428 5514 40476 5516
rect 40532 5514 40580 5516
rect 40448 5462 40476 5514
rect 40572 5462 40580 5514
rect 40428 5460 40476 5462
rect 40532 5460 40580 5462
rect 40636 5514 40684 5516
rect 40740 5514 40788 5516
rect 40636 5462 40644 5514
rect 40740 5462 40768 5514
rect 40636 5460 40684 5462
rect 40740 5460 40788 5462
rect 40844 5460 40892 5516
rect 40268 5450 40948 5460
rect 41132 4676 41188 15092
rect 41468 12850 41524 12862
rect 41468 12798 41470 12850
rect 41522 12798 41524 12850
rect 41244 7588 41300 7598
rect 41244 7586 41412 7588
rect 41244 7534 41246 7586
rect 41298 7534 41412 7586
rect 41244 7532 41412 7534
rect 41244 7522 41300 7532
rect 41132 4610 41188 4620
rect 41244 6580 41300 6590
rect 40124 4498 40180 4508
rect 40236 4340 40292 4350
rect 40236 4246 40292 4284
rect 41132 4228 41188 4238
rect 41020 4116 41076 4126
rect 41132 4116 41188 4172
rect 41020 4114 41188 4116
rect 41020 4062 41022 4114
rect 41074 4062 41188 4114
rect 41020 4060 41188 4062
rect 41020 4050 41076 4060
rect 40268 3948 40948 3958
rect 40324 3892 40372 3948
rect 40428 3946 40476 3948
rect 40532 3946 40580 3948
rect 40448 3894 40476 3946
rect 40572 3894 40580 3946
rect 40428 3892 40476 3894
rect 40532 3892 40580 3894
rect 40636 3946 40684 3948
rect 40740 3946 40788 3948
rect 40636 3894 40644 3946
rect 40740 3894 40768 3946
rect 40636 3892 40684 3894
rect 40740 3892 40788 3894
rect 40844 3892 40892 3948
rect 40268 3882 40948 3892
rect 39228 3726 39230 3778
rect 39282 3726 39284 3778
rect 39228 3714 39284 3726
rect 41020 3780 41076 3790
rect 41020 3686 41076 3724
rect 40908 3668 40964 3678
rect 40908 3574 40964 3612
rect 39116 3502 39118 3554
rect 39170 3502 39172 3554
rect 39116 3490 39172 3502
rect 40348 3556 40404 3566
rect 38556 3378 38612 3388
rect 39004 3444 39060 3454
rect 35768 3164 36448 3174
rect 35824 3108 35872 3164
rect 35928 3162 35976 3164
rect 36032 3162 36080 3164
rect 35948 3110 35976 3162
rect 36072 3110 36080 3162
rect 35928 3108 35976 3110
rect 36032 3108 36080 3110
rect 36136 3162 36184 3164
rect 36240 3162 36288 3164
rect 36136 3110 36144 3162
rect 36240 3110 36268 3162
rect 36136 3108 36184 3110
rect 36240 3108 36288 3110
rect 36344 3108 36392 3164
rect 35768 3098 36448 3108
rect 39004 800 39060 3388
rect 39788 3444 39844 3482
rect 40348 3462 40404 3500
rect 39788 3378 39844 3388
rect 41244 3442 41300 6524
rect 41356 4338 41412 7532
rect 41468 6468 41524 12798
rect 41692 7252 41748 7262
rect 41468 6402 41524 6412
rect 41580 7250 41748 7252
rect 41580 7198 41694 7250
rect 41746 7198 41748 7250
rect 41580 7196 41748 7198
rect 41580 4900 41636 7196
rect 41692 7186 41748 7196
rect 41692 6132 41748 6142
rect 41692 6038 41748 6076
rect 41580 4834 41636 4844
rect 41692 5236 41748 5246
rect 41356 4286 41358 4338
rect 41410 4286 41412 4338
rect 41356 4274 41412 4286
rect 41468 4788 41524 4798
rect 41468 4338 41524 4732
rect 41468 4286 41470 4338
rect 41522 4286 41524 4338
rect 41468 3780 41524 4286
rect 41468 3714 41524 3724
rect 41580 4676 41636 4686
rect 41580 3556 41636 4620
rect 41692 4450 41748 5180
rect 41692 4398 41694 4450
rect 41746 4398 41748 4450
rect 41692 4386 41748 4398
rect 41804 4228 41860 15260
rect 42028 7588 42084 19070
rect 42252 15428 42308 15438
rect 42140 15426 42308 15428
rect 42140 15374 42254 15426
rect 42306 15374 42308 15426
rect 42140 15372 42308 15374
rect 42140 8820 42196 15372
rect 42252 15362 42308 15372
rect 43036 15314 43092 15326
rect 43036 15262 43038 15314
rect 43090 15262 43092 15314
rect 43036 15204 43092 15262
rect 43932 15204 43988 15214
rect 43036 15138 43092 15148
rect 43820 15202 43988 15204
rect 43820 15150 43934 15202
rect 43986 15150 43988 15202
rect 43820 15148 43988 15150
rect 44380 15148 44436 24668
rect 44768 23548 45448 23558
rect 44824 23492 44872 23548
rect 44928 23546 44976 23548
rect 45032 23546 45080 23548
rect 44948 23494 44976 23546
rect 45072 23494 45080 23546
rect 44928 23492 44976 23494
rect 45032 23492 45080 23494
rect 45136 23546 45184 23548
rect 45240 23546 45288 23548
rect 45136 23494 45144 23546
rect 45240 23494 45268 23546
rect 45136 23492 45184 23494
rect 45240 23492 45288 23494
rect 45344 23492 45392 23548
rect 44768 23482 45448 23492
rect 46060 23266 46116 23278
rect 46060 23214 46062 23266
rect 46114 23214 46116 23266
rect 45164 23156 45220 23166
rect 45164 23062 45220 23100
rect 45948 23154 46004 23166
rect 45948 23102 45950 23154
rect 46002 23102 46004 23154
rect 45612 23044 45668 23054
rect 45948 23044 46004 23102
rect 46060 23156 46116 23214
rect 46060 23090 46116 23100
rect 46284 23154 46340 23166
rect 46284 23102 46286 23154
rect 46338 23102 46340 23154
rect 45612 23042 46004 23044
rect 45612 22990 45614 23042
rect 45666 22990 46004 23042
rect 45612 22988 46004 22990
rect 44768 21980 45448 21990
rect 44824 21924 44872 21980
rect 44928 21978 44976 21980
rect 45032 21978 45080 21980
rect 44948 21926 44976 21978
rect 45072 21926 45080 21978
rect 44928 21924 44976 21926
rect 45032 21924 45080 21926
rect 45136 21978 45184 21980
rect 45240 21978 45288 21980
rect 45136 21926 45144 21978
rect 45240 21926 45268 21978
rect 45136 21924 45184 21926
rect 45240 21924 45288 21926
rect 45344 21924 45392 21980
rect 44768 21914 45448 21924
rect 45612 21476 45668 22988
rect 46284 22596 46340 23102
rect 46284 22530 46340 22540
rect 45612 21410 45668 21420
rect 44768 20412 45448 20422
rect 44824 20356 44872 20412
rect 44928 20410 44976 20412
rect 45032 20410 45080 20412
rect 44948 20358 44976 20410
rect 45072 20358 45080 20410
rect 44928 20356 44976 20358
rect 45032 20356 45080 20358
rect 45136 20410 45184 20412
rect 45240 20410 45288 20412
rect 45136 20358 45144 20410
rect 45240 20358 45268 20410
rect 45136 20356 45184 20358
rect 45240 20356 45288 20358
rect 45344 20356 45392 20412
rect 44768 20346 45448 20356
rect 44768 18844 45448 18854
rect 44824 18788 44872 18844
rect 44928 18842 44976 18844
rect 45032 18842 45080 18844
rect 44948 18790 44976 18842
rect 45072 18790 45080 18842
rect 44928 18788 44976 18790
rect 45032 18788 45080 18790
rect 45136 18842 45184 18844
rect 45240 18842 45288 18844
rect 45136 18790 45144 18842
rect 45240 18790 45268 18842
rect 45136 18788 45184 18790
rect 45240 18788 45288 18790
rect 45344 18788 45392 18844
rect 44768 18778 45448 18788
rect 44768 17276 45448 17286
rect 44824 17220 44872 17276
rect 44928 17274 44976 17276
rect 45032 17274 45080 17276
rect 44948 17222 44976 17274
rect 45072 17222 45080 17274
rect 44928 17220 44976 17222
rect 45032 17220 45080 17222
rect 45136 17274 45184 17276
rect 45240 17274 45288 17276
rect 45136 17222 45144 17274
rect 45240 17222 45268 17274
rect 45136 17220 45184 17222
rect 45240 17220 45288 17222
rect 45344 17220 45392 17276
rect 44768 17210 45448 17220
rect 44768 15708 45448 15718
rect 44824 15652 44872 15708
rect 44928 15706 44976 15708
rect 45032 15706 45080 15708
rect 44948 15654 44976 15706
rect 45072 15654 45080 15706
rect 44928 15652 44976 15654
rect 45032 15652 45080 15654
rect 45136 15706 45184 15708
rect 45240 15706 45288 15708
rect 45136 15654 45144 15706
rect 45240 15654 45268 15706
rect 45136 15652 45184 15654
rect 45240 15652 45288 15654
rect 45344 15652 45392 15708
rect 44768 15642 45448 15652
rect 44604 15428 44660 15438
rect 43148 13746 43204 13758
rect 43148 13694 43150 13746
rect 43202 13694 43204 13746
rect 42700 12180 42756 12190
rect 42700 12178 42868 12180
rect 42700 12126 42702 12178
rect 42754 12126 42868 12178
rect 42700 12124 42868 12126
rect 42700 12114 42756 12124
rect 42476 9380 42532 9390
rect 42364 9324 42476 9380
rect 42140 8764 42308 8820
rect 41916 7532 42084 7588
rect 41916 7028 41972 7532
rect 42140 7476 42196 7486
rect 42140 7382 42196 7420
rect 41916 6972 42196 7028
rect 41916 6804 41972 6814
rect 41916 6578 41972 6748
rect 41916 6526 41918 6578
rect 41970 6526 41972 6578
rect 41916 6514 41972 6526
rect 42028 6132 42084 6142
rect 41804 4162 41860 4172
rect 41916 5124 41972 5134
rect 41916 3666 41972 5068
rect 42028 4452 42084 6076
rect 42140 6130 42196 6972
rect 42140 6078 42142 6130
rect 42194 6078 42196 6130
rect 42140 4788 42196 6078
rect 42252 5460 42308 8764
rect 42364 7476 42420 9324
rect 42476 9314 42532 9324
rect 42700 8932 42756 8942
rect 42700 8838 42756 8876
rect 42812 7812 42868 12124
rect 42700 7756 42868 7812
rect 43036 11284 43092 11294
rect 42476 7700 42532 7710
rect 42476 7698 42644 7700
rect 42476 7646 42478 7698
rect 42530 7646 42644 7698
rect 42476 7644 42644 7646
rect 42476 7634 42532 7644
rect 42476 7476 42532 7486
rect 42364 7474 42532 7476
rect 42364 7422 42478 7474
rect 42530 7422 42532 7474
rect 42364 7420 42532 7422
rect 42476 7410 42532 7420
rect 42364 7252 42420 7262
rect 42364 7158 42420 7196
rect 42588 6356 42644 7644
rect 42476 6300 42644 6356
rect 42476 5572 42532 6300
rect 42588 6132 42644 6142
rect 42588 6038 42644 6076
rect 42476 5516 42644 5572
rect 42252 5404 42532 5460
rect 42252 5236 42308 5246
rect 42252 5142 42308 5180
rect 42476 5012 42532 5404
rect 42476 4946 42532 4956
rect 42140 4722 42196 4732
rect 42364 4564 42420 4574
rect 42252 4452 42308 4462
rect 42028 4450 42308 4452
rect 42028 4398 42030 4450
rect 42082 4398 42254 4450
rect 42306 4398 42308 4450
rect 42028 4396 42308 4398
rect 42028 4116 42084 4396
rect 42252 4386 42308 4396
rect 42364 4226 42420 4508
rect 42364 4174 42366 4226
rect 42418 4174 42420 4226
rect 42364 4162 42420 4174
rect 42028 4050 42084 4060
rect 42252 3780 42308 3790
rect 42588 3780 42644 5516
rect 42308 3724 42532 3780
rect 42252 3714 42308 3724
rect 41916 3614 41918 3666
rect 41970 3614 41972 3666
rect 41916 3602 41972 3614
rect 41804 3556 41860 3566
rect 41636 3554 41860 3556
rect 41636 3502 41806 3554
rect 41858 3502 41860 3554
rect 41636 3500 41860 3502
rect 41580 3462 41636 3500
rect 41804 3490 41860 3500
rect 42476 3554 42532 3724
rect 42588 3714 42644 3724
rect 42476 3502 42478 3554
rect 42530 3502 42532 3554
rect 42476 3490 42532 3502
rect 41244 3390 41246 3442
rect 41298 3390 41300 3442
rect 41244 3378 41300 3390
rect 42588 3444 42644 3482
rect 42588 3378 42644 3388
rect 42700 3220 42756 7756
rect 42924 7474 42980 7486
rect 42924 7422 42926 7474
rect 42978 7422 42980 7474
rect 42924 5236 42980 7422
rect 42924 5170 42980 5180
rect 42812 5124 42868 5134
rect 42812 5030 42868 5068
rect 43036 5012 43092 11228
rect 42924 4956 43092 5012
rect 43148 9042 43204 13694
rect 43708 10498 43764 10510
rect 43708 10446 43710 10498
rect 43762 10446 43764 10498
rect 43708 9380 43764 10446
rect 43708 9314 43764 9324
rect 43148 8990 43150 9042
rect 43202 8990 43204 9042
rect 42924 3554 42980 4956
rect 43148 4452 43204 8990
rect 43148 4386 43204 4396
rect 43484 4900 43540 4910
rect 42924 3502 42926 3554
rect 42978 3502 42980 3554
rect 42924 3490 42980 3502
rect 43036 3556 43092 3566
rect 43036 3330 43092 3500
rect 43484 3554 43540 4844
rect 43820 4340 43876 15148
rect 43932 15138 43988 15148
rect 44268 15092 44436 15148
rect 44492 15426 44884 15428
rect 44492 15374 44606 15426
rect 44658 15374 44884 15426
rect 44492 15372 44884 15374
rect 44268 14420 44324 15092
rect 44268 14308 44324 14364
rect 44156 14306 44324 14308
rect 44156 14254 44270 14306
rect 44322 14254 44324 14306
rect 44156 14252 44324 14254
rect 44156 8932 44212 14252
rect 44268 14242 44324 14252
rect 44156 8866 44212 8876
rect 44268 13634 44324 13646
rect 44268 13582 44270 13634
rect 44322 13582 44324 13634
rect 44044 8148 44100 8158
rect 44044 8054 44100 8092
rect 44268 7588 44324 13582
rect 44380 12068 44436 12078
rect 44380 11974 44436 12012
rect 43820 4274 43876 4284
rect 44044 7532 44324 7588
rect 44044 3778 44100 7532
rect 44156 7364 44212 7374
rect 44156 4450 44212 7308
rect 44492 6804 44548 15372
rect 44604 15362 44660 15372
rect 44828 15314 44884 15372
rect 44828 15262 44830 15314
rect 44882 15262 44884 15314
rect 44828 15250 44884 15262
rect 46620 14642 46676 33292
rect 46844 32228 46900 34078
rect 46956 34132 47012 34638
rect 47516 34242 47572 35084
rect 47964 34354 48020 36428
rect 47964 34302 47966 34354
rect 48018 34302 48020 34354
rect 47964 34290 48020 34302
rect 47516 34190 47518 34242
rect 47570 34190 47572 34242
rect 47516 34178 47572 34190
rect 47292 34132 47348 34142
rect 46956 34130 47348 34132
rect 46956 34078 47294 34130
rect 47346 34078 47348 34130
rect 46956 34076 47348 34078
rect 47292 33236 47348 34076
rect 47404 34132 47460 34142
rect 47404 34038 47460 34076
rect 47852 33460 47908 33470
rect 47404 33236 47460 33246
rect 47292 33234 47460 33236
rect 47292 33182 47406 33234
rect 47458 33182 47460 33234
rect 47292 33180 47460 33182
rect 47404 33170 47460 33180
rect 47852 32786 47908 33404
rect 48076 33012 48132 36540
rect 48412 36258 48468 36270
rect 48412 36206 48414 36258
rect 48466 36206 48468 36258
rect 48412 36036 48468 36206
rect 48860 36036 48916 40574
rect 48972 40962 49028 40974
rect 48972 40910 48974 40962
rect 49026 40910 49028 40962
rect 48972 37938 49028 40910
rect 48972 37886 48974 37938
rect 49026 37886 49028 37938
rect 48972 37874 49028 37886
rect 49084 38948 49140 44156
rect 49868 44210 49924 44222
rect 49868 44158 49870 44210
rect 49922 44158 49924 44210
rect 49868 44100 49924 44158
rect 49868 44034 49924 44044
rect 49980 43316 50036 44492
rect 50092 43540 50148 43550
rect 50204 43540 50260 45166
rect 51660 44996 51716 45006
rect 51324 44994 51940 44996
rect 51324 44942 51662 44994
rect 51714 44942 51940 44994
rect 51324 44940 51940 44942
rect 51324 44322 51380 44940
rect 51660 44930 51716 44940
rect 51324 44270 51326 44322
rect 51378 44270 51380 44322
rect 51324 44258 51380 44270
rect 51660 44100 51716 44110
rect 50092 43538 50260 43540
rect 50092 43486 50094 43538
rect 50146 43486 50260 43538
rect 50092 43484 50260 43486
rect 50540 44098 51716 44100
rect 50540 44046 51662 44098
rect 51714 44046 51716 44098
rect 50540 44044 51716 44046
rect 50540 43538 50596 44044
rect 51660 44034 51716 44044
rect 50540 43486 50542 43538
rect 50594 43486 50596 43538
rect 50092 43474 50148 43484
rect 50540 43474 50596 43486
rect 49980 43260 50148 43316
rect 49268 43148 49948 43158
rect 49324 43092 49372 43148
rect 49428 43146 49476 43148
rect 49532 43146 49580 43148
rect 49448 43094 49476 43146
rect 49572 43094 49580 43146
rect 49428 43092 49476 43094
rect 49532 43092 49580 43094
rect 49636 43146 49684 43148
rect 49740 43146 49788 43148
rect 49636 43094 49644 43146
rect 49740 43094 49768 43146
rect 49636 43092 49684 43094
rect 49740 43092 49788 43094
rect 49844 43092 49892 43148
rect 49268 43082 49948 43092
rect 49644 42084 49700 42094
rect 49644 41990 49700 42028
rect 50092 41860 50148 43260
rect 50316 41860 50372 41870
rect 50092 41858 50372 41860
rect 50092 41806 50318 41858
rect 50370 41806 50372 41858
rect 50092 41804 50372 41806
rect 49268 41580 49948 41590
rect 49324 41524 49372 41580
rect 49428 41578 49476 41580
rect 49532 41578 49580 41580
rect 49448 41526 49476 41578
rect 49572 41526 49580 41578
rect 49428 41524 49476 41526
rect 49532 41524 49580 41526
rect 49636 41578 49684 41580
rect 49740 41578 49788 41580
rect 49636 41526 49644 41578
rect 49740 41526 49768 41578
rect 49636 41524 49684 41526
rect 49740 41524 49788 41526
rect 49844 41524 49892 41580
rect 49268 41514 49948 41524
rect 49532 41186 49588 41198
rect 49532 41134 49534 41186
rect 49586 41134 49588 41186
rect 49532 41076 49588 41134
rect 49532 41010 49588 41020
rect 49980 40964 50036 40974
rect 50316 40964 50372 41804
rect 51100 41860 51156 41870
rect 50988 41076 51044 41086
rect 50988 40982 51044 41020
rect 49980 40962 50372 40964
rect 49980 40910 49982 40962
rect 50034 40910 50372 40962
rect 49980 40908 50372 40910
rect 50652 40962 50708 40974
rect 50652 40910 50654 40962
rect 50706 40910 50708 40962
rect 49980 40898 50036 40908
rect 49420 40404 49476 40414
rect 49420 40310 49476 40348
rect 50092 40404 50148 40414
rect 50092 40310 50148 40348
rect 49268 40012 49948 40022
rect 49324 39956 49372 40012
rect 49428 40010 49476 40012
rect 49532 40010 49580 40012
rect 49448 39958 49476 40010
rect 49572 39958 49580 40010
rect 49428 39956 49476 39958
rect 49532 39956 49580 39958
rect 49636 40010 49684 40012
rect 49740 40010 49788 40012
rect 49636 39958 49644 40010
rect 49740 39958 49768 40010
rect 49636 39956 49684 39958
rect 49740 39956 49788 39958
rect 49844 39956 49892 40012
rect 49268 39946 49948 39956
rect 49308 38948 49364 38958
rect 49140 38946 49364 38948
rect 49140 38894 49310 38946
rect 49362 38894 49364 38946
rect 49140 38892 49364 38894
rect 48972 37156 49028 37166
rect 48972 37062 49028 37100
rect 49084 37044 49140 38892
rect 49308 38882 49364 38892
rect 50092 38610 50148 38622
rect 50092 38558 50094 38610
rect 50146 38558 50148 38610
rect 49268 38444 49948 38454
rect 49324 38388 49372 38444
rect 49428 38442 49476 38444
rect 49532 38442 49580 38444
rect 49448 38390 49476 38442
rect 49572 38390 49580 38442
rect 49428 38388 49476 38390
rect 49532 38388 49580 38390
rect 49636 38442 49684 38444
rect 49740 38442 49788 38444
rect 49636 38390 49644 38442
rect 49740 38390 49768 38442
rect 49636 38388 49684 38390
rect 49740 38388 49788 38390
rect 49844 38388 49892 38444
rect 49268 38378 49948 38388
rect 49756 38052 49812 38062
rect 49756 37958 49812 37996
rect 49980 37940 50036 37950
rect 50092 37940 50148 38558
rect 49980 37938 50148 37940
rect 49980 37886 49982 37938
rect 50034 37886 50148 37938
rect 49980 37884 50148 37886
rect 50204 38276 50260 40908
rect 50652 40404 50708 40910
rect 50652 40338 50708 40348
rect 49980 37874 50036 37884
rect 49868 37492 49924 37502
rect 50204 37492 50260 38220
rect 49868 37490 50260 37492
rect 49868 37438 49870 37490
rect 49922 37438 50260 37490
rect 49868 37436 50260 37438
rect 50540 39060 50596 39070
rect 50540 38946 50596 39004
rect 50540 38894 50542 38946
rect 50594 38894 50596 38946
rect 49868 37426 49924 37436
rect 50540 37380 50596 38894
rect 50652 37380 50708 37390
rect 50540 37378 50932 37380
rect 50540 37326 50654 37378
rect 50706 37326 50932 37378
rect 50540 37324 50932 37326
rect 50652 37314 50708 37324
rect 50204 37266 50260 37278
rect 50204 37214 50206 37266
rect 50258 37214 50260 37266
rect 49420 37156 49476 37166
rect 50204 37156 50260 37214
rect 50428 37266 50484 37278
rect 50428 37214 50430 37266
rect 50482 37214 50484 37266
rect 49420 37154 50260 37156
rect 49420 37102 49422 37154
rect 49474 37102 50260 37154
rect 49420 37100 50260 37102
rect 49420 37044 49476 37100
rect 49084 36988 49476 37044
rect 48412 35980 48916 36036
rect 48972 36258 49028 36270
rect 48972 36206 48974 36258
rect 49026 36206 49028 36258
rect 48412 34804 48468 34814
rect 48412 34710 48468 34748
rect 48524 34132 48580 34142
rect 48524 33348 48580 34076
rect 48300 33346 48580 33348
rect 48300 33294 48526 33346
rect 48578 33294 48580 33346
rect 48300 33292 48580 33294
rect 48300 33124 48356 33292
rect 48524 33282 48580 33292
rect 48748 33236 48804 35980
rect 48972 35698 49028 36206
rect 49084 35812 49140 36988
rect 50204 36932 50260 37100
rect 49268 36876 49948 36886
rect 49324 36820 49372 36876
rect 49428 36874 49476 36876
rect 49532 36874 49580 36876
rect 49448 36822 49476 36874
rect 49572 36822 49580 36874
rect 49428 36820 49476 36822
rect 49532 36820 49580 36822
rect 49636 36874 49684 36876
rect 49740 36874 49788 36876
rect 49636 36822 49644 36874
rect 49740 36822 49768 36874
rect 49636 36820 49684 36822
rect 49740 36820 49788 36822
rect 49844 36820 49892 36876
rect 50204 36866 50260 36876
rect 50316 37156 50372 37166
rect 49268 36810 49948 36820
rect 49084 35746 49140 35756
rect 49756 36596 49812 36606
rect 49756 35810 49812 36540
rect 49756 35758 49758 35810
rect 49810 35758 49812 35810
rect 49756 35746 49812 35758
rect 48972 35646 48974 35698
rect 49026 35646 49028 35698
rect 48972 34692 49028 35646
rect 50316 35364 50372 37100
rect 50428 37156 50484 37214
rect 50428 37090 50484 37100
rect 50876 36596 50932 37324
rect 50876 36502 50932 36540
rect 51100 37044 51156 41804
rect 51884 38834 51940 44940
rect 51996 44212 52052 44222
rect 51996 44118 52052 44156
rect 52668 43652 52724 48412
rect 53228 48468 53284 48478
rect 53228 48374 53284 48412
rect 54460 48468 54516 48478
rect 52892 48018 52948 48030
rect 52892 47966 52894 48018
rect 52946 47966 52948 48018
rect 52892 46452 52948 47966
rect 54460 47570 54516 48412
rect 54460 47518 54462 47570
rect 54514 47518 54516 47570
rect 54460 47348 54516 47518
rect 54460 47282 54516 47292
rect 53768 47068 54448 47078
rect 53824 47012 53872 47068
rect 53928 47066 53976 47068
rect 54032 47066 54080 47068
rect 53948 47014 53976 47066
rect 54072 47014 54080 47066
rect 53928 47012 53976 47014
rect 54032 47012 54080 47014
rect 54136 47066 54184 47068
rect 54240 47066 54288 47068
rect 54136 47014 54144 47066
rect 54240 47014 54268 47066
rect 54136 47012 54184 47014
rect 54240 47012 54288 47014
rect 54344 47012 54392 47068
rect 53768 47002 54448 47012
rect 53564 46900 53620 46910
rect 53004 46788 53060 46798
rect 53564 46788 53620 46844
rect 53004 46786 53620 46788
rect 53004 46734 53006 46786
rect 53058 46734 53566 46786
rect 53618 46734 53620 46786
rect 53004 46732 53620 46734
rect 53004 46722 53060 46732
rect 53564 46722 53620 46732
rect 52892 46386 52948 46396
rect 54124 46676 54180 46686
rect 54124 46002 54180 46620
rect 54572 46676 54628 46686
rect 54236 46564 54292 46574
rect 54236 46450 54292 46508
rect 54236 46398 54238 46450
rect 54290 46398 54292 46450
rect 54236 46386 54292 46398
rect 54124 45950 54126 46002
rect 54178 45950 54180 46002
rect 54124 45892 54180 45950
rect 54124 45826 54180 45836
rect 54460 45668 54516 45706
rect 54460 45602 54516 45612
rect 53768 45500 54448 45510
rect 53452 45444 53508 45454
rect 53824 45444 53872 45500
rect 53928 45498 53976 45500
rect 54032 45498 54080 45500
rect 53948 45446 53976 45498
rect 54072 45446 54080 45498
rect 53928 45444 53976 45446
rect 54032 45444 54080 45446
rect 54136 45498 54184 45500
rect 54240 45498 54288 45500
rect 54136 45446 54144 45498
rect 54240 45446 54268 45498
rect 54136 45444 54184 45446
rect 54240 45444 54288 45446
rect 54344 45444 54392 45500
rect 53508 45388 53620 45444
rect 53768 45434 54448 45444
rect 53452 45378 53508 45388
rect 53564 45332 53620 45388
rect 54460 45332 54516 45342
rect 54572 45332 54628 46620
rect 54684 46562 54740 46574
rect 54684 46510 54686 46562
rect 54738 46510 54740 46562
rect 54684 46450 54740 46510
rect 54684 46398 54686 46450
rect 54738 46398 54740 46450
rect 54684 46386 54740 46398
rect 54796 46228 54852 49644
rect 55132 50372 55300 50428
rect 55020 48804 55076 48814
rect 54908 48802 55076 48804
rect 54908 48750 55022 48802
rect 55074 48750 55076 48802
rect 54908 48748 55076 48750
rect 54908 47458 54964 48748
rect 55020 48738 55076 48748
rect 54908 47406 54910 47458
rect 54962 47406 54964 47458
rect 54908 47394 54964 47406
rect 54908 46228 54964 46238
rect 54796 46172 54908 46228
rect 54908 46162 54964 46172
rect 55020 45892 55076 45930
rect 55020 45826 55076 45836
rect 53564 45276 54180 45332
rect 53564 44884 53620 44894
rect 52892 44100 52948 44110
rect 52780 43652 52836 43662
rect 52668 43596 52780 43652
rect 52668 41074 52724 41086
rect 52668 41022 52670 41074
rect 52722 41022 52724 41074
rect 52220 40964 52276 40974
rect 52668 40964 52724 41022
rect 52220 40962 52724 40964
rect 52220 40910 52222 40962
rect 52274 40910 52724 40962
rect 52220 40908 52724 40910
rect 52220 39396 52276 40908
rect 52780 40852 52836 43596
rect 52556 40796 52836 40852
rect 52556 40626 52612 40796
rect 52556 40574 52558 40626
rect 52610 40574 52612 40626
rect 52556 40562 52612 40574
rect 52220 39330 52276 39340
rect 52556 39396 52612 39406
rect 51884 38782 51886 38834
rect 51938 38782 51940 38834
rect 51884 38668 51940 38782
rect 52444 38722 52500 38734
rect 52444 38670 52446 38722
rect 52498 38670 52500 38722
rect 52444 38668 52500 38670
rect 51884 38612 52500 38668
rect 51548 38164 51604 38174
rect 51548 38070 51604 38108
rect 52108 37490 52164 38612
rect 52556 38052 52612 39340
rect 52892 39060 52948 44044
rect 53228 43652 53284 43662
rect 53228 41410 53284 43596
rect 53564 43650 53620 44828
rect 54124 44434 54180 45276
rect 54460 45330 54628 45332
rect 54460 45278 54462 45330
rect 54514 45278 54628 45330
rect 54460 45276 54628 45278
rect 54460 45266 54516 45276
rect 54572 44548 54628 45276
rect 55020 45668 55076 45678
rect 54908 44884 54964 44894
rect 54572 44492 54740 44548
rect 54124 44382 54126 44434
rect 54178 44382 54180 44434
rect 54124 44324 54180 44382
rect 54124 44258 54180 44268
rect 54572 44212 54628 44222
rect 54572 44118 54628 44156
rect 53768 43932 54448 43942
rect 53824 43876 53872 43932
rect 53928 43930 53976 43932
rect 54032 43930 54080 43932
rect 53948 43878 53976 43930
rect 54072 43878 54080 43930
rect 53928 43876 53976 43878
rect 54032 43876 54080 43878
rect 54136 43930 54184 43932
rect 54240 43930 54288 43932
rect 54136 43878 54144 43930
rect 54240 43878 54268 43930
rect 54136 43876 54184 43878
rect 54240 43876 54288 43878
rect 54344 43876 54392 43932
rect 53768 43866 54448 43876
rect 53564 43598 53566 43650
rect 53618 43598 53620 43650
rect 53564 43586 53620 43598
rect 53900 43652 53956 43662
rect 53900 43558 53956 43596
rect 53768 42364 54448 42374
rect 53824 42308 53872 42364
rect 53928 42362 53976 42364
rect 54032 42362 54080 42364
rect 53948 42310 53976 42362
rect 54072 42310 54080 42362
rect 53928 42308 53976 42310
rect 54032 42308 54080 42310
rect 54136 42362 54184 42364
rect 54240 42362 54288 42364
rect 54136 42310 54144 42362
rect 54240 42310 54268 42362
rect 54136 42308 54184 42310
rect 54240 42308 54288 42310
rect 54344 42308 54392 42364
rect 53768 42298 54448 42308
rect 54684 42084 54740 44492
rect 54908 44546 54964 44828
rect 54908 44494 54910 44546
rect 54962 44494 54964 44546
rect 54908 44482 54964 44494
rect 54236 42028 54740 42084
rect 54796 44324 54852 44334
rect 54236 41970 54292 42028
rect 54236 41918 54238 41970
rect 54290 41918 54292 41970
rect 54236 41906 54292 41918
rect 53228 41358 53230 41410
rect 53282 41358 53284 41410
rect 53228 40740 53284 41358
rect 53340 41858 53396 41870
rect 53340 41806 53342 41858
rect 53394 41806 53396 41858
rect 53340 41412 53396 41806
rect 53788 41860 53844 41870
rect 53788 41766 53844 41804
rect 53340 41346 53396 41356
rect 54572 41186 54628 42028
rect 54572 41134 54574 41186
rect 54626 41134 54628 41186
rect 53564 41076 53620 41086
rect 53228 40684 53508 40740
rect 53228 40516 53284 40526
rect 53116 40404 53172 40414
rect 53116 40310 53172 40348
rect 53228 39732 53284 40460
rect 53452 40404 53508 40684
rect 53564 40628 53620 41020
rect 53768 40796 54448 40806
rect 53824 40740 53872 40796
rect 53928 40794 53976 40796
rect 54032 40794 54080 40796
rect 53948 40742 53976 40794
rect 54072 40742 54080 40794
rect 53928 40740 53976 40742
rect 54032 40740 54080 40742
rect 54136 40794 54184 40796
rect 54240 40794 54288 40796
rect 54136 40742 54144 40794
rect 54240 40742 54268 40794
rect 54136 40740 54184 40742
rect 54240 40740 54288 40742
rect 54344 40740 54392 40796
rect 53768 40730 54448 40740
rect 54572 40740 54628 41134
rect 54684 41858 54740 41870
rect 54684 41806 54686 41858
rect 54738 41806 54740 41858
rect 54684 41076 54740 41806
rect 54684 41010 54740 41020
rect 54572 40684 54740 40740
rect 53676 40628 53732 40638
rect 53564 40626 53732 40628
rect 53564 40574 53678 40626
rect 53730 40574 53732 40626
rect 53564 40572 53732 40574
rect 53676 40562 53732 40572
rect 54572 40514 54628 40526
rect 54572 40462 54574 40514
rect 54626 40462 54628 40514
rect 54012 40404 54068 40414
rect 53452 40348 53732 40404
rect 52892 38966 52948 39004
rect 53116 39730 53284 39732
rect 53116 39678 53230 39730
rect 53282 39678 53284 39730
rect 53116 39676 53284 39678
rect 52108 37438 52110 37490
rect 52162 37438 52164 37490
rect 51548 37266 51604 37278
rect 51548 37214 51550 37266
rect 51602 37214 51604 37266
rect 51212 37156 51268 37166
rect 51548 37156 51604 37214
rect 51268 37100 51604 37156
rect 51212 37062 51268 37100
rect 49268 35308 49948 35318
rect 49324 35252 49372 35308
rect 49428 35306 49476 35308
rect 49532 35306 49580 35308
rect 49448 35254 49476 35306
rect 49572 35254 49580 35306
rect 49428 35252 49476 35254
rect 49532 35252 49580 35254
rect 49636 35306 49684 35308
rect 49740 35306 49788 35308
rect 49636 35254 49644 35306
rect 49740 35254 49768 35306
rect 49636 35252 49684 35254
rect 49740 35252 49788 35254
rect 49844 35252 49892 35308
rect 49268 35242 49948 35252
rect 50092 35308 50372 35364
rect 48972 34626 49028 34636
rect 49084 34804 49140 34814
rect 48860 34018 48916 34030
rect 48860 33966 48862 34018
rect 48914 33966 48916 34018
rect 48860 33460 48916 33966
rect 48860 33346 48916 33404
rect 48860 33294 48862 33346
rect 48914 33294 48916 33346
rect 48860 33282 48916 33294
rect 49084 33236 49140 34748
rect 49868 34802 49924 34814
rect 49868 34750 49870 34802
rect 49922 34750 49924 34802
rect 49308 34692 49364 34702
rect 49308 34130 49364 34636
rect 49868 34692 49924 34750
rect 49868 34626 49924 34636
rect 50092 34356 50148 35308
rect 50316 35140 50372 35150
rect 51100 35140 51156 36988
rect 51436 36932 51492 36942
rect 51436 36484 51492 36876
rect 51548 36708 51604 37100
rect 52108 36932 52164 37438
rect 51996 36820 52052 36830
rect 51996 36708 52052 36764
rect 51548 36652 52052 36708
rect 51996 36594 52052 36652
rect 51996 36542 51998 36594
rect 52050 36542 52052 36594
rect 51996 36530 52052 36542
rect 51548 36484 51604 36494
rect 51436 36482 51604 36484
rect 51436 36430 51550 36482
rect 51602 36430 51604 36482
rect 51436 36428 51604 36430
rect 51548 36148 51604 36428
rect 52108 36372 52164 36876
rect 51548 36082 51604 36092
rect 51660 36316 52164 36372
rect 52220 37996 52556 38052
rect 51100 35084 51604 35140
rect 50316 34804 50372 35084
rect 50316 34690 50372 34748
rect 50988 35028 51044 35038
rect 50316 34638 50318 34690
rect 50370 34638 50372 34690
rect 50316 34626 50372 34638
rect 50428 34692 50484 34702
rect 49308 34078 49310 34130
rect 49362 34078 49364 34130
rect 49308 34066 49364 34078
rect 49756 34300 50148 34356
rect 50428 34354 50484 34636
rect 50428 34302 50430 34354
rect 50482 34302 50484 34354
rect 49756 34132 49812 34300
rect 50428 34290 50484 34302
rect 50988 34354 51044 34972
rect 51100 34914 51156 34926
rect 51100 34862 51102 34914
rect 51154 34862 51156 34914
rect 51100 34692 51156 34862
rect 51100 34626 51156 34636
rect 50988 34302 50990 34354
rect 51042 34302 51044 34354
rect 50988 34290 51044 34302
rect 51548 34354 51604 35084
rect 51660 35026 51716 36316
rect 51660 34974 51662 35026
rect 51714 34974 51716 35026
rect 51660 34692 51716 34974
rect 52108 35028 52164 35038
rect 52108 34934 52164 34972
rect 51660 34626 51716 34636
rect 51548 34302 51550 34354
rect 51602 34302 51604 34354
rect 51548 34290 51604 34302
rect 49756 34038 49812 34076
rect 50092 34132 50148 34142
rect 50092 34038 50148 34076
rect 49268 33740 49948 33750
rect 49324 33684 49372 33740
rect 49428 33738 49476 33740
rect 49532 33738 49580 33740
rect 49448 33686 49476 33738
rect 49572 33686 49580 33738
rect 49428 33684 49476 33686
rect 49532 33684 49580 33686
rect 49636 33738 49684 33740
rect 49740 33738 49788 33740
rect 49636 33686 49644 33738
rect 49740 33686 49768 33738
rect 49636 33684 49684 33686
rect 49740 33684 49788 33686
rect 49844 33684 49892 33740
rect 49268 33674 49948 33684
rect 49420 33236 49476 33246
rect 49084 33234 49476 33236
rect 49084 33182 49422 33234
rect 49474 33182 49476 33234
rect 49084 33180 49476 33182
rect 48748 33170 48804 33180
rect 49420 33170 49476 33180
rect 48188 33012 48244 33022
rect 48076 32956 48188 33012
rect 48188 32946 48244 32956
rect 47852 32734 47854 32786
rect 47906 32734 47908 32786
rect 47852 32722 47908 32734
rect 48300 32786 48356 33068
rect 50428 33124 50484 33134
rect 50428 33030 50484 33068
rect 48300 32734 48302 32786
rect 48354 32734 48356 32786
rect 48300 32722 48356 32734
rect 49196 32674 49252 32686
rect 49196 32622 49198 32674
rect 49250 32622 49252 32674
rect 49196 32564 49252 32622
rect 49420 32564 49476 32574
rect 49196 32562 49476 32564
rect 49196 32510 49422 32562
rect 49474 32510 49476 32562
rect 49196 32508 49476 32510
rect 49420 32498 49476 32508
rect 50092 32564 50148 32574
rect 50092 32470 50148 32508
rect 50876 32564 50932 32574
rect 46732 32172 46900 32228
rect 49268 32172 49948 32182
rect 46732 29986 46788 32172
rect 49324 32116 49372 32172
rect 49428 32170 49476 32172
rect 49532 32170 49580 32172
rect 49448 32118 49476 32170
rect 49572 32118 49580 32170
rect 49428 32116 49476 32118
rect 49532 32116 49580 32118
rect 49636 32170 49684 32172
rect 49740 32170 49788 32172
rect 49636 32118 49644 32170
rect 49740 32118 49768 32170
rect 49636 32116 49684 32118
rect 49740 32116 49788 32118
rect 49844 32116 49892 32172
rect 49268 32106 49948 32116
rect 46844 32004 46900 32014
rect 46844 31106 46900 31948
rect 50876 31666 50932 32508
rect 51212 32340 51268 32350
rect 51212 31778 51268 32284
rect 52220 31948 52276 37996
rect 52556 37986 52612 37996
rect 52668 38948 52724 38958
rect 52668 38050 52724 38892
rect 52668 37998 52670 38050
rect 52722 37998 52724 38050
rect 52668 37986 52724 37998
rect 53004 36820 53060 36830
rect 52444 36596 52500 36606
rect 52444 35922 52500 36540
rect 52780 36596 52836 36606
rect 52780 36482 52836 36540
rect 52780 36430 52782 36482
rect 52834 36430 52836 36482
rect 52780 36372 52836 36430
rect 53004 36482 53060 36764
rect 53004 36430 53006 36482
rect 53058 36430 53060 36482
rect 53004 36418 53060 36430
rect 52780 36306 52836 36316
rect 53116 36260 53172 39676
rect 53228 39666 53284 39676
rect 53676 39730 53732 40348
rect 54012 40290 54068 40348
rect 54012 40238 54014 40290
rect 54066 40238 54068 40290
rect 54012 40226 54068 40238
rect 54572 40292 54628 40462
rect 54572 40226 54628 40236
rect 53676 39678 53678 39730
rect 53730 39678 53732 39730
rect 53676 39666 53732 39678
rect 53768 39228 54448 39238
rect 53824 39172 53872 39228
rect 53928 39226 53976 39228
rect 54032 39226 54080 39228
rect 53948 39174 53976 39226
rect 54072 39174 54080 39226
rect 53928 39172 53976 39174
rect 54032 39172 54080 39174
rect 54136 39226 54184 39228
rect 54240 39226 54288 39228
rect 54136 39174 54144 39226
rect 54240 39174 54268 39226
rect 54136 39172 54184 39174
rect 54240 39172 54288 39174
rect 54344 39172 54392 39228
rect 53768 39162 54448 39172
rect 53228 38946 53284 38958
rect 53228 38894 53230 38946
rect 53282 38894 53284 38946
rect 53228 38050 53284 38894
rect 53900 38948 53956 38958
rect 53900 38854 53956 38892
rect 53228 37998 53230 38050
rect 53282 37998 53284 38050
rect 53228 37986 53284 37998
rect 53564 38834 53620 38846
rect 53564 38782 53566 38834
rect 53618 38782 53620 38834
rect 53564 37492 53620 38782
rect 54684 38668 54740 40684
rect 54796 40516 54852 44268
rect 54796 40402 54852 40460
rect 54796 40350 54798 40402
rect 54850 40350 54852 40402
rect 54796 40338 54852 40350
rect 54908 41860 54964 41870
rect 54684 38612 54852 38668
rect 54572 37828 54628 37838
rect 53768 37660 54448 37670
rect 53824 37604 53872 37660
rect 53928 37658 53976 37660
rect 54032 37658 54080 37660
rect 53948 37606 53976 37658
rect 54072 37606 54080 37658
rect 53928 37604 53976 37606
rect 54032 37604 54080 37606
rect 54136 37658 54184 37660
rect 54240 37658 54288 37660
rect 54136 37606 54144 37658
rect 54240 37606 54268 37658
rect 54136 37604 54184 37606
rect 54240 37604 54288 37606
rect 54344 37604 54392 37660
rect 53768 37594 54448 37604
rect 53676 37492 53732 37502
rect 53564 37490 53732 37492
rect 53564 37438 53678 37490
rect 53730 37438 53732 37490
rect 53564 37436 53732 37438
rect 53676 37426 53732 37436
rect 53228 37380 53284 37390
rect 54236 37380 54292 37390
rect 53228 36482 53284 37324
rect 53900 37378 54292 37380
rect 53900 37326 54238 37378
rect 54290 37326 54292 37378
rect 53900 37324 54292 37326
rect 53900 37044 53956 37324
rect 54236 37314 54292 37324
rect 54572 37380 54628 37772
rect 54572 37286 54628 37324
rect 54012 37156 54068 37166
rect 54012 37062 54068 37100
rect 53228 36430 53230 36482
rect 53282 36430 53284 36482
rect 53228 36418 53284 36430
rect 53340 36706 53396 36718
rect 53340 36654 53342 36706
rect 53394 36654 53396 36706
rect 53116 36204 53284 36260
rect 52444 35870 52446 35922
rect 52498 35870 52500 35922
rect 52444 35858 52500 35870
rect 53116 35700 53172 35710
rect 52780 35698 53172 35700
rect 52780 35646 53118 35698
rect 53170 35646 53172 35698
rect 52780 35644 53172 35646
rect 52780 35138 52836 35644
rect 53116 35634 53172 35644
rect 53228 35476 53284 36204
rect 53340 35810 53396 36654
rect 53340 35758 53342 35810
rect 53394 35758 53396 35810
rect 53340 35746 53396 35758
rect 53452 36370 53508 36382
rect 53452 36318 53454 36370
rect 53506 36318 53508 36370
rect 53452 36148 53508 36318
rect 53900 36260 53956 36988
rect 53900 36194 53956 36204
rect 53452 35588 53508 36092
rect 53768 36092 54448 36102
rect 53824 36036 53872 36092
rect 53928 36090 53976 36092
rect 54032 36090 54080 36092
rect 53948 36038 53976 36090
rect 54072 36038 54080 36090
rect 53928 36036 53976 36038
rect 54032 36036 54080 36038
rect 54136 36090 54184 36092
rect 54240 36090 54288 36092
rect 54136 36038 54144 36090
rect 54240 36038 54268 36090
rect 54136 36036 54184 36038
rect 54240 36036 54288 36038
rect 54344 36036 54392 36092
rect 53768 36026 54448 36036
rect 53564 35924 53620 35934
rect 53564 35810 53620 35868
rect 53564 35758 53566 35810
rect 53618 35758 53620 35810
rect 53564 35746 53620 35758
rect 53788 35700 53844 35710
rect 53788 35606 53844 35644
rect 53452 35522 53508 35532
rect 53228 35420 53396 35476
rect 52780 35086 52782 35138
rect 52834 35086 52836 35138
rect 52780 35074 52836 35086
rect 52668 35028 52724 35038
rect 52556 34916 52612 34926
rect 52332 34914 52612 34916
rect 52332 34862 52558 34914
rect 52610 34862 52612 34914
rect 52332 34860 52612 34862
rect 52332 34132 52388 34860
rect 52556 34850 52612 34860
rect 52668 34916 52724 34972
rect 52668 34860 53172 34916
rect 52668 34242 52724 34860
rect 53116 34802 53172 34860
rect 53116 34750 53118 34802
rect 53170 34750 53172 34802
rect 53116 34738 53172 34750
rect 52892 34692 52948 34702
rect 53228 34692 53284 34702
rect 52892 34690 53060 34692
rect 52892 34638 52894 34690
rect 52946 34638 53060 34690
rect 52892 34636 53060 34638
rect 52892 34626 52948 34636
rect 52668 34190 52670 34242
rect 52722 34190 52724 34242
rect 52668 34178 52724 34190
rect 52332 34038 52388 34076
rect 52556 32786 52612 32798
rect 52556 32734 52558 32786
rect 52610 32734 52612 32786
rect 52556 32340 52612 32734
rect 53004 32788 53060 34636
rect 53228 33458 53284 34636
rect 53228 33406 53230 33458
rect 53282 33406 53284 33458
rect 53116 32788 53172 32798
rect 53004 32786 53172 32788
rect 53004 32734 53118 32786
rect 53170 32734 53172 32786
rect 53004 32732 53172 32734
rect 53116 32564 53172 32732
rect 53116 32498 53172 32508
rect 53228 32340 53284 33406
rect 53340 32452 53396 35420
rect 54124 35474 54180 35486
rect 54124 35422 54126 35474
rect 54178 35422 54180 35474
rect 54124 35028 54180 35422
rect 54124 34962 54180 34972
rect 54796 34804 54852 38612
rect 54796 34738 54852 34748
rect 54684 34692 54740 34702
rect 54684 34598 54740 34636
rect 53768 34524 54448 34534
rect 53824 34468 53872 34524
rect 53928 34522 53976 34524
rect 54032 34522 54080 34524
rect 53948 34470 53976 34522
rect 54072 34470 54080 34522
rect 53928 34468 53976 34470
rect 54032 34468 54080 34470
rect 54136 34522 54184 34524
rect 54240 34522 54288 34524
rect 54136 34470 54144 34522
rect 54240 34470 54268 34522
rect 54136 34468 54184 34470
rect 54240 34468 54288 34470
rect 54344 34468 54392 34524
rect 53768 34458 54448 34468
rect 53768 32956 54448 32966
rect 53824 32900 53872 32956
rect 53928 32954 53976 32956
rect 54032 32954 54080 32956
rect 53948 32902 53976 32954
rect 54072 32902 54080 32954
rect 53928 32900 53976 32902
rect 54032 32900 54080 32902
rect 54136 32954 54184 32956
rect 54240 32954 54288 32956
rect 54136 32902 54144 32954
rect 54240 32902 54268 32954
rect 54136 32900 54184 32902
rect 54240 32900 54288 32902
rect 54344 32900 54392 32956
rect 53768 32890 54448 32900
rect 54572 32788 54628 32798
rect 54572 32674 54628 32732
rect 54572 32622 54574 32674
rect 54626 32622 54628 32674
rect 54572 32610 54628 32622
rect 53788 32564 53844 32574
rect 53788 32470 53844 32508
rect 54460 32562 54516 32574
rect 54460 32510 54462 32562
rect 54514 32510 54516 32562
rect 53340 32386 53396 32396
rect 54460 32452 54516 32510
rect 54908 32452 54964 41804
rect 55020 41748 55076 45612
rect 55132 41972 55188 50372
rect 56364 48804 56420 48814
rect 56364 48710 56420 48748
rect 57372 48804 57428 48814
rect 55692 48356 55748 48366
rect 55356 48354 55748 48356
rect 55356 48302 55694 48354
rect 55746 48302 55748 48354
rect 55356 48300 55748 48302
rect 55356 47458 55412 48300
rect 55692 48290 55748 48300
rect 57372 48354 57428 48748
rect 57372 48302 57374 48354
rect 57426 48302 57428 48354
rect 56028 48244 56084 48254
rect 56700 48244 56756 48254
rect 56028 48242 56756 48244
rect 56028 48190 56030 48242
rect 56082 48190 56702 48242
rect 56754 48190 56756 48242
rect 56028 48188 56756 48190
rect 56028 48178 56084 48188
rect 56700 48178 56756 48188
rect 55356 47406 55358 47458
rect 55410 47406 55412 47458
rect 55356 47394 55412 47406
rect 57036 48018 57092 48030
rect 57036 47966 57038 48018
rect 57090 47966 57092 48018
rect 57036 47236 57092 47966
rect 57036 47170 57092 47180
rect 57260 46786 57316 46798
rect 57260 46734 57262 46786
rect 57314 46734 57316 46786
rect 55244 46676 55300 46686
rect 55244 46582 55300 46620
rect 56588 46674 56644 46686
rect 56588 46622 56590 46674
rect 56642 46622 56644 46674
rect 55356 46564 55412 46574
rect 55356 46450 55412 46508
rect 55356 46398 55358 46450
rect 55410 46398 55412 46450
rect 55132 41906 55188 41916
rect 55244 46228 55300 46238
rect 55020 41682 55076 41692
rect 55244 37492 55300 46172
rect 55356 45444 55412 46398
rect 55580 46562 55636 46574
rect 55580 46510 55582 46562
rect 55634 46510 55636 46562
rect 55580 46116 55636 46510
rect 55580 46050 55636 46060
rect 56028 46562 56084 46574
rect 56028 46510 56030 46562
rect 56082 46510 56084 46562
rect 55692 45778 55748 45790
rect 55692 45726 55694 45778
rect 55746 45726 55748 45778
rect 55692 45444 55748 45726
rect 56028 45668 56084 46510
rect 56588 46116 56644 46622
rect 57260 46564 57316 46734
rect 57260 46498 57316 46508
rect 56588 46050 56644 46060
rect 56812 45780 56868 45790
rect 56028 45602 56084 45612
rect 56700 45668 56756 45678
rect 56812 45668 56868 45724
rect 56756 45612 56868 45668
rect 56924 45668 56980 45678
rect 56700 45602 56756 45612
rect 56924 45574 56980 45612
rect 55356 45388 55748 45444
rect 55356 41076 55412 45388
rect 56924 45220 56980 45230
rect 56924 45218 57204 45220
rect 56924 45166 56926 45218
rect 56978 45166 57204 45218
rect 56924 45164 57204 45166
rect 56924 45154 56980 45164
rect 56588 45108 56644 45118
rect 56364 45106 56644 45108
rect 56364 45054 56590 45106
rect 56642 45054 56644 45106
rect 56364 45052 56644 45054
rect 55916 44994 55972 45006
rect 55916 44942 55918 44994
rect 55970 44942 55972 44994
rect 55468 44324 55524 44334
rect 55468 44230 55524 44268
rect 55692 44324 55748 44334
rect 55692 44212 55748 44268
rect 55580 44210 55748 44212
rect 55580 44158 55694 44210
rect 55746 44158 55748 44210
rect 55580 44156 55748 44158
rect 55580 43762 55636 44156
rect 55692 44146 55748 44156
rect 55916 44212 55972 44942
rect 56364 44546 56420 45052
rect 56588 45042 56644 45052
rect 56364 44494 56366 44546
rect 56418 44494 56420 44546
rect 56364 44482 56420 44494
rect 56700 44324 56756 44334
rect 56700 44322 56868 44324
rect 56700 44270 56702 44322
rect 56754 44270 56868 44322
rect 56700 44268 56868 44270
rect 56700 44258 56756 44268
rect 55916 44146 55972 44156
rect 55580 43710 55582 43762
rect 55634 43710 55636 43762
rect 55580 43698 55636 43710
rect 56700 44100 56756 44110
rect 56028 43652 56084 43662
rect 56028 43558 56084 43596
rect 56700 43538 56756 44044
rect 56812 43764 56868 44268
rect 56812 43698 56868 43708
rect 56924 44212 56980 44222
rect 56700 43486 56702 43538
rect 56754 43486 56756 43538
rect 56700 43474 56756 43486
rect 55580 41972 55636 41982
rect 55356 41010 55412 41020
rect 55468 41916 55580 41972
rect 55468 41636 55524 41916
rect 55580 41878 55636 41916
rect 56924 41972 56980 44156
rect 57148 43538 57204 45164
rect 57260 44212 57316 44222
rect 57372 44212 57428 48302
rect 57596 48356 57652 51772
rect 57708 51604 57764 51614
rect 57820 51604 57876 51996
rect 57932 51986 57988 51996
rect 58044 52164 58100 52174
rect 57708 51602 57876 51604
rect 57708 51550 57710 51602
rect 57762 51550 57876 51602
rect 57708 51548 57876 51550
rect 57708 51538 57764 51548
rect 58044 50708 58100 52108
rect 58156 52050 58212 52220
rect 58604 52276 58660 52286
rect 58604 52182 58660 52220
rect 59052 52276 59108 53454
rect 59500 53058 59556 54572
rect 60508 54626 60564 55020
rect 62768 54908 63448 54918
rect 62824 54852 62872 54908
rect 62928 54906 62976 54908
rect 63032 54906 63080 54908
rect 62948 54854 62976 54906
rect 63072 54854 63080 54906
rect 62928 54852 62976 54854
rect 63032 54852 63080 54854
rect 63136 54906 63184 54908
rect 63240 54906 63288 54908
rect 63136 54854 63144 54906
rect 63240 54854 63268 54906
rect 63136 54852 63184 54854
rect 63240 54852 63288 54854
rect 63344 54852 63392 54908
rect 62768 54842 63448 54852
rect 60508 54574 60510 54626
rect 60562 54574 60564 54626
rect 60508 54562 60564 54574
rect 61292 54514 61348 54526
rect 61292 54462 61294 54514
rect 61346 54462 61348 54514
rect 61292 54404 61348 54462
rect 61852 54404 61908 54414
rect 61292 54402 61908 54404
rect 61292 54350 61854 54402
rect 61906 54350 61908 54402
rect 61292 54348 61908 54350
rect 60172 53844 60228 53854
rect 60172 53170 60228 53788
rect 60172 53118 60174 53170
rect 60226 53118 60228 53170
rect 60172 53106 60228 53118
rect 59500 53006 59502 53058
rect 59554 53006 59556 53058
rect 59500 52994 59556 53006
rect 59052 52210 59108 52220
rect 60508 52276 60564 52286
rect 60508 52182 60564 52220
rect 61852 52164 61908 54348
rect 65772 54402 65828 54414
rect 65772 54350 65774 54402
rect 65826 54350 65828 54402
rect 65324 53844 65380 53854
rect 65324 53750 65380 53788
rect 61852 52098 61908 52108
rect 62076 53732 62132 53742
rect 62076 52836 62132 53676
rect 65212 53732 65268 53742
rect 65212 53638 65268 53676
rect 65436 53732 65492 53742
rect 65772 53732 65828 54350
rect 66780 54404 66836 54414
rect 66556 53956 66612 53966
rect 65996 53732 66052 53742
rect 65436 53730 66052 53732
rect 65436 53678 65438 53730
rect 65490 53678 65998 53730
rect 66050 53678 66052 53730
rect 65436 53676 66052 53678
rect 64876 53620 64932 53630
rect 64876 53526 64932 53564
rect 64540 53506 64596 53518
rect 64540 53454 64542 53506
rect 64594 53454 64596 53506
rect 62768 53340 63448 53350
rect 62824 53284 62872 53340
rect 62928 53338 62976 53340
rect 63032 53338 63080 53340
rect 62948 53286 62976 53338
rect 63072 53286 63080 53338
rect 62928 53284 62976 53286
rect 63032 53284 63080 53286
rect 63136 53338 63184 53340
rect 63240 53338 63288 53340
rect 63136 53286 63144 53338
rect 63240 53286 63268 53338
rect 63136 53284 63184 53286
rect 63240 53284 63288 53286
rect 63344 53284 63392 53340
rect 62768 53274 63448 53284
rect 64540 53060 64596 53454
rect 64540 52994 64596 53004
rect 65436 53060 65492 53676
rect 65996 53666 66052 53676
rect 66108 53732 66164 53742
rect 65660 53508 65716 53518
rect 65660 53506 66052 53508
rect 65660 53454 65662 53506
rect 65714 53454 66052 53506
rect 65660 53452 66052 53454
rect 65660 53442 65716 53452
rect 65436 52994 65492 53004
rect 65996 53058 66052 53452
rect 65996 53006 65998 53058
rect 66050 53006 66052 53058
rect 65996 52994 66052 53006
rect 65212 52948 65268 52958
rect 58156 51998 58158 52050
rect 58210 51998 58212 52050
rect 58156 51986 58212 51998
rect 62076 51602 62132 52780
rect 65100 52892 65212 52948
rect 62636 52724 62692 52734
rect 62636 52274 62692 52668
rect 62636 52222 62638 52274
rect 62690 52222 62692 52274
rect 62636 52210 62692 52222
rect 63420 52164 63476 52174
rect 63420 52070 63476 52108
rect 63868 52164 63924 52174
rect 63868 52070 63924 52108
rect 65100 52164 65156 52892
rect 65212 52854 65268 52892
rect 66108 52836 66164 53676
rect 66332 53730 66388 53742
rect 66332 53678 66334 53730
rect 66386 53678 66388 53730
rect 66332 53508 66388 53678
rect 66556 53730 66612 53900
rect 66556 53678 66558 53730
rect 66610 53678 66612 53730
rect 66556 53666 66612 53678
rect 66780 53730 66836 54348
rect 66780 53678 66782 53730
rect 66834 53678 66836 53730
rect 66780 53666 66836 53678
rect 66892 53732 66948 55246
rect 67116 55186 67172 56028
rect 68460 56084 68516 56094
rect 68460 55990 68516 56028
rect 69020 55970 69076 56252
rect 69020 55918 69022 55970
rect 69074 55918 69076 55970
rect 69020 55906 69076 55918
rect 81676 56082 81732 56094
rect 81676 56030 81678 56082
rect 81730 56030 81732 56082
rect 67268 55692 67948 55702
rect 67324 55636 67372 55692
rect 67428 55690 67476 55692
rect 67532 55690 67580 55692
rect 67448 55638 67476 55690
rect 67572 55638 67580 55690
rect 67428 55636 67476 55638
rect 67532 55636 67580 55638
rect 67636 55690 67684 55692
rect 67740 55690 67788 55692
rect 67636 55638 67644 55690
rect 67740 55638 67768 55690
rect 67636 55636 67684 55638
rect 67740 55636 67788 55638
rect 67844 55636 67892 55692
rect 67268 55626 67948 55636
rect 76268 55692 76948 55702
rect 76324 55636 76372 55692
rect 76428 55690 76476 55692
rect 76532 55690 76580 55692
rect 76448 55638 76476 55690
rect 76572 55638 76580 55690
rect 76428 55636 76476 55638
rect 76532 55636 76580 55638
rect 76636 55690 76684 55692
rect 76740 55690 76788 55692
rect 76636 55638 76644 55690
rect 76740 55638 76768 55690
rect 76636 55636 76684 55638
rect 76740 55636 76788 55638
rect 76844 55636 76892 55692
rect 76268 55626 76948 55636
rect 67116 55134 67118 55186
rect 67170 55134 67172 55186
rect 67116 55122 67172 55134
rect 68348 55186 68404 55198
rect 68348 55134 68350 55186
rect 68402 55134 68404 55186
rect 67268 54124 67948 54134
rect 67324 54068 67372 54124
rect 67428 54122 67476 54124
rect 67532 54122 67580 54124
rect 67448 54070 67476 54122
rect 67572 54070 67580 54122
rect 67428 54068 67476 54070
rect 67532 54068 67580 54070
rect 67636 54122 67684 54124
rect 67740 54122 67788 54124
rect 67636 54070 67644 54122
rect 67740 54070 67768 54122
rect 67636 54068 67684 54070
rect 67740 54068 67788 54070
rect 67844 54068 67892 54124
rect 67268 54058 67948 54068
rect 66892 53666 66948 53676
rect 67116 53956 67172 53966
rect 67116 53730 67172 53900
rect 68348 53956 68404 55134
rect 68684 55076 68740 55086
rect 68684 54982 68740 55020
rect 81676 55076 81732 56030
rect 81676 55010 81732 55020
rect 82124 56084 82180 56094
rect 71768 54908 72448 54918
rect 71824 54852 71872 54908
rect 71928 54906 71976 54908
rect 72032 54906 72080 54908
rect 71948 54854 71976 54906
rect 72072 54854 72080 54906
rect 71928 54852 71976 54854
rect 72032 54852 72080 54854
rect 72136 54906 72184 54908
rect 72240 54906 72288 54908
rect 72136 54854 72144 54906
rect 72240 54854 72268 54906
rect 72136 54852 72184 54854
rect 72240 54852 72288 54854
rect 72344 54852 72392 54908
rect 71768 54842 72448 54852
rect 80768 54908 81448 54918
rect 80824 54852 80872 54908
rect 80928 54906 80976 54908
rect 81032 54906 81080 54908
rect 80948 54854 80976 54906
rect 81072 54854 81080 54906
rect 80928 54852 80976 54854
rect 81032 54852 81080 54854
rect 81136 54906 81184 54908
rect 81240 54906 81288 54908
rect 81136 54854 81144 54906
rect 81240 54854 81268 54906
rect 81136 54852 81184 54854
rect 81240 54852 81288 54854
rect 81344 54852 81392 54908
rect 80768 54842 81448 54852
rect 82124 54738 82180 56028
rect 82236 55970 82292 56590
rect 92988 56642 93044 59200
rect 97692 58548 97748 58558
rect 95900 56756 95956 56766
rect 92988 56590 92990 56642
rect 93042 56590 93044 56642
rect 92988 56578 93044 56590
rect 93996 56642 94052 56654
rect 93996 56590 93998 56642
rect 94050 56590 94052 56642
rect 89768 56476 90448 56486
rect 89824 56420 89872 56476
rect 89928 56474 89976 56476
rect 90032 56474 90080 56476
rect 89948 56422 89976 56474
rect 90072 56422 90080 56474
rect 89928 56420 89976 56422
rect 90032 56420 90080 56422
rect 90136 56474 90184 56476
rect 90240 56474 90288 56476
rect 90136 56422 90144 56474
rect 90240 56422 90268 56474
rect 90136 56420 90184 56422
rect 90240 56420 90288 56422
rect 90344 56420 90392 56476
rect 89768 56410 90448 56420
rect 93996 56306 94052 56590
rect 93996 56254 93998 56306
rect 94050 56254 94052 56306
rect 93996 56242 94052 56254
rect 93212 56084 93268 56094
rect 93212 55990 93268 56028
rect 82236 55918 82238 55970
rect 82290 55918 82292 55970
rect 82236 55906 82292 55918
rect 95900 55970 95956 56700
rect 97692 56306 97748 58492
rect 97692 56254 97694 56306
rect 97746 56254 97748 56306
rect 97692 56242 97748 56254
rect 96348 56084 96404 56094
rect 96348 55990 96404 56028
rect 96908 56082 96964 56094
rect 96908 56030 96910 56082
rect 96962 56030 96964 56082
rect 95900 55918 95902 55970
rect 95954 55918 95956 55970
rect 95900 55906 95956 55918
rect 85268 55692 85948 55702
rect 85324 55636 85372 55692
rect 85428 55690 85476 55692
rect 85532 55690 85580 55692
rect 85448 55638 85476 55690
rect 85572 55638 85580 55690
rect 85428 55636 85476 55638
rect 85532 55636 85580 55638
rect 85636 55690 85684 55692
rect 85740 55690 85788 55692
rect 85636 55638 85644 55690
rect 85740 55638 85768 55690
rect 85636 55636 85684 55638
rect 85740 55636 85788 55638
rect 85844 55636 85892 55692
rect 85268 55626 85948 55636
rect 94268 55692 94948 55702
rect 94324 55636 94372 55692
rect 94428 55690 94476 55692
rect 94532 55690 94580 55692
rect 94448 55638 94476 55690
rect 94572 55638 94580 55690
rect 94428 55636 94476 55638
rect 94532 55636 94580 55638
rect 94636 55690 94684 55692
rect 94740 55690 94788 55692
rect 94636 55638 94644 55690
rect 94740 55638 94768 55690
rect 94636 55636 94684 55638
rect 94740 55636 94788 55638
rect 94844 55636 94892 55692
rect 94268 55626 94948 55636
rect 96908 55468 96964 56030
rect 96572 55412 96964 55468
rect 97244 56084 97300 56094
rect 96572 55076 96628 55412
rect 96460 55074 96628 55076
rect 96460 55022 96574 55074
rect 96626 55022 96628 55074
rect 96460 55020 96628 55022
rect 89768 54908 90448 54918
rect 89824 54852 89872 54908
rect 89928 54906 89976 54908
rect 90032 54906 90080 54908
rect 89948 54854 89976 54906
rect 90072 54854 90080 54906
rect 89928 54852 89976 54854
rect 90032 54852 90080 54854
rect 90136 54906 90184 54908
rect 90240 54906 90288 54908
rect 90136 54854 90144 54906
rect 90240 54854 90268 54906
rect 90136 54852 90184 54854
rect 90240 54852 90288 54854
rect 90344 54852 90392 54908
rect 89768 54842 90448 54852
rect 82124 54686 82126 54738
rect 82178 54686 82180 54738
rect 82124 54674 82180 54686
rect 81788 54514 81844 54526
rect 81788 54462 81790 54514
rect 81842 54462 81844 54514
rect 81452 54404 81508 54414
rect 81788 54404 81844 54462
rect 81452 54402 81844 54404
rect 81452 54350 81454 54402
rect 81506 54350 81844 54402
rect 81452 54348 81844 54350
rect 81452 54338 81508 54348
rect 76268 54124 76948 54134
rect 76324 54068 76372 54124
rect 76428 54122 76476 54124
rect 76532 54122 76580 54124
rect 76448 54070 76476 54122
rect 76572 54070 76580 54122
rect 76428 54068 76476 54070
rect 76532 54068 76580 54070
rect 76636 54122 76684 54124
rect 76740 54122 76788 54124
rect 76636 54070 76644 54122
rect 76740 54070 76768 54122
rect 76636 54068 76684 54070
rect 76740 54068 76788 54070
rect 76844 54068 76892 54124
rect 76268 54058 76948 54068
rect 68348 53890 68404 53900
rect 72828 53842 72884 53854
rect 72828 53790 72830 53842
rect 72882 53790 72884 53842
rect 67116 53678 67118 53730
rect 67170 53678 67172 53730
rect 67116 53666 67172 53678
rect 69916 53730 69972 53742
rect 69916 53678 69918 53730
rect 69970 53678 69972 53730
rect 66668 53620 66724 53630
rect 66668 53526 66724 53564
rect 67228 53618 67284 53630
rect 67228 53566 67230 53618
rect 67282 53566 67284 53618
rect 66332 53442 66388 53452
rect 67228 53508 67284 53566
rect 67676 53508 67732 53518
rect 67228 53452 67676 53508
rect 67228 53172 67284 53452
rect 67676 53414 67732 53452
rect 69580 53508 69636 53518
rect 69916 53508 69972 53678
rect 70700 53620 70756 53630
rect 70700 53526 70756 53564
rect 69580 53506 69972 53508
rect 69580 53454 69582 53506
rect 69634 53454 69972 53506
rect 69580 53452 69972 53454
rect 72828 53508 72884 53790
rect 67228 53106 67284 53116
rect 68796 52948 68852 52958
rect 68796 52854 68852 52892
rect 69580 52948 69636 53452
rect 72828 53442 72884 53452
rect 75740 53508 75796 53518
rect 71768 53340 72448 53350
rect 71824 53284 71872 53340
rect 71928 53338 71976 53340
rect 72032 53338 72080 53340
rect 71948 53286 71976 53338
rect 72072 53286 72080 53338
rect 71928 53284 71976 53286
rect 72032 53284 72080 53286
rect 72136 53338 72184 53340
rect 72240 53338 72288 53340
rect 72136 53286 72144 53338
rect 72240 53286 72268 53338
rect 72136 53284 72184 53286
rect 72240 53284 72288 53286
rect 72344 53284 72392 53340
rect 71768 53274 72448 53284
rect 69580 52882 69636 52892
rect 65996 52780 66164 52836
rect 68124 52834 68180 52846
rect 68124 52782 68126 52834
rect 68178 52782 68180 52834
rect 65996 52386 66052 52780
rect 65996 52334 65998 52386
rect 66050 52334 66052 52386
rect 65996 52322 66052 52334
rect 66556 52724 66612 52734
rect 66108 52276 66164 52286
rect 66556 52276 66612 52668
rect 68124 52724 68180 52782
rect 68124 52658 68180 52668
rect 71260 52724 71316 52734
rect 67268 52556 67948 52566
rect 67324 52500 67372 52556
rect 67428 52554 67476 52556
rect 67532 52554 67580 52556
rect 67448 52502 67476 52554
rect 67572 52502 67580 52554
rect 67428 52500 67476 52502
rect 67532 52500 67580 52502
rect 67636 52554 67684 52556
rect 67740 52554 67788 52556
rect 67636 52502 67644 52554
rect 67740 52502 67768 52554
rect 67636 52500 67684 52502
rect 67740 52500 67788 52502
rect 67844 52500 67892 52556
rect 67268 52490 67948 52500
rect 66108 52274 66612 52276
rect 66108 52222 66110 52274
rect 66162 52222 66558 52274
rect 66610 52222 66612 52274
rect 66108 52220 66612 52222
rect 66108 52210 66164 52220
rect 66556 52210 66612 52220
rect 62768 51772 63448 51782
rect 62824 51716 62872 51772
rect 62928 51770 62976 51772
rect 63032 51770 63080 51772
rect 62948 51718 62976 51770
rect 63072 51718 63080 51770
rect 62928 51716 62976 51718
rect 63032 51716 63080 51718
rect 63136 51770 63184 51772
rect 63240 51770 63288 51772
rect 63136 51718 63144 51770
rect 63240 51718 63268 51770
rect 63136 51716 63184 51718
rect 63240 51716 63288 51718
rect 63344 51716 63392 51772
rect 62768 51706 63448 51716
rect 62076 51550 62078 51602
rect 62130 51550 62132 51602
rect 62076 51538 62132 51550
rect 62188 51378 62244 51390
rect 62188 51326 62190 51378
rect 62242 51326 62244 51378
rect 61740 51268 61796 51278
rect 61740 51174 61796 51212
rect 62188 51268 62244 51326
rect 62188 51202 62244 51212
rect 58268 50988 58948 50998
rect 58324 50932 58372 50988
rect 58428 50986 58476 50988
rect 58532 50986 58580 50988
rect 58448 50934 58476 50986
rect 58572 50934 58580 50986
rect 58428 50932 58476 50934
rect 58532 50932 58580 50934
rect 58636 50986 58684 50988
rect 58740 50986 58788 50988
rect 58636 50934 58644 50986
rect 58740 50934 58768 50986
rect 58636 50932 58684 50934
rect 58740 50932 58788 50934
rect 58844 50932 58892 50988
rect 58268 50922 58948 50932
rect 58604 50708 58660 50718
rect 58044 50706 58660 50708
rect 58044 50654 58606 50706
rect 58658 50654 58660 50706
rect 58044 50652 58660 50654
rect 58044 50594 58100 50652
rect 58604 50642 58660 50652
rect 60396 50596 60452 50606
rect 58044 50542 58046 50594
rect 58098 50542 58100 50594
rect 58044 50530 58100 50542
rect 59948 50594 60452 50596
rect 59948 50542 60398 50594
rect 60450 50542 60452 50594
rect 59948 50540 60452 50542
rect 59948 50370 60004 50540
rect 60396 50530 60452 50540
rect 60956 50594 61012 50606
rect 60956 50542 60958 50594
rect 61010 50542 61012 50594
rect 59948 50318 59950 50370
rect 60002 50318 60004 50370
rect 59948 50306 60004 50318
rect 60956 50034 61012 50542
rect 63308 50484 63364 50494
rect 63364 50428 63588 50484
rect 63308 50390 63364 50428
rect 62768 50204 63448 50214
rect 62824 50148 62872 50204
rect 62928 50202 62976 50204
rect 63032 50202 63080 50204
rect 62948 50150 62976 50202
rect 63072 50150 63080 50202
rect 62928 50148 62976 50150
rect 63032 50148 63080 50150
rect 63136 50202 63184 50204
rect 63240 50202 63288 50204
rect 63136 50150 63144 50202
rect 63240 50150 63268 50202
rect 63136 50148 63184 50150
rect 63240 50148 63288 50150
rect 63344 50148 63392 50204
rect 62768 50138 63448 50148
rect 60956 49982 60958 50034
rect 61010 49982 61012 50034
rect 60956 49970 61012 49982
rect 62300 49922 62356 49934
rect 62300 49870 62302 49922
rect 62354 49870 62356 49922
rect 61292 49812 61348 49822
rect 61740 49812 61796 49822
rect 61292 49810 61796 49812
rect 61292 49758 61294 49810
rect 61346 49758 61742 49810
rect 61794 49758 61796 49810
rect 61292 49756 61796 49758
rect 61292 49746 61348 49756
rect 61740 49746 61796 49756
rect 60620 49700 60676 49710
rect 60620 49606 60676 49644
rect 61964 49700 62020 49710
rect 61292 49588 61348 49598
rect 58268 49420 58948 49430
rect 58324 49364 58372 49420
rect 58428 49418 58476 49420
rect 58532 49418 58580 49420
rect 58448 49366 58476 49418
rect 58572 49366 58580 49418
rect 58428 49364 58476 49366
rect 58532 49364 58580 49366
rect 58636 49418 58684 49420
rect 58740 49418 58788 49420
rect 58636 49366 58644 49418
rect 58740 49366 58768 49418
rect 58636 49364 58684 49366
rect 58740 49364 58788 49366
rect 58844 49364 58892 49420
rect 58268 49354 58948 49364
rect 61292 49138 61348 49532
rect 61292 49086 61294 49138
rect 61346 49086 61348 49138
rect 61292 49074 61348 49086
rect 57820 48356 57876 48366
rect 57596 48354 57876 48356
rect 57596 48302 57822 48354
rect 57874 48302 57876 48354
rect 57596 48300 57876 48302
rect 57820 48132 57876 48300
rect 58380 48132 58436 48142
rect 57820 48130 58436 48132
rect 57820 48078 58382 48130
rect 58434 48078 58436 48130
rect 57820 48076 58436 48078
rect 57596 47348 57652 47358
rect 57596 47254 57652 47292
rect 57820 46900 57876 48076
rect 58380 48066 58436 48076
rect 58268 47852 58948 47862
rect 58324 47796 58372 47852
rect 58428 47850 58476 47852
rect 58532 47850 58580 47852
rect 58448 47798 58476 47850
rect 58572 47798 58580 47850
rect 58428 47796 58476 47798
rect 58532 47796 58580 47798
rect 58636 47850 58684 47852
rect 58740 47850 58788 47852
rect 58636 47798 58644 47850
rect 58740 47798 58768 47850
rect 58636 47796 58684 47798
rect 58740 47796 58788 47798
rect 58844 47796 58892 47852
rect 58268 47786 58948 47796
rect 58380 47236 58436 47246
rect 60732 47236 60788 47246
rect 58436 47180 58548 47236
rect 58380 47142 58436 47180
rect 57820 46834 57876 46844
rect 58380 46788 58436 46798
rect 58156 46786 58436 46788
rect 58156 46734 58382 46786
rect 58434 46734 58436 46786
rect 58156 46732 58436 46734
rect 57708 45890 57764 45902
rect 57708 45838 57710 45890
rect 57762 45838 57764 45890
rect 57316 44156 57428 44212
rect 57484 44324 57540 44334
rect 57484 44210 57540 44268
rect 57484 44158 57486 44210
rect 57538 44158 57540 44210
rect 57260 44146 57316 44156
rect 57484 44146 57540 44158
rect 57708 43764 57764 45838
rect 58044 45780 58100 45790
rect 58156 45780 58212 46732
rect 58380 46722 58436 46732
rect 58492 46674 58548 47180
rect 60620 47234 60788 47236
rect 60620 47182 60734 47234
rect 60786 47182 60788 47234
rect 60620 47180 60788 47182
rect 58492 46622 58494 46674
rect 58546 46622 58548 46674
rect 58492 46610 58548 46622
rect 60060 46674 60116 46686
rect 60060 46622 60062 46674
rect 60114 46622 60116 46674
rect 58268 46564 58324 46574
rect 58268 46470 58324 46508
rect 60060 46452 60116 46622
rect 60060 46386 60116 46396
rect 60172 46676 60228 46686
rect 60396 46676 60452 46686
rect 60228 46674 60452 46676
rect 60228 46622 60398 46674
rect 60450 46622 60452 46674
rect 60228 46620 60452 46622
rect 58268 46284 58948 46294
rect 58324 46228 58372 46284
rect 58428 46282 58476 46284
rect 58532 46282 58580 46284
rect 58448 46230 58476 46282
rect 58572 46230 58580 46282
rect 58428 46228 58476 46230
rect 58532 46228 58580 46230
rect 58636 46282 58684 46284
rect 58740 46282 58788 46284
rect 58636 46230 58644 46282
rect 58740 46230 58768 46282
rect 58636 46228 58684 46230
rect 58740 46228 58788 46230
rect 58844 46228 58892 46284
rect 58268 46218 58948 46228
rect 60172 46004 60228 46620
rect 60396 46610 60452 46620
rect 59948 45948 60228 46004
rect 58100 45724 58212 45780
rect 58492 45890 58548 45902
rect 58492 45838 58494 45890
rect 58546 45838 58548 45890
rect 58044 45714 58100 45724
rect 58492 44884 58548 45838
rect 59948 45890 60004 45948
rect 59948 45838 59950 45890
rect 60002 45838 60004 45890
rect 59948 45826 60004 45838
rect 60620 45890 60676 47180
rect 60732 47170 60788 47180
rect 61852 46788 61908 46798
rect 61404 46786 61908 46788
rect 61404 46734 61854 46786
rect 61906 46734 61908 46786
rect 61404 46732 61908 46734
rect 61404 46340 61460 46732
rect 61852 46722 61908 46732
rect 60620 45838 60622 45890
rect 60674 45838 60676 45890
rect 60620 45826 60676 45838
rect 61068 46284 61460 46340
rect 61068 45890 61124 46284
rect 61068 45838 61070 45890
rect 61122 45838 61124 45890
rect 61068 45826 61124 45838
rect 61292 45220 61348 45230
rect 61292 45126 61348 45164
rect 61740 44996 61796 45006
rect 61740 44902 61796 44940
rect 58492 44818 58548 44828
rect 58268 44716 58948 44726
rect 58324 44660 58372 44716
rect 58428 44714 58476 44716
rect 58532 44714 58580 44716
rect 58448 44662 58476 44714
rect 58572 44662 58580 44714
rect 58428 44660 58476 44662
rect 58532 44660 58580 44662
rect 58636 44714 58684 44716
rect 58740 44714 58788 44716
rect 58636 44662 58644 44714
rect 58740 44662 58768 44714
rect 58636 44660 58684 44662
rect 58740 44660 58788 44662
rect 58844 44660 58892 44716
rect 58268 44650 58948 44660
rect 58492 44324 58548 44334
rect 58492 44230 58548 44268
rect 57932 44100 57988 44110
rect 57932 44006 57988 44044
rect 57708 43698 57764 43708
rect 60172 43764 60228 43774
rect 60172 43670 60228 43708
rect 57820 43652 57876 43662
rect 59388 43652 59444 43662
rect 57876 43596 57988 43652
rect 57820 43586 57876 43596
rect 57148 43486 57150 43538
rect 57202 43486 57204 43538
rect 57148 43474 57204 43486
rect 57596 42082 57652 42094
rect 57596 42030 57598 42082
rect 57650 42030 57652 42082
rect 56924 41906 56980 41916
rect 57484 41970 57540 41982
rect 57484 41918 57486 41970
rect 57538 41918 57540 41970
rect 56028 41860 56084 41870
rect 56028 41766 56084 41804
rect 57484 41860 57540 41918
rect 57484 41794 57540 41804
rect 55356 40628 55412 40638
rect 55468 40628 55524 41580
rect 56140 41748 56196 41758
rect 55356 40626 55524 40628
rect 55356 40574 55358 40626
rect 55410 40574 55524 40626
rect 55356 40572 55524 40574
rect 55692 41186 55748 41198
rect 55692 41134 55694 41186
rect 55746 41134 55748 41186
rect 55356 40292 55412 40572
rect 55692 40404 55748 41134
rect 56140 41186 56196 41692
rect 56700 41748 56756 41758
rect 56700 41746 56980 41748
rect 56700 41694 56702 41746
rect 56754 41694 56980 41746
rect 56700 41692 56980 41694
rect 56700 41682 56756 41692
rect 56140 41134 56142 41186
rect 56194 41134 56196 41186
rect 56140 41122 56196 41134
rect 56924 40516 56980 41692
rect 57036 41746 57092 41758
rect 57036 41694 57038 41746
rect 57090 41694 57092 41746
rect 57036 41188 57092 41694
rect 57596 41636 57652 42030
rect 57596 41300 57652 41580
rect 57596 41234 57652 41244
rect 57036 41094 57092 41132
rect 57820 41076 57876 41086
rect 57820 40982 57876 41020
rect 57820 40628 57876 40638
rect 57932 40628 57988 43596
rect 59388 43558 59444 43596
rect 60956 43652 61012 43662
rect 58268 43148 58948 43158
rect 58324 43092 58372 43148
rect 58428 43146 58476 43148
rect 58532 43146 58580 43148
rect 58448 43094 58476 43146
rect 58572 43094 58580 43146
rect 58428 43092 58476 43094
rect 58532 43092 58580 43094
rect 58636 43146 58684 43148
rect 58740 43146 58788 43148
rect 58636 43094 58644 43146
rect 58740 43094 58768 43146
rect 58636 43092 58684 43094
rect 58740 43092 58788 43094
rect 58844 43092 58892 43148
rect 58268 43082 58948 43092
rect 60956 42868 61012 43596
rect 58380 42084 58436 42094
rect 57820 40626 57988 40628
rect 57820 40574 57822 40626
rect 57874 40574 57988 40626
rect 57820 40572 57988 40574
rect 58156 42082 58436 42084
rect 58156 42030 58382 42082
rect 58434 42030 58436 42082
rect 58156 42028 58436 42030
rect 57036 40516 57092 40526
rect 56924 40514 57092 40516
rect 56924 40462 57038 40514
rect 57090 40462 57092 40514
rect 56924 40460 57092 40462
rect 57036 40450 57092 40460
rect 57372 40514 57428 40526
rect 57372 40462 57374 40514
rect 57426 40462 57428 40514
rect 57372 40404 57428 40462
rect 57708 40404 57764 40414
rect 57372 40348 57708 40404
rect 55692 40338 55748 40348
rect 57708 40338 57764 40348
rect 55356 40226 55412 40236
rect 55804 38612 55860 38622
rect 55804 37826 55860 38556
rect 56700 38612 56756 38622
rect 56700 38162 56756 38556
rect 57820 38612 57876 40572
rect 58156 40402 58212 42028
rect 58380 42018 58436 42028
rect 58268 41580 58948 41590
rect 58324 41524 58372 41580
rect 58428 41578 58476 41580
rect 58532 41578 58580 41580
rect 58448 41526 58476 41578
rect 58572 41526 58580 41578
rect 58428 41524 58476 41526
rect 58532 41524 58580 41526
rect 58636 41578 58684 41580
rect 58740 41578 58788 41580
rect 58636 41526 58644 41578
rect 58740 41526 58768 41578
rect 58636 41524 58684 41526
rect 58740 41524 58788 41526
rect 58844 41524 58892 41580
rect 58268 41514 58948 41524
rect 58716 41412 58772 41422
rect 58716 41188 58772 41356
rect 59276 41412 59332 41422
rect 58940 41188 58996 41198
rect 58716 41186 58996 41188
rect 58716 41134 58942 41186
rect 58994 41134 58996 41186
rect 58716 41132 58996 41134
rect 58940 41122 58996 41132
rect 59276 40962 59332 41356
rect 59276 40910 59278 40962
rect 59330 40910 59332 40962
rect 59276 40898 59332 40910
rect 60508 41076 60564 41086
rect 58156 40350 58158 40402
rect 58210 40350 58212 40402
rect 58156 40338 58212 40350
rect 58604 40404 58660 40414
rect 58604 40310 58660 40348
rect 58268 40012 58948 40022
rect 58324 39956 58372 40012
rect 58428 40010 58476 40012
rect 58532 40010 58580 40012
rect 58448 39958 58476 40010
rect 58572 39958 58580 40010
rect 58428 39956 58476 39958
rect 58532 39956 58580 39958
rect 58636 40010 58684 40012
rect 58740 40010 58788 40012
rect 58636 39958 58644 40010
rect 58740 39958 58768 40010
rect 58636 39956 58684 39958
rect 58740 39956 58788 39958
rect 58844 39956 58892 40012
rect 58268 39946 58948 39956
rect 58044 38948 58100 38958
rect 57876 38556 57988 38612
rect 57820 38546 57876 38556
rect 56700 38110 56702 38162
rect 56754 38110 56756 38162
rect 56700 38098 56756 38110
rect 55804 37774 55806 37826
rect 55858 37774 55860 37826
rect 55804 37762 55860 37774
rect 56364 37828 56420 37838
rect 56364 37734 56420 37772
rect 57932 37604 57988 38556
rect 55356 37492 55412 37502
rect 55244 37490 55412 37492
rect 55244 37438 55358 37490
rect 55410 37438 55412 37490
rect 55244 37436 55412 37438
rect 55244 37156 55300 37436
rect 55244 37090 55300 37100
rect 55244 34916 55300 34926
rect 55020 34914 55300 34916
rect 55020 34862 55246 34914
rect 55298 34862 55300 34914
rect 55020 34860 55300 34862
rect 55020 34802 55076 34860
rect 55244 34850 55300 34860
rect 55020 34750 55022 34802
rect 55074 34750 55076 34802
rect 55020 34738 55076 34750
rect 55356 34692 55412 37436
rect 57932 37490 57988 37548
rect 57932 37438 57934 37490
rect 57986 37438 57988 37490
rect 57932 37426 57988 37438
rect 57484 37156 57540 37166
rect 56812 36932 56868 36942
rect 56812 36596 56868 36876
rect 56812 36594 57428 36596
rect 56812 36542 56814 36594
rect 56866 36542 57428 36594
rect 56812 36540 57428 36542
rect 56812 36530 56868 36540
rect 56028 36372 56084 36382
rect 56028 35700 56084 36316
rect 57372 36372 57428 36540
rect 57148 35924 57204 35962
rect 57148 35858 57204 35868
rect 57372 35922 57428 36316
rect 57372 35870 57374 35922
rect 57426 35870 57428 35922
rect 57372 35858 57428 35870
rect 56028 35606 56084 35644
rect 57148 35700 57204 35710
rect 57148 35606 57204 35644
rect 56700 35588 56756 35598
rect 56700 35494 56756 35532
rect 55804 34916 55860 34926
rect 55244 34636 55412 34692
rect 55692 34914 55860 34916
rect 55692 34862 55806 34914
rect 55858 34862 55860 34914
rect 55692 34860 55860 34862
rect 55244 32788 55300 34636
rect 55692 34354 55748 34860
rect 55804 34850 55860 34860
rect 55692 34302 55694 34354
rect 55746 34302 55748 34354
rect 55692 34290 55748 34302
rect 55356 34244 55412 34254
rect 55356 34150 55412 34188
rect 57372 34244 57428 34254
rect 57484 34244 57540 37100
rect 57596 35700 57652 35710
rect 57820 35700 57876 35710
rect 58044 35700 58100 38892
rect 58380 38946 58436 38958
rect 58380 38894 58382 38946
rect 58434 38894 58436 38946
rect 58380 38668 58436 38894
rect 60172 38836 60228 38846
rect 60172 38742 60228 38780
rect 58156 38612 58436 38668
rect 58156 37266 58212 38612
rect 58268 38444 58948 38454
rect 58324 38388 58372 38444
rect 58428 38442 58476 38444
rect 58532 38442 58580 38444
rect 58448 38390 58476 38442
rect 58572 38390 58580 38442
rect 58428 38388 58476 38390
rect 58532 38388 58580 38390
rect 58636 38442 58684 38444
rect 58740 38442 58788 38444
rect 58636 38390 58644 38442
rect 58740 38390 58768 38442
rect 58636 38388 58684 38390
rect 58740 38388 58788 38390
rect 58844 38388 58892 38444
rect 58268 38378 58948 38388
rect 59276 37940 59332 37950
rect 59276 37846 59332 37884
rect 58940 37828 58996 37838
rect 58156 37214 58158 37266
rect 58210 37214 58212 37266
rect 58156 37202 58212 37214
rect 58716 37826 58996 37828
rect 58716 37774 58942 37826
rect 58994 37774 58996 37826
rect 58716 37772 58996 37774
rect 58716 37266 58772 37772
rect 58940 37762 58996 37772
rect 59948 37828 60004 37838
rect 58716 37214 58718 37266
rect 58770 37214 58772 37266
rect 58716 37202 58772 37214
rect 59948 37044 60004 37772
rect 60508 37828 60564 41020
rect 60956 40626 61012 42812
rect 61852 42868 61908 42878
rect 61852 42774 61908 42812
rect 60956 40574 60958 40626
rect 61010 40574 61012 40626
rect 60956 40562 61012 40574
rect 61740 41188 61796 41198
rect 61740 40626 61796 41132
rect 61964 41076 62020 49644
rect 62300 49700 62356 49870
rect 62300 49634 62356 49644
rect 62860 49922 62916 49934
rect 62860 49870 62862 49922
rect 62914 49870 62916 49922
rect 62076 49588 62132 49598
rect 62076 45220 62132 49532
rect 62860 49588 62916 49870
rect 62860 49522 62916 49532
rect 62768 48636 63448 48646
rect 62824 48580 62872 48636
rect 62928 48634 62976 48636
rect 63032 48634 63080 48636
rect 62948 48582 62976 48634
rect 63072 48582 63080 48634
rect 62928 48580 62976 48582
rect 63032 48580 63080 48582
rect 63136 48634 63184 48636
rect 63240 48634 63288 48636
rect 63136 48582 63144 48634
rect 63240 48582 63268 48634
rect 63136 48580 63184 48582
rect 63240 48580 63288 48582
rect 63344 48580 63392 48636
rect 62768 48570 63448 48580
rect 62768 47068 63448 47078
rect 62824 47012 62872 47068
rect 62928 47066 62976 47068
rect 63032 47066 63080 47068
rect 62948 47014 62976 47066
rect 63072 47014 63080 47066
rect 62928 47012 62976 47014
rect 63032 47012 63080 47014
rect 63136 47066 63184 47068
rect 63240 47066 63288 47068
rect 63136 47014 63144 47066
rect 63240 47014 63268 47066
rect 63136 47012 63184 47014
rect 63240 47012 63288 47014
rect 63344 47012 63392 47068
rect 62768 47002 63448 47012
rect 62188 46676 62244 46686
rect 62188 46674 62468 46676
rect 62188 46622 62190 46674
rect 62242 46622 62468 46674
rect 62188 46620 62468 46622
rect 62188 46610 62244 46620
rect 62412 45330 62468 46620
rect 62412 45278 62414 45330
rect 62466 45278 62468 45330
rect 62412 45266 62468 45278
rect 62636 45668 62692 45678
rect 62076 45154 62132 45164
rect 62636 45108 62692 45612
rect 63532 45666 63588 50428
rect 64092 50482 64148 50494
rect 64092 50430 64094 50482
rect 64146 50430 64148 50482
rect 64092 49588 64148 50430
rect 64540 50484 64596 50494
rect 64540 50390 64596 50428
rect 64988 49922 65044 49934
rect 64988 49870 64990 49922
rect 65042 49870 65044 49922
rect 64092 49522 64148 49532
rect 64764 49810 64820 49822
rect 64764 49758 64766 49810
rect 64818 49758 64820 49810
rect 63644 49476 63700 49486
rect 63644 49138 63700 49420
rect 64764 49250 64820 49758
rect 64988 49812 65044 49870
rect 64988 49746 65044 49756
rect 64764 49198 64766 49250
rect 64818 49198 64820 49250
rect 64764 49186 64820 49198
rect 64876 49588 64932 49598
rect 63644 49086 63646 49138
rect 63698 49086 63700 49138
rect 63644 49028 63700 49086
rect 63644 48962 63700 48972
rect 64204 48916 64260 48926
rect 64204 48822 64260 48860
rect 63868 48468 63924 48478
rect 63868 47236 63924 48412
rect 64540 48356 64596 48366
rect 64540 47572 64596 48300
rect 64876 48354 64932 49532
rect 65100 49252 65156 52108
rect 70588 51490 70644 51502
rect 71036 51492 71092 51502
rect 70588 51438 70590 51490
rect 70642 51438 70644 51490
rect 67268 50988 67948 50998
rect 67324 50932 67372 50988
rect 67428 50986 67476 50988
rect 67532 50986 67580 50988
rect 67448 50934 67476 50986
rect 67572 50934 67580 50986
rect 67428 50932 67476 50934
rect 67532 50932 67580 50934
rect 67636 50986 67684 50988
rect 67740 50986 67788 50988
rect 67636 50934 67644 50986
rect 67740 50934 67768 50986
rect 67636 50932 67684 50934
rect 67740 50932 67788 50934
rect 67844 50932 67892 50988
rect 67268 50922 67948 50932
rect 70476 50596 70532 50606
rect 70588 50596 70644 51438
rect 70476 50594 70644 50596
rect 70476 50542 70478 50594
rect 70530 50542 70644 50594
rect 70476 50540 70644 50542
rect 70924 51490 71092 51492
rect 70924 51438 71038 51490
rect 71090 51438 71092 51490
rect 70924 51436 71092 51438
rect 70924 50594 70980 51436
rect 71036 51426 71092 51436
rect 70924 50542 70926 50594
rect 70978 50542 70980 50594
rect 70476 50530 70532 50540
rect 70924 50530 70980 50542
rect 65548 50372 65604 50382
rect 65436 50370 65604 50372
rect 65436 50318 65550 50370
rect 65602 50318 65604 50370
rect 65436 50316 65604 50318
rect 65436 49810 65492 50316
rect 65548 50306 65604 50316
rect 68124 50372 68180 50382
rect 68124 50034 68180 50316
rect 68124 49982 68126 50034
rect 68178 49982 68180 50034
rect 68124 49970 68180 49982
rect 69244 50372 69300 50382
rect 69244 50034 69300 50316
rect 69244 49982 69246 50034
rect 69298 49982 69300 50034
rect 69244 49970 69300 49982
rect 65436 49758 65438 49810
rect 65490 49758 65492 49810
rect 65436 49746 65492 49758
rect 65772 49812 65828 49822
rect 65772 49718 65828 49756
rect 71260 49698 71316 52668
rect 71768 51772 72448 51782
rect 71824 51716 71872 51772
rect 71928 51770 71976 51772
rect 72032 51770 72080 51772
rect 71948 51718 71976 51770
rect 72072 51718 72080 51770
rect 71928 51716 71976 51718
rect 72032 51716 72080 51718
rect 72136 51770 72184 51772
rect 72240 51770 72288 51772
rect 72136 51718 72144 51770
rect 72240 51718 72268 51770
rect 72136 51716 72184 51718
rect 72240 51716 72288 51718
rect 72344 51716 72392 51772
rect 71768 51706 72448 51716
rect 71372 51492 71428 51502
rect 71372 51398 71428 51436
rect 72492 51492 72548 51502
rect 72548 51436 72660 51492
rect 72492 51426 72548 51436
rect 71768 50204 72448 50214
rect 71824 50148 71872 50204
rect 71928 50202 71976 50204
rect 72032 50202 72080 50204
rect 71948 50150 71976 50202
rect 72072 50150 72080 50202
rect 71928 50148 71976 50150
rect 72032 50148 72080 50150
rect 72136 50202 72184 50204
rect 72240 50202 72288 50204
rect 72136 50150 72144 50202
rect 72240 50150 72268 50202
rect 72136 50148 72184 50150
rect 72240 50148 72288 50150
rect 72344 50148 72392 50204
rect 71768 50138 72448 50148
rect 72380 50036 72436 50046
rect 72604 50036 72660 51436
rect 74284 51268 74340 51278
rect 74284 50706 74340 51212
rect 74284 50654 74286 50706
rect 74338 50654 74340 50706
rect 73164 50484 73220 50494
rect 73164 50390 73220 50428
rect 73948 50482 74004 50494
rect 73948 50430 73950 50482
rect 74002 50430 74004 50482
rect 72380 50034 72660 50036
rect 72380 49982 72382 50034
rect 72434 49982 72660 50034
rect 72380 49980 72660 49982
rect 72380 49970 72436 49980
rect 72940 49922 72996 49934
rect 72940 49870 72942 49922
rect 72994 49870 72996 49922
rect 71260 49646 71262 49698
rect 71314 49646 71316 49698
rect 64876 48302 64878 48354
rect 64930 48302 64932 48354
rect 64876 48290 64932 48302
rect 64988 49196 65156 49252
rect 65884 49588 65940 49598
rect 64988 48020 65044 49196
rect 65100 49028 65156 49038
rect 65100 48934 65156 48972
rect 65324 48916 65380 48926
rect 65884 48916 65940 49532
rect 68908 49588 68964 49598
rect 68908 49494 68964 49532
rect 67268 49420 67948 49430
rect 67324 49364 67372 49420
rect 67428 49418 67476 49420
rect 67532 49418 67580 49420
rect 67448 49366 67476 49418
rect 67572 49366 67580 49418
rect 67428 49364 67476 49366
rect 67532 49364 67580 49366
rect 67636 49418 67684 49420
rect 67740 49418 67788 49420
rect 67636 49366 67644 49418
rect 67740 49366 67768 49418
rect 67636 49364 67684 49366
rect 67740 49364 67788 49366
rect 67844 49364 67892 49420
rect 67268 49354 67948 49364
rect 65324 48822 65380 48860
rect 65436 48914 65940 48916
rect 65436 48862 65886 48914
rect 65938 48862 65940 48914
rect 65436 48860 65940 48862
rect 65324 48468 65380 48478
rect 65436 48468 65492 48860
rect 65884 48850 65940 48860
rect 71260 49028 71316 49646
rect 71708 49700 71764 49710
rect 71708 49606 71764 49644
rect 72940 49700 72996 49870
rect 73500 49924 73556 49934
rect 73500 49922 73892 49924
rect 73500 49870 73502 49922
rect 73554 49870 73892 49922
rect 73500 49868 73892 49870
rect 73500 49858 73556 49868
rect 72940 49634 72996 49644
rect 72716 49586 72772 49598
rect 72716 49534 72718 49586
rect 72770 49534 72772 49586
rect 65324 48466 65492 48468
rect 65324 48414 65326 48466
rect 65378 48414 65492 48466
rect 65324 48412 65492 48414
rect 65548 48468 65604 48478
rect 65324 48402 65380 48412
rect 65100 48356 65156 48366
rect 65100 48262 65156 48300
rect 65548 48242 65604 48412
rect 65548 48190 65550 48242
rect 65602 48190 65604 48242
rect 65548 48178 65604 48190
rect 71036 48354 71092 48366
rect 71036 48302 71038 48354
rect 71090 48302 71092 48354
rect 64540 47506 64596 47516
rect 64764 47964 65044 48020
rect 65212 48130 65268 48142
rect 65212 48078 65214 48130
rect 65266 48078 65268 48130
rect 63868 47170 63924 47180
rect 64652 45892 64708 45902
rect 64540 45836 64652 45892
rect 64540 45778 64596 45836
rect 64652 45826 64708 45836
rect 64540 45726 64542 45778
rect 64594 45726 64596 45778
rect 64540 45714 64596 45726
rect 63532 45614 63534 45666
rect 63586 45614 63588 45666
rect 62768 45500 63448 45510
rect 62824 45444 62872 45500
rect 62928 45498 62976 45500
rect 63032 45498 63080 45500
rect 62948 45446 62976 45498
rect 63072 45446 63080 45498
rect 62928 45444 62976 45446
rect 63032 45444 63080 45446
rect 63136 45498 63184 45500
rect 63240 45498 63288 45500
rect 63136 45446 63144 45498
rect 63240 45446 63268 45498
rect 63136 45444 63184 45446
rect 63240 45444 63288 45446
rect 63344 45444 63392 45500
rect 62768 45434 63448 45444
rect 63532 45444 63588 45614
rect 64092 45668 64148 45678
rect 64092 45574 64148 45612
rect 64652 45668 64708 45678
rect 64652 45574 64708 45612
rect 63532 45378 63588 45388
rect 64540 45444 64596 45454
rect 64540 45330 64596 45388
rect 64540 45278 64542 45330
rect 64594 45278 64596 45330
rect 64540 45266 64596 45278
rect 63308 45220 63364 45230
rect 63084 45164 63308 45220
rect 62748 45108 62804 45118
rect 62636 45106 62804 45108
rect 62636 45054 62750 45106
rect 62802 45054 62804 45106
rect 62636 45052 62804 45054
rect 62748 45042 62804 45052
rect 61964 41010 62020 41020
rect 62076 44996 62132 45006
rect 61740 40574 61742 40626
rect 61794 40574 61796 40626
rect 61740 40562 61796 40574
rect 62076 40964 62132 44940
rect 63084 44548 63140 45164
rect 63308 45126 63364 45164
rect 63532 45106 63588 45118
rect 63532 45054 63534 45106
rect 63586 45054 63588 45106
rect 63532 44996 63588 45054
rect 63532 44930 63588 44940
rect 63084 44434 63140 44492
rect 64428 44548 64484 44558
rect 64428 44454 64484 44492
rect 63084 44382 63086 44434
rect 63138 44382 63140 44434
rect 63084 44370 63140 44382
rect 64652 44210 64708 44222
rect 64652 44158 64654 44210
rect 64706 44158 64708 44210
rect 63532 44100 63588 44110
rect 63532 44006 63588 44044
rect 64092 44098 64148 44110
rect 64092 44046 64094 44098
rect 64146 44046 64148 44098
rect 62768 43932 63448 43942
rect 62824 43876 62872 43932
rect 62928 43930 62976 43932
rect 63032 43930 63080 43932
rect 62948 43878 62976 43930
rect 63072 43878 63080 43930
rect 62928 43876 62976 43878
rect 63032 43876 63080 43878
rect 63136 43930 63184 43932
rect 63240 43930 63288 43932
rect 63136 43878 63144 43930
rect 63240 43878 63268 43930
rect 63136 43876 63184 43878
rect 63240 43876 63288 43878
rect 63344 43876 63392 43932
rect 62768 43866 63448 43876
rect 63420 43764 63476 43774
rect 62412 43650 62468 43662
rect 63084 43652 63140 43662
rect 62412 43598 62414 43650
rect 62466 43598 62468 43650
rect 62300 42756 62356 42766
rect 62412 42756 62468 43598
rect 62300 42754 62468 42756
rect 62300 42702 62302 42754
rect 62354 42702 62468 42754
rect 62300 42700 62468 42702
rect 62748 43650 63140 43652
rect 62748 43598 63086 43650
rect 63138 43598 63140 43650
rect 62748 43596 63140 43598
rect 62748 42754 62804 43596
rect 63084 43586 63140 43596
rect 63420 43650 63476 43708
rect 64092 43764 64148 44046
rect 64092 43698 64148 43708
rect 64652 44100 64708 44158
rect 63420 43598 63422 43650
rect 63474 43598 63476 43650
rect 63420 43586 63476 43598
rect 64540 43428 64596 43438
rect 64540 43334 64596 43372
rect 62748 42702 62750 42754
rect 62802 42702 62804 42754
rect 62300 42690 62356 42700
rect 62748 42690 62804 42702
rect 62768 42364 63448 42374
rect 62824 42308 62872 42364
rect 62928 42362 62976 42364
rect 63032 42362 63080 42364
rect 62948 42310 62976 42362
rect 63072 42310 63080 42362
rect 62928 42308 62976 42310
rect 63032 42308 63080 42310
rect 63136 42362 63184 42364
rect 63240 42362 63288 42364
rect 63136 42310 63144 42362
rect 63240 42310 63268 42362
rect 63136 42308 63184 42310
rect 63240 42308 63288 42310
rect 63344 42308 63392 42364
rect 64652 42308 64708 44044
rect 62768 42298 63448 42308
rect 64428 42252 64708 42308
rect 63980 41188 64036 41198
rect 63756 41186 64036 41188
rect 63756 41134 63982 41186
rect 64034 41134 64036 41186
rect 63756 41132 64036 41134
rect 63756 41074 63812 41132
rect 63980 41122 64036 41132
rect 63756 41022 63758 41074
rect 63810 41022 63812 41074
rect 63756 41010 63812 41022
rect 60956 39060 61012 39070
rect 60956 38836 61012 39004
rect 60956 38274 61012 38780
rect 60956 38222 60958 38274
rect 61010 38222 61012 38274
rect 60956 38210 61012 38222
rect 60620 37940 60676 37950
rect 60620 37846 60676 37884
rect 61180 37938 61236 37950
rect 61180 37886 61182 37938
rect 61234 37886 61236 37938
rect 60508 37762 60564 37772
rect 61180 37828 61236 37886
rect 61180 37762 61236 37772
rect 61740 37940 61796 37950
rect 60956 37604 61012 37614
rect 60956 37490 61012 37548
rect 60956 37438 60958 37490
rect 61010 37438 61012 37490
rect 60956 37426 61012 37438
rect 61740 37490 61796 37884
rect 61740 37438 61742 37490
rect 61794 37438 61796 37490
rect 61740 37426 61796 37438
rect 59948 36978 60004 36988
rect 58268 36876 58948 36886
rect 58324 36820 58372 36876
rect 58428 36874 58476 36876
rect 58532 36874 58580 36876
rect 58448 36822 58476 36874
rect 58572 36822 58580 36874
rect 58428 36820 58476 36822
rect 58532 36820 58580 36822
rect 58636 36874 58684 36876
rect 58740 36874 58788 36876
rect 58636 36822 58644 36874
rect 58740 36822 58768 36874
rect 58636 36820 58684 36822
rect 58740 36820 58788 36822
rect 58844 36820 58892 36876
rect 58268 36810 58948 36820
rect 57596 35698 57764 35700
rect 57596 35646 57598 35698
rect 57650 35646 57764 35698
rect 57596 35644 57764 35646
rect 57596 35634 57652 35644
rect 57428 34188 57540 34244
rect 57708 34916 57764 35644
rect 57820 35698 58100 35700
rect 57820 35646 57822 35698
rect 57874 35646 58100 35698
rect 57820 35644 58100 35646
rect 57820 35588 57876 35644
rect 57820 35522 57876 35532
rect 58268 35308 58948 35318
rect 58324 35252 58372 35308
rect 58428 35306 58476 35308
rect 58532 35306 58580 35308
rect 58448 35254 58476 35306
rect 58572 35254 58580 35306
rect 58428 35252 58476 35254
rect 58532 35252 58580 35254
rect 58636 35306 58684 35308
rect 58740 35306 58788 35308
rect 58636 35254 58644 35306
rect 58740 35254 58768 35306
rect 58636 35252 58684 35254
rect 58740 35252 58788 35254
rect 58844 35252 58892 35308
rect 58268 35242 58948 35252
rect 57708 34242 57764 34860
rect 58940 34916 58996 34926
rect 58940 34822 58996 34860
rect 61628 34916 61684 34926
rect 61964 34916 62020 34926
rect 61628 34914 62020 34916
rect 61628 34862 61630 34914
rect 61682 34862 61966 34914
rect 62018 34862 62020 34914
rect 61628 34860 62020 34862
rect 61628 34850 61684 34860
rect 61516 34804 61572 34814
rect 58156 34690 58212 34702
rect 58156 34638 58158 34690
rect 58210 34638 58212 34690
rect 58156 34468 58212 34638
rect 58156 34402 58212 34412
rect 60732 34580 60788 34590
rect 57708 34190 57710 34242
rect 57762 34190 57764 34242
rect 57372 34150 57428 34188
rect 57708 34178 57764 34190
rect 56028 34132 56084 34142
rect 56812 34132 56868 34142
rect 56028 34130 56868 34132
rect 56028 34078 56030 34130
rect 56082 34078 56814 34130
rect 56866 34078 56868 34130
rect 56028 34076 56868 34078
rect 56028 34066 56084 34076
rect 56812 34066 56868 34076
rect 57148 33906 57204 33918
rect 57148 33854 57150 33906
rect 57202 33854 57204 33906
rect 56364 33122 56420 33134
rect 56364 33070 56366 33122
rect 56418 33070 56420 33122
rect 55244 32694 55300 32732
rect 55692 32788 55748 32798
rect 55692 32694 55748 32732
rect 56364 32788 56420 33070
rect 56364 32722 56420 32732
rect 57148 32788 57204 33854
rect 58268 33740 58948 33750
rect 58324 33684 58372 33740
rect 58428 33738 58476 33740
rect 58532 33738 58580 33740
rect 58448 33686 58476 33738
rect 58572 33686 58580 33738
rect 58428 33684 58476 33686
rect 58532 33684 58580 33686
rect 58636 33738 58684 33740
rect 58740 33738 58788 33740
rect 58636 33686 58644 33738
rect 58740 33686 58768 33738
rect 58636 33684 58684 33686
rect 58740 33684 58788 33686
rect 58844 33684 58892 33740
rect 58268 33674 58948 33684
rect 59836 33236 59892 33246
rect 57148 32722 57204 32732
rect 57820 32788 57876 32798
rect 56028 32676 56084 32686
rect 56028 32582 56084 32620
rect 57260 32676 57316 32686
rect 57260 32582 57316 32620
rect 57820 32674 57876 32732
rect 57820 32622 57822 32674
rect 57874 32622 57876 32674
rect 57820 32610 57876 32622
rect 59836 32786 59892 33180
rect 59836 32734 59838 32786
rect 59890 32734 59892 32786
rect 59836 32676 59892 32734
rect 59836 32610 59892 32620
rect 60284 33124 60340 33134
rect 57036 32564 57092 32574
rect 57036 32470 57092 32508
rect 59164 32564 59220 32574
rect 54460 32396 54964 32452
rect 52556 32284 53284 32340
rect 53116 32116 53172 32126
rect 52220 31892 52836 31948
rect 51212 31726 51214 31778
rect 51266 31726 51268 31778
rect 51212 31714 51268 31726
rect 50876 31614 50878 31666
rect 50930 31614 50932 31666
rect 50876 31602 50932 31614
rect 46844 31054 46846 31106
rect 46898 31054 46900 31106
rect 46844 31042 46900 31054
rect 47180 30996 47236 31006
rect 46956 30884 47012 30894
rect 46956 30790 47012 30828
rect 46732 29934 46734 29986
rect 46786 29934 46788 29986
rect 46732 29922 46788 29934
rect 46844 30212 46900 30222
rect 47068 30212 47124 30222
rect 46844 28642 46900 30156
rect 46956 30156 47068 30212
rect 46956 29428 47012 30156
rect 47068 30118 47124 30156
rect 47180 30100 47236 30940
rect 49268 30604 49948 30614
rect 49324 30548 49372 30604
rect 49428 30602 49476 30604
rect 49532 30602 49580 30604
rect 49448 30550 49476 30602
rect 49572 30550 49580 30602
rect 49428 30548 49476 30550
rect 49532 30548 49580 30550
rect 49636 30602 49684 30604
rect 49740 30602 49788 30604
rect 49636 30550 49644 30602
rect 49740 30550 49768 30602
rect 49636 30548 49684 30550
rect 49740 30548 49788 30550
rect 49844 30548 49892 30604
rect 49268 30538 49948 30548
rect 49756 30212 49812 30222
rect 47628 30100 47684 30110
rect 47180 30098 47684 30100
rect 47180 30046 47630 30098
rect 47682 30046 47684 30098
rect 47180 30044 47684 30046
rect 47628 30034 47684 30044
rect 49196 30100 49252 30110
rect 49196 30006 49252 30044
rect 49308 29986 49364 29998
rect 49308 29934 49310 29986
rect 49362 29934 49364 29986
rect 49308 29764 49364 29934
rect 49308 29698 49364 29708
rect 46956 29334 47012 29372
rect 49756 29204 49812 30156
rect 52668 30210 52724 30222
rect 52668 30158 52670 30210
rect 52722 30158 52724 30210
rect 50204 29986 50260 29998
rect 50204 29934 50206 29986
rect 50258 29934 50260 29986
rect 50204 29426 50260 29934
rect 52108 29988 52164 29998
rect 52668 29988 52724 30158
rect 52108 29986 52724 29988
rect 52108 29934 52110 29986
rect 52162 29934 52724 29986
rect 52108 29932 52724 29934
rect 50204 29374 50206 29426
rect 50258 29374 50260 29426
rect 50204 29362 50260 29374
rect 50540 29764 50596 29774
rect 50540 29426 50596 29708
rect 50540 29374 50542 29426
rect 50594 29374 50596 29426
rect 50540 29362 50596 29374
rect 49756 29138 49812 29148
rect 49268 29036 49948 29046
rect 49324 28980 49372 29036
rect 49428 29034 49476 29036
rect 49532 29034 49580 29036
rect 49448 28982 49476 29034
rect 49572 28982 49580 29034
rect 49428 28980 49476 28982
rect 49532 28980 49580 28982
rect 49636 29034 49684 29036
rect 49740 29034 49788 29036
rect 49636 28982 49644 29034
rect 49740 28982 49768 29034
rect 49636 28980 49684 28982
rect 49740 28980 49788 28982
rect 49844 28980 49892 29036
rect 49268 28970 49948 28980
rect 46844 28590 46846 28642
rect 46898 28590 46900 28642
rect 46844 28578 46900 28590
rect 47404 28644 47460 28654
rect 47740 28644 47796 28654
rect 47404 28642 47796 28644
rect 47404 28590 47406 28642
rect 47458 28590 47742 28642
rect 47794 28590 47796 28642
rect 47404 28588 47796 28590
rect 47404 28578 47460 28588
rect 47740 28578 47796 28588
rect 48076 28418 48132 28430
rect 48076 28366 48078 28418
rect 48130 28366 48132 28418
rect 48076 27860 48132 28366
rect 48524 28420 48580 28430
rect 48524 28418 48692 28420
rect 48524 28366 48526 28418
rect 48578 28366 48692 28418
rect 48524 28364 48692 28366
rect 48524 28354 48580 28364
rect 48076 27794 48132 27804
rect 48636 27858 48692 28364
rect 51772 28082 51828 28094
rect 51772 28030 51774 28082
rect 51826 28030 51828 28082
rect 51772 27972 51828 28030
rect 51772 27906 51828 27916
rect 48636 27806 48638 27858
rect 48690 27806 48692 27858
rect 48636 27794 48692 27806
rect 49196 27860 49252 27870
rect 49196 27766 49252 27804
rect 46844 27748 46900 27758
rect 46844 27654 46900 27692
rect 49268 27468 49948 27478
rect 49324 27412 49372 27468
rect 49428 27466 49476 27468
rect 49532 27466 49580 27468
rect 49448 27414 49476 27466
rect 49572 27414 49580 27466
rect 49428 27412 49476 27414
rect 49532 27412 49580 27414
rect 49636 27466 49684 27468
rect 49740 27466 49788 27468
rect 49636 27414 49644 27466
rect 49740 27414 49768 27466
rect 49636 27412 49684 27414
rect 49740 27412 49788 27414
rect 49844 27412 49892 27468
rect 49268 27402 49948 27412
rect 49644 26402 49700 26414
rect 49644 26350 49646 26402
rect 49698 26350 49700 26402
rect 48412 26292 48468 26302
rect 49644 26292 49700 26350
rect 49868 26292 49924 26302
rect 49644 26290 49924 26292
rect 49644 26238 49870 26290
rect 49922 26238 49924 26290
rect 49644 26236 49924 26238
rect 48412 25730 48468 26236
rect 49868 26226 49924 26236
rect 50428 26292 50484 26302
rect 50428 26198 50484 26236
rect 49268 25900 49948 25910
rect 49324 25844 49372 25900
rect 49428 25898 49476 25900
rect 49532 25898 49580 25900
rect 49448 25846 49476 25898
rect 49572 25846 49580 25898
rect 49428 25844 49476 25846
rect 49532 25844 49580 25846
rect 49636 25898 49684 25900
rect 49740 25898 49788 25900
rect 49636 25846 49644 25898
rect 49740 25846 49768 25898
rect 49636 25844 49684 25846
rect 49740 25844 49788 25846
rect 49844 25844 49892 25900
rect 49268 25834 49948 25844
rect 48412 25678 48414 25730
rect 48466 25678 48468 25730
rect 48412 25666 48468 25678
rect 47628 25284 47684 25294
rect 47628 25190 47684 25228
rect 49268 24332 49948 24342
rect 49324 24276 49372 24332
rect 49428 24330 49476 24332
rect 49532 24330 49580 24332
rect 49448 24278 49476 24330
rect 49572 24278 49580 24330
rect 49428 24276 49476 24278
rect 49532 24276 49580 24278
rect 49636 24330 49684 24332
rect 49740 24330 49788 24332
rect 49636 24278 49644 24330
rect 49740 24278 49768 24330
rect 49636 24276 49684 24278
rect 49740 24276 49788 24278
rect 49844 24276 49892 24332
rect 49268 24266 49948 24276
rect 49268 22764 49948 22774
rect 49324 22708 49372 22764
rect 49428 22762 49476 22764
rect 49532 22762 49580 22764
rect 49448 22710 49476 22762
rect 49572 22710 49580 22762
rect 49428 22708 49476 22710
rect 49532 22708 49580 22710
rect 49636 22762 49684 22764
rect 49740 22762 49788 22764
rect 49636 22710 49644 22762
rect 49740 22710 49768 22762
rect 49636 22708 49684 22710
rect 49740 22708 49788 22710
rect 49844 22708 49892 22764
rect 49268 22698 49948 22708
rect 46956 21476 47012 21486
rect 46956 20692 47012 21420
rect 49268 21196 49948 21206
rect 49324 21140 49372 21196
rect 49428 21194 49476 21196
rect 49532 21194 49580 21196
rect 49448 21142 49476 21194
rect 49572 21142 49580 21194
rect 49428 21140 49476 21142
rect 49532 21140 49580 21142
rect 49636 21194 49684 21196
rect 49740 21194 49788 21196
rect 49636 21142 49644 21194
rect 49740 21142 49768 21194
rect 49636 21140 49684 21142
rect 49740 21140 49788 21142
rect 49844 21140 49892 21196
rect 49268 21130 49948 21140
rect 46956 20626 47012 20636
rect 49268 19628 49948 19638
rect 49324 19572 49372 19628
rect 49428 19626 49476 19628
rect 49532 19626 49580 19628
rect 49448 19574 49476 19626
rect 49572 19574 49580 19626
rect 49428 19572 49476 19574
rect 49532 19572 49580 19574
rect 49636 19626 49684 19628
rect 49740 19626 49788 19628
rect 49636 19574 49644 19626
rect 49740 19574 49768 19626
rect 49636 19572 49684 19574
rect 49740 19572 49788 19574
rect 49844 19572 49892 19628
rect 49268 19562 49948 19572
rect 49268 18060 49948 18070
rect 49324 18004 49372 18060
rect 49428 18058 49476 18060
rect 49532 18058 49580 18060
rect 49448 18006 49476 18058
rect 49572 18006 49580 18058
rect 49428 18004 49476 18006
rect 49532 18004 49580 18006
rect 49636 18058 49684 18060
rect 49740 18058 49788 18060
rect 49636 18006 49644 18058
rect 49740 18006 49768 18058
rect 49636 18004 49684 18006
rect 49740 18004 49788 18006
rect 49844 18004 49892 18060
rect 49268 17994 49948 18004
rect 49268 16492 49948 16502
rect 49324 16436 49372 16492
rect 49428 16490 49476 16492
rect 49532 16490 49580 16492
rect 49448 16438 49476 16490
rect 49572 16438 49580 16490
rect 49428 16436 49476 16438
rect 49532 16436 49580 16438
rect 49636 16490 49684 16492
rect 49740 16490 49788 16492
rect 49636 16438 49644 16490
rect 49740 16438 49768 16490
rect 49636 16436 49684 16438
rect 49740 16436 49788 16438
rect 49844 16436 49892 16492
rect 49268 16426 49948 16436
rect 49268 14924 49948 14934
rect 49324 14868 49372 14924
rect 49428 14922 49476 14924
rect 49532 14922 49580 14924
rect 49448 14870 49476 14922
rect 49572 14870 49580 14922
rect 49428 14868 49476 14870
rect 49532 14868 49580 14870
rect 49636 14922 49684 14924
rect 49740 14922 49788 14924
rect 49636 14870 49644 14922
rect 49740 14870 49768 14922
rect 49636 14868 49684 14870
rect 49740 14868 49788 14870
rect 49844 14868 49892 14924
rect 49268 14858 49948 14868
rect 46620 14590 46622 14642
rect 46674 14590 46676 14642
rect 46620 14578 46676 14590
rect 44940 14532 44996 14542
rect 44604 14530 44996 14532
rect 44604 14478 44942 14530
rect 44994 14478 44996 14530
rect 44604 14476 44996 14478
rect 44604 11508 44660 14476
rect 44940 14466 44996 14476
rect 45388 14532 45444 14542
rect 45948 14532 46004 14542
rect 45388 14530 45668 14532
rect 45388 14478 45390 14530
rect 45442 14478 45668 14530
rect 45388 14476 45668 14478
rect 45388 14466 45444 14476
rect 44768 14140 45448 14150
rect 44824 14084 44872 14140
rect 44928 14138 44976 14140
rect 45032 14138 45080 14140
rect 44948 14086 44976 14138
rect 45072 14086 45080 14138
rect 44928 14084 44976 14086
rect 45032 14084 45080 14086
rect 45136 14138 45184 14140
rect 45240 14138 45288 14140
rect 45136 14086 45144 14138
rect 45240 14086 45268 14138
rect 45136 14084 45184 14086
rect 45240 14084 45288 14086
rect 45344 14084 45392 14140
rect 44768 14074 45448 14084
rect 45388 13748 45444 13758
rect 45388 13074 45444 13692
rect 45388 13022 45390 13074
rect 45442 13022 45444 13074
rect 45388 13010 45444 13022
rect 44768 12572 45448 12582
rect 44824 12516 44872 12572
rect 44928 12570 44976 12572
rect 45032 12570 45080 12572
rect 44948 12518 44976 12570
rect 45072 12518 45080 12570
rect 44928 12516 44976 12518
rect 45032 12516 45080 12518
rect 45136 12570 45184 12572
rect 45240 12570 45288 12572
rect 45136 12518 45144 12570
rect 45240 12518 45268 12570
rect 45136 12516 45184 12518
rect 45240 12516 45288 12518
rect 45344 12516 45392 12572
rect 44768 12506 45448 12516
rect 45612 11732 45668 14476
rect 44604 11442 44660 11452
rect 45500 11676 45668 11732
rect 45500 11172 45556 11676
rect 45612 11508 45668 11518
rect 45668 11452 45780 11508
rect 45612 11442 45668 11452
rect 45500 11116 45668 11172
rect 44768 11004 45448 11014
rect 44824 10948 44872 11004
rect 44928 11002 44976 11004
rect 45032 11002 45080 11004
rect 44948 10950 44976 11002
rect 45072 10950 45080 11002
rect 44928 10948 44976 10950
rect 45032 10948 45080 10950
rect 45136 11002 45184 11004
rect 45240 11002 45288 11004
rect 45136 10950 45144 11002
rect 45240 10950 45268 11002
rect 45136 10948 45184 10950
rect 45240 10948 45288 10950
rect 45344 10948 45392 11004
rect 44768 10938 45448 10948
rect 45052 9940 45108 9950
rect 45052 9846 45108 9884
rect 45164 9604 45220 9642
rect 45164 9538 45220 9548
rect 44768 9436 45448 9446
rect 44824 9380 44872 9436
rect 44928 9434 44976 9436
rect 45032 9434 45080 9436
rect 44948 9382 44976 9434
rect 45072 9382 45080 9434
rect 44928 9380 44976 9382
rect 45032 9380 45080 9382
rect 45136 9434 45184 9436
rect 45240 9434 45288 9436
rect 45136 9382 45144 9434
rect 45240 9382 45268 9434
rect 45136 9380 45184 9382
rect 45240 9380 45288 9382
rect 45344 9380 45392 9436
rect 44768 9370 45448 9380
rect 45388 9268 45444 9278
rect 45388 8258 45444 9212
rect 45388 8206 45390 8258
rect 45442 8206 45444 8258
rect 45388 8194 45444 8206
rect 44828 8148 44884 8158
rect 44828 8054 44884 8092
rect 44768 7868 45448 7878
rect 44824 7812 44872 7868
rect 44928 7866 44976 7868
rect 45032 7866 45080 7868
rect 44948 7814 44976 7866
rect 45072 7814 45080 7866
rect 44928 7812 44976 7814
rect 45032 7812 45080 7814
rect 45136 7866 45184 7868
rect 45240 7866 45288 7868
rect 45136 7814 45144 7866
rect 45240 7814 45268 7866
rect 45136 7812 45184 7814
rect 45240 7812 45288 7814
rect 45344 7812 45392 7868
rect 44768 7802 45448 7812
rect 45388 7362 45444 7374
rect 45388 7310 45390 7362
rect 45442 7310 45444 7362
rect 44492 6748 44660 6804
rect 44268 6692 44324 6702
rect 44268 6690 44548 6692
rect 44268 6638 44270 6690
rect 44322 6638 44548 6690
rect 44268 6636 44548 6638
rect 44268 6626 44324 6636
rect 44156 4398 44158 4450
rect 44210 4398 44212 4450
rect 44156 4386 44212 4398
rect 44380 5236 44436 5246
rect 44044 3726 44046 3778
rect 44098 3726 44100 3778
rect 44044 3714 44100 3726
rect 44268 3668 44324 3678
rect 44380 3668 44436 5180
rect 44492 4564 44548 6636
rect 44604 4788 44660 6748
rect 45388 6692 45444 7310
rect 45388 6626 45444 6636
rect 45612 6690 45668 11116
rect 45724 8370 45780 11452
rect 45948 9602 46004 14476
rect 46732 14532 46788 14542
rect 46732 14438 46788 14476
rect 47068 14530 47124 14542
rect 47068 14478 47070 14530
rect 47122 14478 47124 14530
rect 47068 14420 47124 14478
rect 47068 14354 47124 14364
rect 52108 14308 52164 29932
rect 52108 14242 52164 14252
rect 52444 27858 52500 27870
rect 52444 27806 52446 27858
rect 52498 27806 52500 27858
rect 52444 27748 52500 27806
rect 48972 13972 49028 13982
rect 46172 13748 46228 13758
rect 46060 13636 46116 13646
rect 46060 9938 46116 13580
rect 46060 9886 46062 9938
rect 46114 9886 46116 9938
rect 46060 9874 46116 9886
rect 46172 9940 46228 13692
rect 46956 12964 47012 12974
rect 47180 12964 47236 12974
rect 46956 12962 47180 12964
rect 46956 12910 46958 12962
rect 47010 12910 47180 12962
rect 46956 12908 47180 12910
rect 46956 12898 47012 12908
rect 47180 12850 47236 12908
rect 48076 12962 48132 12974
rect 48076 12910 48078 12962
rect 48130 12910 48132 12962
rect 47180 12798 47182 12850
rect 47234 12798 47236 12850
rect 47180 12786 47236 12798
rect 47740 12852 47796 12862
rect 46844 12292 46900 12302
rect 46508 12180 46564 12190
rect 45948 9550 45950 9602
rect 46002 9550 46004 9602
rect 45948 9538 46004 9550
rect 45724 8318 45726 8370
rect 45778 8318 45780 8370
rect 45724 8306 45780 8318
rect 45836 8932 45892 8942
rect 45836 8258 45892 8876
rect 45836 8206 45838 8258
rect 45890 8206 45892 8258
rect 45836 8194 45892 8206
rect 45948 8930 46004 8942
rect 45948 8878 45950 8930
rect 46002 8878 46004 8930
rect 45948 6916 46004 8878
rect 46172 8372 46228 9884
rect 45612 6638 45614 6690
rect 45666 6638 45668 6690
rect 45612 6626 45668 6638
rect 45724 6860 46004 6916
rect 46060 8316 46228 8372
rect 46396 11394 46452 11406
rect 46396 11342 46398 11394
rect 46450 11342 46452 11394
rect 45388 6468 45444 6506
rect 45388 6402 45444 6412
rect 44768 6300 45448 6310
rect 44824 6244 44872 6300
rect 44928 6298 44976 6300
rect 45032 6298 45080 6300
rect 44948 6246 44976 6298
rect 45072 6246 45080 6298
rect 44928 6244 44976 6246
rect 45032 6244 45080 6246
rect 45136 6298 45184 6300
rect 45240 6298 45288 6300
rect 45136 6246 45144 6298
rect 45240 6246 45268 6298
rect 45136 6244 45184 6246
rect 45240 6244 45288 6246
rect 45344 6244 45392 6300
rect 44768 6234 45448 6244
rect 44940 6132 44996 6142
rect 44940 5236 44996 6076
rect 44940 5142 44996 5180
rect 45276 5794 45332 5806
rect 45276 5742 45278 5794
rect 45330 5742 45332 5794
rect 45276 5012 45332 5742
rect 45724 5348 45780 6860
rect 45276 4946 45332 4956
rect 45612 5292 45780 5348
rect 45836 6692 45892 6702
rect 44604 4722 44660 4732
rect 44768 4732 45448 4742
rect 44824 4676 44872 4732
rect 44928 4730 44976 4732
rect 45032 4730 45080 4732
rect 44948 4678 44976 4730
rect 45072 4678 45080 4730
rect 44928 4676 44976 4678
rect 45032 4676 45080 4678
rect 45136 4730 45184 4732
rect 45240 4730 45288 4732
rect 45136 4678 45144 4730
rect 45240 4678 45268 4730
rect 45136 4676 45184 4678
rect 45240 4676 45288 4678
rect 45344 4676 45392 4732
rect 44768 4666 45448 4676
rect 45612 4564 45668 5292
rect 45836 5122 45892 6636
rect 46060 6690 46116 8316
rect 46284 8260 46340 8270
rect 46284 8166 46340 8204
rect 46060 6638 46062 6690
rect 46114 6638 46116 6690
rect 46060 6468 46116 6638
rect 46060 6402 46116 6412
rect 46172 8148 46228 8158
rect 45836 5070 45838 5122
rect 45890 5070 45892 5122
rect 45836 5058 45892 5070
rect 46172 5122 46228 8092
rect 46284 8036 46340 8046
rect 46284 6802 46340 7980
rect 46284 6750 46286 6802
rect 46338 6750 46340 6802
rect 46284 6738 46340 6750
rect 46396 6020 46452 11342
rect 46396 5954 46452 5964
rect 46284 5684 46340 5694
rect 46284 5234 46340 5628
rect 46284 5182 46286 5234
rect 46338 5182 46340 5234
rect 46284 5170 46340 5182
rect 46172 5070 46174 5122
rect 46226 5070 46228 5122
rect 46172 5058 46228 5070
rect 46508 4900 46564 12124
rect 44492 4508 44884 4564
rect 44828 3778 44884 4508
rect 44828 3726 44830 3778
rect 44882 3726 44884 3778
rect 44828 3714 44884 3726
rect 45164 4508 45668 4564
rect 45948 4844 46564 4900
rect 46620 4900 46676 4910
rect 45164 3778 45220 4508
rect 45164 3726 45166 3778
rect 45218 3726 45220 3778
rect 45164 3714 45220 3726
rect 45276 3780 45332 3790
rect 45276 3686 45332 3724
rect 45948 3778 46004 4844
rect 46620 4806 46676 4844
rect 45948 3726 45950 3778
rect 46002 3726 46004 3778
rect 45948 3714 46004 3726
rect 46844 3778 46900 12236
rect 47180 12068 47236 12078
rect 47068 11284 47124 11294
rect 47068 11190 47124 11228
rect 47180 10610 47236 12012
rect 47180 10558 47182 10610
rect 47234 10558 47236 10610
rect 47180 10546 47236 10558
rect 47068 9826 47124 9838
rect 47068 9774 47070 9826
rect 47122 9774 47124 9826
rect 47068 6804 47124 9774
rect 47068 6738 47124 6748
rect 46844 3726 46846 3778
rect 46898 3726 46900 3778
rect 46844 3714 46900 3726
rect 44268 3666 44436 3668
rect 44268 3614 44270 3666
rect 44322 3614 44436 3666
rect 44268 3612 44436 3614
rect 44268 3602 44324 3612
rect 43484 3502 43486 3554
rect 43538 3502 43540 3554
rect 43484 3490 43540 3502
rect 44380 3556 44436 3612
rect 47740 3666 47796 12796
rect 47852 12738 47908 12750
rect 47852 12686 47854 12738
rect 47906 12686 47908 12738
rect 47852 6690 47908 12686
rect 48076 7364 48132 12910
rect 48860 12292 48916 12302
rect 48860 12198 48916 12236
rect 48748 12180 48804 12190
rect 48748 12086 48804 12124
rect 48188 12068 48244 12078
rect 48188 11974 48244 12012
rect 48972 10052 49028 13916
rect 51660 13860 51716 13870
rect 51660 13746 51716 13804
rect 52444 13860 52500 27692
rect 52780 27076 52836 31892
rect 53116 31890 53172 32060
rect 53116 31838 53118 31890
rect 53170 31838 53172 31890
rect 53116 31826 53172 31838
rect 53116 29652 53172 29662
rect 53228 29652 53284 32284
rect 53452 32340 53508 32350
rect 53452 32246 53508 32284
rect 54460 32116 54516 32396
rect 54460 32050 54516 32060
rect 56700 32338 56756 32350
rect 56700 32286 56702 32338
rect 56754 32286 56756 32338
rect 56700 31948 56756 32286
rect 58268 32172 58948 32182
rect 58324 32116 58372 32172
rect 58428 32170 58476 32172
rect 58532 32170 58580 32172
rect 58448 32118 58476 32170
rect 58572 32118 58580 32170
rect 58428 32116 58476 32118
rect 58532 32116 58580 32118
rect 58636 32170 58684 32172
rect 58740 32170 58788 32172
rect 58636 32118 58644 32170
rect 58740 32118 58768 32170
rect 58636 32116 58684 32118
rect 58740 32116 58788 32118
rect 58844 32116 58892 32172
rect 58268 32106 58948 32116
rect 56140 31892 56756 31948
rect 56140 31778 56196 31892
rect 56140 31726 56142 31778
rect 56194 31726 56196 31778
rect 56140 31714 56196 31726
rect 55356 31556 55412 31566
rect 53768 31388 54448 31398
rect 53824 31332 53872 31388
rect 53928 31386 53976 31388
rect 54032 31386 54080 31388
rect 53948 31334 53976 31386
rect 54072 31334 54080 31386
rect 53928 31332 53976 31334
rect 54032 31332 54080 31334
rect 54136 31386 54184 31388
rect 54240 31386 54288 31388
rect 54136 31334 54144 31386
rect 54240 31334 54268 31386
rect 54136 31332 54184 31334
rect 54240 31332 54288 31334
rect 54344 31332 54392 31388
rect 53768 31322 54448 31332
rect 53768 29820 54448 29830
rect 53824 29764 53872 29820
rect 53928 29818 53976 29820
rect 54032 29818 54080 29820
rect 53948 29766 53976 29818
rect 54072 29766 54080 29818
rect 53928 29764 53976 29766
rect 54032 29764 54080 29766
rect 54136 29818 54184 29820
rect 54240 29818 54288 29820
rect 54136 29766 54144 29818
rect 54240 29766 54268 29818
rect 54136 29764 54184 29766
rect 54240 29764 54288 29766
rect 54344 29764 54392 29820
rect 53768 29754 54448 29764
rect 52892 29650 53284 29652
rect 52892 29598 53118 29650
rect 53170 29598 53284 29650
rect 52892 29596 53284 29598
rect 52892 28082 52948 29596
rect 53116 29586 53172 29596
rect 53228 29540 53284 29596
rect 53228 29474 53284 29484
rect 54236 29540 54292 29550
rect 54236 29446 54292 29484
rect 55244 29540 55300 29550
rect 54908 29428 54964 29438
rect 53676 29204 53732 29214
rect 53676 28756 53732 29148
rect 54908 28866 54964 29372
rect 54908 28814 54910 28866
rect 54962 28814 54964 28866
rect 54908 28802 54964 28814
rect 52892 28030 52894 28082
rect 52946 28030 52948 28082
rect 52892 27972 52948 28030
rect 53340 28700 53732 28756
rect 52948 27916 53060 27972
rect 52892 27906 52948 27916
rect 52780 27020 52948 27076
rect 52892 26404 52948 27020
rect 53004 26514 53060 27916
rect 53004 26462 53006 26514
rect 53058 26462 53060 26514
rect 53004 26450 53060 26462
rect 52892 26338 52948 26348
rect 53340 20188 53396 28700
rect 55020 28532 55076 28542
rect 55020 28438 55076 28476
rect 54572 28420 54628 28430
rect 54908 28420 54964 28430
rect 54572 28418 54964 28420
rect 54572 28366 54574 28418
rect 54626 28366 54910 28418
rect 54962 28366 54964 28418
rect 54572 28364 54964 28366
rect 53768 28252 54448 28262
rect 53824 28196 53872 28252
rect 53928 28250 53976 28252
rect 54032 28250 54080 28252
rect 53948 28198 53976 28250
rect 54072 28198 54080 28250
rect 53928 28196 53976 28198
rect 54032 28196 54080 28198
rect 54136 28250 54184 28252
rect 54240 28250 54288 28252
rect 54136 28198 54144 28250
rect 54240 28198 54268 28250
rect 54136 28196 54184 28198
rect 54240 28196 54288 28198
rect 54344 28196 54392 28252
rect 53768 28186 54448 28196
rect 53676 27972 53732 27982
rect 53676 27186 53732 27916
rect 53676 27134 53678 27186
rect 53730 27134 53732 27186
rect 53676 27122 53732 27134
rect 54572 27188 54628 28364
rect 54908 28354 54964 28364
rect 55020 28084 55076 28094
rect 55244 28084 55300 29484
rect 55356 28642 55412 31500
rect 55356 28590 55358 28642
rect 55410 28590 55412 28642
rect 55356 28578 55412 28590
rect 55804 31554 55860 31566
rect 55804 31502 55806 31554
rect 55858 31502 55860 31554
rect 55804 28642 55860 31502
rect 56476 31556 56532 31566
rect 56476 31462 56532 31500
rect 58268 30604 58948 30614
rect 58324 30548 58372 30604
rect 58428 30602 58476 30604
rect 58532 30602 58580 30604
rect 58448 30550 58476 30602
rect 58572 30550 58580 30602
rect 58428 30548 58476 30550
rect 58532 30548 58580 30550
rect 58636 30602 58684 30604
rect 58740 30602 58788 30604
rect 58636 30550 58644 30602
rect 58740 30550 58768 30602
rect 58636 30548 58684 30550
rect 58740 30548 58788 30550
rect 58844 30548 58892 30604
rect 58268 30538 58948 30548
rect 59052 29988 59108 29998
rect 59052 29894 59108 29932
rect 56028 29540 56084 29550
rect 56924 29540 56980 29550
rect 56028 29538 56196 29540
rect 56028 29486 56030 29538
rect 56082 29486 56196 29538
rect 56028 29484 56196 29486
rect 56028 29474 56084 29484
rect 55804 28590 55806 28642
rect 55858 28590 55860 28642
rect 55804 28578 55860 28590
rect 54572 27122 54628 27132
rect 54796 28082 56084 28084
rect 54796 28030 55022 28082
rect 55074 28030 56084 28082
rect 54796 28028 56084 28030
rect 53564 26852 53620 26862
rect 53564 26514 53620 26796
rect 54236 26852 54292 26862
rect 54236 26850 54628 26852
rect 54236 26798 54238 26850
rect 54290 26798 54628 26850
rect 54236 26796 54628 26798
rect 54236 26786 54292 26796
rect 53768 26684 54448 26694
rect 53824 26628 53872 26684
rect 53928 26682 53976 26684
rect 54032 26682 54080 26684
rect 53948 26630 53976 26682
rect 54072 26630 54080 26682
rect 53928 26628 53976 26630
rect 54032 26628 54080 26630
rect 54136 26682 54184 26684
rect 54240 26682 54288 26684
rect 54136 26630 54144 26682
rect 54240 26630 54268 26682
rect 54136 26628 54184 26630
rect 54240 26628 54288 26630
rect 54344 26628 54392 26684
rect 53768 26618 54448 26628
rect 53564 26462 53566 26514
rect 53618 26462 53620 26514
rect 53564 26450 53620 26462
rect 53452 26404 53508 26414
rect 53452 25618 53508 26348
rect 53788 26404 53844 26414
rect 53788 26310 53844 26348
rect 54572 26292 54628 26796
rect 53452 25566 53454 25618
rect 53506 25566 53508 25618
rect 53452 25554 53508 25566
rect 54236 26236 54628 26292
rect 54236 25506 54292 26236
rect 54796 26178 54852 28028
rect 55020 28018 55076 28028
rect 56028 27746 56084 28028
rect 56140 27860 56196 29484
rect 56924 29446 56980 29484
rect 57596 29540 57652 29550
rect 57596 29446 57652 29484
rect 56812 29428 56868 29438
rect 56812 29334 56868 29372
rect 57148 29426 57204 29438
rect 57148 29374 57150 29426
rect 57202 29374 57204 29426
rect 56924 28532 56980 28542
rect 56476 27860 56532 27870
rect 56140 27858 56532 27860
rect 56140 27806 56478 27858
rect 56530 27806 56532 27858
rect 56140 27804 56532 27806
rect 56476 27794 56532 27804
rect 56028 27694 56030 27746
rect 56082 27694 56084 27746
rect 56028 26740 56084 27694
rect 56924 27298 56980 28476
rect 57148 27858 57204 29374
rect 58268 29036 58948 29046
rect 58324 28980 58372 29036
rect 58428 29034 58476 29036
rect 58532 29034 58580 29036
rect 58448 28982 58476 29034
rect 58572 28982 58580 29034
rect 58428 28980 58476 28982
rect 58532 28980 58580 28982
rect 58636 29034 58684 29036
rect 58740 29034 58788 29036
rect 58636 28982 58644 29034
rect 58740 28982 58768 29034
rect 58636 28980 58684 28982
rect 58740 28980 58788 28982
rect 58844 28980 58892 29036
rect 59164 28980 59220 32508
rect 60284 32452 60340 33068
rect 60732 32788 60788 34524
rect 61516 34356 61572 34748
rect 61628 34356 61684 34366
rect 61516 34354 61684 34356
rect 61516 34302 61630 34354
rect 61682 34302 61684 34354
rect 61516 34300 61684 34302
rect 61628 34244 61684 34300
rect 61628 34178 61684 34188
rect 61068 34018 61124 34030
rect 61068 33966 61070 34018
rect 61122 33966 61124 34018
rect 61068 33572 61124 33966
rect 61740 33796 61796 34860
rect 61964 34850 62020 34860
rect 60844 33460 60900 33470
rect 60844 33366 60900 33404
rect 61068 32788 61124 33516
rect 61628 33740 61796 33796
rect 61516 33122 61572 33134
rect 61516 33070 61518 33122
rect 61570 33070 61572 33122
rect 61180 32788 61236 32798
rect 60732 32786 61012 32788
rect 60732 32734 60734 32786
rect 60786 32734 61012 32786
rect 60732 32732 61012 32734
rect 60732 32722 60788 32732
rect 60956 32564 61012 32732
rect 61124 32786 61236 32788
rect 61124 32734 61182 32786
rect 61234 32734 61236 32786
rect 61124 32732 61236 32734
rect 61068 32694 61124 32732
rect 61180 32722 61236 32732
rect 61404 32674 61460 32686
rect 61404 32622 61406 32674
rect 61458 32622 61460 32674
rect 61404 32564 61460 32622
rect 60956 32508 61460 32564
rect 60284 32358 60340 32396
rect 60396 31780 60452 31790
rect 59948 31778 60452 31780
rect 59948 31726 60398 31778
rect 60450 31726 60452 31778
rect 59948 31724 60452 31726
rect 59948 31666 60004 31724
rect 60396 31714 60452 31724
rect 61068 31780 61124 31790
rect 61068 31778 61236 31780
rect 61068 31726 61070 31778
rect 61122 31726 61236 31778
rect 61068 31724 61236 31726
rect 61068 31714 61124 31724
rect 59948 31614 59950 31666
rect 60002 31614 60004 31666
rect 59948 31602 60004 31614
rect 61180 31218 61236 31724
rect 61180 31166 61182 31218
rect 61234 31166 61236 31218
rect 61180 31154 61236 31166
rect 61516 30994 61572 33070
rect 61516 30942 61518 30994
rect 61570 30942 61572 30994
rect 61516 30930 61572 30942
rect 61628 29988 61684 33740
rect 62076 33460 62132 40908
rect 62768 40796 63448 40806
rect 62824 40740 62872 40796
rect 62928 40794 62976 40796
rect 63032 40794 63080 40796
rect 62948 40742 62976 40794
rect 63072 40742 63080 40794
rect 62928 40740 62976 40742
rect 63032 40740 63080 40742
rect 63136 40794 63184 40796
rect 63240 40794 63288 40796
rect 63136 40742 63144 40794
rect 63240 40742 63268 40794
rect 63136 40740 63184 40742
rect 63240 40740 63288 40742
rect 63344 40740 63392 40796
rect 62768 40730 63448 40740
rect 62768 39228 63448 39238
rect 62824 39172 62872 39228
rect 62928 39226 62976 39228
rect 63032 39226 63080 39228
rect 62948 39174 62976 39226
rect 63072 39174 63080 39226
rect 62928 39172 62976 39174
rect 63032 39172 63080 39174
rect 63136 39226 63184 39228
rect 63240 39226 63288 39228
rect 63136 39174 63144 39226
rect 63240 39174 63268 39226
rect 63136 39172 63184 39174
rect 63240 39172 63288 39174
rect 63344 39172 63392 39228
rect 62768 39162 63448 39172
rect 63868 38388 63924 38398
rect 63308 38052 63364 38062
rect 63084 38050 63364 38052
rect 63084 37998 63310 38050
rect 63362 37998 63364 38050
rect 63084 37996 63364 37998
rect 63084 37938 63140 37996
rect 63308 37986 63364 37996
rect 63084 37886 63086 37938
rect 63138 37886 63140 37938
rect 63084 37874 63140 37886
rect 62768 37660 63448 37670
rect 62824 37604 62872 37660
rect 62928 37658 62976 37660
rect 63032 37658 63080 37660
rect 62948 37606 62976 37658
rect 63072 37606 63080 37658
rect 62928 37604 62976 37606
rect 63032 37604 63080 37606
rect 63136 37658 63184 37660
rect 63240 37658 63288 37660
rect 63136 37606 63144 37658
rect 63240 37606 63268 37658
rect 63136 37604 63184 37606
rect 63240 37604 63288 37606
rect 63344 37604 63392 37660
rect 62768 37594 63448 37604
rect 63868 37490 63924 38332
rect 64428 38388 64484 42252
rect 64652 41188 64708 41198
rect 64652 41094 64708 41132
rect 64652 39844 64708 39854
rect 64428 38322 64484 38332
rect 64540 38836 64596 38846
rect 63980 38052 64036 38062
rect 63980 38050 64484 38052
rect 63980 37998 63982 38050
rect 64034 37998 64484 38050
rect 63980 37996 64484 37998
rect 63980 37986 64036 37996
rect 63868 37438 63870 37490
rect 63922 37438 63924 37490
rect 63868 37156 63924 37438
rect 64428 37490 64484 37996
rect 64428 37438 64430 37490
rect 64482 37438 64484 37490
rect 64428 37426 64484 37438
rect 63868 37090 63924 37100
rect 62768 36092 63448 36102
rect 62824 36036 62872 36092
rect 62928 36090 62976 36092
rect 63032 36090 63080 36092
rect 62948 36038 62976 36090
rect 63072 36038 63080 36090
rect 62928 36036 62976 36038
rect 63032 36036 63080 36038
rect 63136 36090 63184 36092
rect 63240 36090 63288 36092
rect 63136 36038 63144 36090
rect 63240 36038 63268 36090
rect 63136 36036 63184 36038
rect 63240 36036 63288 36038
rect 63344 36036 63392 36092
rect 62768 36026 63448 36036
rect 62972 35810 63028 35822
rect 62972 35758 62974 35810
rect 63026 35758 63028 35810
rect 62636 35700 62692 35710
rect 62188 35698 62692 35700
rect 62188 35646 62638 35698
rect 62690 35646 62692 35698
rect 62188 35644 62692 35646
rect 62188 34354 62244 35644
rect 62636 35634 62692 35644
rect 62972 34692 63028 35758
rect 64540 35700 64596 38780
rect 64540 35634 64596 35644
rect 64316 35028 64372 35038
rect 64652 35028 64708 39788
rect 64764 38668 64820 47964
rect 64988 46788 65044 46798
rect 64988 46694 65044 46732
rect 64876 46676 64932 46686
rect 64876 45890 64932 46620
rect 65212 46674 65268 48078
rect 67268 47852 67948 47862
rect 67324 47796 67372 47852
rect 67428 47850 67476 47852
rect 67532 47850 67580 47852
rect 67448 47798 67476 47850
rect 67572 47798 67580 47850
rect 67428 47796 67476 47798
rect 67532 47796 67580 47798
rect 67636 47850 67684 47852
rect 67740 47850 67788 47852
rect 67636 47798 67644 47850
rect 67740 47798 67768 47850
rect 67636 47796 67684 47798
rect 67740 47796 67788 47798
rect 67844 47796 67892 47852
rect 67268 47786 67948 47796
rect 71036 47458 71092 48302
rect 71036 47406 71038 47458
rect 71090 47406 71092 47458
rect 71036 47394 71092 47406
rect 65436 46788 65492 46798
rect 65436 46694 65492 46732
rect 67564 46786 67620 46798
rect 67564 46734 67566 46786
rect 67618 46734 67620 46786
rect 65212 46622 65214 46674
rect 65266 46622 65268 46674
rect 65212 46610 65268 46622
rect 65772 46676 65828 46686
rect 65772 46582 65828 46620
rect 66444 46674 66500 46686
rect 66444 46622 66446 46674
rect 66498 46622 66500 46674
rect 64876 45838 64878 45890
rect 64930 45838 64932 45890
rect 64876 45826 64932 45838
rect 65324 45892 65380 45902
rect 65324 45666 65380 45836
rect 65324 45614 65326 45666
rect 65378 45614 65380 45666
rect 65212 44212 65268 44222
rect 65212 44118 65268 44156
rect 64988 43426 65044 43438
rect 64988 43374 64990 43426
rect 65042 43374 65044 43426
rect 64988 42868 65044 43374
rect 64988 42802 65044 42812
rect 64988 42532 65044 42542
rect 64988 42438 65044 42476
rect 65212 41188 65268 41198
rect 65212 40626 65268 41132
rect 65212 40574 65214 40626
rect 65266 40574 65268 40626
rect 65212 40562 65268 40574
rect 65324 39844 65380 45614
rect 65884 44212 65940 44222
rect 65884 43652 65940 44156
rect 65996 43652 66052 43662
rect 65884 43650 66052 43652
rect 65884 43598 65998 43650
rect 66050 43598 66052 43650
rect 65884 43596 66052 43598
rect 65436 43540 65492 43550
rect 65772 43540 65828 43550
rect 65436 43446 65492 43484
rect 65660 43538 65828 43540
rect 65660 43486 65774 43538
rect 65826 43486 65828 43538
rect 65660 43484 65828 43486
rect 65548 43428 65604 43438
rect 65548 42084 65604 43372
rect 65660 42868 65716 43484
rect 65772 43474 65828 43484
rect 65772 42980 65828 42990
rect 65884 42980 65940 43596
rect 65996 43586 66052 43596
rect 65772 42978 65940 42980
rect 65772 42926 65774 42978
rect 65826 42926 65940 42978
rect 65772 42924 65940 42926
rect 66332 43538 66388 43550
rect 66332 43486 66334 43538
rect 66386 43486 66388 43538
rect 66332 43428 66388 43486
rect 65772 42914 65828 42924
rect 65660 42802 65716 42812
rect 66332 42756 66388 43372
rect 66444 43314 66500 46622
rect 67564 46564 67620 46734
rect 67564 46508 68068 46564
rect 66780 46452 66836 46462
rect 66780 46358 66836 46396
rect 67268 46284 67948 46294
rect 67324 46228 67372 46284
rect 67428 46282 67476 46284
rect 67532 46282 67580 46284
rect 67448 46230 67476 46282
rect 67572 46230 67580 46282
rect 67428 46228 67476 46230
rect 67532 46228 67580 46230
rect 67636 46282 67684 46284
rect 67740 46282 67788 46284
rect 67636 46230 67644 46282
rect 67740 46230 67768 46282
rect 67636 46228 67684 46230
rect 67740 46228 67788 46230
rect 67844 46228 67892 46284
rect 67268 46218 67948 46228
rect 68012 45892 68068 46508
rect 68236 45892 68292 45902
rect 68796 45892 68852 45902
rect 68012 45890 68292 45892
rect 68012 45838 68238 45890
rect 68290 45838 68292 45890
rect 68012 45836 68292 45838
rect 68236 45826 68292 45836
rect 68572 45890 68852 45892
rect 68572 45838 68798 45890
rect 68850 45838 68852 45890
rect 68572 45836 68852 45838
rect 67788 45666 67844 45678
rect 67788 45614 67790 45666
rect 67842 45614 67844 45666
rect 67788 45444 67844 45614
rect 67844 45388 68068 45444
rect 67788 45378 67844 45388
rect 67268 44716 67948 44726
rect 67324 44660 67372 44716
rect 67428 44714 67476 44716
rect 67532 44714 67580 44716
rect 67448 44662 67476 44714
rect 67572 44662 67580 44714
rect 67428 44660 67476 44662
rect 67532 44660 67580 44662
rect 67636 44714 67684 44716
rect 67740 44714 67788 44716
rect 67636 44662 67644 44714
rect 67740 44662 67768 44714
rect 67636 44660 67684 44662
rect 67740 44660 67788 44662
rect 67844 44660 67892 44716
rect 67268 44650 67948 44660
rect 66444 43262 66446 43314
rect 66498 43262 66500 43314
rect 66444 43250 66500 43262
rect 67004 43540 67060 43550
rect 66668 42868 66724 42878
rect 66444 42756 66500 42766
rect 66332 42700 66444 42756
rect 66444 42690 66500 42700
rect 65324 39778 65380 39788
rect 65436 42028 65604 42084
rect 64764 38612 65380 38668
rect 64764 37268 64820 37278
rect 65212 37268 65268 37278
rect 64764 37266 65268 37268
rect 64764 37214 64766 37266
rect 64818 37214 65214 37266
rect 65266 37214 65268 37266
rect 64764 37212 65268 37214
rect 64764 37202 64820 37212
rect 65212 37202 65268 37212
rect 64876 36596 64932 36606
rect 64876 36502 64932 36540
rect 62972 34636 63588 34692
rect 62768 34524 63448 34534
rect 62824 34468 62872 34524
rect 62928 34522 62976 34524
rect 63032 34522 63080 34524
rect 62948 34470 62976 34522
rect 63072 34470 63080 34522
rect 62928 34468 62976 34470
rect 63032 34468 63080 34470
rect 63136 34522 63184 34524
rect 63240 34522 63288 34524
rect 63136 34470 63144 34522
rect 63240 34470 63268 34522
rect 63136 34468 63184 34470
rect 63240 34468 63288 34470
rect 63344 34468 63392 34524
rect 62768 34458 63448 34468
rect 63532 34468 63588 34636
rect 63532 34412 63924 34468
rect 62188 34302 62190 34354
rect 62242 34302 62244 34354
rect 62188 34290 62244 34302
rect 62972 34244 63028 34254
rect 62972 34130 63028 34188
rect 62972 34078 62974 34130
rect 63026 34078 63028 34130
rect 62972 34066 63028 34078
rect 63084 34242 63140 34254
rect 63084 34190 63086 34242
rect 63138 34190 63140 34242
rect 61852 33348 61908 33358
rect 61852 33254 61908 33292
rect 62076 33234 62132 33404
rect 62524 33906 62580 33918
rect 62524 33854 62526 33906
rect 62578 33854 62580 33906
rect 62524 33572 62580 33854
rect 62076 33182 62078 33234
rect 62130 33182 62132 33234
rect 62076 33170 62132 33182
rect 62412 33348 62468 33358
rect 61740 32564 61796 32574
rect 62412 32564 62468 33292
rect 62524 33234 62580 33516
rect 62524 33182 62526 33234
rect 62578 33182 62580 33234
rect 62524 33170 62580 33182
rect 63084 33124 63140 34190
rect 63756 34242 63812 34254
rect 63756 34190 63758 34242
rect 63810 34190 63812 34242
rect 63756 34132 63812 34190
rect 63196 34076 63812 34132
rect 63196 33346 63252 34076
rect 63868 34020 63924 34412
rect 64316 34130 64372 34972
rect 64316 34078 64318 34130
rect 64370 34078 64372 34130
rect 64316 34066 64372 34078
rect 64540 34972 64708 35028
rect 63196 33294 63198 33346
rect 63250 33294 63252 33346
rect 63196 33282 63252 33294
rect 63532 33964 63924 34020
rect 63532 33346 63588 33964
rect 63532 33294 63534 33346
rect 63586 33294 63588 33346
rect 63532 33282 63588 33294
rect 63644 33684 63700 33694
rect 63196 33124 63252 33134
rect 63084 33068 63196 33124
rect 63196 33058 63252 33068
rect 62768 32956 63448 32966
rect 62824 32900 62872 32956
rect 62928 32954 62976 32956
rect 63032 32954 63080 32956
rect 62948 32902 62976 32954
rect 63072 32902 63080 32954
rect 62928 32900 62976 32902
rect 63032 32900 63080 32902
rect 63136 32954 63184 32956
rect 63240 32954 63288 32956
rect 63136 32902 63144 32954
rect 63240 32902 63268 32954
rect 63136 32900 63184 32902
rect 63240 32900 63288 32902
rect 63344 32900 63392 32956
rect 62768 32890 63448 32900
rect 63308 32676 63364 32686
rect 63308 32582 63364 32620
rect 62524 32564 62580 32574
rect 62412 32562 62580 32564
rect 62412 32510 62526 32562
rect 62578 32510 62580 32562
rect 62412 32508 62580 32510
rect 61740 32470 61796 32508
rect 62524 32004 62580 32508
rect 62972 32564 63028 32574
rect 62972 32470 63028 32508
rect 63084 32452 63140 32462
rect 63644 32452 63700 33628
rect 63756 33124 63812 33134
rect 63756 32786 63812 33068
rect 63756 32734 63758 32786
rect 63810 32734 63812 32786
rect 63756 32722 63812 32734
rect 64540 32564 64596 34972
rect 64652 34804 64708 34814
rect 65324 34804 65380 38612
rect 65436 36372 65492 42028
rect 65996 40964 66052 40974
rect 65996 40626 66052 40908
rect 65996 40574 65998 40626
rect 66050 40574 66052 40626
rect 65996 40562 66052 40574
rect 66108 40516 66164 40526
rect 65548 40404 65604 40414
rect 65548 40310 65604 40348
rect 66108 39394 66164 40460
rect 66556 40404 66612 40414
rect 66556 40310 66612 40348
rect 66108 39342 66110 39394
rect 66162 39342 66164 39394
rect 65548 39060 65604 39070
rect 66108 39060 66164 39342
rect 65604 39004 66164 39060
rect 66668 39060 66724 42812
rect 67004 42196 67060 43484
rect 67268 43148 67948 43158
rect 67324 43092 67372 43148
rect 67428 43146 67476 43148
rect 67532 43146 67580 43148
rect 67448 43094 67476 43146
rect 67572 43094 67580 43146
rect 67428 43092 67476 43094
rect 67532 43092 67580 43094
rect 67636 43146 67684 43148
rect 67740 43146 67788 43148
rect 67636 43094 67644 43146
rect 67740 43094 67768 43146
rect 67636 43092 67684 43094
rect 67740 43092 67788 43094
rect 67844 43092 67892 43148
rect 67268 43082 67948 43092
rect 68012 42980 68068 45388
rect 68572 45330 68628 45836
rect 68796 45826 68852 45836
rect 68572 45278 68574 45330
rect 68626 45278 68628 45330
rect 68572 45266 68628 45278
rect 70476 45668 70532 45678
rect 68908 45108 68964 45118
rect 68908 45014 68964 45052
rect 70140 45108 70196 45118
rect 70140 45014 70196 45052
rect 70476 45106 70532 45612
rect 71260 45444 71316 48972
rect 72156 49028 72212 49038
rect 72156 48934 72212 48972
rect 72716 49028 72772 49534
rect 71820 48916 71876 48926
rect 71820 48822 71876 48860
rect 71768 48636 72448 48646
rect 71824 48580 71872 48636
rect 71928 48634 71976 48636
rect 72032 48634 72080 48636
rect 71948 48582 71976 48634
rect 72072 48582 72080 48634
rect 71928 48580 71976 48582
rect 72032 48580 72080 48582
rect 72136 48634 72184 48636
rect 72240 48634 72288 48636
rect 72136 48582 72144 48634
rect 72240 48582 72268 48634
rect 72136 48580 72184 48582
rect 72240 48580 72288 48582
rect 72344 48580 72392 48636
rect 71768 48570 72448 48580
rect 71372 48354 71428 48366
rect 71372 48302 71374 48354
rect 71426 48302 71428 48354
rect 71372 47460 71428 48302
rect 71708 48244 71764 48254
rect 71708 48150 71764 48188
rect 72380 48244 72436 48254
rect 72380 48150 72436 48188
rect 72716 48242 72772 48972
rect 73836 49476 73892 49868
rect 73948 49476 74004 50430
rect 74284 50484 74340 50654
rect 74284 50418 74340 50428
rect 74956 50484 75012 50494
rect 73836 49420 74004 49476
rect 73500 48804 73556 48814
rect 73500 48802 73668 48804
rect 73500 48750 73502 48802
rect 73554 48750 73668 48802
rect 73500 48748 73668 48750
rect 73500 48738 73556 48748
rect 72716 48190 72718 48242
rect 72770 48190 72772 48242
rect 72716 48178 72772 48190
rect 72940 48692 72996 48702
rect 72940 48354 72996 48636
rect 72940 48302 72942 48354
rect 72994 48302 72996 48354
rect 72940 48020 72996 48302
rect 73500 48354 73556 48366
rect 73500 48302 73502 48354
rect 73554 48302 73556 48354
rect 73500 48244 73556 48302
rect 73612 48356 73668 48748
rect 73836 48580 73892 49420
rect 73948 48804 74004 48814
rect 73948 48802 74116 48804
rect 73948 48750 73950 48802
rect 74002 48750 74116 48802
rect 73948 48748 74116 48750
rect 73948 48738 74004 48748
rect 73836 48524 74004 48580
rect 73612 48290 73668 48300
rect 73948 48354 74004 48524
rect 74060 48468 74116 48748
rect 74060 48402 74116 48412
rect 74620 48468 74676 48478
rect 73948 48302 73950 48354
rect 74002 48302 74004 48354
rect 73948 48290 74004 48302
rect 74172 48356 74228 48366
rect 74172 48262 74228 48300
rect 73500 48178 73556 48188
rect 74396 48244 74452 48254
rect 72940 47954 72996 47964
rect 74284 48130 74340 48142
rect 74284 48078 74286 48130
rect 74338 48078 74340 48130
rect 71484 47460 71540 47470
rect 71372 47458 71540 47460
rect 71372 47406 71486 47458
rect 71538 47406 71540 47458
rect 71372 47404 71540 47406
rect 71484 47394 71540 47404
rect 74060 47236 74116 47246
rect 74060 47142 74116 47180
rect 71768 47068 72448 47078
rect 71824 47012 71872 47068
rect 71928 47066 71976 47068
rect 72032 47066 72080 47068
rect 71948 47014 71976 47066
rect 72072 47014 72080 47066
rect 71928 47012 71976 47014
rect 72032 47012 72080 47014
rect 72136 47066 72184 47068
rect 72240 47066 72288 47068
rect 72136 47014 72144 47066
rect 72240 47014 72268 47066
rect 72136 47012 72184 47014
rect 72240 47012 72288 47014
rect 72344 47012 72392 47068
rect 71768 47002 72448 47012
rect 74284 47012 74340 48078
rect 74396 47684 74452 48188
rect 74620 48242 74676 48412
rect 74620 48190 74622 48242
rect 74674 48190 74676 48242
rect 74620 48132 74676 48190
rect 74620 48066 74676 48076
rect 74620 47684 74676 47694
rect 74396 47682 74676 47684
rect 74396 47630 74622 47682
rect 74674 47630 74676 47682
rect 74396 47628 74676 47630
rect 74620 47618 74676 47628
rect 74956 47570 75012 50428
rect 75740 50034 75796 53452
rect 80768 53340 81448 53350
rect 80824 53284 80872 53340
rect 80928 53338 80976 53340
rect 81032 53338 81080 53340
rect 80948 53286 80976 53338
rect 81072 53286 81080 53338
rect 80928 53284 80976 53286
rect 81032 53284 81080 53286
rect 81136 53338 81184 53340
rect 81240 53338 81288 53340
rect 81136 53286 81144 53338
rect 81240 53286 81268 53338
rect 81136 53284 81184 53286
rect 81240 53284 81288 53286
rect 81344 53284 81392 53340
rect 80768 53274 81448 53284
rect 81452 52836 81508 52846
rect 81564 52836 81620 54348
rect 85268 54124 85948 54134
rect 85324 54068 85372 54124
rect 85428 54122 85476 54124
rect 85532 54122 85580 54124
rect 85448 54070 85476 54122
rect 85572 54070 85580 54122
rect 85428 54068 85476 54070
rect 85532 54068 85580 54070
rect 85636 54122 85684 54124
rect 85740 54122 85788 54124
rect 85636 54070 85644 54122
rect 85740 54070 85768 54122
rect 85636 54068 85684 54070
rect 85740 54068 85788 54070
rect 85844 54068 85892 54124
rect 85268 54058 85948 54068
rect 94268 54124 94948 54134
rect 94324 54068 94372 54124
rect 94428 54122 94476 54124
rect 94532 54122 94580 54124
rect 94448 54070 94476 54122
rect 94572 54070 94580 54122
rect 94428 54068 94476 54070
rect 94532 54068 94580 54070
rect 94636 54122 94684 54124
rect 94740 54122 94788 54124
rect 94636 54070 94644 54122
rect 94740 54070 94768 54122
rect 94636 54068 94684 54070
rect 94740 54068 94788 54070
rect 94844 54068 94892 54124
rect 94268 54058 94948 54068
rect 89768 53340 90448 53350
rect 89824 53284 89872 53340
rect 89928 53338 89976 53340
rect 90032 53338 90080 53340
rect 89948 53286 89976 53338
rect 90072 53286 90080 53338
rect 89928 53284 89976 53286
rect 90032 53284 90080 53286
rect 90136 53338 90184 53340
rect 90240 53338 90288 53340
rect 90136 53286 90144 53338
rect 90240 53286 90268 53338
rect 90136 53284 90184 53286
rect 90240 53284 90288 53286
rect 90344 53284 90392 53340
rect 89768 53274 90448 53284
rect 81508 52780 81620 52836
rect 81452 52770 81508 52780
rect 76268 52556 76948 52566
rect 76324 52500 76372 52556
rect 76428 52554 76476 52556
rect 76532 52554 76580 52556
rect 76448 52502 76476 52554
rect 76572 52502 76580 52554
rect 76428 52500 76476 52502
rect 76532 52500 76580 52502
rect 76636 52554 76684 52556
rect 76740 52554 76788 52556
rect 76636 52502 76644 52554
rect 76740 52502 76768 52554
rect 76636 52500 76684 52502
rect 76740 52500 76788 52502
rect 76844 52500 76892 52556
rect 76268 52490 76948 52500
rect 85268 52556 85948 52566
rect 85324 52500 85372 52556
rect 85428 52554 85476 52556
rect 85532 52554 85580 52556
rect 85448 52502 85476 52554
rect 85572 52502 85580 52554
rect 85428 52500 85476 52502
rect 85532 52500 85580 52502
rect 85636 52554 85684 52556
rect 85740 52554 85788 52556
rect 85636 52502 85644 52554
rect 85740 52502 85768 52554
rect 85636 52500 85684 52502
rect 85740 52500 85788 52502
rect 85844 52500 85892 52556
rect 85268 52490 85948 52500
rect 94268 52556 94948 52566
rect 94324 52500 94372 52556
rect 94428 52554 94476 52556
rect 94532 52554 94580 52556
rect 94448 52502 94476 52554
rect 94572 52502 94580 52554
rect 94428 52500 94476 52502
rect 94532 52500 94580 52502
rect 94636 52554 94684 52556
rect 94740 52554 94788 52556
rect 94636 52502 94644 52554
rect 94740 52502 94768 52554
rect 94636 52500 94684 52502
rect 94740 52500 94788 52502
rect 94844 52500 94892 52556
rect 94268 52490 94948 52500
rect 80768 51772 81448 51782
rect 80824 51716 80872 51772
rect 80928 51770 80976 51772
rect 81032 51770 81080 51772
rect 80948 51718 80976 51770
rect 81072 51718 81080 51770
rect 80928 51716 80976 51718
rect 81032 51716 81080 51718
rect 81136 51770 81184 51772
rect 81240 51770 81288 51772
rect 81136 51718 81144 51770
rect 81240 51718 81268 51770
rect 81136 51716 81184 51718
rect 81240 51716 81288 51718
rect 81344 51716 81392 51772
rect 80768 51706 81448 51716
rect 89768 51772 90448 51782
rect 89824 51716 89872 51772
rect 89928 51770 89976 51772
rect 90032 51770 90080 51772
rect 89948 51718 89976 51770
rect 90072 51718 90080 51770
rect 89928 51716 89976 51718
rect 90032 51716 90080 51718
rect 90136 51770 90184 51772
rect 90240 51770 90288 51772
rect 90136 51718 90144 51770
rect 90240 51718 90268 51770
rect 90136 51716 90184 51718
rect 90240 51716 90288 51718
rect 90344 51716 90392 51772
rect 89768 51706 90448 51716
rect 90972 51604 91028 51614
rect 90972 51510 91028 51548
rect 77084 51490 77140 51502
rect 77084 51438 77086 51490
rect 77138 51438 77140 51490
rect 76636 51268 76692 51278
rect 76636 51174 76692 51212
rect 76268 50988 76948 50998
rect 76324 50932 76372 50988
rect 76428 50986 76476 50988
rect 76532 50986 76580 50988
rect 76448 50934 76476 50986
rect 76572 50934 76580 50986
rect 76428 50932 76476 50934
rect 76532 50932 76580 50934
rect 76636 50986 76684 50988
rect 76740 50986 76788 50988
rect 76636 50934 76644 50986
rect 76740 50934 76768 50986
rect 76636 50932 76684 50934
rect 76740 50932 76788 50934
rect 76844 50932 76892 50988
rect 76268 50922 76948 50932
rect 76300 50596 76356 50606
rect 76524 50596 76580 50606
rect 76300 50594 76468 50596
rect 76300 50542 76302 50594
rect 76354 50542 76468 50594
rect 76300 50540 76468 50542
rect 76300 50530 76356 50540
rect 76412 50148 76468 50540
rect 76524 50482 76580 50540
rect 76972 50596 77028 50606
rect 77084 50596 77140 51438
rect 90748 51378 90804 51390
rect 90748 51326 90750 51378
rect 90802 51326 90804 51378
rect 79660 51268 79716 51278
rect 76972 50594 77140 50596
rect 76972 50542 76974 50594
rect 77026 50542 77140 50594
rect 76972 50540 77140 50542
rect 77308 50596 77364 50606
rect 76972 50530 77028 50540
rect 77308 50502 77364 50540
rect 76524 50430 76526 50482
rect 76578 50430 76580 50482
rect 76524 50418 76580 50430
rect 77980 50484 78036 50494
rect 77756 50372 78036 50428
rect 79660 50482 79716 51212
rect 85268 50988 85948 50998
rect 85324 50932 85372 50988
rect 85428 50986 85476 50988
rect 85532 50986 85580 50988
rect 85448 50934 85476 50986
rect 85572 50934 85580 50986
rect 85428 50932 85476 50934
rect 85532 50932 85580 50934
rect 85636 50986 85684 50988
rect 85740 50986 85788 50988
rect 85636 50934 85644 50986
rect 85740 50934 85768 50986
rect 85636 50932 85684 50934
rect 85740 50932 85788 50934
rect 85844 50932 85892 50988
rect 85268 50922 85948 50932
rect 79660 50430 79662 50482
rect 79714 50430 79716 50482
rect 79660 50428 79716 50430
rect 80444 50484 80500 50494
rect 79660 50372 79828 50428
rect 80444 50390 80500 50428
rect 86828 50372 86884 50382
rect 76412 50092 76916 50148
rect 75740 49982 75742 50034
rect 75794 49982 75796 50034
rect 75740 49812 75796 49982
rect 76860 50034 76916 50092
rect 76860 49982 76862 50034
rect 76914 49982 76916 50034
rect 76860 49970 76916 49982
rect 77420 49922 77476 49934
rect 77420 49870 77422 49922
rect 77474 49870 77476 49922
rect 75740 49746 75796 49756
rect 77196 49812 77252 49822
rect 77196 49718 77252 49756
rect 76188 49700 76244 49710
rect 76188 49606 76244 49644
rect 77420 49700 77476 49870
rect 77756 49922 77812 50372
rect 77756 49870 77758 49922
rect 77810 49870 77812 49922
rect 77420 49634 77476 49644
rect 77644 49812 77700 49822
rect 76268 49420 76948 49430
rect 76324 49364 76372 49420
rect 76428 49418 76476 49420
rect 76532 49418 76580 49420
rect 76448 49366 76476 49418
rect 76572 49366 76580 49418
rect 76428 49364 76476 49366
rect 76532 49364 76580 49366
rect 76636 49418 76684 49420
rect 76740 49418 76788 49420
rect 76636 49366 76644 49418
rect 76740 49366 76768 49418
rect 76636 49364 76684 49366
rect 76740 49364 76788 49366
rect 76844 49364 76892 49420
rect 76268 49354 76948 49364
rect 77644 49140 77700 49756
rect 77644 49046 77700 49084
rect 77196 48356 77252 48366
rect 77196 48262 77252 48300
rect 77644 48356 77700 48366
rect 77756 48356 77812 49870
rect 77644 48354 77812 48356
rect 77644 48302 77646 48354
rect 77698 48302 77812 48354
rect 77644 48300 77812 48302
rect 77980 49140 78036 49150
rect 77644 48290 77700 48300
rect 76412 48244 76468 48254
rect 76412 48150 76468 48188
rect 76972 48242 77028 48254
rect 76972 48190 76974 48242
rect 77026 48190 77028 48242
rect 75964 48132 76020 48142
rect 74956 47518 74958 47570
rect 75010 47518 75012 47570
rect 74956 47236 75012 47518
rect 75292 47684 75348 47694
rect 75012 47180 75236 47236
rect 74956 47170 75012 47180
rect 74284 46956 75012 47012
rect 73724 46786 73780 46798
rect 73724 46734 73726 46786
rect 73778 46734 73780 46786
rect 73052 46676 73108 46686
rect 73052 46114 73108 46620
rect 73052 46062 73054 46114
rect 73106 46062 73108 46114
rect 73052 46050 73108 46062
rect 73388 46564 73444 46574
rect 73724 46564 73780 46734
rect 73948 46676 74004 46686
rect 74508 46676 74564 46686
rect 73948 46674 74116 46676
rect 73948 46622 73950 46674
rect 74002 46622 74116 46674
rect 73948 46620 74116 46622
rect 73948 46610 74004 46620
rect 73388 46562 73780 46564
rect 73388 46510 73390 46562
rect 73442 46510 73780 46562
rect 73388 46508 73780 46510
rect 72716 45892 72772 45902
rect 72940 45892 72996 45902
rect 72716 45890 72940 45892
rect 72716 45838 72718 45890
rect 72770 45838 72940 45890
rect 72716 45836 72940 45838
rect 72716 45826 72772 45836
rect 72940 45798 72996 45836
rect 73388 45780 73444 46508
rect 73388 45714 73444 45724
rect 70476 45054 70478 45106
rect 70530 45054 70532 45106
rect 70476 45042 70532 45054
rect 71148 45388 71316 45444
rect 71372 45666 71428 45678
rect 71372 45614 71374 45666
rect 71426 45614 71428 45666
rect 71372 45444 71428 45614
rect 71932 45668 71988 45706
rect 71932 45602 71988 45612
rect 73052 45668 73108 45678
rect 73052 45574 73108 45612
rect 71768 45500 72448 45510
rect 71824 45444 71872 45500
rect 71928 45498 71976 45500
rect 72032 45498 72080 45500
rect 71948 45446 71976 45498
rect 72072 45446 72080 45498
rect 71928 45444 71976 45446
rect 72032 45444 72080 45446
rect 72136 45498 72184 45500
rect 72240 45498 72288 45500
rect 72136 45446 72144 45498
rect 72240 45446 72268 45498
rect 72136 45444 72184 45446
rect 72240 45444 72288 45446
rect 72344 45444 72392 45500
rect 71768 45434 72448 45444
rect 71148 45218 71204 45388
rect 71372 45378 71428 45388
rect 71148 45166 71150 45218
rect 71202 45166 71204 45218
rect 69468 44996 69524 45006
rect 69468 44902 69524 44940
rect 69692 44324 69748 44334
rect 71148 44324 71204 45166
rect 71260 45108 71316 45118
rect 71260 45014 71316 45052
rect 73612 44996 73668 45006
rect 73612 44902 73668 44940
rect 74060 44546 74116 46620
rect 74508 46582 74564 46620
rect 74956 46674 75012 46956
rect 74956 46622 74958 46674
rect 75010 46622 75012 46674
rect 74956 46610 75012 46622
rect 74060 44494 74062 44546
rect 74114 44494 74116 44546
rect 74060 44482 74116 44494
rect 74508 44996 74564 45006
rect 71260 44324 71316 44334
rect 71148 44268 71260 44324
rect 69692 44230 69748 44268
rect 71260 43762 71316 44268
rect 73612 44324 73668 44334
rect 73612 44230 73668 44268
rect 73836 44322 73892 44334
rect 73836 44270 73838 44322
rect 73890 44270 73892 44322
rect 73052 44100 73108 44110
rect 73276 44100 73332 44110
rect 73052 44006 73108 44044
rect 73164 44044 73276 44100
rect 71768 43932 72448 43942
rect 71824 43876 71872 43932
rect 71928 43930 71976 43932
rect 72032 43930 72080 43932
rect 71948 43878 71976 43930
rect 72072 43878 72080 43930
rect 71928 43876 71976 43878
rect 72032 43876 72080 43878
rect 72136 43930 72184 43932
rect 72240 43930 72288 43932
rect 72136 43878 72144 43930
rect 72240 43878 72268 43930
rect 72136 43876 72184 43878
rect 72240 43876 72288 43878
rect 72344 43876 72392 43932
rect 71768 43866 72448 43876
rect 71260 43710 71262 43762
rect 71314 43710 71316 43762
rect 67788 42924 68068 42980
rect 69916 43650 69972 43662
rect 70364 43652 70420 43662
rect 69916 43598 69918 43650
rect 69970 43598 69972 43650
rect 67060 42140 67172 42196
rect 67004 42130 67060 42140
rect 67004 41972 67060 41982
rect 67004 40962 67060 41916
rect 67116 41412 67172 42140
rect 67788 41972 67844 42924
rect 67900 42756 67956 42766
rect 69804 42756 69860 42766
rect 69916 42756 69972 43598
rect 67956 42700 68068 42756
rect 67900 42690 67956 42700
rect 67788 41878 67844 41916
rect 67268 41580 67948 41590
rect 67324 41524 67372 41580
rect 67428 41578 67476 41580
rect 67532 41578 67580 41580
rect 67448 41526 67476 41578
rect 67572 41526 67580 41578
rect 67428 41524 67476 41526
rect 67532 41524 67580 41526
rect 67636 41578 67684 41580
rect 67740 41578 67788 41580
rect 67636 41526 67644 41578
rect 67740 41526 67768 41578
rect 67636 41524 67684 41526
rect 67740 41524 67788 41526
rect 67844 41524 67892 41580
rect 67268 41514 67948 41524
rect 67116 41356 67284 41412
rect 67004 40910 67006 40962
rect 67058 40910 67060 40962
rect 66892 40180 66948 40190
rect 66892 39508 66948 40124
rect 67004 39732 67060 40910
rect 67116 40964 67172 40974
rect 67116 40514 67172 40908
rect 67116 40462 67118 40514
rect 67170 40462 67172 40514
rect 67116 40450 67172 40462
rect 67228 40180 67284 41356
rect 67676 40962 67732 40974
rect 67676 40910 67678 40962
rect 67730 40910 67732 40962
rect 67452 40516 67508 40526
rect 67452 40422 67508 40460
rect 67116 40124 67284 40180
rect 67676 40180 67732 40910
rect 67116 39844 67172 40124
rect 67676 40114 67732 40124
rect 67268 40012 67948 40022
rect 67324 39956 67372 40012
rect 67428 40010 67476 40012
rect 67532 40010 67580 40012
rect 67448 39958 67476 40010
rect 67572 39958 67580 40010
rect 67428 39956 67476 39958
rect 67532 39956 67580 39958
rect 67636 40010 67684 40012
rect 67740 40010 67788 40012
rect 67636 39958 67644 40010
rect 67740 39958 67768 40010
rect 67636 39956 67684 39958
rect 67740 39956 67788 39958
rect 67844 39956 67892 40012
rect 67268 39946 67948 39956
rect 68012 39844 68068 42700
rect 69804 42754 69972 42756
rect 69804 42702 69806 42754
rect 69858 42702 69972 42754
rect 69804 42700 69972 42702
rect 70252 43650 70420 43652
rect 70252 43598 70366 43650
rect 70418 43598 70420 43650
rect 70252 43596 70420 43598
rect 70252 42754 70308 43596
rect 70364 43586 70420 43596
rect 70700 43540 70756 43550
rect 70700 43446 70756 43484
rect 71260 43428 71316 43710
rect 71708 43652 71764 43662
rect 71708 43558 71764 43596
rect 72492 43652 72548 43662
rect 73164 43652 73220 44044
rect 73276 44034 73332 44044
rect 73836 43988 73892 44270
rect 74508 44322 74564 44940
rect 74508 44270 74510 44322
rect 74562 44270 74564 44322
rect 74060 44210 74116 44222
rect 74060 44158 74062 44210
rect 74114 44158 74116 44210
rect 73948 43988 74004 43998
rect 73836 43932 73948 43988
rect 73948 43922 74004 43932
rect 74060 43708 74116 44158
rect 73500 43652 74116 43708
rect 72548 43596 72660 43652
rect 72492 43586 72548 43596
rect 72380 43540 72436 43550
rect 72380 43446 72436 43484
rect 71260 43362 71316 43372
rect 70252 42702 70254 42754
rect 70306 42702 70308 42754
rect 69804 42690 69860 42700
rect 70252 42690 70308 42702
rect 69356 42532 69412 42542
rect 69356 42438 69412 42476
rect 72492 42532 72548 42570
rect 72492 42466 72548 42476
rect 71768 42364 72448 42374
rect 71824 42308 71872 42364
rect 71928 42362 71976 42364
rect 72032 42362 72080 42364
rect 71948 42310 71976 42362
rect 72072 42310 72080 42362
rect 71928 42308 71976 42310
rect 72032 42308 72080 42310
rect 72136 42362 72184 42364
rect 72240 42362 72288 42364
rect 72136 42310 72144 42362
rect 72240 42310 72268 42362
rect 72136 42308 72184 42310
rect 72240 42308 72288 42310
rect 72344 42308 72392 42364
rect 71768 42298 72448 42308
rect 72268 41860 72324 41870
rect 72268 41300 72324 41804
rect 72268 41234 72324 41244
rect 71036 41188 71092 41198
rect 70812 41186 71092 41188
rect 70812 41134 71038 41186
rect 71090 41134 71092 41186
rect 70812 41132 71092 41134
rect 70812 41074 70868 41132
rect 71036 41122 71092 41132
rect 71596 41186 71652 41198
rect 71596 41134 71598 41186
rect 71650 41134 71652 41186
rect 70812 41022 70814 41074
rect 70866 41022 70868 41074
rect 70812 41010 70868 41022
rect 71372 41076 71428 41086
rect 68572 40962 68628 40974
rect 68572 40910 68574 40962
rect 68626 40910 68628 40962
rect 68124 40628 68180 40638
rect 68572 40628 68628 40910
rect 68180 40572 68628 40628
rect 68124 40514 68180 40572
rect 68124 40462 68126 40514
rect 68178 40462 68180 40514
rect 68124 40450 68180 40462
rect 67116 39788 67284 39844
rect 67004 39676 67172 39732
rect 66892 39442 66948 39452
rect 65548 37266 65604 39004
rect 66668 38966 66724 39004
rect 67116 39058 67172 39676
rect 67116 39006 67118 39058
rect 67170 39006 67172 39058
rect 67004 38948 67060 38958
rect 65548 37214 65550 37266
rect 65602 37214 65604 37266
rect 65548 36596 65604 37214
rect 66108 38388 66164 38398
rect 66108 37716 66164 38332
rect 66444 37828 66500 37838
rect 66444 37734 66500 37772
rect 67004 37826 67060 38892
rect 67004 37774 67006 37826
rect 67058 37774 67060 37826
rect 66108 37266 66164 37660
rect 66332 37380 66388 37390
rect 67004 37380 67060 37774
rect 67116 37828 67172 39006
rect 67228 39730 67284 39788
rect 67228 39678 67230 39730
rect 67282 39678 67284 39730
rect 67228 38836 67284 39678
rect 67228 38770 67284 38780
rect 67676 39788 68068 39844
rect 68236 40402 68292 40414
rect 68908 40404 68964 40414
rect 69356 40404 69412 40414
rect 68236 40350 68238 40402
rect 68290 40350 68292 40402
rect 67676 39730 67732 39788
rect 67676 39678 67678 39730
rect 67730 39678 67732 39730
rect 67676 38668 67732 39678
rect 68236 39508 68292 40350
rect 68684 40402 68964 40404
rect 68684 40350 68910 40402
rect 68962 40350 68964 40402
rect 68684 40348 68964 40350
rect 68348 39844 68404 39854
rect 68348 39618 68404 39788
rect 68348 39566 68350 39618
rect 68402 39566 68404 39618
rect 68348 39554 68404 39566
rect 68684 39618 68740 40348
rect 68908 40338 68964 40348
rect 69020 40402 69412 40404
rect 69020 40350 69358 40402
rect 69410 40350 69412 40402
rect 69020 40348 69412 40350
rect 71372 40404 71428 41020
rect 71596 40628 71652 41134
rect 71768 40796 72448 40806
rect 71824 40740 71872 40796
rect 71928 40794 71976 40796
rect 72032 40794 72080 40796
rect 71948 40742 71976 40794
rect 72072 40742 72080 40794
rect 71928 40740 71976 40742
rect 72032 40740 72080 40742
rect 72136 40794 72184 40796
rect 72240 40794 72288 40796
rect 72136 40742 72144 40794
rect 72240 40742 72268 40794
rect 72136 40740 72184 40742
rect 72240 40740 72288 40742
rect 72344 40740 72392 40796
rect 71768 40730 72448 40740
rect 71596 40562 71652 40572
rect 72268 40628 72324 40638
rect 72604 40628 72660 43596
rect 73164 43538 73220 43596
rect 73164 43486 73166 43538
rect 73218 43486 73220 43538
rect 73164 43474 73220 43486
rect 73276 43650 73556 43652
rect 73276 43598 73502 43650
rect 73554 43598 73556 43650
rect 73276 43596 73556 43598
rect 72716 43428 72772 43438
rect 72716 43334 72772 43372
rect 73276 42978 73332 43596
rect 73500 43586 73556 43596
rect 73276 42926 73278 42978
rect 73330 42926 73332 42978
rect 73276 42914 73332 42926
rect 74508 42532 74564 44270
rect 74508 42466 74564 42476
rect 74620 44324 74676 44334
rect 74620 42196 74676 44268
rect 75068 44324 75124 44334
rect 75068 44230 75124 44268
rect 74956 43988 75012 43998
rect 74956 43426 75012 43932
rect 74956 43374 74958 43426
rect 75010 43374 75012 43426
rect 74956 43314 75012 43374
rect 74956 43262 74958 43314
rect 75010 43262 75012 43314
rect 74956 43250 75012 43262
rect 72268 40534 72324 40572
rect 72492 40572 72660 40628
rect 73500 41860 73556 41870
rect 71708 40404 71764 40414
rect 71372 40348 71708 40404
rect 69020 40180 69076 40348
rect 69356 40338 69412 40348
rect 71708 40310 71764 40348
rect 68684 39566 68686 39618
rect 68738 39566 68740 39618
rect 68684 39554 68740 39566
rect 68796 40124 69076 40180
rect 69692 40180 69748 40190
rect 67900 39452 68292 39508
rect 68460 39508 68516 39518
rect 67788 39060 67844 39070
rect 67788 38834 67844 39004
rect 67900 39058 67956 39452
rect 68460 39414 68516 39452
rect 67900 39006 67902 39058
rect 67954 39006 67956 39058
rect 67900 38994 67956 39006
rect 68012 38948 68068 38958
rect 68012 38854 68068 38892
rect 68348 38836 68404 38846
rect 67788 38782 67790 38834
rect 67842 38782 67844 38834
rect 67788 38770 67844 38782
rect 68124 38834 68404 38836
rect 68124 38782 68350 38834
rect 68402 38782 68404 38834
rect 68124 38780 68404 38782
rect 68124 38724 68180 38780
rect 68348 38770 68404 38780
rect 67900 38668 68180 38724
rect 67676 38612 67956 38668
rect 67268 38444 67948 38454
rect 67324 38388 67372 38444
rect 67428 38442 67476 38444
rect 67532 38442 67580 38444
rect 67448 38390 67476 38442
rect 67572 38390 67580 38442
rect 67428 38388 67476 38390
rect 67532 38388 67580 38390
rect 67636 38442 67684 38444
rect 67740 38442 67788 38444
rect 67636 38390 67644 38442
rect 67740 38390 67768 38442
rect 67636 38388 67684 38390
rect 67740 38388 67788 38390
rect 67844 38388 67892 38444
rect 67268 38378 67948 38388
rect 67788 38276 67844 38286
rect 67676 38162 67732 38174
rect 67676 38110 67678 38162
rect 67730 38110 67732 38162
rect 67116 37762 67172 37772
rect 67228 38052 67284 38062
rect 67228 37826 67284 37996
rect 67228 37774 67230 37826
rect 67282 37774 67284 37826
rect 66332 37378 67060 37380
rect 66332 37326 66334 37378
rect 66386 37326 67060 37378
rect 66332 37324 67060 37326
rect 66332 37314 66388 37324
rect 66108 37214 66110 37266
rect 66162 37214 66164 37266
rect 66108 37202 66164 37214
rect 66892 37154 66948 37166
rect 66892 37102 66894 37154
rect 66946 37102 66948 37154
rect 66892 37044 66948 37102
rect 66892 36978 66948 36988
rect 67228 37044 67284 37774
rect 67676 37828 67732 38110
rect 67676 37762 67732 37772
rect 67788 37490 67844 38220
rect 68572 38276 68628 38286
rect 68572 38052 68628 38220
rect 68796 38162 68852 40124
rect 69692 40086 69748 40124
rect 69020 39844 69076 39854
rect 69020 39730 69076 39788
rect 69020 39678 69022 39730
rect 69074 39678 69076 39730
rect 69020 39666 69076 39678
rect 72492 39396 72548 40572
rect 72604 40404 72660 40414
rect 73164 40404 73220 40414
rect 72604 40402 73220 40404
rect 72604 40350 72606 40402
rect 72658 40350 73166 40402
rect 73218 40350 73220 40402
rect 72604 40348 73220 40350
rect 72604 40338 72660 40348
rect 73164 40338 73220 40348
rect 73500 40290 73556 41804
rect 74172 41076 74228 41086
rect 74060 40962 74116 40974
rect 74060 40910 74062 40962
rect 74114 40910 74116 40962
rect 73948 40404 74004 40414
rect 73948 40310 74004 40348
rect 73500 40238 73502 40290
rect 73554 40238 73556 40290
rect 72492 39340 72660 39396
rect 71768 39228 72448 39238
rect 71824 39172 71872 39228
rect 71928 39226 71976 39228
rect 72032 39226 72080 39228
rect 71948 39174 71976 39226
rect 72072 39174 72080 39226
rect 71928 39172 71976 39174
rect 72032 39172 72080 39174
rect 72136 39226 72184 39228
rect 72240 39226 72288 39228
rect 72136 39174 72144 39226
rect 72240 39174 72268 39226
rect 72136 39172 72184 39174
rect 72240 39172 72288 39174
rect 72344 39172 72392 39228
rect 71768 39162 72448 39172
rect 72492 39060 72548 39070
rect 72604 39060 72660 39340
rect 72492 39058 72660 39060
rect 72492 39006 72494 39058
rect 72546 39006 72660 39058
rect 72492 39004 72660 39006
rect 72716 39394 72772 39406
rect 72716 39342 72718 39394
rect 72770 39342 72772 39394
rect 72716 39060 72772 39342
rect 72940 39060 72996 39070
rect 73500 39060 73556 40238
rect 74060 40292 74116 40910
rect 74172 40514 74228 41020
rect 74620 40852 74676 42140
rect 75068 41188 75124 41198
rect 75180 41188 75236 47180
rect 75292 46786 75348 47628
rect 75292 46734 75294 46786
rect 75346 46734 75348 46786
rect 75292 46722 75348 46734
rect 75852 45892 75908 45902
rect 75404 44324 75460 44334
rect 75404 43764 75460 44268
rect 75404 43762 75572 43764
rect 75404 43710 75406 43762
rect 75458 43710 75572 43762
rect 75404 43708 75572 43710
rect 75404 43698 75460 43708
rect 75516 43540 75572 43708
rect 75740 43540 75796 43550
rect 75516 43538 75796 43540
rect 75516 43486 75742 43538
rect 75794 43486 75796 43538
rect 75516 43484 75796 43486
rect 75740 43474 75796 43484
rect 75068 41186 75236 41188
rect 75068 41134 75070 41186
rect 75122 41134 75236 41186
rect 75068 41132 75236 41134
rect 75292 43316 75348 43326
rect 74732 41076 74788 41086
rect 74732 40982 74788 41020
rect 74620 40796 75012 40852
rect 74172 40462 74174 40514
rect 74226 40462 74228 40514
rect 74172 40450 74228 40462
rect 74172 40292 74228 40302
rect 74060 40236 74172 40292
rect 74172 40226 74228 40236
rect 72716 39058 73556 39060
rect 72716 39006 72942 39058
rect 72994 39006 73556 39058
rect 72716 39004 73556 39006
rect 69020 38836 69076 38846
rect 69020 38742 69076 38780
rect 72492 38668 72548 39004
rect 72940 38994 72996 39004
rect 68796 38110 68798 38162
rect 68850 38110 68852 38162
rect 68796 38098 68852 38110
rect 72380 38612 72548 38668
rect 68572 37958 68628 37996
rect 68348 37940 68404 37950
rect 68348 37846 68404 37884
rect 72380 37940 72436 38612
rect 72492 38052 72548 38062
rect 73164 38052 73220 38062
rect 72492 38050 73220 38052
rect 72492 37998 72494 38050
rect 72546 37998 73166 38050
rect 73218 37998 73220 38050
rect 72492 37996 73220 37998
rect 72492 37986 72548 37996
rect 73164 37986 73220 37996
rect 73500 38050 73556 39004
rect 74844 38836 74900 38846
rect 73500 37998 73502 38050
rect 73554 37998 73556 38050
rect 72380 37874 72436 37884
rect 68796 37826 68852 37838
rect 68796 37774 68798 37826
rect 68850 37774 68852 37826
rect 67788 37438 67790 37490
rect 67842 37438 67844 37490
rect 67788 37426 67844 37438
rect 68236 37604 68292 37614
rect 68236 37490 68292 37548
rect 68236 37438 68238 37490
rect 68290 37438 68292 37490
rect 68236 37426 68292 37438
rect 67228 36978 67284 36988
rect 68684 37044 68740 37054
rect 67268 36876 67948 36886
rect 67324 36820 67372 36876
rect 67428 36874 67476 36876
rect 67532 36874 67580 36876
rect 67448 36822 67476 36874
rect 67572 36822 67580 36874
rect 67428 36820 67476 36822
rect 67532 36820 67580 36822
rect 67636 36874 67684 36876
rect 67740 36874 67788 36876
rect 67636 36822 67644 36874
rect 67740 36822 67768 36874
rect 67636 36820 67684 36822
rect 67740 36820 67788 36822
rect 67844 36820 67892 36876
rect 67268 36810 67948 36820
rect 65548 36530 65604 36540
rect 67452 36596 67508 36606
rect 67452 36502 67508 36540
rect 65436 36306 65492 36316
rect 67788 36372 67844 36382
rect 68684 36372 68740 36988
rect 68796 36820 68852 37774
rect 68908 37826 68964 37838
rect 68908 37774 68910 37826
rect 68962 37774 68964 37826
rect 68908 37604 68964 37774
rect 71932 37828 71988 37866
rect 71932 37762 71988 37772
rect 72604 37828 72660 37838
rect 71768 37660 72448 37670
rect 71824 37604 71872 37660
rect 71928 37658 71976 37660
rect 72032 37658 72080 37660
rect 71948 37606 71976 37658
rect 72072 37606 72080 37658
rect 71928 37604 71976 37606
rect 72032 37604 72080 37606
rect 72136 37658 72184 37660
rect 72240 37658 72288 37660
rect 72136 37606 72144 37658
rect 72240 37606 72268 37658
rect 72136 37604 72184 37606
rect 72240 37604 72288 37606
rect 72344 37604 72392 37660
rect 71768 37594 72448 37604
rect 68908 37538 68964 37548
rect 72380 37268 72436 37278
rect 72604 37268 72660 37772
rect 72380 37266 72660 37268
rect 72380 37214 72382 37266
rect 72434 37214 72660 37266
rect 72380 37212 72660 37214
rect 72716 37826 72772 37838
rect 72716 37774 72718 37826
rect 72770 37774 72772 37826
rect 72716 37266 72772 37774
rect 72716 37214 72718 37266
rect 72770 37214 72772 37266
rect 72380 37202 72436 37212
rect 72716 37202 72772 37214
rect 68796 36754 68852 36764
rect 69468 36932 69524 36942
rect 68796 36596 68852 36606
rect 68796 36502 68852 36540
rect 69468 36482 69524 36876
rect 69468 36430 69470 36482
rect 69522 36430 69524 36482
rect 69468 36372 69524 36430
rect 67844 36316 68068 36372
rect 68684 36316 68852 36372
rect 67788 36278 67844 36316
rect 67268 35308 67948 35318
rect 67324 35252 67372 35308
rect 67428 35306 67476 35308
rect 67532 35306 67580 35308
rect 67448 35254 67476 35306
rect 67572 35254 67580 35306
rect 67428 35252 67476 35254
rect 67532 35252 67580 35254
rect 67636 35306 67684 35308
rect 67740 35306 67788 35308
rect 67636 35254 67644 35306
rect 67740 35254 67768 35306
rect 67636 35252 67684 35254
rect 67740 35252 67788 35254
rect 67844 35252 67892 35308
rect 67268 35242 67948 35252
rect 65436 34804 65492 34814
rect 65324 34802 65492 34804
rect 65324 34750 65438 34802
rect 65490 34750 65492 34802
rect 65324 34748 65492 34750
rect 64652 34354 64708 34748
rect 64652 34302 64654 34354
rect 64706 34302 64708 34354
rect 64652 34290 64708 34302
rect 65436 34356 65492 34748
rect 67004 34692 67060 34702
rect 65436 34300 65604 34356
rect 64652 34130 64708 34142
rect 64876 34132 64932 34142
rect 65436 34132 65492 34142
rect 64652 34078 64654 34130
rect 64706 34078 64708 34130
rect 64652 33684 64708 34078
rect 64652 33618 64708 33628
rect 64764 34130 65492 34132
rect 64764 34078 64878 34130
rect 64930 34078 65438 34130
rect 65490 34078 65492 34130
rect 64764 34076 65492 34078
rect 64540 32498 64596 32508
rect 63084 32450 63700 32452
rect 63084 32398 63086 32450
rect 63138 32398 63700 32450
rect 63084 32396 63700 32398
rect 63084 32386 63140 32396
rect 62524 31938 62580 31948
rect 64092 32004 64148 32014
rect 64092 31910 64148 31948
rect 63532 31892 63588 31902
rect 63532 31554 63588 31836
rect 64428 31892 64484 31902
rect 64428 31798 64484 31836
rect 63532 31502 63534 31554
rect 63586 31502 63588 31554
rect 63532 31490 63588 31502
rect 64652 31556 64708 31566
rect 62768 31388 63448 31398
rect 62824 31332 62872 31388
rect 62928 31386 62976 31388
rect 63032 31386 63080 31388
rect 62948 31334 62976 31386
rect 63072 31334 63080 31386
rect 62928 31332 62976 31334
rect 63032 31332 63080 31334
rect 63136 31386 63184 31388
rect 63240 31386 63288 31388
rect 63136 31334 63144 31386
rect 63240 31334 63268 31386
rect 63136 31332 63184 31334
rect 63240 31332 63288 31334
rect 63344 31332 63392 31388
rect 62768 31322 63448 31332
rect 61628 29876 61684 29932
rect 58268 28970 58948 28980
rect 59052 28924 59220 28980
rect 61516 29820 61684 29876
rect 62768 29820 63448 29830
rect 58940 28868 58996 28878
rect 59052 28868 59108 28924
rect 58940 28866 59108 28868
rect 58940 28814 58942 28866
rect 58994 28814 59108 28866
rect 58940 28812 59108 28814
rect 60732 28868 60788 28878
rect 58940 28802 58996 28812
rect 60732 28754 60788 28812
rect 61180 28868 61236 28878
rect 61180 28866 61348 28868
rect 61180 28814 61182 28866
rect 61234 28814 61348 28866
rect 61180 28812 61348 28814
rect 61180 28802 61236 28812
rect 60732 28702 60734 28754
rect 60786 28702 60788 28754
rect 60732 28644 60788 28702
rect 60732 28578 60788 28588
rect 61292 28644 61348 28812
rect 61292 28578 61348 28588
rect 61068 28530 61124 28542
rect 61068 28478 61070 28530
rect 61122 28478 61124 28530
rect 58156 28420 58212 28430
rect 58044 28418 58212 28420
rect 58044 28366 58158 28418
rect 58210 28366 58212 28418
rect 58044 28364 58212 28366
rect 57148 27806 57150 27858
rect 57202 27806 57204 27858
rect 57148 27794 57204 27806
rect 57260 27972 57316 27982
rect 56924 27246 56926 27298
rect 56978 27246 56980 27298
rect 56924 27076 56980 27246
rect 57260 27300 57316 27916
rect 57932 27748 57988 27758
rect 57260 27298 57652 27300
rect 57260 27246 57262 27298
rect 57314 27246 57652 27298
rect 57260 27244 57652 27246
rect 57260 27234 57316 27244
rect 56924 27010 56980 27020
rect 57036 26852 57092 26862
rect 57036 26758 57092 26796
rect 56028 26674 56084 26684
rect 57596 26514 57652 27244
rect 57932 27298 57988 27692
rect 57932 27246 57934 27298
rect 57986 27246 57988 27298
rect 57932 27234 57988 27246
rect 57820 27076 57876 27086
rect 57820 26982 57876 27020
rect 57932 26962 57988 26974
rect 57932 26910 57934 26962
rect 57986 26910 57988 26962
rect 57932 26516 57988 26910
rect 57596 26462 57598 26514
rect 57650 26462 57652 26514
rect 57596 26450 57652 26462
rect 57708 26460 57988 26516
rect 58044 26740 58100 28364
rect 58156 28354 58212 28364
rect 61068 28420 61124 28478
rect 61180 28532 61236 28542
rect 61516 28532 61572 29820
rect 62824 29764 62872 29820
rect 62928 29818 62976 29820
rect 63032 29818 63080 29820
rect 62948 29766 62976 29818
rect 63072 29766 63080 29818
rect 62928 29764 62976 29766
rect 63032 29764 63080 29766
rect 63136 29818 63184 29820
rect 63240 29818 63288 29820
rect 63136 29766 63144 29818
rect 63240 29766 63268 29818
rect 63136 29764 63184 29766
rect 63240 29764 63288 29766
rect 63344 29764 63392 29820
rect 62768 29754 63448 29764
rect 61628 29652 61684 29662
rect 61628 28644 61684 29596
rect 64652 29540 64708 31500
rect 64652 29474 64708 29484
rect 61740 28868 61796 28878
rect 61740 28774 61796 28812
rect 62300 28644 62356 28654
rect 61628 28642 62356 28644
rect 61628 28590 62302 28642
rect 62354 28590 62356 28642
rect 61628 28588 62356 28590
rect 61180 28438 61236 28476
rect 61404 28476 61572 28532
rect 61740 28530 61796 28588
rect 62300 28578 62356 28588
rect 62972 28644 63028 28654
rect 59612 28082 59668 28094
rect 59612 28030 59614 28082
rect 59666 28030 59668 28082
rect 58268 27468 58948 27478
rect 58324 27412 58372 27468
rect 58428 27466 58476 27468
rect 58532 27466 58580 27468
rect 58448 27414 58476 27466
rect 58572 27414 58580 27466
rect 58428 27412 58476 27414
rect 58532 27412 58580 27414
rect 58636 27466 58684 27468
rect 58740 27466 58788 27468
rect 58636 27414 58644 27466
rect 58740 27414 58768 27466
rect 58636 27412 58684 27414
rect 58740 27412 58788 27414
rect 58844 27412 58892 27468
rect 58268 27402 58948 27412
rect 57036 26292 57092 26302
rect 54796 26126 54798 26178
rect 54850 26126 54852 26178
rect 54796 26114 54852 26126
rect 56700 26236 57036 26292
rect 54236 25454 54238 25506
rect 54290 25454 54292 25506
rect 54236 25442 54292 25454
rect 54572 25508 54628 25518
rect 54572 25414 54628 25452
rect 53768 25116 54448 25126
rect 53824 25060 53872 25116
rect 53928 25114 53976 25116
rect 54032 25114 54080 25116
rect 53948 25062 53976 25114
rect 54072 25062 54080 25114
rect 53928 25060 53976 25062
rect 54032 25060 54080 25062
rect 54136 25114 54184 25116
rect 54240 25114 54288 25116
rect 54136 25062 54144 25114
rect 54240 25062 54268 25114
rect 54136 25060 54184 25062
rect 54240 25060 54288 25062
rect 54344 25060 54392 25116
rect 53768 25050 54448 25060
rect 53768 23548 54448 23558
rect 53824 23492 53872 23548
rect 53928 23546 53976 23548
rect 54032 23546 54080 23548
rect 53948 23494 53976 23546
rect 54072 23494 54080 23546
rect 53928 23492 53976 23494
rect 54032 23492 54080 23494
rect 54136 23546 54184 23548
rect 54240 23546 54288 23548
rect 54136 23494 54144 23546
rect 54240 23494 54268 23546
rect 54136 23492 54184 23494
rect 54240 23492 54288 23494
rect 54344 23492 54392 23548
rect 53768 23482 54448 23492
rect 53768 21980 54448 21990
rect 53824 21924 53872 21980
rect 53928 21978 53976 21980
rect 54032 21978 54080 21980
rect 53948 21926 53976 21978
rect 54072 21926 54080 21978
rect 53928 21924 53976 21926
rect 54032 21924 54080 21926
rect 54136 21978 54184 21980
rect 54240 21978 54288 21980
rect 54136 21926 54144 21978
rect 54240 21926 54268 21978
rect 54136 21924 54184 21926
rect 54240 21924 54288 21926
rect 54344 21924 54392 21980
rect 53768 21914 54448 21924
rect 56028 21028 56084 21038
rect 55468 20916 55524 20926
rect 55468 20822 55524 20860
rect 56028 20804 56084 20972
rect 56700 21028 56756 26236
rect 57036 26198 57092 26236
rect 57708 25730 57764 26460
rect 57932 26292 57988 26302
rect 57932 26198 57988 26236
rect 57708 25678 57710 25730
rect 57762 25678 57764 25730
rect 57708 25666 57764 25678
rect 57148 25620 57204 25630
rect 57148 25282 57204 25564
rect 58044 25620 58100 26684
rect 59612 26740 59668 28030
rect 60172 27972 60228 27982
rect 60172 27878 60228 27916
rect 59948 27300 60004 27310
rect 59948 27186 60004 27244
rect 59948 27134 59950 27186
rect 60002 27134 60004 27186
rect 59948 27122 60004 27134
rect 60620 27300 60676 27310
rect 60508 26964 60564 26974
rect 59612 26674 59668 26684
rect 59948 26852 60004 26862
rect 59612 26516 59668 26526
rect 59612 26422 59668 26460
rect 58492 26404 58548 26414
rect 58492 26310 58548 26348
rect 59948 26404 60004 26796
rect 60060 26516 60116 26526
rect 60060 26422 60116 26460
rect 59948 26310 60004 26348
rect 60060 26068 60116 26078
rect 60060 25974 60116 26012
rect 58268 25900 58948 25910
rect 58324 25844 58372 25900
rect 58428 25898 58476 25900
rect 58532 25898 58580 25900
rect 58448 25846 58476 25898
rect 58572 25846 58580 25898
rect 58428 25844 58476 25846
rect 58532 25844 58580 25846
rect 58636 25898 58684 25900
rect 58740 25898 58788 25900
rect 58636 25846 58644 25898
rect 58740 25846 58768 25898
rect 58636 25844 58684 25846
rect 58740 25844 58788 25846
rect 58844 25844 58892 25900
rect 58268 25834 58948 25844
rect 58044 25526 58100 25564
rect 57148 25230 57150 25282
rect 57202 25230 57204 25282
rect 57148 25218 57204 25230
rect 60172 24948 60228 24958
rect 60172 24854 60228 24892
rect 60508 24834 60564 26908
rect 60620 26962 60676 27244
rect 60844 27076 60900 27086
rect 60844 26982 60900 27020
rect 61068 27074 61124 28364
rect 61404 28196 61460 28476
rect 61292 28140 61460 28196
rect 61628 28474 61684 28486
rect 61628 28422 61630 28474
rect 61682 28422 61684 28474
rect 61740 28478 61742 28530
rect 61794 28478 61796 28530
rect 61740 28466 61796 28478
rect 62972 28530 63028 28588
rect 63196 28644 63252 28654
rect 63196 28550 63252 28588
rect 63532 28644 63588 28654
rect 62972 28478 62974 28530
rect 63026 28478 63028 28530
rect 62972 28466 63028 28478
rect 61628 28420 61684 28422
rect 61068 27022 61070 27074
rect 61122 27022 61124 27074
rect 60620 26910 60622 26962
rect 60674 26910 60676 26962
rect 60620 26898 60676 26910
rect 61068 26852 61124 27022
rect 61068 26786 61124 26796
rect 61180 28084 61236 28094
rect 61180 26962 61236 28028
rect 61180 26910 61182 26962
rect 61234 26910 61236 26962
rect 60844 26516 60900 26526
rect 61180 26516 61236 26910
rect 60844 26514 61236 26516
rect 60844 26462 60846 26514
rect 60898 26462 61236 26514
rect 60844 26460 61236 26462
rect 60844 26450 60900 26460
rect 60620 24948 60676 24958
rect 60620 24854 60676 24892
rect 60508 24782 60510 24834
rect 60562 24782 60564 24834
rect 59388 24724 59444 24734
rect 58268 24332 58948 24342
rect 58324 24276 58372 24332
rect 58428 24330 58476 24332
rect 58532 24330 58580 24332
rect 58448 24278 58476 24330
rect 58572 24278 58580 24330
rect 58428 24276 58476 24278
rect 58532 24276 58580 24278
rect 58636 24330 58684 24332
rect 58740 24330 58788 24332
rect 58636 24278 58644 24330
rect 58740 24278 58768 24330
rect 58636 24276 58684 24278
rect 58740 24276 58788 24278
rect 58844 24276 58892 24332
rect 58268 24266 58948 24276
rect 59388 24052 59444 24668
rect 59388 24050 59892 24052
rect 59388 23998 59390 24050
rect 59442 23998 59892 24050
rect 59388 23996 59892 23998
rect 59388 23986 59444 23996
rect 59724 23828 59780 23838
rect 59724 23734 59780 23772
rect 59836 23826 59892 23996
rect 59836 23774 59838 23826
rect 59890 23774 59892 23826
rect 59836 23762 59892 23774
rect 60508 23938 60564 24782
rect 60620 24500 60676 24510
rect 60620 24406 60676 24444
rect 60508 23886 60510 23938
rect 60562 23886 60564 23938
rect 60508 23828 60564 23886
rect 61180 24052 61236 24062
rect 60508 23762 60564 23772
rect 61068 23828 61124 23838
rect 61068 23734 61124 23772
rect 61180 23826 61236 23996
rect 61180 23774 61182 23826
rect 61234 23774 61236 23826
rect 60060 23714 60116 23726
rect 60060 23662 60062 23714
rect 60114 23662 60116 23714
rect 58268 22764 58948 22774
rect 58324 22708 58372 22764
rect 58428 22762 58476 22764
rect 58532 22762 58580 22764
rect 58448 22710 58476 22762
rect 58572 22710 58580 22762
rect 58428 22708 58476 22710
rect 58532 22708 58580 22710
rect 58636 22762 58684 22764
rect 58740 22762 58788 22764
rect 58636 22710 58644 22762
rect 58740 22710 58768 22762
rect 58636 22708 58684 22710
rect 58740 22708 58788 22710
rect 58844 22708 58892 22764
rect 58268 22698 58948 22708
rect 60060 22372 60116 23662
rect 60284 23716 60340 23726
rect 60284 23604 60340 23660
rect 60620 23714 60676 23726
rect 60844 23716 60900 23726
rect 60620 23662 60622 23714
rect 60674 23662 60676 23714
rect 60620 23604 60676 23662
rect 60284 23548 60676 23604
rect 60732 23714 60900 23716
rect 60732 23662 60846 23714
rect 60898 23662 60900 23714
rect 60732 23660 60900 23662
rect 60284 23378 60340 23548
rect 60284 23326 60286 23378
rect 60338 23326 60340 23378
rect 60284 23314 60340 23326
rect 60732 23380 60788 23660
rect 60844 23650 60900 23660
rect 61180 23492 61236 23774
rect 60732 23314 60788 23324
rect 60844 23436 61236 23492
rect 60844 23378 60900 23436
rect 60844 23326 60846 23378
rect 60898 23326 60900 23378
rect 60844 23314 60900 23326
rect 60060 22306 60116 22316
rect 58268 21196 58948 21206
rect 58324 21140 58372 21196
rect 58428 21194 58476 21196
rect 58532 21194 58580 21196
rect 58448 21142 58476 21194
rect 58572 21142 58580 21194
rect 58428 21140 58476 21142
rect 58532 21140 58580 21142
rect 58636 21194 58684 21196
rect 58740 21194 58788 21196
rect 58636 21142 58644 21194
rect 58740 21142 58768 21194
rect 58636 21140 58684 21142
rect 58740 21140 58788 21142
rect 58844 21140 58892 21196
rect 58268 21130 58948 21140
rect 56028 20710 56084 20748
rect 56140 20916 56196 20926
rect 56140 20690 56196 20860
rect 56700 20914 56756 20972
rect 56700 20862 56702 20914
rect 56754 20862 56756 20914
rect 56700 20850 56756 20862
rect 56364 20804 56420 20814
rect 56364 20710 56420 20748
rect 56140 20638 56142 20690
rect 56194 20638 56196 20690
rect 56140 20626 56196 20638
rect 53768 20412 54448 20422
rect 53824 20356 53872 20412
rect 53928 20410 53976 20412
rect 54032 20410 54080 20412
rect 53948 20358 53976 20410
rect 54072 20358 54080 20410
rect 53928 20356 53976 20358
rect 54032 20356 54080 20358
rect 54136 20410 54184 20412
rect 54240 20410 54288 20412
rect 54136 20358 54144 20410
rect 54240 20358 54268 20410
rect 54136 20356 54184 20358
rect 54240 20356 54288 20358
rect 54344 20356 54392 20412
rect 53768 20346 54448 20356
rect 53116 20132 53396 20188
rect 53116 15148 53172 20132
rect 58268 19628 58948 19638
rect 58324 19572 58372 19628
rect 58428 19626 58476 19628
rect 58532 19626 58580 19628
rect 58448 19574 58476 19626
rect 58572 19574 58580 19626
rect 58428 19572 58476 19574
rect 58532 19572 58580 19574
rect 58636 19626 58684 19628
rect 58740 19626 58788 19628
rect 58636 19574 58644 19626
rect 58740 19574 58768 19626
rect 58636 19572 58684 19574
rect 58740 19572 58788 19574
rect 58844 19572 58892 19628
rect 58268 19562 58948 19572
rect 53768 18844 54448 18854
rect 53824 18788 53872 18844
rect 53928 18842 53976 18844
rect 54032 18842 54080 18844
rect 53948 18790 53976 18842
rect 54072 18790 54080 18842
rect 53928 18788 53976 18790
rect 54032 18788 54080 18790
rect 54136 18842 54184 18844
rect 54240 18842 54288 18844
rect 54136 18790 54144 18842
rect 54240 18790 54268 18842
rect 54136 18788 54184 18790
rect 54240 18788 54288 18790
rect 54344 18788 54392 18844
rect 53768 18778 54448 18788
rect 58268 18060 58948 18070
rect 58324 18004 58372 18060
rect 58428 18058 58476 18060
rect 58532 18058 58580 18060
rect 58448 18006 58476 18058
rect 58572 18006 58580 18058
rect 58428 18004 58476 18006
rect 58532 18004 58580 18006
rect 58636 18058 58684 18060
rect 58740 18058 58788 18060
rect 58636 18006 58644 18058
rect 58740 18006 58768 18058
rect 58636 18004 58684 18006
rect 58740 18004 58788 18006
rect 58844 18004 58892 18060
rect 58268 17994 58948 18004
rect 53768 17276 54448 17286
rect 53824 17220 53872 17276
rect 53928 17274 53976 17276
rect 54032 17274 54080 17276
rect 53948 17222 53976 17274
rect 54072 17222 54080 17274
rect 53928 17220 53976 17222
rect 54032 17220 54080 17222
rect 54136 17274 54184 17276
rect 54240 17274 54288 17276
rect 54136 17222 54144 17274
rect 54240 17222 54268 17274
rect 54136 17220 54184 17222
rect 54240 17220 54288 17222
rect 54344 17220 54392 17276
rect 53768 17210 54448 17220
rect 58268 16492 58948 16502
rect 58324 16436 58372 16492
rect 58428 16490 58476 16492
rect 58532 16490 58580 16492
rect 58448 16438 58476 16490
rect 58572 16438 58580 16490
rect 58428 16436 58476 16438
rect 58532 16436 58580 16438
rect 58636 16490 58684 16492
rect 58740 16490 58788 16492
rect 58636 16438 58644 16490
rect 58740 16438 58768 16490
rect 58636 16436 58684 16438
rect 58740 16436 58788 16438
rect 58844 16436 58892 16492
rect 58268 16426 58948 16436
rect 53768 15708 54448 15718
rect 53824 15652 53872 15708
rect 53928 15706 53976 15708
rect 54032 15706 54080 15708
rect 53948 15654 53976 15706
rect 54072 15654 54080 15706
rect 53928 15652 53976 15654
rect 54032 15652 54080 15654
rect 54136 15706 54184 15708
rect 54240 15706 54288 15708
rect 54136 15654 54144 15706
rect 54240 15654 54268 15706
rect 54136 15652 54184 15654
rect 54240 15652 54288 15654
rect 54344 15652 54392 15708
rect 53768 15642 54448 15652
rect 52444 13794 52500 13804
rect 53004 15092 53172 15148
rect 53004 13972 53060 15092
rect 58268 14924 58948 14934
rect 58324 14868 58372 14924
rect 58428 14922 58476 14924
rect 58532 14922 58580 14924
rect 58448 14870 58476 14922
rect 58572 14870 58580 14922
rect 58428 14868 58476 14870
rect 58532 14868 58580 14870
rect 58636 14922 58684 14924
rect 58740 14922 58788 14924
rect 58636 14870 58644 14922
rect 58740 14870 58768 14922
rect 58636 14868 58684 14870
rect 58740 14868 58788 14870
rect 58844 14868 58892 14924
rect 58268 14858 58948 14868
rect 53768 14140 54448 14150
rect 53824 14084 53872 14140
rect 53928 14138 53976 14140
rect 54032 14138 54080 14140
rect 53948 14086 53976 14138
rect 54072 14086 54080 14138
rect 53928 14084 53976 14086
rect 54032 14084 54080 14086
rect 54136 14138 54184 14140
rect 54240 14138 54288 14140
rect 54136 14086 54144 14138
rect 54240 14086 54268 14138
rect 54136 14084 54184 14086
rect 54240 14084 54288 14086
rect 54344 14084 54392 14140
rect 53768 14074 54448 14084
rect 51660 13694 51662 13746
rect 51714 13694 51716 13746
rect 51660 13682 51716 13694
rect 52108 13746 52164 13758
rect 52108 13694 52110 13746
rect 52162 13694 52164 13746
rect 51212 13634 51268 13646
rect 51212 13582 51214 13634
rect 51266 13582 51268 13634
rect 49268 13356 49948 13366
rect 49324 13300 49372 13356
rect 49428 13354 49476 13356
rect 49532 13354 49580 13356
rect 49448 13302 49476 13354
rect 49572 13302 49580 13354
rect 49428 13300 49476 13302
rect 49532 13300 49580 13302
rect 49636 13354 49684 13356
rect 49740 13354 49788 13356
rect 49636 13302 49644 13354
rect 49740 13302 49768 13354
rect 49636 13300 49684 13302
rect 49740 13300 49788 13302
rect 49844 13300 49892 13356
rect 49268 13290 49948 13300
rect 50092 12962 50148 12974
rect 50092 12910 50094 12962
rect 50146 12910 50148 12962
rect 49532 12852 49588 12862
rect 49532 12758 49588 12796
rect 49268 11788 49948 11798
rect 49324 11732 49372 11788
rect 49428 11786 49476 11788
rect 49532 11786 49580 11788
rect 49448 11734 49476 11786
rect 49572 11734 49580 11786
rect 49428 11732 49476 11734
rect 49532 11732 49580 11734
rect 49636 11786 49684 11788
rect 49740 11786 49788 11788
rect 49636 11734 49644 11786
rect 49740 11734 49768 11786
rect 49636 11732 49684 11734
rect 49740 11732 49788 11734
rect 49844 11732 49892 11788
rect 49268 11722 49948 11732
rect 49268 10220 49948 10230
rect 49324 10164 49372 10220
rect 49428 10218 49476 10220
rect 49532 10218 49580 10220
rect 49448 10166 49476 10218
rect 49572 10166 49580 10218
rect 49428 10164 49476 10166
rect 49532 10164 49580 10166
rect 49636 10218 49684 10220
rect 49740 10218 49788 10220
rect 49636 10166 49644 10218
rect 49740 10166 49768 10218
rect 49636 10164 49684 10166
rect 49740 10164 49788 10166
rect 49844 10164 49892 10220
rect 49268 10154 49948 10164
rect 50092 10052 50148 12910
rect 50428 12740 50484 12750
rect 50428 11956 50484 12684
rect 50876 12740 50932 12750
rect 50876 12646 50932 12684
rect 48860 9996 49028 10052
rect 49756 9996 50148 10052
rect 50316 11900 50484 11956
rect 51100 12178 51156 12190
rect 51100 12126 51102 12178
rect 51154 12126 51156 12178
rect 48860 9154 48916 9996
rect 48860 9102 48862 9154
rect 48914 9102 48916 9154
rect 48748 8818 48804 8830
rect 48748 8766 48750 8818
rect 48802 8766 48804 8818
rect 48748 8260 48804 8766
rect 48748 8194 48804 8204
rect 48076 7298 48132 7308
rect 48636 8146 48692 8158
rect 48636 8094 48638 8146
rect 48690 8094 48692 8146
rect 48636 6916 48692 8094
rect 48860 7812 48916 9102
rect 48972 9714 49028 9726
rect 48972 9662 48974 9714
rect 49026 9662 49028 9714
rect 48972 8036 49028 9662
rect 49196 9156 49252 9166
rect 49084 9154 49252 9156
rect 49084 9102 49198 9154
rect 49250 9102 49252 9154
rect 49084 9100 49252 9102
rect 49084 8484 49140 9100
rect 49196 9090 49252 9100
rect 49756 8930 49812 9996
rect 49756 8878 49758 8930
rect 49810 8878 49812 8930
rect 49756 8866 49812 8878
rect 50204 9042 50260 9054
rect 50204 8990 50206 9042
rect 50258 8990 50260 9042
rect 50092 8818 50148 8830
rect 50092 8766 50094 8818
rect 50146 8766 50148 8818
rect 49268 8652 49948 8662
rect 49324 8596 49372 8652
rect 49428 8650 49476 8652
rect 49532 8650 49580 8652
rect 49448 8598 49476 8650
rect 49572 8598 49580 8650
rect 49428 8596 49476 8598
rect 49532 8596 49580 8598
rect 49636 8650 49684 8652
rect 49740 8650 49788 8652
rect 49636 8598 49644 8650
rect 49740 8598 49768 8650
rect 49636 8596 49684 8598
rect 49740 8596 49788 8598
rect 49844 8596 49892 8652
rect 49268 8586 49948 8596
rect 49084 8428 49252 8484
rect 48972 7970 49028 7980
rect 48860 7756 49028 7812
rect 48972 7698 49028 7756
rect 48972 7646 48974 7698
rect 49026 7646 49028 7698
rect 48972 7634 49028 7646
rect 49196 7364 49252 8428
rect 49868 8372 49924 8382
rect 49868 7700 49924 8316
rect 49868 7606 49924 7644
rect 48636 6850 48692 6860
rect 48860 7308 49252 7364
rect 47852 6638 47854 6690
rect 47906 6638 47908 6690
rect 47852 6626 47908 6638
rect 48188 5908 48244 5918
rect 48188 5814 48244 5852
rect 48860 5460 48916 7308
rect 49268 7084 49948 7094
rect 49324 7028 49372 7084
rect 49428 7082 49476 7084
rect 49532 7082 49580 7084
rect 49448 7030 49476 7082
rect 49572 7030 49580 7082
rect 49428 7028 49476 7030
rect 49532 7028 49580 7030
rect 49636 7082 49684 7084
rect 49740 7082 49788 7084
rect 49636 7030 49644 7082
rect 49740 7030 49768 7082
rect 49636 7028 49684 7030
rect 49740 7028 49788 7030
rect 49844 7028 49892 7084
rect 49268 7018 49948 7028
rect 49084 6916 49140 6926
rect 49084 5906 49140 6860
rect 50092 6692 50148 8766
rect 50204 7812 50260 8990
rect 50316 8372 50372 11900
rect 50316 8306 50372 8316
rect 50428 10498 50484 10510
rect 50428 10446 50430 10498
rect 50482 10446 50484 10498
rect 50204 7746 50260 7756
rect 50092 6626 50148 6636
rect 50316 7474 50372 7486
rect 50316 7422 50318 7474
rect 50370 7422 50372 7474
rect 49980 6580 50036 6590
rect 49308 6468 49364 6478
rect 49084 5854 49086 5906
rect 49138 5854 49140 5906
rect 49084 5842 49140 5854
rect 49196 6412 49308 6468
rect 48972 5684 49028 5694
rect 49196 5684 49252 6412
rect 49308 6402 49364 6412
rect 49980 6018 50036 6524
rect 49980 5966 49982 6018
rect 50034 5966 50036 6018
rect 49980 5954 50036 5966
rect 50092 6132 50148 6142
rect 49308 5908 49364 5918
rect 49868 5908 49924 5918
rect 49308 5906 49924 5908
rect 49308 5854 49310 5906
rect 49362 5854 49870 5906
rect 49922 5854 49924 5906
rect 49308 5852 49924 5854
rect 49308 5842 49364 5852
rect 49868 5842 49924 5852
rect 49420 5684 49476 5694
rect 49196 5682 49476 5684
rect 49196 5630 49422 5682
rect 49474 5630 49476 5682
rect 49196 5628 49476 5630
rect 48972 5590 49028 5628
rect 49420 5618 49476 5628
rect 49268 5516 49948 5526
rect 49324 5460 49372 5516
rect 49428 5514 49476 5516
rect 49532 5514 49580 5516
rect 49448 5462 49476 5514
rect 49572 5462 49580 5514
rect 49428 5460 49476 5462
rect 49532 5460 49580 5462
rect 49636 5514 49684 5516
rect 49740 5514 49788 5516
rect 49636 5462 49644 5514
rect 49740 5462 49768 5514
rect 49636 5460 49684 5462
rect 49740 5460 49788 5462
rect 49844 5460 49892 5516
rect 48860 5404 49140 5460
rect 49268 5450 49948 5460
rect 48300 5124 48356 5134
rect 48300 5030 48356 5068
rect 48188 4340 48244 4350
rect 48188 4246 48244 4284
rect 49084 4338 49140 5404
rect 49868 5124 49924 5134
rect 49420 5012 49476 5022
rect 49420 4450 49476 4956
rect 49868 4562 49924 5068
rect 49868 4510 49870 4562
rect 49922 4510 49924 4562
rect 49868 4498 49924 4510
rect 49420 4398 49422 4450
rect 49474 4398 49476 4450
rect 49420 4386 49476 4398
rect 49756 4452 49812 4462
rect 49756 4358 49812 4396
rect 49980 4452 50036 4462
rect 49980 4358 50036 4396
rect 49084 4286 49086 4338
rect 49138 4286 49140 4338
rect 49084 4274 49140 4286
rect 48524 4116 48580 4126
rect 48524 3668 48580 4060
rect 49196 4116 49252 4154
rect 49196 4050 49252 4060
rect 49268 3948 49948 3958
rect 49324 3892 49372 3948
rect 49428 3946 49476 3948
rect 49532 3946 49580 3948
rect 49448 3894 49476 3946
rect 49572 3894 49580 3946
rect 49428 3892 49476 3894
rect 49532 3892 49580 3894
rect 49636 3946 49684 3948
rect 49740 3946 49788 3948
rect 49636 3894 49644 3946
rect 49740 3894 49768 3946
rect 49636 3892 49684 3894
rect 49740 3892 49788 3894
rect 49844 3892 49892 3948
rect 49268 3882 49948 3892
rect 50092 3780 50148 6076
rect 50316 5796 50372 7422
rect 50428 6132 50484 10446
rect 51100 10164 51156 12126
rect 51100 10098 51156 10108
rect 50428 6066 50484 6076
rect 50540 9042 50596 9054
rect 50540 8990 50542 9042
rect 50594 8990 50596 9042
rect 50428 5796 50484 5806
rect 50316 5794 50484 5796
rect 50316 5742 50430 5794
rect 50482 5742 50484 5794
rect 50316 5740 50484 5742
rect 50428 5236 50484 5740
rect 50204 5180 50484 5236
rect 50204 4452 50260 5180
rect 50540 4788 50596 8990
rect 51212 7700 51268 13582
rect 51324 12740 51380 12750
rect 51324 12646 51380 12684
rect 51212 7634 51268 7644
rect 51324 12066 51380 12078
rect 51324 12014 51326 12066
rect 51378 12014 51380 12066
rect 50764 5906 50820 5918
rect 50764 5854 50766 5906
rect 50818 5854 50820 5906
rect 50764 4900 50820 5854
rect 50764 4834 50820 4844
rect 50204 4386 50260 4396
rect 50316 4732 50596 4788
rect 47740 3614 47742 3666
rect 47794 3614 47796 3666
rect 47740 3602 47796 3614
rect 47964 3666 48580 3668
rect 47964 3614 48526 3666
rect 48578 3614 48580 3666
rect 47964 3612 48580 3614
rect 44492 3556 44548 3566
rect 44380 3554 44548 3556
rect 44380 3502 44494 3554
rect 44546 3502 44548 3554
rect 44380 3500 44548 3502
rect 44492 3490 44548 3500
rect 44940 3556 44996 3566
rect 43820 3444 43876 3482
rect 44940 3462 44996 3500
rect 46396 3556 46452 3566
rect 43820 3378 43876 3388
rect 43036 3278 43038 3330
rect 43090 3278 43092 3330
rect 43036 3266 43092 3278
rect 43932 3332 43988 3342
rect 43932 3238 43988 3276
rect 46396 3330 46452 3500
rect 47964 3554 48020 3612
rect 48524 3602 48580 3612
rect 49756 3724 50148 3780
rect 50204 3780 50260 3790
rect 47964 3502 47966 3554
rect 48018 3502 48020 3554
rect 47964 3490 48020 3502
rect 49308 3556 49364 3566
rect 46732 3444 46788 3482
rect 46732 3378 46788 3388
rect 48860 3444 48916 3482
rect 49308 3462 49364 3500
rect 49420 3554 49476 3566
rect 49420 3502 49422 3554
rect 49474 3502 49476 3554
rect 48860 3378 48916 3388
rect 49420 3444 49476 3502
rect 49420 3378 49476 3388
rect 49756 3442 49812 3724
rect 49980 3556 50036 3566
rect 50204 3556 50260 3724
rect 50316 3666 50372 4732
rect 51324 4338 51380 12014
rect 52108 10052 52164 13694
rect 53004 13746 53060 13916
rect 55580 13972 55636 13982
rect 55580 13878 55636 13916
rect 55132 13860 55188 13870
rect 55132 13766 55188 13804
rect 59052 13858 59108 13870
rect 59052 13806 59054 13858
rect 59106 13806 59108 13858
rect 53004 13694 53006 13746
rect 53058 13694 53060 13746
rect 53004 13682 53060 13694
rect 53452 13746 53508 13758
rect 53452 13694 53454 13746
rect 53506 13694 53508 13746
rect 52332 13636 52388 13646
rect 52332 13542 52388 13580
rect 52780 12290 52836 12302
rect 52780 12238 52782 12290
rect 52834 12238 52836 12290
rect 52108 9986 52164 9996
rect 52444 12180 52500 12190
rect 52780 12180 52836 12238
rect 52444 12178 52836 12180
rect 52444 12126 52446 12178
rect 52498 12126 52836 12178
rect 52444 12124 52836 12126
rect 51884 8258 51940 8270
rect 51884 8206 51886 8258
rect 51938 8206 51940 8258
rect 51884 7588 51940 8206
rect 51884 7522 51940 7532
rect 51996 7476 52052 7486
rect 51884 6804 51940 6814
rect 51996 6804 52052 7420
rect 51884 6802 52052 6804
rect 51884 6750 51886 6802
rect 51938 6750 52052 6802
rect 51884 6748 52052 6750
rect 51884 6738 51940 6748
rect 51772 5236 51828 5246
rect 51772 5142 51828 5180
rect 51324 4286 51326 4338
rect 51378 4286 51380 4338
rect 51324 4274 51380 4286
rect 52332 4564 52388 4574
rect 50316 3614 50318 3666
rect 50370 3614 50372 3666
rect 50316 3602 50372 3614
rect 51436 4116 51492 4126
rect 51436 3666 51492 4060
rect 51436 3614 51438 3666
rect 51490 3614 51492 3666
rect 51436 3602 51492 3614
rect 51884 3668 51940 3678
rect 52332 3668 52388 4508
rect 51884 3666 52388 3668
rect 51884 3614 51886 3666
rect 51938 3614 52334 3666
rect 52386 3614 52388 3666
rect 51884 3612 52388 3614
rect 51884 3602 51940 3612
rect 52332 3602 52388 3612
rect 52444 3668 52500 12124
rect 53228 10610 53284 10622
rect 53228 10558 53230 10610
rect 53282 10558 53284 10610
rect 52780 9826 52836 9838
rect 52780 9774 52782 9826
rect 52834 9774 52836 9826
rect 52668 8258 52724 8270
rect 52668 8206 52670 8258
rect 52722 8206 52724 8258
rect 52668 4452 52724 8206
rect 52780 7476 52836 9774
rect 52780 7410 52836 7420
rect 53228 5236 53284 10558
rect 53452 5348 53508 13694
rect 54572 13748 54628 13758
rect 54572 13654 54628 13692
rect 58828 13746 58884 13758
rect 58828 13694 58830 13746
rect 58882 13694 58884 13746
rect 58828 13524 58884 13694
rect 58940 13524 58996 13534
rect 58828 13468 58940 13524
rect 58940 13458 58996 13468
rect 58268 13356 58948 13366
rect 58324 13300 58372 13356
rect 58428 13354 58476 13356
rect 58532 13354 58580 13356
rect 58448 13302 58476 13354
rect 58572 13302 58580 13354
rect 58428 13300 58476 13302
rect 58532 13300 58580 13302
rect 58636 13354 58684 13356
rect 58740 13354 58788 13356
rect 58636 13302 58644 13354
rect 58740 13302 58768 13354
rect 58636 13300 58684 13302
rect 58740 13300 58788 13302
rect 58844 13300 58892 13356
rect 58268 13290 58948 13300
rect 53768 12572 54448 12582
rect 53824 12516 53872 12572
rect 53928 12570 53976 12572
rect 54032 12570 54080 12572
rect 53948 12518 53976 12570
rect 54072 12518 54080 12570
rect 53928 12516 53976 12518
rect 54032 12516 54080 12518
rect 54136 12570 54184 12572
rect 54240 12570 54288 12572
rect 54136 12518 54144 12570
rect 54240 12518 54268 12570
rect 54136 12516 54184 12518
rect 54240 12516 54288 12518
rect 54344 12516 54392 12572
rect 53768 12506 54448 12516
rect 57820 12404 57876 12414
rect 57708 12348 57820 12404
rect 56140 11394 56196 11406
rect 56140 11342 56142 11394
rect 56194 11342 56196 11394
rect 53768 11004 54448 11014
rect 53824 10948 53872 11004
rect 53928 11002 53976 11004
rect 54032 11002 54080 11004
rect 53948 10950 53976 11002
rect 54072 10950 54080 11002
rect 53928 10948 53976 10950
rect 54032 10948 54080 10950
rect 54136 11002 54184 11004
rect 54240 11002 54288 11004
rect 54136 10950 54144 11002
rect 54240 10950 54268 11002
rect 54136 10948 54184 10950
rect 54240 10948 54288 10950
rect 54344 10948 54392 11004
rect 53768 10938 54448 10948
rect 54684 10164 54740 10174
rect 54684 9938 54740 10108
rect 54684 9886 54686 9938
rect 54738 9886 54740 9938
rect 54684 9874 54740 9886
rect 53768 9436 54448 9446
rect 53824 9380 53872 9436
rect 53928 9434 53976 9436
rect 54032 9434 54080 9436
rect 53948 9382 53976 9434
rect 54072 9382 54080 9434
rect 53928 9380 53976 9382
rect 54032 9380 54080 9382
rect 54136 9434 54184 9436
rect 54240 9434 54288 9436
rect 54136 9382 54144 9434
rect 54240 9382 54268 9434
rect 54136 9380 54184 9382
rect 54240 9380 54288 9382
rect 54344 9380 54392 9436
rect 53768 9370 54448 9380
rect 54572 8930 54628 8942
rect 54572 8878 54574 8930
rect 54626 8878 54628 8930
rect 53768 7868 54448 7878
rect 53824 7812 53872 7868
rect 53928 7866 53976 7868
rect 54032 7866 54080 7868
rect 53948 7814 53976 7866
rect 54072 7814 54080 7866
rect 53928 7812 53976 7814
rect 54032 7812 54080 7814
rect 54136 7866 54184 7868
rect 54240 7866 54288 7868
rect 54136 7814 54144 7866
rect 54240 7814 54268 7866
rect 54136 7812 54184 7814
rect 54240 7812 54288 7814
rect 54344 7812 54392 7868
rect 53768 7802 54448 7812
rect 53788 7362 53844 7374
rect 53788 7310 53790 7362
rect 53842 7310 53844 7362
rect 53788 6468 53844 7310
rect 54348 6692 54404 6702
rect 54572 6692 54628 8878
rect 56140 8372 56196 11342
rect 56140 8306 56196 8316
rect 56700 11282 56756 11294
rect 56700 11230 56702 11282
rect 56754 11230 56756 11282
rect 54684 8148 54740 8158
rect 54684 8054 54740 8092
rect 54348 6690 54628 6692
rect 54348 6638 54350 6690
rect 54402 6638 54628 6690
rect 54348 6636 54628 6638
rect 54348 6626 54404 6636
rect 53788 6402 53844 6412
rect 53768 6300 54448 6310
rect 53824 6244 53872 6300
rect 53928 6298 53976 6300
rect 54032 6298 54080 6300
rect 53948 6246 53976 6298
rect 54072 6246 54080 6298
rect 53928 6244 53976 6246
rect 54032 6244 54080 6246
rect 54136 6298 54184 6300
rect 54240 6298 54288 6300
rect 54136 6246 54144 6298
rect 54240 6246 54268 6298
rect 54136 6244 54184 6246
rect 54240 6244 54288 6246
rect 54344 6244 54392 6300
rect 53768 6234 54448 6244
rect 54572 5908 54628 6636
rect 54572 5842 54628 5852
rect 54684 7700 54740 7710
rect 53452 5282 53508 5292
rect 53228 5170 53284 5180
rect 54684 5234 54740 7644
rect 55356 7476 55412 7486
rect 54908 6580 54964 6590
rect 54908 6486 54964 6524
rect 55356 6018 55412 7420
rect 56588 7476 56644 7486
rect 56588 7382 56644 7420
rect 55356 5966 55358 6018
rect 55410 5966 55412 6018
rect 55356 5954 55412 5966
rect 54684 5182 54686 5234
rect 54738 5182 54740 5234
rect 54684 5170 54740 5182
rect 53768 4732 54448 4742
rect 53824 4676 53872 4732
rect 53928 4730 53976 4732
rect 54032 4730 54080 4732
rect 53948 4678 53976 4730
rect 54072 4678 54080 4730
rect 53928 4676 53976 4678
rect 54032 4676 54080 4678
rect 54136 4730 54184 4732
rect 54240 4730 54288 4732
rect 54136 4678 54144 4730
rect 54240 4678 54268 4730
rect 54136 4676 54184 4678
rect 54240 4676 54288 4678
rect 54344 4676 54392 4732
rect 53768 4666 54448 4676
rect 52780 4452 52836 4462
rect 52668 4396 52780 4452
rect 52780 4358 52836 4396
rect 56700 3780 56756 11230
rect 57148 5906 57204 5918
rect 57148 5854 57150 5906
rect 57202 5854 57204 5906
rect 57148 5236 57204 5854
rect 57148 5170 57204 5180
rect 56700 3714 56756 3724
rect 57484 4116 57540 4126
rect 52444 3602 52500 3612
rect 55468 3668 55524 3678
rect 55468 3574 55524 3612
rect 57484 3666 57540 4060
rect 57708 3892 57764 12348
rect 57820 12338 57876 12348
rect 59052 12404 59108 13806
rect 60508 13748 60564 13758
rect 60396 13746 60564 13748
rect 60396 13694 60510 13746
rect 60562 13694 60564 13746
rect 60396 13692 60564 13694
rect 59052 12338 59108 12348
rect 60284 13524 60340 13534
rect 58268 11788 58948 11798
rect 58324 11732 58372 11788
rect 58428 11786 58476 11788
rect 58532 11786 58580 11788
rect 58448 11734 58476 11786
rect 58572 11734 58580 11786
rect 58428 11732 58476 11734
rect 58532 11732 58580 11734
rect 58636 11786 58684 11788
rect 58740 11786 58788 11788
rect 58636 11734 58644 11786
rect 58740 11734 58768 11786
rect 58636 11732 58684 11734
rect 58740 11732 58788 11734
rect 58844 11732 58892 11788
rect 58268 11722 58948 11732
rect 58156 11396 58212 11406
rect 58156 11302 58212 11340
rect 59388 11394 59444 11406
rect 59388 11342 59390 11394
rect 59442 11342 59444 11394
rect 58044 11282 58100 11294
rect 58044 11230 58046 11282
rect 58098 11230 58100 11282
rect 57820 8372 57876 8382
rect 57876 8316 57988 8372
rect 57820 8306 57876 8316
rect 57932 5572 57988 8316
rect 58044 6692 58100 11230
rect 59164 11284 59220 11294
rect 59388 11284 59444 11342
rect 59164 11282 59444 11284
rect 59164 11230 59166 11282
rect 59218 11230 59444 11282
rect 59164 11228 59444 11230
rect 59164 11218 59220 11228
rect 59388 11172 59444 11228
rect 58268 10220 58948 10230
rect 58324 10164 58372 10220
rect 58428 10218 58476 10220
rect 58532 10218 58580 10220
rect 58448 10166 58476 10218
rect 58572 10166 58580 10218
rect 58428 10164 58476 10166
rect 58532 10164 58580 10166
rect 58636 10218 58684 10220
rect 58740 10218 58788 10220
rect 58636 10166 58644 10218
rect 58740 10166 58768 10218
rect 58636 10164 58684 10166
rect 58740 10164 58788 10166
rect 58844 10164 58892 10220
rect 58268 10154 58948 10164
rect 59276 10052 59332 10062
rect 58268 8652 58948 8662
rect 58324 8596 58372 8652
rect 58428 8650 58476 8652
rect 58532 8650 58580 8652
rect 58448 8598 58476 8650
rect 58572 8598 58580 8650
rect 58428 8596 58476 8598
rect 58532 8596 58580 8598
rect 58636 8650 58684 8652
rect 58740 8650 58788 8652
rect 58636 8598 58644 8650
rect 58740 8598 58768 8650
rect 58636 8596 58684 8598
rect 58740 8596 58788 8598
rect 58844 8596 58892 8652
rect 58268 8586 58948 8596
rect 58828 8372 58884 8382
rect 58828 8278 58884 8316
rect 58940 8258 58996 8270
rect 58940 8206 58942 8258
rect 58994 8206 58996 8258
rect 58828 8034 58884 8046
rect 58828 7982 58830 8034
rect 58882 7982 58884 8034
rect 58828 7252 58884 7982
rect 58940 7364 58996 8206
rect 59164 8258 59220 8270
rect 59164 8206 59166 8258
rect 59218 8206 59220 8258
rect 59164 7588 59220 8206
rect 59164 7522 59220 7532
rect 59276 7586 59332 9996
rect 59276 7534 59278 7586
rect 59330 7534 59332 7586
rect 59276 7522 59332 7534
rect 58940 7308 59220 7364
rect 58828 7196 59108 7252
rect 58268 7084 58948 7094
rect 58324 7028 58372 7084
rect 58428 7082 58476 7084
rect 58532 7082 58580 7084
rect 58448 7030 58476 7082
rect 58572 7030 58580 7082
rect 58428 7028 58476 7030
rect 58532 7028 58580 7030
rect 58636 7082 58684 7084
rect 58740 7082 58788 7084
rect 58636 7030 58644 7082
rect 58740 7030 58768 7082
rect 58636 7028 58684 7030
rect 58740 7028 58788 7030
rect 58844 7028 58892 7084
rect 58268 7018 58948 7028
rect 58044 6626 58100 6636
rect 58828 6804 58884 6814
rect 58828 6018 58884 6748
rect 59052 6580 59108 7196
rect 59164 6916 59220 7308
rect 59276 6916 59332 6926
rect 59164 6914 59332 6916
rect 59164 6862 59278 6914
rect 59330 6862 59332 6914
rect 59164 6860 59332 6862
rect 59276 6850 59332 6860
rect 59052 6514 59108 6524
rect 59388 6468 59444 11116
rect 59948 10610 60004 10622
rect 59948 10558 59950 10610
rect 60002 10558 60004 10610
rect 59836 8930 59892 8942
rect 59836 8878 59838 8930
rect 59890 8878 59892 8930
rect 59500 6916 59556 6926
rect 59724 6916 59780 6926
rect 59500 6914 59780 6916
rect 59500 6862 59502 6914
rect 59554 6862 59726 6914
rect 59778 6862 59780 6914
rect 59500 6860 59780 6862
rect 59500 6850 59556 6860
rect 59724 6850 59780 6860
rect 59836 6690 59892 8878
rect 59836 6638 59838 6690
rect 59890 6638 59892 6690
rect 59836 6626 59892 6638
rect 58828 5966 58830 6018
rect 58882 5966 58884 6018
rect 58828 5954 58884 5966
rect 59276 6466 59444 6468
rect 59276 6414 59390 6466
rect 59442 6414 59444 6466
rect 59276 6412 59444 6414
rect 57932 5516 58100 5572
rect 57932 5348 57988 5358
rect 58044 5348 58100 5516
rect 58268 5516 58948 5526
rect 58324 5460 58372 5516
rect 58428 5514 58476 5516
rect 58532 5514 58580 5516
rect 58448 5462 58476 5514
rect 58572 5462 58580 5514
rect 58428 5460 58476 5462
rect 58532 5460 58580 5462
rect 58636 5514 58684 5516
rect 58740 5514 58788 5516
rect 58636 5462 58644 5514
rect 58740 5462 58768 5514
rect 58636 5460 58684 5462
rect 58740 5460 58788 5462
rect 58844 5460 58892 5516
rect 58268 5450 58948 5460
rect 58268 5348 58324 5358
rect 58044 5346 58324 5348
rect 58044 5294 58270 5346
rect 58322 5294 58324 5346
rect 58044 5292 58324 5294
rect 57932 5122 57988 5292
rect 58268 5282 58324 5292
rect 58716 5348 58772 5358
rect 57932 5070 57934 5122
rect 57986 5070 57988 5122
rect 57932 5058 57988 5070
rect 58716 4450 58772 5292
rect 59164 5124 59220 5134
rect 59164 5030 59220 5068
rect 59052 5010 59108 5022
rect 59052 4958 59054 5010
rect 59106 4958 59108 5010
rect 59052 4900 59108 4958
rect 59276 5010 59332 6412
rect 59388 6402 59444 6412
rect 59836 6356 59892 6366
rect 59836 5348 59892 6300
rect 59948 5572 60004 10558
rect 59948 5516 60116 5572
rect 59948 5348 60004 5358
rect 59836 5346 60004 5348
rect 59836 5294 59950 5346
rect 60002 5294 60004 5346
rect 59836 5292 60004 5294
rect 59948 5282 60004 5292
rect 59836 5122 59892 5134
rect 59836 5070 59838 5122
rect 59890 5070 59892 5122
rect 59276 4958 59278 5010
rect 59330 4958 59332 5010
rect 59276 4900 59332 4958
rect 59612 5012 59668 5022
rect 59612 4918 59668 4956
rect 59052 4844 59332 4900
rect 58716 4398 58718 4450
rect 58770 4398 58772 4450
rect 58716 4386 58772 4398
rect 59276 4340 59332 4844
rect 59276 4274 59332 4284
rect 59388 4900 59444 4910
rect 59388 4116 59444 4844
rect 58268 3948 58948 3958
rect 58324 3892 58372 3948
rect 58428 3946 58476 3948
rect 58532 3946 58580 3948
rect 58448 3894 58476 3946
rect 58572 3894 58580 3946
rect 58428 3892 58476 3894
rect 58532 3892 58580 3894
rect 58636 3946 58684 3948
rect 58740 3946 58788 3948
rect 58636 3894 58644 3946
rect 58740 3894 58768 3946
rect 58636 3892 58684 3894
rect 58740 3892 58788 3894
rect 58844 3892 58892 3948
rect 57708 3836 58212 3892
rect 58268 3882 58948 3892
rect 58156 3780 58212 3836
rect 58268 3780 58324 3790
rect 58156 3778 58324 3780
rect 58156 3726 58270 3778
rect 58322 3726 58324 3778
rect 58156 3724 58324 3726
rect 58268 3714 58324 3724
rect 59052 3780 59108 3790
rect 57484 3614 57486 3666
rect 57538 3614 57540 3666
rect 57484 3602 57540 3614
rect 59052 3666 59108 3724
rect 59052 3614 59054 3666
rect 59106 3614 59108 3666
rect 59052 3602 59108 3614
rect 49980 3554 50260 3556
rect 49980 3502 49982 3554
rect 50034 3502 50206 3554
rect 50258 3502 50260 3554
rect 49980 3500 50260 3502
rect 49980 3490 50036 3500
rect 50204 3490 50260 3500
rect 50428 3556 50484 3566
rect 50428 3444 50484 3500
rect 54572 3556 54628 3566
rect 49756 3390 49758 3442
rect 49810 3390 49812 3442
rect 49756 3378 49812 3390
rect 50316 3388 50484 3444
rect 52668 3444 52724 3482
rect 54572 3462 54628 3500
rect 55020 3556 55076 3566
rect 55020 3462 55076 3500
rect 57820 3556 57876 3566
rect 58156 3556 58212 3566
rect 57820 3554 58156 3556
rect 57820 3502 57822 3554
rect 57874 3502 58156 3554
rect 57820 3500 58156 3502
rect 57820 3490 57876 3500
rect 58156 3462 58212 3500
rect 59388 3554 59444 4060
rect 59836 3668 59892 5070
rect 59836 3602 59892 3612
rect 59388 3502 59390 3554
rect 59442 3502 59444 3554
rect 59388 3490 59444 3502
rect 60060 3554 60116 5516
rect 60284 4228 60340 13468
rect 60396 12290 60452 13692
rect 60508 13682 60564 13692
rect 61068 13634 61124 13646
rect 61068 13582 61070 13634
rect 61122 13582 61124 13634
rect 61068 13076 61124 13582
rect 61068 13020 61236 13076
rect 61068 12852 61124 12862
rect 60396 12238 60398 12290
rect 60450 12238 60452 12290
rect 60396 12226 60452 12238
rect 60732 12850 61124 12852
rect 60732 12798 61070 12850
rect 61122 12798 61124 12850
rect 60732 12796 61124 12798
rect 60620 11172 60676 11182
rect 60620 11078 60676 11116
rect 60508 6692 60564 6702
rect 60508 6598 60564 6636
rect 60732 6020 60788 12796
rect 61068 12786 61124 12796
rect 61068 11172 61124 11182
rect 61068 11078 61124 11116
rect 61180 7140 61236 13020
rect 61292 11508 61348 28140
rect 61628 27074 61684 28364
rect 62636 28420 62692 28430
rect 62636 27748 62692 28364
rect 63084 28420 63140 28458
rect 63084 28354 63140 28364
rect 62768 28252 63448 28262
rect 62824 28196 62872 28252
rect 62928 28250 62976 28252
rect 63032 28250 63080 28252
rect 62948 28198 62976 28250
rect 63072 28198 63080 28250
rect 62928 28196 62976 28198
rect 63032 28196 63080 28198
rect 63136 28250 63184 28252
rect 63240 28250 63288 28252
rect 63136 28198 63144 28250
rect 63240 28198 63268 28250
rect 63136 28196 63184 28198
rect 63240 28196 63288 28198
rect 63344 28196 63392 28252
rect 62768 28186 63448 28196
rect 62636 27692 63140 27748
rect 61628 27022 61630 27074
rect 61682 27022 61684 27074
rect 61628 27010 61684 27022
rect 61740 27636 61796 27646
rect 61740 26964 61796 27580
rect 62748 27076 62804 27086
rect 61740 26870 61796 26908
rect 61964 26964 62020 26974
rect 62300 26964 62356 27002
rect 62748 26982 62804 27020
rect 63084 27074 63140 27692
rect 63084 27022 63086 27074
rect 63138 27022 63140 27074
rect 63084 27010 63140 27022
rect 61964 26962 62244 26964
rect 61964 26910 61966 26962
rect 62018 26910 62244 26962
rect 61964 26908 62244 26910
rect 61964 26898 62020 26908
rect 61404 26852 61460 26862
rect 61404 26758 61460 26796
rect 62188 25508 62244 26908
rect 62300 26898 62356 26908
rect 62300 26740 62356 26750
rect 62300 26292 62356 26684
rect 62768 26684 63448 26694
rect 62824 26628 62872 26684
rect 62928 26682 62976 26684
rect 63032 26682 63080 26684
rect 62948 26630 62976 26682
rect 63072 26630 63080 26682
rect 62928 26628 62976 26630
rect 63032 26628 63080 26630
rect 63136 26682 63184 26684
rect 63240 26682 63288 26684
rect 63136 26630 63144 26682
rect 63240 26630 63268 26682
rect 63136 26628 63184 26630
rect 63240 26628 63288 26630
rect 63344 26628 63392 26684
rect 62768 26618 63448 26628
rect 62300 26198 62356 26236
rect 62300 25508 62356 25518
rect 62188 25506 62356 25508
rect 62188 25454 62302 25506
rect 62354 25454 62356 25506
rect 62188 25452 62356 25454
rect 62300 25442 62356 25452
rect 62972 25508 63028 25518
rect 62972 25414 63028 25452
rect 61852 25284 61908 25294
rect 61740 25282 61908 25284
rect 61740 25230 61854 25282
rect 61906 25230 61908 25282
rect 61740 25228 61908 25230
rect 61740 23938 61796 25228
rect 61852 25218 61908 25228
rect 62412 25282 62468 25294
rect 62412 25230 62414 25282
rect 62466 25230 62468 25282
rect 61740 23886 61742 23938
rect 61794 23886 61796 23938
rect 61740 23874 61796 23886
rect 62076 24500 62132 24510
rect 61404 23716 61460 23726
rect 62076 23716 62132 24444
rect 62188 23940 62244 23950
rect 62412 23940 62468 25230
rect 62524 25284 62580 25294
rect 62524 25190 62580 25228
rect 63308 25284 63364 25322
rect 63532 25284 63588 28588
rect 63644 28642 63700 28654
rect 63644 28590 63646 28642
rect 63698 28590 63700 28642
rect 63644 27636 63700 28590
rect 64428 28644 64484 28654
rect 64428 28550 64484 28588
rect 64764 28644 64820 34076
rect 64876 34066 64932 34076
rect 65436 34066 65492 34076
rect 65548 33908 65604 34300
rect 65436 33852 65604 33908
rect 64876 32450 64932 32462
rect 64876 32398 64878 32450
rect 64930 32398 64932 32450
rect 64876 31668 64932 32398
rect 65100 31668 65156 31678
rect 64876 31612 65100 31668
rect 65100 31574 65156 31612
rect 65212 31554 65268 31566
rect 65212 31502 65214 31554
rect 65266 31502 65268 31554
rect 65100 31220 65156 31230
rect 65100 30994 65156 31164
rect 65100 30942 65102 30994
rect 65154 30942 65156 30994
rect 65100 30930 65156 30942
rect 65212 30996 65268 31502
rect 65324 31556 65380 31566
rect 65324 31462 65380 31500
rect 65436 31332 65492 33852
rect 66108 33684 66164 33694
rect 66108 33122 66164 33628
rect 67004 33684 67060 34636
rect 67900 34692 67956 34702
rect 67900 34598 67956 34636
rect 68012 34244 68068 36316
rect 68460 36258 68516 36270
rect 68460 36206 68462 36258
rect 68514 36206 68516 36258
rect 68124 36036 68180 36046
rect 68124 35698 68180 35980
rect 68460 36036 68516 36206
rect 68460 35970 68516 35980
rect 68348 35866 68404 35878
rect 68348 35814 68350 35866
rect 68402 35814 68404 35866
rect 68124 35646 68126 35698
rect 68178 35646 68180 35698
rect 68124 35634 68180 35646
rect 68236 35700 68292 35710
rect 68012 34178 68068 34188
rect 67268 33740 67948 33750
rect 67324 33684 67372 33740
rect 67428 33738 67476 33740
rect 67532 33738 67580 33740
rect 67448 33686 67476 33738
rect 67572 33686 67580 33738
rect 67428 33684 67476 33686
rect 67532 33684 67580 33686
rect 67636 33738 67684 33740
rect 67740 33738 67788 33740
rect 67636 33686 67644 33738
rect 67740 33686 67768 33738
rect 67636 33684 67684 33686
rect 67740 33684 67788 33686
rect 67844 33684 67892 33740
rect 67268 33674 67948 33684
rect 67004 33458 67060 33628
rect 67004 33406 67006 33458
rect 67058 33406 67060 33458
rect 66108 33070 66110 33122
rect 66162 33070 66164 33122
rect 66108 33058 66164 33070
rect 66668 33124 66724 33134
rect 66668 33030 66724 33068
rect 67004 31892 67060 33406
rect 68236 32676 68292 35644
rect 68348 35364 68404 35814
rect 68684 35812 68740 35822
rect 68348 35298 68404 35308
rect 68460 35810 68740 35812
rect 68460 35758 68686 35810
rect 68738 35758 68740 35810
rect 68460 35756 68740 35758
rect 68460 34914 68516 35756
rect 68684 35746 68740 35756
rect 68460 34862 68462 34914
rect 68514 34862 68516 34914
rect 68460 34850 68516 34862
rect 68796 34692 68852 36316
rect 69468 36306 69524 36316
rect 69580 36820 69636 36830
rect 69580 36370 69636 36764
rect 73500 36596 73556 37998
rect 73948 38050 74004 38062
rect 73948 37998 73950 38050
rect 74002 37998 74004 38050
rect 73948 37940 74004 37998
rect 73948 37874 74004 37884
rect 74284 37940 74340 37950
rect 74284 37846 74340 37884
rect 73500 36530 73556 36540
rect 69580 36318 69582 36370
rect 69634 36318 69636 36370
rect 69580 35924 69636 36318
rect 71768 36092 72448 36102
rect 71824 36036 71872 36092
rect 71928 36090 71976 36092
rect 72032 36090 72080 36092
rect 71948 36038 71976 36090
rect 72072 36038 72080 36090
rect 71928 36036 71976 36038
rect 72032 36036 72080 36038
rect 72136 36090 72184 36092
rect 72240 36090 72288 36092
rect 72136 36038 72144 36090
rect 72240 36038 72268 36090
rect 72136 36036 72184 36038
rect 72240 36036 72288 36038
rect 72344 36036 72392 36092
rect 71768 36026 72448 36036
rect 69580 35858 69636 35868
rect 71932 35924 71988 35934
rect 68908 35364 68964 35374
rect 68908 34914 68964 35308
rect 71932 35138 71988 35868
rect 73724 35924 73780 35934
rect 72380 35812 72436 35822
rect 71932 35086 71934 35138
rect 71986 35086 71988 35138
rect 71932 35074 71988 35086
rect 72156 35810 72436 35812
rect 72156 35758 72382 35810
rect 72434 35758 72436 35810
rect 72156 35756 72436 35758
rect 68908 34862 68910 34914
rect 68962 34862 68964 34914
rect 68908 34850 68964 34862
rect 72156 34914 72212 35756
rect 72380 35746 72436 35756
rect 72156 34862 72158 34914
rect 72210 34862 72212 34914
rect 72156 34850 72212 34862
rect 72716 34914 72772 34926
rect 72716 34862 72718 34914
rect 72770 34862 72772 34914
rect 68236 32610 68292 32620
rect 68460 34636 68852 34692
rect 71148 34692 71204 34702
rect 67268 32172 67948 32182
rect 67324 32116 67372 32172
rect 67428 32170 67476 32172
rect 67532 32170 67580 32172
rect 67448 32118 67476 32170
rect 67572 32118 67580 32170
rect 67428 32116 67476 32118
rect 67532 32116 67580 32118
rect 67636 32170 67684 32172
rect 67740 32170 67788 32172
rect 67636 32118 67644 32170
rect 67740 32118 67768 32170
rect 67636 32116 67684 32118
rect 67740 32116 67788 32118
rect 67844 32116 67892 32172
rect 67268 32106 67948 32116
rect 67004 31826 67060 31836
rect 67900 31892 67956 31902
rect 65772 31780 65828 31790
rect 65772 31778 66500 31780
rect 65772 31726 65774 31778
rect 65826 31726 66500 31778
rect 65772 31724 66500 31726
rect 65772 31714 65828 31724
rect 65212 30930 65268 30940
rect 65324 31276 65492 31332
rect 65996 31554 66052 31566
rect 65996 31502 65998 31554
rect 66050 31502 66052 31554
rect 64764 28578 64820 28588
rect 63644 27570 63700 27580
rect 63868 28418 63924 28430
rect 63868 28366 63870 28418
rect 63922 28366 63924 28418
rect 63868 27076 63924 28366
rect 63868 27010 63924 27020
rect 63364 25228 63588 25284
rect 63308 25218 63364 25228
rect 62768 25116 63448 25126
rect 62824 25060 62872 25116
rect 62928 25114 62976 25116
rect 63032 25114 63080 25116
rect 62948 25062 62976 25114
rect 63072 25062 63080 25114
rect 62928 25060 62976 25062
rect 63032 25060 63080 25062
rect 63136 25114 63184 25116
rect 63240 25114 63288 25116
rect 63136 25062 63144 25114
rect 63240 25062 63268 25114
rect 63136 25060 63184 25062
rect 63240 25060 63288 25062
rect 63344 25060 63392 25116
rect 62768 25050 63448 25060
rect 62188 23938 62468 23940
rect 62188 23886 62190 23938
rect 62242 23886 62468 23938
rect 62188 23884 62468 23886
rect 62188 23874 62244 23884
rect 62076 23660 62356 23716
rect 61404 23622 61460 23660
rect 62300 23378 62356 23660
rect 62768 23548 63448 23558
rect 62824 23492 62872 23548
rect 62928 23546 62976 23548
rect 63032 23546 63080 23548
rect 62948 23494 62976 23546
rect 63072 23494 63080 23546
rect 62928 23492 62976 23494
rect 63032 23492 63080 23494
rect 63136 23546 63184 23548
rect 63240 23546 63288 23548
rect 63136 23494 63144 23546
rect 63240 23494 63268 23546
rect 63136 23492 63184 23494
rect 63240 23492 63288 23494
rect 63344 23492 63392 23548
rect 62768 23482 63448 23492
rect 62300 23326 62302 23378
rect 62354 23326 62356 23378
rect 62300 23314 62356 23326
rect 62524 23380 62580 23390
rect 63308 23380 63364 23390
rect 63532 23380 63588 25228
rect 62524 23378 63588 23380
rect 62524 23326 62526 23378
rect 62578 23326 63310 23378
rect 63362 23326 63588 23378
rect 62524 23324 63588 23326
rect 64540 26292 64596 26302
rect 62524 23314 62580 23324
rect 63308 23314 63364 23324
rect 62972 23156 63028 23166
rect 62972 23062 63028 23100
rect 64204 23156 64260 23166
rect 62412 23042 62468 23054
rect 62412 22990 62414 23042
rect 62466 22990 62468 23042
rect 61852 22148 61908 22158
rect 61740 22146 61908 22148
rect 61740 22094 61854 22146
rect 61906 22094 61908 22146
rect 61740 22092 61908 22094
rect 61740 20802 61796 22092
rect 61852 22082 61908 22092
rect 61740 20750 61742 20802
rect 61794 20750 61796 20802
rect 61740 20738 61796 20750
rect 62188 20804 62244 20814
rect 62412 20804 62468 22990
rect 62768 21980 63448 21990
rect 62824 21924 62872 21980
rect 62928 21978 62976 21980
rect 63032 21978 63080 21980
rect 62948 21926 62976 21978
rect 63072 21926 63080 21978
rect 62928 21924 62976 21926
rect 63032 21924 63080 21926
rect 63136 21978 63184 21980
rect 63240 21978 63288 21980
rect 63136 21926 63144 21978
rect 63240 21926 63268 21978
rect 63136 21924 63184 21926
rect 63240 21924 63288 21926
rect 63344 21924 63392 21980
rect 62768 21914 63448 21924
rect 64204 21812 64260 23100
rect 64316 22372 64372 22382
rect 64540 22372 64596 26236
rect 65324 26068 65380 31276
rect 65996 31220 66052 31502
rect 65996 31154 66052 31164
rect 65436 30996 65492 31006
rect 65436 30902 65492 30940
rect 66444 30210 66500 31724
rect 66556 31556 66612 31566
rect 66556 31462 66612 31500
rect 67900 31220 67956 31836
rect 67900 31218 68068 31220
rect 67900 31166 67902 31218
rect 67954 31166 68068 31218
rect 67900 31164 68068 31166
rect 67900 31154 67956 31164
rect 67268 30604 67948 30614
rect 67324 30548 67372 30604
rect 67428 30602 67476 30604
rect 67532 30602 67580 30604
rect 67448 30550 67476 30602
rect 67572 30550 67580 30602
rect 67428 30548 67476 30550
rect 67532 30548 67580 30550
rect 67636 30602 67684 30604
rect 67740 30602 67788 30604
rect 67636 30550 67644 30602
rect 67740 30550 67768 30602
rect 67636 30548 67684 30550
rect 67740 30548 67788 30550
rect 67844 30548 67892 30604
rect 67268 30538 67948 30548
rect 66444 30158 66446 30210
rect 66498 30158 66500 30210
rect 66444 30146 66500 30158
rect 66668 30212 66724 30222
rect 66668 30098 66724 30156
rect 66668 30046 66670 30098
rect 66722 30046 66724 30098
rect 66668 30034 66724 30046
rect 66780 30100 66836 30110
rect 67228 30100 67284 30110
rect 66780 30098 67284 30100
rect 66780 30046 66782 30098
rect 66834 30046 67230 30098
rect 67282 30046 67284 30098
rect 66780 30044 67284 30046
rect 66780 28308 66836 30044
rect 67228 30034 67284 30044
rect 67268 29036 67948 29046
rect 67324 28980 67372 29036
rect 67428 29034 67476 29036
rect 67532 29034 67580 29036
rect 67448 28982 67476 29034
rect 67572 28982 67580 29034
rect 67428 28980 67476 28982
rect 67532 28980 67580 28982
rect 67636 29034 67684 29036
rect 67740 29034 67788 29036
rect 67636 28982 67644 29034
rect 67740 28982 67768 29034
rect 67636 28980 67684 28982
rect 67740 28980 67788 28982
rect 67844 28980 67892 29036
rect 67268 28970 67948 28980
rect 68012 28868 68068 31164
rect 67340 28812 68068 28868
rect 68348 29316 68404 29326
rect 67340 28756 67396 28812
rect 66220 28252 66836 28308
rect 66220 28082 66276 28252
rect 66220 28030 66222 28082
rect 66274 28030 66276 28082
rect 65660 27972 65716 27982
rect 65660 27878 65716 27916
rect 65772 27860 65828 27870
rect 66220 27860 66276 28030
rect 65772 27858 66276 27860
rect 65772 27806 65774 27858
rect 65826 27806 66276 27858
rect 65772 27804 66276 27806
rect 66332 27972 66388 27982
rect 65660 27636 65716 27646
rect 65660 27542 65716 27580
rect 65436 26962 65492 26974
rect 65436 26910 65438 26962
rect 65490 26910 65492 26962
rect 65436 26292 65492 26910
rect 65436 26226 65492 26236
rect 65324 26012 65492 26068
rect 65324 25620 65380 25630
rect 64988 25508 65044 25518
rect 64988 25414 65044 25452
rect 65324 25506 65380 25564
rect 65324 25454 65326 25506
rect 65378 25454 65380 25506
rect 65324 25442 65380 25454
rect 65212 25282 65268 25294
rect 65212 25230 65214 25282
rect 65266 25230 65268 25282
rect 64652 23828 64708 23838
rect 64652 23714 64708 23772
rect 64652 23662 64654 23714
rect 64706 23662 64708 23714
rect 64652 23650 64708 23662
rect 65212 23714 65268 25230
rect 65212 23662 65214 23714
rect 65266 23662 65268 23714
rect 65212 23604 65268 23662
rect 65212 23538 65268 23548
rect 64652 22372 64708 22382
rect 64316 22370 64708 22372
rect 64316 22318 64318 22370
rect 64370 22318 64654 22370
rect 64706 22318 64708 22370
rect 64316 22316 64708 22318
rect 64316 22306 64372 22316
rect 64652 22306 64708 22316
rect 64316 21812 64372 21822
rect 64204 21810 64372 21812
rect 64204 21758 64318 21810
rect 64370 21758 64372 21810
rect 64204 21756 64372 21758
rect 64316 21746 64372 21756
rect 64540 21698 64596 21710
rect 64540 21646 64542 21698
rect 64594 21646 64596 21698
rect 64540 21028 64596 21646
rect 64652 21700 64708 21710
rect 64652 21606 64708 21644
rect 65100 21700 65156 21710
rect 65100 21606 65156 21644
rect 64540 20962 64596 20972
rect 65212 21028 65268 21038
rect 65212 20934 65268 20972
rect 62188 20802 62468 20804
rect 62188 20750 62190 20802
rect 62242 20750 62468 20802
rect 62188 20748 62468 20750
rect 64652 20916 64708 20926
rect 62188 20738 62244 20748
rect 64652 20578 64708 20860
rect 64652 20526 64654 20578
rect 64706 20526 64708 20578
rect 64652 20514 64708 20526
rect 62768 20412 63448 20422
rect 62824 20356 62872 20412
rect 62928 20410 62976 20412
rect 63032 20410 63080 20412
rect 62948 20358 62976 20410
rect 63072 20358 63080 20410
rect 62928 20356 62976 20358
rect 63032 20356 63080 20358
rect 63136 20410 63184 20412
rect 63240 20410 63288 20412
rect 63136 20358 63144 20410
rect 63240 20358 63268 20410
rect 63136 20356 63184 20358
rect 63240 20356 63288 20358
rect 63344 20356 63392 20412
rect 62768 20346 63448 20356
rect 62768 18844 63448 18854
rect 62824 18788 62872 18844
rect 62928 18842 62976 18844
rect 63032 18842 63080 18844
rect 62948 18790 62976 18842
rect 63072 18790 63080 18842
rect 62928 18788 62976 18790
rect 63032 18788 63080 18790
rect 63136 18842 63184 18844
rect 63240 18842 63288 18844
rect 63136 18790 63144 18842
rect 63240 18790 63268 18842
rect 63136 18788 63184 18790
rect 63240 18788 63288 18790
rect 63344 18788 63392 18844
rect 62768 18778 63448 18788
rect 62768 17276 63448 17286
rect 62824 17220 62872 17276
rect 62928 17274 62976 17276
rect 63032 17274 63080 17276
rect 62948 17222 62976 17274
rect 63072 17222 63080 17274
rect 62928 17220 62976 17222
rect 63032 17220 63080 17222
rect 63136 17274 63184 17276
rect 63240 17274 63288 17276
rect 63136 17222 63144 17274
rect 63240 17222 63268 17274
rect 63136 17220 63184 17222
rect 63240 17220 63288 17222
rect 63344 17220 63392 17276
rect 62768 17210 63448 17220
rect 62768 15708 63448 15718
rect 62824 15652 62872 15708
rect 62928 15706 62976 15708
rect 63032 15706 63080 15708
rect 62948 15654 62976 15706
rect 63072 15654 63080 15706
rect 62928 15652 62976 15654
rect 63032 15652 63080 15654
rect 63136 15706 63184 15708
rect 63240 15706 63288 15708
rect 63136 15654 63144 15706
rect 63240 15654 63268 15706
rect 63136 15652 63184 15654
rect 63240 15652 63288 15654
rect 63344 15652 63392 15708
rect 62768 15642 63448 15652
rect 65436 15148 65492 26012
rect 65772 25620 65828 27804
rect 66220 27300 66276 27310
rect 66332 27300 66388 27916
rect 66220 27298 66332 27300
rect 66220 27246 66222 27298
rect 66274 27246 66332 27298
rect 66220 27244 66332 27246
rect 66220 27234 66276 27244
rect 66332 27206 66388 27244
rect 66780 26740 66836 28252
rect 67228 28754 67396 28756
rect 67228 28702 67342 28754
rect 67394 28702 67396 28754
rect 67228 28700 67396 28702
rect 67228 27748 67284 28700
rect 67340 28690 67396 28700
rect 68348 28756 68404 29260
rect 68348 28690 68404 28700
rect 68236 28644 68292 28654
rect 67788 28642 68292 28644
rect 67788 28590 68238 28642
rect 68290 28590 68292 28642
rect 67788 28588 68292 28590
rect 67788 28530 67844 28588
rect 68236 28578 68292 28588
rect 67788 28478 67790 28530
rect 67842 28478 67844 28530
rect 67788 28466 67844 28478
rect 66780 26674 66836 26684
rect 67004 27692 67284 27748
rect 65772 25526 65828 25564
rect 66668 26402 66724 26414
rect 66668 26350 66670 26402
rect 66722 26350 66724 26402
rect 66332 24948 66388 24958
rect 66332 24854 66388 24892
rect 66668 24722 66724 26350
rect 66668 24670 66670 24722
rect 66722 24670 66724 24722
rect 66668 24658 66724 24670
rect 67004 24948 67060 27692
rect 67268 27468 67948 27478
rect 67324 27412 67372 27468
rect 67428 27466 67476 27468
rect 67532 27466 67580 27468
rect 67448 27414 67476 27466
rect 67572 27414 67580 27466
rect 67428 27412 67476 27414
rect 67532 27412 67580 27414
rect 67636 27466 67684 27468
rect 67740 27466 67788 27468
rect 67636 27414 67644 27466
rect 67740 27414 67768 27466
rect 67636 27412 67684 27414
rect 67740 27412 67788 27414
rect 67844 27412 67892 27468
rect 67268 27402 67948 27412
rect 67228 27300 67284 27310
rect 67228 27074 67284 27244
rect 67228 27022 67230 27074
rect 67282 27022 67284 27074
rect 67228 27010 67284 27022
rect 67564 27300 67620 27310
rect 67564 26962 67620 27244
rect 67564 26910 67566 26962
rect 67618 26910 67620 26962
rect 67564 26898 67620 26910
rect 68460 26908 68516 34636
rect 71148 34598 71204 34636
rect 71768 34524 72448 34534
rect 71824 34468 71872 34524
rect 71928 34522 71976 34524
rect 72032 34522 72080 34524
rect 71948 34470 71976 34522
rect 72072 34470 72080 34522
rect 71928 34468 71976 34470
rect 72032 34468 72080 34470
rect 72136 34522 72184 34524
rect 72240 34522 72288 34524
rect 72136 34470 72144 34522
rect 72240 34470 72268 34522
rect 72136 34468 72184 34470
rect 72240 34468 72288 34470
rect 72344 34468 72392 34524
rect 71768 34458 72448 34468
rect 72492 34356 72548 34366
rect 72716 34356 72772 34862
rect 72828 34356 72884 34366
rect 72716 34354 72884 34356
rect 72716 34302 72830 34354
rect 72882 34302 72884 34354
rect 72716 34300 72884 34302
rect 72492 34132 72548 34300
rect 72828 34290 72884 34300
rect 72716 34132 72772 34142
rect 72492 34130 72772 34132
rect 72492 34078 72718 34130
rect 72770 34078 72772 34130
rect 72492 34076 72772 34078
rect 72716 34066 72772 34076
rect 72940 34130 72996 34142
rect 72940 34078 72942 34130
rect 72994 34078 72996 34130
rect 72940 33908 72996 34078
rect 73388 34132 73444 34142
rect 73388 34038 73444 34076
rect 73724 34018 73780 35868
rect 74732 35476 74788 35486
rect 74508 34356 74564 34366
rect 74508 34262 74564 34300
rect 74284 34132 74340 34142
rect 74620 34132 74676 34142
rect 74284 34038 74340 34076
rect 74508 34130 74676 34132
rect 74508 34078 74622 34130
rect 74674 34078 74676 34130
rect 74508 34076 74676 34078
rect 74732 34132 74788 35420
rect 74844 34244 74900 38780
rect 74956 37828 75012 40796
rect 75068 40292 75124 41132
rect 75068 38668 75124 40236
rect 75292 39060 75348 43260
rect 75404 42532 75460 42542
rect 75404 42438 75460 42476
rect 75740 41972 75796 41982
rect 75628 40964 75684 41002
rect 75404 39060 75460 39070
rect 75292 39004 75404 39060
rect 75068 38612 75348 38668
rect 74956 37734 75012 37772
rect 75292 38610 75348 38612
rect 75292 38558 75294 38610
rect 75346 38558 75348 38610
rect 75292 37490 75348 38558
rect 75404 38276 75460 39004
rect 75404 38162 75460 38220
rect 75404 38110 75406 38162
rect 75458 38110 75460 38162
rect 75404 38098 75460 38110
rect 75628 38052 75684 40908
rect 75628 37986 75684 37996
rect 75292 37438 75294 37490
rect 75346 37438 75348 37490
rect 75292 37156 75348 37438
rect 75292 37090 75348 37100
rect 75740 36932 75796 41916
rect 75852 40964 75908 45836
rect 75964 41858 76020 48076
rect 76972 48132 77028 48190
rect 77420 48244 77476 48254
rect 77420 48150 77476 48188
rect 76972 48066 77028 48076
rect 77308 48130 77364 48142
rect 77308 48078 77310 48130
rect 77362 48078 77364 48130
rect 76268 47852 76948 47862
rect 76324 47796 76372 47852
rect 76428 47850 76476 47852
rect 76532 47850 76580 47852
rect 76448 47798 76476 47850
rect 76572 47798 76580 47850
rect 76428 47796 76476 47798
rect 76532 47796 76580 47798
rect 76636 47850 76684 47852
rect 76740 47850 76788 47852
rect 76636 47798 76644 47850
rect 76740 47798 76768 47850
rect 76636 47796 76684 47798
rect 76740 47796 76788 47798
rect 76844 47796 76892 47852
rect 76268 47786 76948 47796
rect 77308 47348 77364 48078
rect 77420 48020 77476 48030
rect 77420 47570 77476 47964
rect 77420 47518 77422 47570
rect 77474 47518 77476 47570
rect 77420 47506 77476 47518
rect 77308 47282 77364 47292
rect 76860 46788 76916 46798
rect 76636 46786 76916 46788
rect 76636 46734 76862 46786
rect 76914 46734 76916 46786
rect 76636 46732 76916 46734
rect 76636 46564 76692 46732
rect 76860 46722 76916 46732
rect 77084 46676 77140 46686
rect 77084 46674 77252 46676
rect 77084 46622 77086 46674
rect 77138 46622 77252 46674
rect 77084 46620 77252 46622
rect 77084 46610 77140 46620
rect 76636 46470 76692 46508
rect 76268 46284 76948 46294
rect 76324 46228 76372 46284
rect 76428 46282 76476 46284
rect 76532 46282 76580 46284
rect 76448 46230 76476 46282
rect 76572 46230 76580 46282
rect 76428 46228 76476 46230
rect 76532 46228 76580 46230
rect 76636 46282 76684 46284
rect 76740 46282 76788 46284
rect 76636 46230 76644 46282
rect 76740 46230 76768 46282
rect 76636 46228 76684 46230
rect 76740 46228 76788 46230
rect 76844 46228 76892 46284
rect 76268 46218 76948 46228
rect 77084 45892 77140 45902
rect 77084 45798 77140 45836
rect 77196 45444 77252 46620
rect 77644 46674 77700 46686
rect 77644 46622 77646 46674
rect 77698 46622 77700 46674
rect 77308 45892 77364 45902
rect 77308 45798 77364 45836
rect 77644 45890 77700 46622
rect 77980 46004 78036 49084
rect 78876 49140 78932 49150
rect 78428 48916 78484 48926
rect 78316 48356 78372 48366
rect 78316 48262 78372 48300
rect 78092 48242 78148 48254
rect 78092 48190 78094 48242
rect 78146 48190 78148 48242
rect 78092 48020 78148 48190
rect 78148 47964 78260 48020
rect 78092 47954 78148 47964
rect 78092 47348 78148 47358
rect 78092 46674 78148 47292
rect 78092 46622 78094 46674
rect 78146 46622 78148 46674
rect 78092 46610 78148 46622
rect 77644 45838 77646 45890
rect 77698 45838 77700 45890
rect 77644 45826 77700 45838
rect 77756 46002 78036 46004
rect 77756 45950 77982 46002
rect 78034 45950 78036 46002
rect 77756 45948 78036 45950
rect 77420 45668 77476 45678
rect 77420 45574 77476 45612
rect 77084 45388 77252 45444
rect 76748 45220 76804 45230
rect 76748 45126 76804 45164
rect 76300 44996 76356 45006
rect 76300 44902 76356 44940
rect 76268 44716 76948 44726
rect 76324 44660 76372 44716
rect 76428 44714 76476 44716
rect 76532 44714 76580 44716
rect 76448 44662 76476 44714
rect 76572 44662 76580 44714
rect 76428 44660 76476 44662
rect 76532 44660 76580 44662
rect 76636 44714 76684 44716
rect 76740 44714 76788 44716
rect 76636 44662 76644 44714
rect 76740 44662 76768 44714
rect 76636 44660 76684 44662
rect 76740 44660 76788 44662
rect 76844 44660 76892 44716
rect 76268 44650 76948 44660
rect 76636 44100 76692 44110
rect 76636 44006 76692 44044
rect 77084 43762 77140 45388
rect 77756 45220 77812 45948
rect 77980 45938 78036 45948
rect 77812 45164 78036 45220
rect 77756 45126 77812 45164
rect 77532 45106 77588 45118
rect 77532 45054 77534 45106
rect 77586 45054 77588 45106
rect 77532 44996 77588 45054
rect 77308 44322 77364 44334
rect 77308 44270 77310 44322
rect 77362 44270 77364 44322
rect 77308 44100 77364 44270
rect 77308 44034 77364 44044
rect 77420 44210 77476 44222
rect 77420 44158 77422 44210
rect 77474 44158 77476 44210
rect 77084 43710 77086 43762
rect 77138 43710 77140 43762
rect 77084 43698 77140 43710
rect 76972 43652 77028 43662
rect 76972 43558 77028 43596
rect 77420 43652 77476 44158
rect 77420 43586 77476 43596
rect 76636 43538 76692 43550
rect 76636 43486 76638 43538
rect 76690 43486 76692 43538
rect 76636 43316 76692 43486
rect 77196 43538 77252 43550
rect 77196 43486 77198 43538
rect 77250 43486 77252 43538
rect 77196 43316 77252 43486
rect 76636 43260 77140 43316
rect 76268 43148 76948 43158
rect 76324 43092 76372 43148
rect 76428 43146 76476 43148
rect 76532 43146 76580 43148
rect 76448 43094 76476 43146
rect 76572 43094 76580 43146
rect 76428 43092 76476 43094
rect 76532 43092 76580 43094
rect 76636 43146 76684 43148
rect 76740 43146 76788 43148
rect 76636 43094 76644 43146
rect 76740 43094 76768 43146
rect 76636 43092 76684 43094
rect 76740 43092 76788 43094
rect 76844 43092 76892 43148
rect 76268 43082 76948 43092
rect 77084 42532 77140 43260
rect 77196 43250 77252 43260
rect 77532 43092 77588 44940
rect 77980 44546 78036 45164
rect 77980 44494 77982 44546
rect 78034 44494 78036 44546
rect 77980 44482 78036 44494
rect 76860 41972 76916 41982
rect 76860 41878 76916 41916
rect 75964 41806 75966 41858
rect 76018 41806 76020 41858
rect 75964 41188 76020 41806
rect 76412 41860 76468 41870
rect 76412 41766 76468 41804
rect 76268 41580 76948 41590
rect 76324 41524 76372 41580
rect 76428 41578 76476 41580
rect 76532 41578 76580 41580
rect 76448 41526 76476 41578
rect 76572 41526 76580 41578
rect 76428 41524 76476 41526
rect 76532 41524 76580 41526
rect 76636 41578 76684 41580
rect 76740 41578 76788 41580
rect 76636 41526 76644 41578
rect 76740 41526 76768 41578
rect 76636 41524 76684 41526
rect 76740 41524 76788 41526
rect 76844 41524 76892 41580
rect 76268 41514 76948 41524
rect 76748 41412 76804 41422
rect 76188 41188 76244 41198
rect 75964 41132 76188 41188
rect 76188 41122 76244 41132
rect 76748 41186 76804 41356
rect 76860 41300 76916 41310
rect 76860 41298 77028 41300
rect 76860 41246 76862 41298
rect 76914 41246 77028 41298
rect 76860 41244 77028 41246
rect 76860 41234 76916 41244
rect 76748 41134 76750 41186
rect 76802 41134 76804 41186
rect 76748 41122 76804 41134
rect 76300 41076 76356 41086
rect 76300 40982 76356 41020
rect 76524 41074 76580 41086
rect 76524 41022 76526 41074
rect 76578 41022 76580 41074
rect 76412 40964 76468 40974
rect 76524 40964 76580 41022
rect 76860 41076 76916 41086
rect 76860 40982 76916 41020
rect 75852 40908 76132 40964
rect 76076 40404 76132 40908
rect 76468 40908 76580 40964
rect 76412 40898 76468 40908
rect 76300 40852 76356 40862
rect 76300 40628 76356 40796
rect 76300 40626 76580 40628
rect 76300 40574 76302 40626
rect 76354 40574 76580 40626
rect 76300 40572 76580 40574
rect 76300 40562 76356 40572
rect 76524 40514 76580 40572
rect 76524 40462 76526 40514
rect 76578 40462 76580 40514
rect 76524 40450 76580 40462
rect 75964 40348 76132 40404
rect 76636 40402 76692 40414
rect 76636 40350 76638 40402
rect 76690 40350 76692 40402
rect 75964 39844 76020 40348
rect 76636 40292 76692 40350
rect 76972 40404 77028 41244
rect 76972 40338 77028 40348
rect 75964 39778 76020 39788
rect 76076 40236 76692 40292
rect 76076 38274 76132 40236
rect 76268 40012 76948 40022
rect 76324 39956 76372 40012
rect 76428 40010 76476 40012
rect 76532 40010 76580 40012
rect 76448 39958 76476 40010
rect 76572 39958 76580 40010
rect 76428 39956 76476 39958
rect 76532 39956 76580 39958
rect 76636 40010 76684 40012
rect 76740 40010 76788 40012
rect 76636 39958 76644 40010
rect 76740 39958 76768 40010
rect 76636 39956 76684 39958
rect 76740 39956 76788 39958
rect 76844 39956 76892 40012
rect 76268 39946 76948 39956
rect 76412 38948 76468 38958
rect 77084 38948 77140 42476
rect 77196 43036 77588 43092
rect 77196 39060 77252 43036
rect 77756 42644 77812 42654
rect 77532 42642 77812 42644
rect 77532 42590 77758 42642
rect 77810 42590 77812 42642
rect 77532 42588 77812 42590
rect 77532 42194 77588 42588
rect 77756 42578 77812 42588
rect 77532 42142 77534 42194
rect 77586 42142 77588 42194
rect 77532 42130 77588 42142
rect 78092 42530 78148 42542
rect 78092 42478 78094 42530
rect 78146 42478 78148 42530
rect 77980 42084 78036 42094
rect 77868 41860 77924 41870
rect 77868 41766 77924 41804
rect 77980 41186 78036 42028
rect 77980 41134 77982 41186
rect 78034 41134 78036 41186
rect 77980 41122 78036 41134
rect 78092 41188 78148 42478
rect 78204 42082 78260 47964
rect 78428 46786 78484 48860
rect 78876 48242 78932 49084
rect 79772 49138 79828 50372
rect 86716 50370 86884 50372
rect 86716 50318 86830 50370
rect 86882 50318 86884 50370
rect 86716 50316 86884 50318
rect 80768 50204 81448 50214
rect 80824 50148 80872 50204
rect 80928 50202 80976 50204
rect 81032 50202 81080 50204
rect 80948 50150 80976 50202
rect 81072 50150 81080 50202
rect 80928 50148 80976 50150
rect 81032 50148 81080 50150
rect 81136 50202 81184 50204
rect 81240 50202 81288 50204
rect 81136 50150 81144 50202
rect 81240 50150 81268 50202
rect 81136 50148 81184 50150
rect 81240 50148 81288 50150
rect 81344 50148 81392 50204
rect 80768 50138 81448 50148
rect 86268 49922 86324 49934
rect 86268 49870 86270 49922
rect 86322 49870 86324 49922
rect 86044 49810 86100 49822
rect 86044 49758 86046 49810
rect 86098 49758 86100 49810
rect 85268 49420 85948 49430
rect 85324 49364 85372 49420
rect 85428 49418 85476 49420
rect 85532 49418 85580 49420
rect 85448 49366 85476 49418
rect 85572 49366 85580 49418
rect 85428 49364 85476 49366
rect 85532 49364 85580 49366
rect 85636 49418 85684 49420
rect 85740 49418 85788 49420
rect 85636 49366 85644 49418
rect 85740 49366 85768 49418
rect 85636 49364 85684 49366
rect 85740 49364 85788 49366
rect 85844 49364 85892 49420
rect 85268 49354 85948 49364
rect 86044 49252 86100 49758
rect 86156 49252 86212 49262
rect 86044 49250 86212 49252
rect 86044 49198 86158 49250
rect 86210 49198 86212 49250
rect 86044 49196 86212 49198
rect 86156 49186 86212 49196
rect 79772 49086 79774 49138
rect 79826 49086 79828 49138
rect 79772 49074 79828 49086
rect 85148 49026 85204 49038
rect 85148 48974 85150 49026
rect 85202 48974 85204 49026
rect 85036 48916 85092 48926
rect 85036 48822 85092 48860
rect 80220 48802 80276 48814
rect 80220 48750 80222 48802
rect 80274 48750 80276 48802
rect 78876 48190 78878 48242
rect 78930 48190 78932 48242
rect 78876 48178 78932 48190
rect 79548 48244 79604 48254
rect 79212 48018 79268 48030
rect 79212 47966 79214 48018
rect 79266 47966 79268 48018
rect 79212 47458 79268 47966
rect 79212 47406 79214 47458
rect 79266 47406 79268 47458
rect 79212 47394 79268 47406
rect 79548 47346 79604 48188
rect 80220 48242 80276 48750
rect 84700 48802 84756 48814
rect 84700 48750 84702 48802
rect 84754 48750 84756 48802
rect 84700 48692 84756 48750
rect 85148 48692 85204 48974
rect 85820 49028 85876 49038
rect 85820 48934 85876 48972
rect 86268 48804 86324 49870
rect 86716 49026 86772 50316
rect 86828 50306 86884 50316
rect 89768 50204 90448 50214
rect 89824 50148 89872 50204
rect 89928 50202 89976 50204
rect 90032 50202 90080 50204
rect 89948 50150 89976 50202
rect 90072 50150 90080 50202
rect 89928 50148 89976 50150
rect 90032 50148 90080 50150
rect 90136 50202 90184 50204
rect 90240 50202 90288 50204
rect 90136 50150 90144 50202
rect 90240 50150 90268 50202
rect 90136 50148 90184 50150
rect 90240 50148 90288 50150
rect 90344 50148 90392 50204
rect 89768 50138 90448 50148
rect 90524 49700 90580 49710
rect 90524 49138 90580 49644
rect 90748 49252 90804 51326
rect 94268 50988 94948 50998
rect 94324 50932 94372 50988
rect 94428 50986 94476 50988
rect 94532 50986 94580 50988
rect 94448 50934 94476 50986
rect 94572 50934 94580 50986
rect 94428 50932 94476 50934
rect 94532 50932 94580 50934
rect 94636 50986 94684 50988
rect 94740 50986 94788 50988
rect 94636 50934 94644 50986
rect 94740 50934 94768 50986
rect 94636 50932 94684 50934
rect 94740 50932 94788 50934
rect 94844 50932 94892 50988
rect 94268 50922 94948 50932
rect 96236 50482 96292 50494
rect 96236 50430 96238 50482
rect 96290 50430 96292 50482
rect 92428 49700 92484 49710
rect 92428 49606 92484 49644
rect 95452 49700 95508 49710
rect 94268 49420 94948 49430
rect 94324 49364 94372 49420
rect 94428 49418 94476 49420
rect 94532 49418 94580 49420
rect 94448 49366 94476 49418
rect 94572 49366 94580 49418
rect 94428 49364 94476 49366
rect 94532 49364 94580 49366
rect 94636 49418 94684 49420
rect 94740 49418 94788 49420
rect 94636 49366 94644 49418
rect 94740 49366 94768 49418
rect 94636 49364 94684 49366
rect 94740 49364 94788 49366
rect 94844 49364 94892 49420
rect 94268 49354 94948 49364
rect 90748 49186 90804 49196
rect 90524 49086 90526 49138
rect 90578 49086 90580 49138
rect 86716 48974 86718 49026
rect 86770 48974 86772 49026
rect 86716 48962 86772 48974
rect 87052 49026 87108 49038
rect 87052 48974 87054 49026
rect 87106 48974 87108 49026
rect 87052 48804 87108 48974
rect 90188 49028 90244 49038
rect 90188 48934 90244 48972
rect 86268 48748 87108 48804
rect 89628 48916 89684 48926
rect 89628 48802 89684 48860
rect 90524 48916 90580 49086
rect 92540 49028 92596 49038
rect 93100 49028 93156 49038
rect 90524 48850 90580 48860
rect 92316 49026 92596 49028
rect 92316 48974 92542 49026
rect 92594 48974 92596 49026
rect 92316 48972 92596 48974
rect 92316 48914 92372 48972
rect 92540 48962 92596 48972
rect 92876 49026 93156 49028
rect 92876 48974 93102 49026
rect 93154 48974 93156 49026
rect 92876 48972 93156 48974
rect 92316 48862 92318 48914
rect 92370 48862 92372 48914
rect 92316 48850 92372 48862
rect 89628 48750 89630 48802
rect 89682 48750 89684 48802
rect 80768 48636 81448 48646
rect 84700 48636 85204 48692
rect 80824 48580 80872 48636
rect 80928 48634 80976 48636
rect 81032 48634 81080 48636
rect 80948 48582 80976 48634
rect 81072 48582 81080 48634
rect 80928 48580 80976 48582
rect 81032 48580 81080 48582
rect 81136 48634 81184 48636
rect 81240 48634 81288 48636
rect 81136 48582 81144 48634
rect 81240 48582 81268 48634
rect 81136 48580 81184 48582
rect 81240 48580 81288 48582
rect 81344 48580 81392 48636
rect 80768 48570 81448 48580
rect 83132 48468 83188 48478
rect 83132 48466 83524 48468
rect 83132 48414 83134 48466
rect 83186 48414 83524 48466
rect 83132 48412 83524 48414
rect 83132 48402 83188 48412
rect 80220 48190 80222 48242
rect 80274 48190 80276 48242
rect 80220 48178 80276 48190
rect 80556 48244 80612 48254
rect 80556 48150 80612 48188
rect 79548 47294 79550 47346
rect 79602 47294 79604 47346
rect 79548 47282 79604 47294
rect 80768 47068 81448 47078
rect 80824 47012 80872 47068
rect 80928 47066 80976 47068
rect 81032 47066 81080 47068
rect 80948 47014 80976 47066
rect 81072 47014 81080 47066
rect 80928 47012 80976 47014
rect 81032 47012 81080 47014
rect 81136 47066 81184 47068
rect 81240 47066 81288 47068
rect 81136 47014 81144 47066
rect 81240 47014 81268 47066
rect 81136 47012 81184 47014
rect 81240 47012 81288 47014
rect 81344 47012 81392 47068
rect 80768 47002 81448 47012
rect 78428 46734 78430 46786
rect 78482 46734 78484 46786
rect 78428 46722 78484 46734
rect 79100 46004 79156 46014
rect 79100 45910 79156 45948
rect 79548 46004 79604 46014
rect 78652 45780 78708 45790
rect 78316 45668 78372 45678
rect 78316 45106 78372 45612
rect 78652 45330 78708 45724
rect 79324 45780 79380 45790
rect 79324 45686 79380 45724
rect 78652 45278 78654 45330
rect 78706 45278 78708 45330
rect 78652 45266 78708 45278
rect 78316 45054 78318 45106
rect 78370 45054 78372 45106
rect 78316 45042 78372 45054
rect 78316 44212 78372 44222
rect 78316 44118 78372 44156
rect 78204 42030 78206 42082
rect 78258 42030 78260 42082
rect 78204 41972 78260 42030
rect 78204 41906 78260 41916
rect 78652 42082 78708 42094
rect 78652 42030 78654 42082
rect 78706 42030 78708 42082
rect 78652 41412 78708 42030
rect 79100 42084 79156 42094
rect 79100 41990 79156 42028
rect 78652 41346 78708 41356
rect 78428 41188 78484 41198
rect 78092 41186 78484 41188
rect 78092 41134 78430 41186
rect 78482 41134 78484 41186
rect 78092 41132 78484 41134
rect 78428 41122 78484 41132
rect 77644 40964 77700 40974
rect 77644 40870 77700 40908
rect 78540 40964 78596 40974
rect 77420 40404 77476 40414
rect 77756 40404 77812 40414
rect 77420 40402 77700 40404
rect 77420 40350 77422 40402
rect 77474 40350 77700 40402
rect 77420 40348 77700 40350
rect 77420 40338 77476 40348
rect 77196 38994 77252 39004
rect 77308 39058 77364 39070
rect 77308 39006 77310 39058
rect 77362 39006 77364 39058
rect 76412 38946 77140 38948
rect 76412 38894 76414 38946
rect 76466 38894 77140 38946
rect 76412 38892 77140 38894
rect 76412 38882 76468 38892
rect 76860 38724 76916 38762
rect 76860 38658 76916 38668
rect 76972 38668 77028 38892
rect 77196 38834 77252 38846
rect 77196 38782 77198 38834
rect 77250 38782 77252 38834
rect 77196 38724 77252 38782
rect 76972 38612 77140 38668
rect 77196 38658 77252 38668
rect 76268 38444 76948 38454
rect 76324 38388 76372 38444
rect 76428 38442 76476 38444
rect 76532 38442 76580 38444
rect 76448 38390 76476 38442
rect 76572 38390 76580 38442
rect 76428 38388 76476 38390
rect 76532 38388 76580 38390
rect 76636 38442 76684 38444
rect 76740 38442 76788 38444
rect 76636 38390 76644 38442
rect 76740 38390 76768 38442
rect 76636 38388 76684 38390
rect 76740 38388 76788 38390
rect 76844 38388 76892 38444
rect 76268 38378 76948 38388
rect 76076 38222 76078 38274
rect 76130 38222 76132 38274
rect 76076 38210 76132 38222
rect 76188 38050 76244 38062
rect 76188 37998 76190 38050
rect 76242 37998 76244 38050
rect 76188 37828 76244 37998
rect 76972 38052 77028 38062
rect 77084 38052 77140 38612
rect 76972 38050 77140 38052
rect 76972 37998 76974 38050
rect 77026 37998 77140 38050
rect 76972 37996 77140 37998
rect 77196 38276 77252 38286
rect 77308 38276 77364 39006
rect 77420 38948 77476 38958
rect 77420 38668 77476 38892
rect 77532 38948 77588 38958
rect 77644 38948 77700 40348
rect 77756 40310 77812 40348
rect 78092 40292 78148 40302
rect 78092 40198 78148 40236
rect 77756 39844 77812 39854
rect 77812 39788 77924 39844
rect 77756 39778 77812 39788
rect 77532 38946 77700 38948
rect 77532 38894 77534 38946
rect 77586 38894 77700 38946
rect 77532 38892 77700 38894
rect 77756 39060 77812 39070
rect 77532 38882 77588 38892
rect 77420 38612 77700 38668
rect 77308 38220 77588 38276
rect 77196 38052 77252 38220
rect 77420 38052 77476 38062
rect 77196 38050 77476 38052
rect 77196 37998 77422 38050
rect 77474 37998 77476 38050
rect 77196 37996 77476 37998
rect 76972 37986 77028 37996
rect 77420 37986 77476 37996
rect 76188 37762 76244 37772
rect 76300 37940 76356 37950
rect 75852 37492 75908 37502
rect 76300 37492 76356 37884
rect 77532 37828 77588 38220
rect 77532 37762 77588 37772
rect 77644 37604 77700 38612
rect 77532 37548 77700 37604
rect 75852 37490 76356 37492
rect 75852 37438 75854 37490
rect 75906 37438 76356 37490
rect 75852 37436 76356 37438
rect 76860 37492 76916 37502
rect 75852 37426 75908 37436
rect 76860 37398 76916 37436
rect 77532 37492 77588 37548
rect 77532 37266 77588 37436
rect 77532 37214 77534 37266
rect 77586 37214 77588 37266
rect 77532 37202 77588 37214
rect 77644 37378 77700 37390
rect 77644 37326 77646 37378
rect 77698 37326 77700 37378
rect 76188 37156 76244 37166
rect 76188 37062 76244 37100
rect 77644 37044 77700 37326
rect 77196 36988 77700 37044
rect 77756 37156 77812 39004
rect 77868 39058 77924 39788
rect 77868 39006 77870 39058
rect 77922 39006 77924 39058
rect 77868 38724 77924 39006
rect 78540 39060 78596 40908
rect 78540 38966 78596 39004
rect 78988 38946 79044 38958
rect 78988 38894 78990 38946
rect 79042 38894 79044 38946
rect 78988 38668 79044 38894
rect 77868 38658 77924 38668
rect 78876 38612 79044 38668
rect 79548 38724 79604 45948
rect 82796 46004 82852 46014
rect 79884 45892 79940 45902
rect 80444 45892 80500 45902
rect 79884 45798 79940 45836
rect 79996 45890 80500 45892
rect 79996 45838 80446 45890
rect 80498 45838 80500 45890
rect 79996 45836 80500 45838
rect 79660 45668 79716 45678
rect 79996 45668 80052 45836
rect 80444 45826 80500 45836
rect 80556 45892 80612 45902
rect 79660 45666 80052 45668
rect 79660 45614 79662 45666
rect 79714 45614 80052 45666
rect 79660 45612 80052 45614
rect 79660 45602 79716 45612
rect 80556 45332 80612 45836
rect 82796 45778 82852 45948
rect 82796 45726 82798 45778
rect 82850 45726 82852 45778
rect 82796 45714 82852 45726
rect 80768 45500 81448 45510
rect 80824 45444 80872 45500
rect 80928 45498 80976 45500
rect 81032 45498 81080 45500
rect 80948 45446 80976 45498
rect 81072 45446 81080 45498
rect 80928 45444 80976 45446
rect 81032 45444 81080 45446
rect 81136 45498 81184 45500
rect 81240 45498 81288 45500
rect 81136 45446 81144 45498
rect 81240 45446 81268 45498
rect 81136 45444 81184 45446
rect 81240 45444 81288 45446
rect 81344 45444 81392 45500
rect 80768 45434 81448 45444
rect 81004 45332 81060 45342
rect 80556 45330 81060 45332
rect 80556 45278 81006 45330
rect 81058 45278 81060 45330
rect 80556 45276 81060 45278
rect 81004 45266 81060 45276
rect 79772 44212 79828 44222
rect 79772 44118 79828 44156
rect 80108 44098 80164 44110
rect 81116 44100 81172 44110
rect 80108 44046 80110 44098
rect 80162 44046 80164 44098
rect 80108 43764 80164 44046
rect 80556 44098 81172 44100
rect 80556 44046 81118 44098
rect 81170 44046 81172 44098
rect 80556 44044 81172 44046
rect 80556 43764 80612 44044
rect 81116 44034 81172 44044
rect 80768 43932 81448 43942
rect 80824 43876 80872 43932
rect 80928 43930 80976 43932
rect 81032 43930 81080 43932
rect 80948 43878 80976 43930
rect 81072 43878 81080 43930
rect 80928 43876 80976 43878
rect 81032 43876 81080 43878
rect 81136 43930 81184 43932
rect 81240 43930 81288 43932
rect 81136 43878 81144 43930
rect 81240 43878 81268 43930
rect 81136 43876 81184 43878
rect 81240 43876 81288 43878
rect 81344 43876 81392 43932
rect 80768 43866 81448 43876
rect 81340 43764 81396 43774
rect 80556 43708 80836 43764
rect 80108 43698 80164 43708
rect 80780 43538 80836 43708
rect 80780 43486 80782 43538
rect 80834 43486 80836 43538
rect 80780 43474 80836 43486
rect 81340 43538 81396 43708
rect 81340 43486 81342 43538
rect 81394 43486 81396 43538
rect 81340 43474 81396 43486
rect 83468 43708 83524 48412
rect 83692 48356 83748 48366
rect 83692 48262 83748 48300
rect 85148 48244 85204 48636
rect 85036 46900 85092 46910
rect 85148 46900 85204 48188
rect 85268 47852 85948 47862
rect 85324 47796 85372 47852
rect 85428 47850 85476 47852
rect 85532 47850 85580 47852
rect 85448 47798 85476 47850
rect 85572 47798 85580 47850
rect 85428 47796 85476 47798
rect 85532 47796 85580 47798
rect 85636 47850 85684 47852
rect 85740 47850 85788 47852
rect 85636 47798 85644 47850
rect 85740 47798 85768 47850
rect 85636 47796 85684 47798
rect 85740 47796 85788 47798
rect 85844 47796 85892 47852
rect 85268 47786 85948 47796
rect 85036 46898 85204 46900
rect 85036 46846 85038 46898
rect 85090 46846 85204 46898
rect 85036 46844 85204 46846
rect 86268 47516 86884 47572
rect 85036 46834 85092 46844
rect 85484 46562 85540 46574
rect 85484 46510 85486 46562
rect 85538 46510 85540 46562
rect 85484 46452 85540 46510
rect 85484 46386 85540 46396
rect 85268 46284 85948 46294
rect 85324 46228 85372 46284
rect 85428 46282 85476 46284
rect 85532 46282 85580 46284
rect 85448 46230 85476 46282
rect 85572 46230 85580 46282
rect 85428 46228 85476 46230
rect 85532 46228 85580 46230
rect 85636 46282 85684 46284
rect 85740 46282 85788 46284
rect 85636 46230 85644 46282
rect 85740 46230 85768 46282
rect 85636 46228 85684 46230
rect 85740 46228 85788 46230
rect 85844 46228 85892 46284
rect 85268 46218 85948 46228
rect 86156 45892 86212 45902
rect 86268 45892 86324 47516
rect 86828 47460 86884 47516
rect 86828 47404 87108 47460
rect 86716 47348 86772 47358
rect 86716 47346 86996 47348
rect 86716 47294 86718 47346
rect 86770 47294 86996 47346
rect 86716 47292 86996 47294
rect 86716 47282 86772 47292
rect 86380 47236 86436 47246
rect 86380 47234 86548 47236
rect 86380 47182 86382 47234
rect 86434 47182 86548 47234
rect 86380 47180 86548 47182
rect 86380 47170 86436 47180
rect 86380 46786 86436 46798
rect 86380 46734 86382 46786
rect 86434 46734 86436 46786
rect 86380 46452 86436 46734
rect 86380 46386 86436 46396
rect 86156 45890 86324 45892
rect 86156 45838 86158 45890
rect 86210 45838 86324 45890
rect 86156 45836 86324 45838
rect 86492 45890 86548 47180
rect 86940 47012 86996 47292
rect 87052 47346 87108 47404
rect 87052 47294 87054 47346
rect 87106 47294 87108 47346
rect 87052 47282 87108 47294
rect 86940 46956 87332 47012
rect 87276 46898 87332 46956
rect 87276 46846 87278 46898
rect 87330 46846 87332 46898
rect 87276 46834 87332 46846
rect 89628 46900 89684 48750
rect 89768 48636 90448 48646
rect 89824 48580 89872 48636
rect 89928 48634 89976 48636
rect 90032 48634 90080 48636
rect 89948 48582 89976 48634
rect 90072 48582 90080 48634
rect 89928 48580 89976 48582
rect 90032 48580 90080 48582
rect 90136 48634 90184 48636
rect 90240 48634 90288 48636
rect 90136 48582 90144 48634
rect 90240 48582 90268 48634
rect 90136 48580 90184 48582
rect 90240 48580 90288 48582
rect 90344 48580 90392 48636
rect 89768 48570 90448 48580
rect 92540 48354 92596 48366
rect 92540 48302 92542 48354
rect 92594 48302 92596 48354
rect 91196 48244 91252 48254
rect 91084 48188 91196 48244
rect 89768 47068 90448 47078
rect 89824 47012 89872 47068
rect 89928 47066 89976 47068
rect 90032 47066 90080 47068
rect 89948 47014 89976 47066
rect 90072 47014 90080 47066
rect 89928 47012 89976 47014
rect 90032 47012 90080 47014
rect 90136 47066 90184 47068
rect 90240 47066 90288 47068
rect 90136 47014 90144 47066
rect 90240 47014 90268 47066
rect 90136 47012 90184 47014
rect 90240 47012 90288 47014
rect 90344 47012 90392 47068
rect 89768 47002 90448 47012
rect 89628 46844 90020 46900
rect 86492 45838 86494 45890
rect 86546 45838 86548 45890
rect 86156 45826 86212 45836
rect 86492 45826 86548 45838
rect 86716 46786 86772 46798
rect 86716 46734 86718 46786
rect 86770 46734 86772 46786
rect 83580 45668 83636 45678
rect 83580 45574 83636 45612
rect 86716 45220 86772 46734
rect 86940 46452 86996 46462
rect 86940 46358 86996 46396
rect 89628 46452 89684 46462
rect 89628 46114 89684 46396
rect 89628 46062 89630 46114
rect 89682 46062 89684 46114
rect 89628 45780 89684 46062
rect 89628 45714 89684 45724
rect 89964 46002 90020 46844
rect 89964 45950 89966 46002
rect 90018 45950 90020 46002
rect 89068 45668 89124 45678
rect 89068 45574 89124 45612
rect 89964 45668 90020 45950
rect 89964 45602 90020 45612
rect 89768 45500 90448 45510
rect 89824 45444 89872 45500
rect 89928 45498 89976 45500
rect 90032 45498 90080 45500
rect 89948 45446 89976 45498
rect 90072 45446 90080 45498
rect 89928 45444 89976 45446
rect 90032 45444 90080 45446
rect 90136 45498 90184 45500
rect 90240 45498 90288 45500
rect 90136 45446 90144 45498
rect 90240 45446 90268 45498
rect 90136 45444 90184 45446
rect 90240 45444 90288 45446
rect 90344 45444 90392 45500
rect 89768 45434 90448 45444
rect 86716 45154 86772 45164
rect 90636 45220 90692 45230
rect 91084 45220 91140 48188
rect 91196 48150 91252 48188
rect 92316 48244 92372 48254
rect 92316 48150 92372 48188
rect 91644 48130 91700 48142
rect 91644 48078 91646 48130
rect 91698 48078 91700 48130
rect 91644 47684 91700 48078
rect 91644 47618 91700 47628
rect 92540 47684 92596 48302
rect 92540 47618 92596 47628
rect 92652 47460 92708 47470
rect 92652 47366 92708 47404
rect 92876 47346 92932 48972
rect 93100 48962 93156 48972
rect 95452 48914 95508 49644
rect 95452 48862 95454 48914
rect 95506 48862 95508 48914
rect 95452 48850 95508 48862
rect 96236 48802 96292 50430
rect 96236 48750 96238 48802
rect 96290 48750 96292 48802
rect 93100 48692 93156 48702
rect 93100 48242 93156 48636
rect 96236 48692 96292 48750
rect 96236 48626 96292 48636
rect 96236 48244 96292 48254
rect 93100 48190 93102 48242
rect 93154 48190 93156 48242
rect 93100 48178 93156 48190
rect 96124 48242 96292 48244
rect 96124 48190 96238 48242
rect 96290 48190 96292 48242
rect 96124 48188 96292 48190
rect 93436 48018 93492 48030
rect 93436 47966 93438 48018
rect 93490 47966 93492 48018
rect 93436 47460 93492 47966
rect 94268 47852 94948 47862
rect 94324 47796 94372 47852
rect 94428 47850 94476 47852
rect 94532 47850 94580 47852
rect 94448 47798 94476 47850
rect 94572 47798 94580 47850
rect 94428 47796 94476 47798
rect 94532 47796 94580 47798
rect 94636 47850 94684 47852
rect 94740 47850 94788 47852
rect 94636 47798 94644 47850
rect 94740 47798 94768 47850
rect 94636 47796 94684 47798
rect 94740 47796 94788 47798
rect 94844 47796 94892 47852
rect 94268 47786 94948 47796
rect 93436 47394 93492 47404
rect 92876 47294 92878 47346
rect 92930 47294 92932 47346
rect 92876 47282 92932 47294
rect 91980 46788 92036 46798
rect 91868 46676 91924 46686
rect 91868 46582 91924 46620
rect 91980 45890 92036 46732
rect 91980 45838 91982 45890
rect 92034 45838 92036 45890
rect 91980 45826 92036 45838
rect 92204 46786 92260 46798
rect 92204 46734 92206 46786
rect 92258 46734 92260 46786
rect 92204 45892 92260 46734
rect 92540 46788 92596 46798
rect 92540 46694 92596 46732
rect 92876 46676 92932 46686
rect 96012 46676 96068 46686
rect 92540 45892 92596 45902
rect 92204 45890 92596 45892
rect 92204 45838 92542 45890
rect 92594 45838 92596 45890
rect 92204 45836 92596 45838
rect 92540 45826 92596 45836
rect 91308 45666 91364 45678
rect 91308 45614 91310 45666
rect 91362 45614 91364 45666
rect 91308 45556 91364 45614
rect 91308 45490 91364 45500
rect 92540 45668 92596 45678
rect 91196 45332 91252 45342
rect 91196 45238 91252 45276
rect 91980 45332 92036 45342
rect 90692 45164 90916 45220
rect 90636 45126 90692 45164
rect 85268 44716 85948 44726
rect 85324 44660 85372 44716
rect 85428 44714 85476 44716
rect 85532 44714 85580 44716
rect 85448 44662 85476 44714
rect 85572 44662 85580 44714
rect 85428 44660 85476 44662
rect 85532 44660 85580 44662
rect 85636 44714 85684 44716
rect 85740 44714 85788 44716
rect 85636 44662 85644 44714
rect 85740 44662 85768 44714
rect 85636 44660 85684 44662
rect 85740 44660 85788 44662
rect 85844 44660 85892 44716
rect 85268 44650 85948 44660
rect 89768 43932 90448 43942
rect 89824 43876 89872 43932
rect 89928 43930 89976 43932
rect 90032 43930 90080 43932
rect 89948 43878 89976 43930
rect 90072 43878 90080 43930
rect 89928 43876 89976 43878
rect 90032 43876 90080 43878
rect 90136 43930 90184 43932
rect 90240 43930 90288 43932
rect 90136 43878 90144 43930
rect 90240 43878 90268 43930
rect 90136 43876 90184 43878
rect 90240 43876 90288 43878
rect 90344 43876 90392 43932
rect 89768 43866 90448 43876
rect 88396 43764 88452 43774
rect 83468 43652 83748 43708
rect 80556 43426 80612 43438
rect 80556 43374 80558 43426
rect 80610 43374 80612 43426
rect 80556 41972 80612 43374
rect 80768 42364 81448 42374
rect 80824 42308 80872 42364
rect 80928 42362 80976 42364
rect 81032 42362 81080 42364
rect 80948 42310 80976 42362
rect 81072 42310 81080 42362
rect 80928 42308 80976 42310
rect 81032 42308 81080 42310
rect 81136 42362 81184 42364
rect 81240 42362 81288 42364
rect 81136 42310 81144 42362
rect 81240 42310 81268 42362
rect 81136 42308 81184 42310
rect 81240 42308 81288 42310
rect 81344 42308 81392 42364
rect 80768 42298 81448 42308
rect 80556 41906 80612 41916
rect 80892 41972 80948 41982
rect 80892 40964 80948 41916
rect 81676 41972 81732 41982
rect 81564 41412 81620 41422
rect 81564 41318 81620 41356
rect 80892 40898 80948 40908
rect 80768 40796 81448 40806
rect 80824 40740 80872 40796
rect 80928 40794 80976 40796
rect 81032 40794 81080 40796
rect 80948 40742 80976 40794
rect 81072 40742 81080 40794
rect 80928 40740 80976 40742
rect 81032 40740 81080 40742
rect 81136 40794 81184 40796
rect 81240 40794 81288 40796
rect 81136 40742 81144 40794
rect 81240 40742 81268 40794
rect 81136 40740 81184 40742
rect 81240 40740 81288 40742
rect 81344 40740 81392 40796
rect 80768 40730 81448 40740
rect 80768 39228 81448 39238
rect 80824 39172 80872 39228
rect 80928 39226 80976 39228
rect 81032 39226 81080 39228
rect 80948 39174 80976 39226
rect 81072 39174 81080 39226
rect 80928 39172 80976 39174
rect 81032 39172 81080 39174
rect 81136 39226 81184 39228
rect 81240 39226 81288 39228
rect 81136 39174 81144 39226
rect 81240 39174 81268 39226
rect 81136 39172 81184 39174
rect 81240 39172 81288 39174
rect 81344 39172 81392 39228
rect 80768 39162 81448 39172
rect 79548 38658 79604 38668
rect 78316 38052 78372 38062
rect 78540 38052 78596 38062
rect 78316 38050 78484 38052
rect 78316 37998 78318 38050
rect 78370 37998 78484 38050
rect 78316 37996 78484 37998
rect 78316 37986 78372 37996
rect 78316 37828 78372 37838
rect 78316 37266 78372 37772
rect 78428 37604 78484 37996
rect 78540 37938 78596 37996
rect 78876 38050 78932 38612
rect 78876 37998 78878 38050
rect 78930 37998 78932 38050
rect 78876 37986 78932 37998
rect 79324 38052 79380 38062
rect 79324 37958 79380 37996
rect 78540 37886 78542 37938
rect 78594 37886 78596 37938
rect 78540 37874 78596 37886
rect 81676 37938 81732 41916
rect 83468 41972 83524 43652
rect 83692 43650 83748 43652
rect 83692 43598 83694 43650
rect 83746 43598 83748 43650
rect 83692 43586 83748 43598
rect 84476 43652 84532 43662
rect 84476 43558 84532 43596
rect 86604 43650 86660 43662
rect 86604 43598 86606 43650
rect 86658 43598 86660 43650
rect 85268 43148 85948 43158
rect 85324 43092 85372 43148
rect 85428 43146 85476 43148
rect 85532 43146 85580 43148
rect 85448 43094 85476 43146
rect 85572 43094 85580 43146
rect 85428 43092 85476 43094
rect 85532 43092 85580 43094
rect 85636 43146 85684 43148
rect 85740 43146 85788 43148
rect 85636 43094 85644 43146
rect 85740 43094 85768 43146
rect 85636 43092 85684 43094
rect 85740 43092 85788 43094
rect 85844 43092 85892 43148
rect 85268 43082 85948 43092
rect 86604 42754 86660 43598
rect 86940 42756 86996 42766
rect 86604 42702 86606 42754
rect 86658 42702 86660 42754
rect 86604 42690 86660 42702
rect 86828 42754 86996 42756
rect 86828 42702 86942 42754
rect 86994 42702 86996 42754
rect 86828 42700 86996 42702
rect 86828 42194 86884 42700
rect 86940 42690 86996 42700
rect 86828 42142 86830 42194
rect 86882 42142 86884 42194
rect 86828 42130 86884 42142
rect 87500 42140 88228 42196
rect 83468 41906 83524 41916
rect 87164 41972 87220 41982
rect 87164 41878 87220 41916
rect 85268 41580 85948 41590
rect 85324 41524 85372 41580
rect 85428 41578 85476 41580
rect 85532 41578 85580 41580
rect 85448 41526 85476 41578
rect 85572 41526 85580 41578
rect 85428 41524 85476 41526
rect 85532 41524 85580 41526
rect 85636 41578 85684 41580
rect 85740 41578 85788 41580
rect 85636 41526 85644 41578
rect 85740 41526 85768 41578
rect 85636 41524 85684 41526
rect 85740 41524 85788 41526
rect 85844 41524 85892 41580
rect 85268 41514 85948 41524
rect 82572 40964 82628 40974
rect 82460 40962 82628 40964
rect 82460 40910 82574 40962
rect 82626 40910 82628 40962
rect 82460 40908 82628 40910
rect 82460 40402 82516 40908
rect 82572 40898 82628 40908
rect 84588 40964 84644 40974
rect 84588 40962 85092 40964
rect 84588 40910 84590 40962
rect 84642 40910 85092 40962
rect 84588 40908 85092 40910
rect 84588 40898 84644 40908
rect 84140 40740 84196 40750
rect 82796 40404 82852 40414
rect 82460 40350 82462 40402
rect 82514 40350 82516 40402
rect 82460 40338 82516 40350
rect 82572 40402 82852 40404
rect 82572 40350 82798 40402
rect 82850 40350 82852 40402
rect 82572 40348 82852 40350
rect 82124 39732 82180 39742
rect 82180 39676 82516 39732
rect 82124 39638 82180 39676
rect 82460 39618 82516 39676
rect 82572 39730 82628 40348
rect 82796 40338 82852 40348
rect 82572 39678 82574 39730
rect 82626 39678 82628 39730
rect 82572 39666 82628 39678
rect 82460 39566 82462 39618
rect 82514 39566 82516 39618
rect 82460 39554 82516 39566
rect 83020 39620 83076 39630
rect 83020 39526 83076 39564
rect 83916 39620 83972 39630
rect 83916 39526 83972 39564
rect 84140 39506 84196 40684
rect 84924 39620 84980 39630
rect 84924 39526 84980 39564
rect 85036 39620 85092 40908
rect 85372 40628 85428 40638
rect 85372 40534 85428 40572
rect 85932 40628 85988 40638
rect 85932 40534 85988 40572
rect 86268 40516 86324 40526
rect 86268 40422 86324 40460
rect 86828 40516 86884 40526
rect 85268 40012 85948 40022
rect 85324 39956 85372 40012
rect 85428 40010 85476 40012
rect 85532 40010 85580 40012
rect 85448 39958 85476 40010
rect 85572 39958 85580 40010
rect 85428 39956 85476 39958
rect 85532 39956 85580 39958
rect 85636 40010 85684 40012
rect 85740 40010 85788 40012
rect 85636 39958 85644 40010
rect 85740 39958 85768 40010
rect 85636 39956 85684 39958
rect 85740 39956 85788 39958
rect 85844 39956 85892 40012
rect 85268 39946 85948 39956
rect 85372 39620 85428 39630
rect 85596 39620 85652 39630
rect 86604 39620 86660 39630
rect 85036 39618 85316 39620
rect 85036 39566 85038 39618
rect 85090 39566 85316 39618
rect 85036 39564 85316 39566
rect 85036 39554 85092 39564
rect 84140 39454 84142 39506
rect 84194 39454 84196 39506
rect 84140 39442 84196 39454
rect 84252 39506 84308 39518
rect 84252 39454 84254 39506
rect 84306 39454 84308 39506
rect 82684 39394 82740 39406
rect 82684 39342 82686 39394
rect 82738 39342 82740 39394
rect 82684 39060 82740 39342
rect 82684 38994 82740 39004
rect 83468 39394 83524 39406
rect 83468 39342 83470 39394
rect 83522 39342 83524 39394
rect 83468 39060 83524 39342
rect 83468 38994 83524 39004
rect 83916 38948 83972 38958
rect 83692 38722 83748 38734
rect 83692 38670 83694 38722
rect 83746 38670 83748 38722
rect 83692 38610 83748 38670
rect 83692 38558 83694 38610
rect 83746 38558 83748 38610
rect 83692 38546 83748 38558
rect 81676 37886 81678 37938
rect 81730 37886 81732 37938
rect 81676 37874 81732 37886
rect 82460 37828 82516 37838
rect 82460 37734 82516 37772
rect 83468 37828 83524 37838
rect 80768 37660 81448 37670
rect 80824 37604 80872 37660
rect 80928 37658 80976 37660
rect 81032 37658 81080 37660
rect 80948 37606 80976 37658
rect 81072 37606 81080 37658
rect 80928 37604 80976 37606
rect 81032 37604 81080 37606
rect 81136 37658 81184 37660
rect 81240 37658 81288 37660
rect 81136 37606 81144 37658
rect 81240 37606 81268 37658
rect 81136 37604 81184 37606
rect 81240 37604 81288 37606
rect 81344 37604 81392 37660
rect 78428 37548 78708 37604
rect 80768 37594 81448 37604
rect 78652 37490 78708 37548
rect 78652 37438 78654 37490
rect 78706 37438 78708 37490
rect 78652 37426 78708 37438
rect 83468 37380 83524 37772
rect 83468 37314 83524 37324
rect 78316 37214 78318 37266
rect 78370 37214 78372 37266
rect 78316 37202 78372 37214
rect 83916 37266 83972 38892
rect 84252 38668 84308 39454
rect 84364 39508 84420 39518
rect 84364 39058 84420 39452
rect 84812 39508 84868 39518
rect 84812 39414 84868 39452
rect 84364 39006 84366 39058
rect 84418 39006 84420 39058
rect 84364 38994 84420 39006
rect 84476 39060 84532 39070
rect 84140 38612 84308 38668
rect 84140 38610 84196 38612
rect 84140 38558 84142 38610
rect 84194 38558 84196 38610
rect 84140 37940 84196 38558
rect 84140 37874 84196 37884
rect 84252 37828 84308 37838
rect 84252 37734 84308 37772
rect 84364 37826 84420 37838
rect 84364 37774 84366 37826
rect 84418 37774 84420 37826
rect 83916 37214 83918 37266
rect 83970 37214 83972 37266
rect 83916 37202 83972 37214
rect 84364 37266 84420 37774
rect 84476 37828 84532 39004
rect 85260 39060 85316 39564
rect 85372 39618 85652 39620
rect 85372 39566 85374 39618
rect 85426 39566 85598 39618
rect 85650 39566 85652 39618
rect 85372 39564 85652 39566
rect 85372 39554 85428 39564
rect 85596 39554 85652 39564
rect 86380 39618 86660 39620
rect 86380 39566 86606 39618
rect 86658 39566 86660 39618
rect 86380 39564 86660 39566
rect 85932 39506 85988 39518
rect 85932 39454 85934 39506
rect 85986 39454 85988 39506
rect 85820 39396 85876 39406
rect 85820 39302 85876 39340
rect 85260 38966 85316 39004
rect 84700 38948 84756 38958
rect 84700 38854 84756 38892
rect 85708 38722 85764 38734
rect 85708 38670 85710 38722
rect 85762 38670 85764 38722
rect 85708 38612 85764 38670
rect 85932 38612 85988 39454
rect 86380 39506 86436 39564
rect 86604 39554 86660 39564
rect 86380 39454 86382 39506
rect 86434 39454 86436 39506
rect 86380 39442 86436 39454
rect 85708 38556 86100 38612
rect 85268 38444 85948 38454
rect 85324 38388 85372 38444
rect 85428 38442 85476 38444
rect 85532 38442 85580 38444
rect 85448 38390 85476 38442
rect 85572 38390 85580 38442
rect 85428 38388 85476 38390
rect 85532 38388 85580 38390
rect 85636 38442 85684 38444
rect 85740 38442 85788 38444
rect 85636 38390 85644 38442
rect 85740 38390 85768 38442
rect 85636 38388 85684 38390
rect 85740 38388 85788 38390
rect 85844 38388 85892 38444
rect 85268 38378 85948 38388
rect 84924 38052 84980 38062
rect 85148 38052 85204 38062
rect 84924 38050 85204 38052
rect 84924 37998 84926 38050
rect 84978 37998 85150 38050
rect 85202 37998 85204 38050
rect 84924 37996 85204 37998
rect 84924 37986 84980 37996
rect 85148 37986 85204 37996
rect 85484 37938 85540 37950
rect 85484 37886 85486 37938
rect 85538 37886 85540 37938
rect 84924 37828 84980 37838
rect 84476 37826 84868 37828
rect 84476 37774 84478 37826
rect 84530 37774 84868 37826
rect 84476 37772 84868 37774
rect 84476 37762 84532 37772
rect 84364 37214 84366 37266
rect 84418 37214 84420 37266
rect 84364 37202 84420 37214
rect 75740 36866 75796 36876
rect 76268 36876 76948 36886
rect 76324 36820 76372 36876
rect 76428 36874 76476 36876
rect 76532 36874 76580 36876
rect 76448 36822 76476 36874
rect 76572 36822 76580 36874
rect 76428 36820 76476 36822
rect 76532 36820 76580 36822
rect 76636 36874 76684 36876
rect 76740 36874 76788 36876
rect 76636 36822 76644 36874
rect 76740 36822 76768 36874
rect 76636 36820 76684 36822
rect 76740 36820 76788 36822
rect 76844 36820 76892 36876
rect 76268 36810 76948 36820
rect 77196 36596 77252 36988
rect 77196 36502 77252 36540
rect 76268 35308 76948 35318
rect 76324 35252 76372 35308
rect 76428 35306 76476 35308
rect 76532 35306 76580 35308
rect 76448 35254 76476 35306
rect 76572 35254 76580 35306
rect 76428 35252 76476 35254
rect 76532 35252 76580 35254
rect 76636 35306 76684 35308
rect 76740 35306 76788 35308
rect 76636 35254 76644 35306
rect 76740 35254 76768 35306
rect 76636 35252 76684 35254
rect 76740 35252 76788 35254
rect 76844 35252 76892 35308
rect 76268 35242 76948 35252
rect 77644 34804 77700 34814
rect 77756 34804 77812 37100
rect 84252 36708 84308 36718
rect 77980 36484 78036 36494
rect 77980 35924 78036 36428
rect 81564 36372 81620 36382
rect 78428 36260 78484 36270
rect 78204 35924 78260 35934
rect 77980 35922 78260 35924
rect 77980 35870 77982 35922
rect 78034 35870 78206 35922
rect 78258 35870 78260 35922
rect 77980 35868 78260 35870
rect 77980 35858 78036 35868
rect 78204 35858 78260 35868
rect 78428 35924 78484 36204
rect 78988 36260 79044 36270
rect 78988 36166 79044 36204
rect 80768 36092 81448 36102
rect 80824 36036 80872 36092
rect 80928 36090 80976 36092
rect 81032 36090 81080 36092
rect 80948 36038 80976 36090
rect 81072 36038 81080 36090
rect 80928 36036 80976 36038
rect 81032 36036 81080 36038
rect 81136 36090 81184 36092
rect 81240 36090 81288 36092
rect 81136 36038 81144 36090
rect 81240 36038 81268 36090
rect 81136 36036 81184 36038
rect 81240 36036 81288 36038
rect 81344 36036 81392 36092
rect 80768 36026 81448 36036
rect 78428 35830 78484 35868
rect 79100 35810 79156 35822
rect 79100 35758 79102 35810
rect 79154 35758 79156 35810
rect 78876 35700 78932 35710
rect 78876 35606 78932 35644
rect 78316 35586 78372 35598
rect 78316 35534 78318 35586
rect 78370 35534 78372 35586
rect 78092 35364 78148 35374
rect 78092 34914 78148 35308
rect 78092 34862 78094 34914
rect 78146 34862 78148 34914
rect 78092 34850 78148 34862
rect 78316 34916 78372 35534
rect 79100 35364 79156 35758
rect 80220 35812 80276 35822
rect 80220 35718 80276 35756
rect 81564 35812 81620 36316
rect 84252 35924 84308 36652
rect 84812 36260 84868 37772
rect 84588 35924 84644 35934
rect 84252 35922 84644 35924
rect 84252 35870 84254 35922
rect 84306 35870 84590 35922
rect 84642 35870 84644 35922
rect 84252 35868 84644 35870
rect 84252 35858 84308 35868
rect 84588 35858 84644 35868
rect 79996 35700 80052 35710
rect 79996 35606 80052 35644
rect 80332 35698 80388 35710
rect 80332 35646 80334 35698
rect 80386 35646 80388 35698
rect 80332 35588 80388 35646
rect 80780 35588 80836 35598
rect 80332 35586 80836 35588
rect 80332 35534 80782 35586
rect 80834 35534 80836 35586
rect 80332 35532 80836 35534
rect 80332 35476 80388 35532
rect 80332 35410 80388 35420
rect 79100 35298 79156 35308
rect 80780 35364 80836 35532
rect 80780 35298 80836 35308
rect 81564 35138 81620 35756
rect 81564 35086 81566 35138
rect 81618 35086 81620 35138
rect 81564 35074 81620 35086
rect 84588 35700 84644 35710
rect 78428 34916 78484 34926
rect 78316 34914 78484 34916
rect 78316 34862 78430 34914
rect 78482 34862 78484 34914
rect 78316 34860 78484 34862
rect 78428 34850 78484 34860
rect 84588 34914 84644 35644
rect 84588 34862 84590 34914
rect 84642 34862 84644 34914
rect 84588 34850 84644 34862
rect 84700 35698 84756 35710
rect 84700 35646 84702 35698
rect 84754 35646 84756 35698
rect 84700 34916 84756 35646
rect 84812 35698 84868 36204
rect 84812 35646 84814 35698
rect 84866 35646 84868 35698
rect 84812 35364 84868 35646
rect 84924 35588 84980 37772
rect 85372 37826 85428 37838
rect 85372 37774 85374 37826
rect 85426 37774 85428 37826
rect 85372 37044 85428 37774
rect 85484 37828 85540 37886
rect 85484 37762 85540 37772
rect 85932 37828 85988 37838
rect 86044 37828 86100 38556
rect 85988 37772 86100 37828
rect 85932 37734 85988 37772
rect 86828 37492 86884 40460
rect 87500 40292 87556 42140
rect 88172 42082 88228 42140
rect 88172 42030 88174 42082
rect 88226 42030 88228 42082
rect 88172 42018 88228 42030
rect 88396 41972 88452 43708
rect 90860 43764 90916 45164
rect 91084 45154 91140 45164
rect 91756 45220 91812 45230
rect 91756 45106 91812 45164
rect 91980 45218 92036 45276
rect 91980 45166 91982 45218
rect 92034 45166 92036 45218
rect 91980 45154 92036 45166
rect 91756 45054 91758 45106
rect 91810 45054 91812 45106
rect 91756 45042 91812 45054
rect 92540 45106 92596 45612
rect 92876 45330 92932 46620
rect 95900 46620 96012 46676
rect 94268 46284 94948 46294
rect 94324 46228 94372 46284
rect 94428 46282 94476 46284
rect 94532 46282 94580 46284
rect 94448 46230 94476 46282
rect 94572 46230 94580 46282
rect 94428 46228 94476 46230
rect 94532 46228 94580 46230
rect 94636 46282 94684 46284
rect 94740 46282 94788 46284
rect 94636 46230 94644 46282
rect 94740 46230 94768 46282
rect 94636 46228 94684 46230
rect 94740 46228 94788 46230
rect 94844 46228 94892 46284
rect 94268 46218 94948 46228
rect 92876 45278 92878 45330
rect 92930 45278 92932 45330
rect 92876 45266 92932 45278
rect 95004 45666 95060 45678
rect 95004 45614 95006 45666
rect 95058 45614 95060 45666
rect 95004 45556 95060 45614
rect 95676 45668 95732 45678
rect 95676 45574 95732 45612
rect 92540 45054 92542 45106
rect 92594 45054 92596 45106
rect 92540 45042 92596 45054
rect 94268 44716 94948 44726
rect 94324 44660 94372 44716
rect 94428 44714 94476 44716
rect 94532 44714 94580 44716
rect 94448 44662 94476 44714
rect 94572 44662 94580 44714
rect 94428 44660 94476 44662
rect 94532 44660 94580 44662
rect 94636 44714 94684 44716
rect 94740 44714 94788 44716
rect 94636 44662 94644 44714
rect 94740 44662 94768 44714
rect 94636 44660 94684 44662
rect 94740 44660 94788 44662
rect 94844 44660 94892 44716
rect 94268 44650 94948 44660
rect 90412 42756 90468 42766
rect 89964 42754 90692 42756
rect 89964 42702 90414 42754
rect 90466 42702 90692 42754
rect 89964 42700 90692 42702
rect 88284 41970 88452 41972
rect 88284 41918 88398 41970
rect 88450 41918 88452 41970
rect 88284 41916 88452 41918
rect 88284 41748 88340 41916
rect 88396 41906 88452 41916
rect 88844 42532 88900 42542
rect 88844 41970 88900 42476
rect 89516 42532 89572 42542
rect 89964 42532 90020 42700
rect 90412 42690 90468 42700
rect 89516 42530 90020 42532
rect 89516 42478 89518 42530
rect 89570 42478 90020 42530
rect 89516 42476 90020 42478
rect 90076 42532 90132 42570
rect 89516 42466 89572 42476
rect 90076 42466 90132 42476
rect 89768 42364 90448 42374
rect 89824 42308 89872 42364
rect 89928 42362 89976 42364
rect 90032 42362 90080 42364
rect 89948 42310 89976 42362
rect 90072 42310 90080 42362
rect 89928 42308 89976 42310
rect 90032 42308 90080 42310
rect 90136 42362 90184 42364
rect 90240 42362 90288 42364
rect 90136 42310 90144 42362
rect 90240 42310 90268 42362
rect 90136 42308 90184 42310
rect 90240 42308 90288 42310
rect 90344 42308 90392 42364
rect 89768 42298 90448 42308
rect 88844 41918 88846 41970
rect 88898 41918 88900 41970
rect 88844 41906 88900 41918
rect 89180 41972 89236 41982
rect 89180 41878 89236 41916
rect 87612 41692 88340 41748
rect 87612 41298 87668 41692
rect 87612 41246 87614 41298
rect 87666 41246 87668 41298
rect 87612 41234 87668 41246
rect 89768 40796 90448 40806
rect 89824 40740 89872 40796
rect 89928 40794 89976 40796
rect 90032 40794 90080 40796
rect 89948 40742 89976 40794
rect 90072 40742 90080 40794
rect 89928 40740 89976 40742
rect 90032 40740 90080 40742
rect 90136 40794 90184 40796
rect 90240 40794 90288 40796
rect 90136 40742 90144 40794
rect 90240 40742 90268 40794
rect 90136 40740 90184 40742
rect 90240 40740 90288 40742
rect 90344 40740 90392 40796
rect 89768 40730 90448 40740
rect 90636 40628 90692 42700
rect 90860 42530 90916 43708
rect 92316 43764 92372 43774
rect 91420 43650 91476 43662
rect 91420 43598 91422 43650
rect 91474 43598 91476 43650
rect 91420 43540 91476 43598
rect 91644 43540 91700 43550
rect 92204 43540 92260 43550
rect 91420 43538 91700 43540
rect 91420 43486 91646 43538
rect 91698 43486 91700 43538
rect 91420 43484 91700 43486
rect 91644 43474 91700 43484
rect 92092 43538 92260 43540
rect 92092 43486 92206 43538
rect 92258 43486 92260 43538
rect 92092 43484 92260 43486
rect 90860 42478 90862 42530
rect 90914 42478 90916 42530
rect 90748 40628 90804 40638
rect 90636 40626 90804 40628
rect 90636 40574 90750 40626
rect 90802 40574 90804 40626
rect 90636 40572 90804 40574
rect 87500 40226 87556 40236
rect 89516 40516 89572 40526
rect 87164 39620 87220 39630
rect 87164 39526 87220 39564
rect 89516 39394 89572 40460
rect 90636 39730 90692 40572
rect 90748 40516 90804 40572
rect 90748 40450 90804 40460
rect 90636 39678 90638 39730
rect 90690 39678 90692 39730
rect 90636 39666 90692 39678
rect 89516 39342 89518 39394
rect 89570 39342 89572 39394
rect 89068 38948 89124 38958
rect 87164 38612 87220 38622
rect 87164 38164 87220 38556
rect 89068 38164 89124 38892
rect 87164 38162 87556 38164
rect 87164 38110 87166 38162
rect 87218 38110 87556 38162
rect 87164 38108 87556 38110
rect 87164 38098 87220 38108
rect 87500 38052 87556 38108
rect 89068 38098 89124 38108
rect 87500 37958 87556 37996
rect 86828 37398 86884 37436
rect 88060 37826 88116 37838
rect 88060 37774 88062 37826
rect 88114 37774 88116 37826
rect 88060 37492 88116 37774
rect 88060 37398 88116 37436
rect 89516 37492 89572 39342
rect 90300 39396 90356 39434
rect 90300 39330 90356 39340
rect 89768 39228 90448 39238
rect 89824 39172 89872 39228
rect 89928 39226 89976 39228
rect 90032 39226 90080 39228
rect 89948 39174 89976 39226
rect 90072 39174 90080 39226
rect 89928 39172 89976 39174
rect 90032 39172 90080 39174
rect 90136 39226 90184 39228
rect 90240 39226 90288 39228
rect 90136 39174 90144 39226
rect 90240 39174 90268 39226
rect 90136 39172 90184 39174
rect 90240 39172 90288 39174
rect 90344 39172 90392 39228
rect 89768 39162 90448 39172
rect 89740 39060 89796 39070
rect 89740 38966 89796 39004
rect 90860 39060 90916 42478
rect 90972 43428 91028 43438
rect 90972 39956 91028 43372
rect 91980 42642 92036 42654
rect 91980 42590 91982 42642
rect 92034 42590 92036 42642
rect 91420 42532 91476 42542
rect 91980 42532 92036 42590
rect 91420 42530 92036 42532
rect 91420 42478 91422 42530
rect 91474 42478 92036 42530
rect 91420 42476 92036 42478
rect 91420 41748 91476 42476
rect 91980 42196 92036 42206
rect 92092 42196 92148 43484
rect 92204 43474 92260 43484
rect 92316 42754 92372 43708
rect 94556 43650 94612 43662
rect 94556 43598 94558 43650
rect 94610 43598 94612 43650
rect 94556 43428 94612 43598
rect 94556 43362 94612 43372
rect 94268 43148 94948 43158
rect 94324 43092 94372 43148
rect 94428 43146 94476 43148
rect 94532 43146 94580 43148
rect 94448 43094 94476 43146
rect 94572 43094 94580 43146
rect 94428 43092 94476 43094
rect 94532 43092 94580 43094
rect 94636 43146 94684 43148
rect 94740 43146 94788 43148
rect 94636 43094 94644 43146
rect 94740 43094 94768 43146
rect 94636 43092 94684 43094
rect 94740 43092 94788 43094
rect 94844 43092 94892 43148
rect 94268 43082 94948 43092
rect 92764 42980 92820 42990
rect 92764 42886 92820 42924
rect 92316 42702 92318 42754
rect 92370 42702 92372 42754
rect 92316 42690 92372 42702
rect 91980 42194 92148 42196
rect 91980 42142 91982 42194
rect 92034 42142 92148 42194
rect 91980 42140 92148 42142
rect 92316 42532 92372 42542
rect 91980 42130 92036 42140
rect 92316 41970 92372 42476
rect 93100 42532 93156 42542
rect 93100 42438 93156 42476
rect 92316 41918 92318 41970
rect 92370 41918 92372 41970
rect 92316 41906 92372 41918
rect 91084 41692 91476 41748
rect 91084 40180 91140 41692
rect 94268 41580 94948 41590
rect 94324 41524 94372 41580
rect 94428 41578 94476 41580
rect 94532 41578 94580 41580
rect 94448 41526 94476 41578
rect 94572 41526 94580 41578
rect 94428 41524 94476 41526
rect 94532 41524 94580 41526
rect 94636 41578 94684 41580
rect 94740 41578 94788 41580
rect 94636 41526 94644 41578
rect 94740 41526 94768 41578
rect 94636 41524 94684 41526
rect 94740 41524 94788 41526
rect 94844 41524 94892 41580
rect 94268 41514 94948 41524
rect 95004 41076 95060 45500
rect 95564 44210 95620 44222
rect 95564 44158 95566 44210
rect 95618 44158 95620 44210
rect 95564 43708 95620 44158
rect 95900 44210 95956 46620
rect 96012 46610 96068 46620
rect 96124 45780 96180 48188
rect 96236 48178 96292 48188
rect 96124 45714 96180 45724
rect 96236 46674 96292 46686
rect 96236 46622 96238 46674
rect 96290 46622 96292 46674
rect 96236 45668 96292 46622
rect 96236 45602 96292 45612
rect 95900 44158 95902 44210
rect 95954 44158 95956 44210
rect 95900 44146 95956 44158
rect 96236 44210 96292 44222
rect 96236 44158 96238 44210
rect 96290 44158 96292 44210
rect 95340 43652 95620 43708
rect 95340 43314 95396 43652
rect 95340 43262 95342 43314
rect 95394 43262 95396 43314
rect 95340 42980 95396 43262
rect 95340 42914 95396 42924
rect 96236 42868 96292 44158
rect 96460 43708 96516 55020
rect 96572 55010 96628 55020
rect 97020 55298 97076 55310
rect 97020 55246 97022 55298
rect 97074 55246 97076 55298
rect 96908 53732 96964 53742
rect 96572 53730 96964 53732
rect 96572 53678 96910 53730
rect 96962 53678 96964 53730
rect 96572 53676 96964 53678
rect 96572 50482 96628 53676
rect 96908 53666 96964 53676
rect 96572 50430 96574 50482
rect 96626 50430 96628 50482
rect 96572 50418 96628 50430
rect 96908 51938 96964 51950
rect 96908 51886 96910 51938
rect 96962 51886 96964 51938
rect 96908 50036 96964 51886
rect 97020 51604 97076 55246
rect 97020 51538 97076 51548
rect 96908 49980 97076 50036
rect 96908 49812 96964 49822
rect 96572 49810 96964 49812
rect 96572 49758 96910 49810
rect 96962 49758 96964 49810
rect 96572 49756 96964 49758
rect 96572 48466 96628 49756
rect 96908 49746 96964 49756
rect 96572 48414 96574 48466
rect 96626 48414 96628 48466
rect 96572 48402 96628 48414
rect 96908 48244 96964 48254
rect 96572 48242 96964 48244
rect 96572 48190 96910 48242
rect 96962 48190 96964 48242
rect 96572 48188 96964 48190
rect 96572 46898 96628 48188
rect 96908 48178 96964 48188
rect 96572 46846 96574 46898
rect 96626 46846 96628 46898
rect 96572 46834 96628 46846
rect 96908 46676 96964 46686
rect 96908 46582 96964 46620
rect 97020 46452 97076 49980
rect 96572 46396 97076 46452
rect 96572 44210 96628 46396
rect 96572 44158 96574 44210
rect 96626 44158 96628 44210
rect 96572 44146 96628 44158
rect 96908 44322 96964 44334
rect 96908 44270 96910 44322
rect 96962 44270 96964 44322
rect 96908 43708 96964 44270
rect 97244 43708 97300 56028
rect 98140 56084 98196 56094
rect 98140 55990 98196 56028
rect 98028 55186 98084 55198
rect 98028 55134 98030 55186
rect 98082 55134 98084 55186
rect 98028 54964 98084 55134
rect 98028 54898 98084 54908
rect 98028 53618 98084 53630
rect 98028 53566 98030 53618
rect 98082 53566 98084 53618
rect 98028 53172 98084 53566
rect 98028 53106 98084 53116
rect 97692 52162 97748 52174
rect 97692 52110 97694 52162
rect 97746 52110 97748 52162
rect 97692 51380 97748 52110
rect 97692 51314 97748 51324
rect 98028 49698 98084 49710
rect 98028 49646 98030 49698
rect 98082 49646 98084 49698
rect 98028 49588 98084 49646
rect 98028 49522 98084 49532
rect 98028 48130 98084 48142
rect 98028 48078 98030 48130
rect 98082 48078 98084 48130
rect 98028 47796 98084 48078
rect 98028 47730 98084 47740
rect 98028 46562 98084 46574
rect 98028 46510 98030 46562
rect 98082 46510 98084 46562
rect 98028 46004 98084 46510
rect 98028 45938 98084 45948
rect 98028 44212 98084 44222
rect 98028 44118 98084 44156
rect 96236 42802 96292 42812
rect 96348 43652 96516 43708
rect 96572 43652 96964 43708
rect 97020 43652 97300 43708
rect 96236 42644 96292 42654
rect 94780 41020 95060 41076
rect 96124 42642 96292 42644
rect 96124 42590 96238 42642
rect 96290 42590 96292 42642
rect 96124 42588 96292 42590
rect 91420 40628 91476 40638
rect 91420 40626 92260 40628
rect 91420 40574 91422 40626
rect 91474 40574 92260 40626
rect 91420 40572 92260 40574
rect 91420 40562 91476 40572
rect 91196 40404 91252 40414
rect 91196 40402 91812 40404
rect 91196 40350 91198 40402
rect 91250 40350 91812 40402
rect 91196 40348 91812 40350
rect 91196 40338 91252 40348
rect 91084 40114 91140 40124
rect 91644 40180 91700 40190
rect 90972 39900 91140 39956
rect 90860 38994 90916 39004
rect 90188 38948 90244 38958
rect 90188 38854 90244 38892
rect 90972 38948 91028 38958
rect 90972 38854 91028 38892
rect 90972 38052 91028 38062
rect 91084 38052 91140 39900
rect 91028 37996 91140 38052
rect 91308 38948 91364 38958
rect 90972 37986 91028 37996
rect 89768 37660 90448 37670
rect 89824 37604 89872 37660
rect 89928 37658 89976 37660
rect 90032 37658 90080 37660
rect 89948 37606 89976 37658
rect 90072 37606 90080 37658
rect 89928 37604 89976 37606
rect 90032 37604 90080 37606
rect 90136 37658 90184 37660
rect 90240 37658 90288 37660
rect 90136 37606 90144 37658
rect 90240 37606 90268 37658
rect 90136 37604 90184 37606
rect 90240 37604 90288 37606
rect 90344 37604 90392 37660
rect 89768 37594 90448 37604
rect 85372 36978 85428 36988
rect 87500 37044 87556 37054
rect 87500 36950 87556 36988
rect 85268 36876 85948 36886
rect 85324 36820 85372 36876
rect 85428 36874 85476 36876
rect 85532 36874 85580 36876
rect 85448 36822 85476 36874
rect 85572 36822 85580 36874
rect 85428 36820 85476 36822
rect 85532 36820 85580 36822
rect 85636 36874 85684 36876
rect 85740 36874 85788 36876
rect 85636 36822 85644 36874
rect 85740 36822 85768 36874
rect 85636 36820 85684 36822
rect 85740 36820 85788 36822
rect 85844 36820 85892 36876
rect 85268 36810 85948 36820
rect 89292 36260 89348 36270
rect 85484 35812 85540 35822
rect 85484 35718 85540 35756
rect 89292 35810 89348 36204
rect 89516 35924 89572 37436
rect 90412 37380 90468 37390
rect 90412 37378 90692 37380
rect 90412 37326 90414 37378
rect 90466 37326 90692 37378
rect 90412 37324 90692 37326
rect 90412 37314 90468 37324
rect 90524 36370 90580 36382
rect 90524 36318 90526 36370
rect 90578 36318 90580 36370
rect 89768 36092 90448 36102
rect 89824 36036 89872 36092
rect 89928 36090 89976 36092
rect 90032 36090 90080 36092
rect 89948 36038 89976 36090
rect 90072 36038 90080 36090
rect 89928 36036 89976 36038
rect 90032 36036 90080 36038
rect 90136 36090 90184 36092
rect 90240 36090 90288 36092
rect 90136 36038 90144 36090
rect 90240 36038 90268 36090
rect 90136 36036 90184 36038
rect 90240 36036 90288 36038
rect 90344 36036 90392 36092
rect 89768 36026 90448 36036
rect 89516 35858 89572 35868
rect 89852 35924 89908 35934
rect 90524 35924 90580 36318
rect 89852 35922 90580 35924
rect 89852 35870 89854 35922
rect 89906 35870 90580 35922
rect 89852 35868 90580 35870
rect 89852 35858 89908 35868
rect 89292 35758 89294 35810
rect 89346 35758 89348 35810
rect 89292 35746 89348 35758
rect 85260 35700 85316 35710
rect 85260 35606 85316 35644
rect 86044 35698 86100 35710
rect 86044 35646 86046 35698
rect 86098 35646 86100 35698
rect 84924 35522 84980 35532
rect 85148 35476 85204 35486
rect 85148 35364 85204 35420
rect 86044 35476 86100 35646
rect 86044 35410 86100 35420
rect 86156 35700 86212 35710
rect 84812 35308 85204 35364
rect 85036 34916 85092 34926
rect 84700 34914 85092 34916
rect 84700 34862 85038 34914
rect 85090 34862 85092 34914
rect 84700 34860 85092 34862
rect 85036 34850 85092 34860
rect 77700 34748 77812 34804
rect 80780 34804 80836 34814
rect 77644 34710 77700 34748
rect 80780 34710 80836 34748
rect 75180 34692 75236 34702
rect 75180 34598 75236 34636
rect 75740 34690 75796 34702
rect 75740 34638 75742 34690
rect 75794 34638 75796 34690
rect 75740 34356 75796 34638
rect 75740 34290 75796 34300
rect 75852 34692 75908 34702
rect 74844 34188 75236 34244
rect 74732 34076 75012 34132
rect 73724 33966 73726 34018
rect 73778 33966 73780 34018
rect 73724 33908 73780 33966
rect 72940 33852 73780 33908
rect 71768 32956 72448 32966
rect 71824 32900 71872 32956
rect 71928 32954 71976 32956
rect 72032 32954 72080 32956
rect 71948 32902 71976 32954
rect 72072 32902 72080 32954
rect 71928 32900 71976 32902
rect 72032 32900 72080 32902
rect 72136 32954 72184 32956
rect 72240 32954 72288 32956
rect 72136 32902 72144 32954
rect 72240 32902 72268 32954
rect 72136 32900 72184 32902
rect 72240 32900 72288 32902
rect 72344 32900 72392 32956
rect 71768 32890 72448 32900
rect 68572 31892 68628 31902
rect 70700 31892 70756 31902
rect 68628 31836 68964 31892
rect 68572 31798 68628 31836
rect 68908 31556 68964 31836
rect 69244 31780 69300 31790
rect 69020 31778 69300 31780
rect 69020 31726 69246 31778
rect 69298 31726 69300 31778
rect 69020 31724 69300 31726
rect 69020 31666 69076 31724
rect 69244 31714 69300 31724
rect 69804 31778 69860 31790
rect 69804 31726 69806 31778
rect 69858 31726 69860 31778
rect 69020 31614 69022 31666
rect 69074 31614 69076 31666
rect 69020 31602 69076 31614
rect 68908 31218 68964 31500
rect 68908 31166 68910 31218
rect 68962 31166 68964 31218
rect 68908 31154 68964 31166
rect 69020 31444 69076 31454
rect 68572 30770 68628 30782
rect 68572 30718 68574 30770
rect 68626 30718 68628 30770
rect 68572 30212 68628 30718
rect 68572 30146 68628 30156
rect 68796 29652 68852 29662
rect 69020 29652 69076 31388
rect 69804 31218 69860 31726
rect 69804 31166 69806 31218
rect 69858 31166 69860 31218
rect 69804 31154 69860 31166
rect 69916 31444 69972 31454
rect 69916 31218 69972 31388
rect 69916 31166 69918 31218
rect 69970 31166 69972 31218
rect 69916 31154 69972 31166
rect 70700 31444 70756 31836
rect 72940 31892 72996 33852
rect 72940 31826 72996 31836
rect 73052 33348 73108 33358
rect 72940 31668 72996 31678
rect 72604 31612 72940 31668
rect 70700 31218 70756 31388
rect 70700 31166 70702 31218
rect 70754 31166 70756 31218
rect 70700 31154 70756 31166
rect 71148 31556 71204 31566
rect 69468 31108 69524 31118
rect 69692 31108 69748 31118
rect 69524 31106 69748 31108
rect 69524 31054 69694 31106
rect 69746 31054 69748 31106
rect 69524 31052 69748 31054
rect 69468 31014 69524 31052
rect 69692 31042 69748 31052
rect 70364 30996 70420 31006
rect 70364 30902 70420 30940
rect 68796 29650 69020 29652
rect 68796 29598 68798 29650
rect 68850 29598 69020 29650
rect 68796 29596 69020 29598
rect 68796 29586 68852 29596
rect 69020 29558 69076 29596
rect 69692 29652 69748 29662
rect 69692 29558 69748 29596
rect 68572 29426 68628 29438
rect 68572 29374 68574 29426
rect 68626 29374 68628 29426
rect 68572 29316 68628 29374
rect 69244 29428 69300 29438
rect 69244 29334 69300 29372
rect 70476 29428 70532 29438
rect 68572 29250 68628 29260
rect 68684 29314 68740 29326
rect 68684 29262 68686 29314
rect 68738 29262 68740 29314
rect 68684 28644 68740 29262
rect 68796 28644 68852 28654
rect 68684 28642 68852 28644
rect 68684 28590 68798 28642
rect 68850 28590 68852 28642
rect 68684 28588 68852 28590
rect 68796 28578 68852 28588
rect 70476 28082 70532 29372
rect 70476 28030 70478 28082
rect 70530 28030 70532 28082
rect 70476 28018 70532 28030
rect 70700 28644 70756 28654
rect 70700 28082 70756 28588
rect 71148 28530 71204 31500
rect 72156 31556 72212 31594
rect 72156 31490 72212 31500
rect 71768 31388 72448 31398
rect 71824 31332 71872 31388
rect 71928 31386 71976 31388
rect 72032 31386 72080 31388
rect 71948 31334 71976 31386
rect 72072 31334 72080 31386
rect 71928 31332 71976 31334
rect 72032 31332 72080 31334
rect 72136 31386 72184 31388
rect 72240 31386 72288 31388
rect 72136 31334 72144 31386
rect 72240 31334 72268 31386
rect 72136 31332 72184 31334
rect 72240 31332 72288 31334
rect 72344 31332 72392 31388
rect 71768 31322 72448 31332
rect 72380 31220 72436 31230
rect 72604 31220 72660 31612
rect 72940 31574 72996 31612
rect 72940 31220 72996 31230
rect 73052 31220 73108 33292
rect 74508 33348 74564 34076
rect 74620 34066 74676 34076
rect 74508 33282 74564 33292
rect 74060 31668 74116 31678
rect 74060 31574 74116 31612
rect 74396 31556 74452 31566
rect 74396 31462 74452 31500
rect 72380 31218 72660 31220
rect 72380 31166 72382 31218
rect 72434 31166 72660 31218
rect 72380 31164 72660 31166
rect 72716 31218 73108 31220
rect 72716 31166 72942 31218
rect 72994 31166 73108 31218
rect 72716 31164 73108 31166
rect 72380 31154 72436 31164
rect 72268 30996 72324 31006
rect 72268 30772 72324 30940
rect 72492 30996 72548 31006
rect 72716 30996 72772 31164
rect 72940 31154 72996 31164
rect 72492 30994 72772 30996
rect 72492 30942 72494 30994
rect 72546 30942 72772 30994
rect 72492 30940 72772 30942
rect 72492 30930 72548 30940
rect 72380 30772 72436 30782
rect 72268 30770 72436 30772
rect 72268 30718 72382 30770
rect 72434 30718 72436 30770
rect 72268 30716 72436 30718
rect 72380 30706 72436 30716
rect 72492 30212 72548 30222
rect 72492 30118 72548 30156
rect 72828 30100 72884 30110
rect 72828 30006 72884 30044
rect 71768 29820 72448 29830
rect 71824 29764 71872 29820
rect 71928 29818 71976 29820
rect 72032 29818 72080 29820
rect 71948 29766 71976 29818
rect 72072 29766 72080 29818
rect 71928 29764 71976 29766
rect 72032 29764 72080 29766
rect 72136 29818 72184 29820
rect 72240 29818 72288 29820
rect 72136 29766 72144 29818
rect 72240 29766 72268 29818
rect 72136 29764 72184 29766
rect 72240 29764 72288 29766
rect 72344 29764 72392 29820
rect 71768 29754 72448 29764
rect 71932 28644 71988 28654
rect 71932 28550 71988 28588
rect 72380 28644 72436 28654
rect 72380 28550 72436 28588
rect 72716 28644 72772 28654
rect 71148 28478 71150 28530
rect 71202 28478 71204 28530
rect 71148 28466 71204 28478
rect 72716 28530 72772 28588
rect 72716 28478 72718 28530
rect 72770 28478 72772 28530
rect 72716 28466 72772 28478
rect 71768 28252 72448 28262
rect 71824 28196 71872 28252
rect 71928 28250 71976 28252
rect 72032 28250 72080 28252
rect 71948 28198 71976 28250
rect 72072 28198 72080 28250
rect 71928 28196 71976 28198
rect 72032 28196 72080 28198
rect 72136 28250 72184 28252
rect 72240 28250 72288 28252
rect 72136 28198 72144 28250
rect 72240 28198 72268 28250
rect 72136 28196 72184 28198
rect 72240 28196 72288 28198
rect 72344 28196 72392 28252
rect 71768 28186 72448 28196
rect 70700 28030 70702 28082
rect 70754 28030 70756 28082
rect 70700 28018 70756 28030
rect 70812 27972 70868 27982
rect 70812 26908 70868 27916
rect 71260 27972 71316 27982
rect 71260 27878 71316 27916
rect 73052 27972 73108 31164
rect 74172 28532 74228 28542
rect 74396 28532 74452 28542
rect 74172 28530 74452 28532
rect 74172 28478 74174 28530
rect 74226 28478 74398 28530
rect 74450 28478 74452 28530
rect 74172 28476 74452 28478
rect 74172 28466 74228 28476
rect 67116 26852 67172 26862
rect 68460 26852 68628 26908
rect 67116 26514 67172 26796
rect 67116 26462 67118 26514
rect 67170 26462 67172 26514
rect 67116 26450 67172 26462
rect 67340 26404 67396 26414
rect 67340 26310 67396 26348
rect 68124 26404 68180 26414
rect 68124 26310 68180 26348
rect 67788 26292 67844 26302
rect 67788 26290 68068 26292
rect 67788 26238 67790 26290
rect 67842 26238 68068 26290
rect 67788 26236 68068 26238
rect 67788 26226 67844 26236
rect 67228 26178 67284 26190
rect 67228 26126 67230 26178
rect 67282 26126 67284 26178
rect 67228 26068 67284 26126
rect 67116 26012 67284 26068
rect 67116 25732 67172 26012
rect 67268 25900 67948 25910
rect 67324 25844 67372 25900
rect 67428 25898 67476 25900
rect 67532 25898 67580 25900
rect 67448 25846 67476 25898
rect 67572 25846 67580 25898
rect 67428 25844 67476 25846
rect 67532 25844 67580 25846
rect 67636 25898 67684 25900
rect 67740 25898 67788 25900
rect 67636 25846 67644 25898
rect 67740 25846 67768 25898
rect 67636 25844 67684 25846
rect 67740 25844 67788 25846
rect 67844 25844 67892 25900
rect 67268 25834 67948 25844
rect 68012 25844 68068 26236
rect 68572 25956 68628 26852
rect 70476 26852 70868 26908
rect 72604 27188 72660 27198
rect 68908 26740 68964 26750
rect 68572 25900 68740 25956
rect 68012 25788 68628 25844
rect 67116 25676 67284 25732
rect 65548 23828 65604 23838
rect 65548 23714 65604 23772
rect 65548 23662 65550 23714
rect 65602 23662 65604 23714
rect 65548 23380 65604 23662
rect 66332 23604 66388 23614
rect 65996 23380 66052 23390
rect 65548 23324 65996 23380
rect 65660 22594 65716 23324
rect 65996 23286 66052 23324
rect 66332 23266 66388 23548
rect 67004 23380 67060 24892
rect 67228 24722 67284 25676
rect 68572 25506 68628 25788
rect 68572 25454 68574 25506
rect 68626 25454 68628 25506
rect 68572 25442 68628 25454
rect 67228 24670 67230 24722
rect 67282 24670 67284 24722
rect 67228 24658 67284 24670
rect 67268 24332 67948 24342
rect 67324 24276 67372 24332
rect 67428 24330 67476 24332
rect 67532 24330 67580 24332
rect 67448 24278 67476 24330
rect 67572 24278 67580 24330
rect 67428 24276 67476 24278
rect 67532 24276 67580 24278
rect 67636 24330 67684 24332
rect 67740 24330 67788 24332
rect 67636 24278 67644 24330
rect 67740 24278 67768 24330
rect 67636 24276 67684 24278
rect 67740 24276 67788 24278
rect 67844 24276 67892 24332
rect 67268 24266 67948 24276
rect 67004 23314 67060 23324
rect 66332 23214 66334 23266
rect 66386 23214 66388 23266
rect 66332 23202 66388 23214
rect 66668 23266 66724 23278
rect 66668 23214 66670 23266
rect 66722 23214 66724 23266
rect 65660 22542 65662 22594
rect 65714 22542 65716 22594
rect 65548 20916 65604 20926
rect 65660 20916 65716 22542
rect 66668 21812 66724 23214
rect 67116 23154 67172 23166
rect 67116 23102 67118 23154
rect 67170 23102 67172 23154
rect 67116 22258 67172 23102
rect 67564 23156 67620 23166
rect 67564 23154 68516 23156
rect 67564 23102 67566 23154
rect 67618 23102 68516 23154
rect 67564 23100 68516 23102
rect 67564 23090 67620 23100
rect 67268 22764 67948 22774
rect 67324 22708 67372 22764
rect 67428 22762 67476 22764
rect 67532 22762 67580 22764
rect 67448 22710 67476 22762
rect 67572 22710 67580 22762
rect 67428 22708 67476 22710
rect 67532 22708 67580 22710
rect 67636 22762 67684 22764
rect 67740 22762 67788 22764
rect 67636 22710 67644 22762
rect 67740 22710 67768 22762
rect 67636 22708 67684 22710
rect 67740 22708 67788 22710
rect 67844 22708 67892 22764
rect 67268 22698 67948 22708
rect 68460 22482 68516 23100
rect 68460 22430 68462 22482
rect 68514 22430 68516 22482
rect 68460 22418 68516 22430
rect 68572 22484 68628 22494
rect 68348 22372 68404 22382
rect 68348 22278 68404 22316
rect 68572 22370 68628 22428
rect 68572 22318 68574 22370
rect 68626 22318 68628 22370
rect 68572 22306 68628 22318
rect 67116 22206 67118 22258
rect 67170 22206 67172 22258
rect 67116 22194 67172 22206
rect 66668 21746 66724 21756
rect 67268 21196 67948 21206
rect 67324 21140 67372 21196
rect 67428 21194 67476 21196
rect 67532 21194 67580 21196
rect 67448 21142 67476 21194
rect 67572 21142 67580 21194
rect 67428 21140 67476 21142
rect 67532 21140 67580 21142
rect 67636 21194 67684 21196
rect 67740 21194 67788 21196
rect 67636 21142 67644 21194
rect 67740 21142 67768 21194
rect 67636 21140 67684 21142
rect 67740 21140 67788 21142
rect 67844 21140 67892 21196
rect 67268 21130 67948 21140
rect 65604 20860 65716 20916
rect 65884 21028 65940 21038
rect 65548 20822 65604 20860
rect 65884 20130 65940 20972
rect 68684 20916 68740 25900
rect 68908 25620 68964 26684
rect 70476 26740 70532 26852
rect 70476 26674 70532 26684
rect 71768 26684 72448 26694
rect 71824 26628 71872 26684
rect 71928 26682 71976 26684
rect 72032 26682 72080 26684
rect 71948 26630 71976 26682
rect 72072 26630 72080 26682
rect 71928 26628 71976 26630
rect 72032 26628 72080 26630
rect 72136 26682 72184 26684
rect 72240 26682 72288 26684
rect 72136 26630 72144 26682
rect 72240 26630 72268 26682
rect 72136 26628 72184 26630
rect 72240 26628 72288 26630
rect 72344 26628 72392 26684
rect 71768 26618 72448 26628
rect 72492 26516 72548 26526
rect 72604 26516 72660 27132
rect 73052 26964 73108 27916
rect 73612 27858 73668 27870
rect 73612 27806 73614 27858
rect 73666 27806 73668 27858
rect 73164 27748 73220 27758
rect 73164 27654 73220 27692
rect 73612 27748 73668 27806
rect 73668 27692 73780 27748
rect 73612 27682 73668 27692
rect 73724 27188 73780 27692
rect 73836 27188 73892 27198
rect 74284 27188 74340 28476
rect 74396 28466 74452 28476
rect 74620 27748 74676 27758
rect 74956 27748 75012 34076
rect 75068 34018 75124 34030
rect 75068 33966 75070 34018
rect 75122 33966 75124 34018
rect 75068 33348 75124 33966
rect 75068 33282 75124 33292
rect 75180 28644 75236 34188
rect 75852 32228 75908 34636
rect 76412 34692 76468 34702
rect 76188 34356 76244 34366
rect 76188 34242 76244 34300
rect 76412 34356 76468 34636
rect 84364 34690 84420 34702
rect 84364 34638 84366 34690
rect 84418 34638 84420 34690
rect 80768 34524 81448 34534
rect 80824 34468 80872 34524
rect 80928 34522 80976 34524
rect 81032 34522 81080 34524
rect 80948 34470 80976 34522
rect 81072 34470 81080 34522
rect 80928 34468 80976 34470
rect 81032 34468 81080 34470
rect 81136 34522 81184 34524
rect 81240 34522 81288 34524
rect 81136 34470 81144 34522
rect 81240 34470 81268 34522
rect 81136 34468 81184 34470
rect 81240 34468 81288 34470
rect 81344 34468 81392 34524
rect 80768 34458 81448 34468
rect 76412 34290 76468 34300
rect 84364 34356 84420 34638
rect 84364 34290 84420 34300
rect 76188 34190 76190 34242
rect 76242 34190 76244 34242
rect 76188 34178 76244 34190
rect 76524 34244 76580 34254
rect 76524 34150 76580 34188
rect 76268 33740 76948 33750
rect 76324 33684 76372 33740
rect 76428 33738 76476 33740
rect 76532 33738 76580 33740
rect 76448 33686 76476 33738
rect 76572 33686 76580 33738
rect 76428 33684 76476 33686
rect 76532 33684 76580 33686
rect 76636 33738 76684 33740
rect 76740 33738 76788 33740
rect 76636 33686 76644 33738
rect 76740 33686 76768 33738
rect 76636 33684 76684 33686
rect 76740 33684 76788 33686
rect 76844 33684 76892 33740
rect 76268 33674 76948 33684
rect 80768 32956 81448 32966
rect 80824 32900 80872 32956
rect 80928 32954 80976 32956
rect 81032 32954 81080 32956
rect 80948 32902 80976 32954
rect 81072 32902 81080 32954
rect 80928 32900 80976 32902
rect 81032 32900 81080 32902
rect 81136 32954 81184 32956
rect 81240 32954 81288 32956
rect 81136 32902 81144 32954
rect 81240 32902 81268 32954
rect 81136 32900 81184 32902
rect 81240 32900 81288 32902
rect 81344 32900 81392 32956
rect 80768 32890 81448 32900
rect 75740 32172 75908 32228
rect 76268 32172 76948 32182
rect 75404 29428 75460 29438
rect 75404 28866 75460 29372
rect 75404 28814 75406 28866
rect 75458 28814 75460 28866
rect 75404 28802 75460 28814
rect 75180 28588 75460 28644
rect 74620 27746 75236 27748
rect 74620 27694 74622 27746
rect 74674 27694 75236 27746
rect 74620 27692 75236 27694
rect 74620 27682 74676 27692
rect 73724 27186 74340 27188
rect 73724 27134 73838 27186
rect 73890 27134 74340 27186
rect 73724 27132 74340 27134
rect 73836 27094 73892 27132
rect 74284 27076 74340 27132
rect 74284 27074 74788 27076
rect 74284 27022 74286 27074
rect 74338 27022 74788 27074
rect 74284 27020 74788 27022
rect 74284 27010 74340 27020
rect 73052 26898 73108 26908
rect 72492 26514 72660 26516
rect 72492 26462 72494 26514
rect 72546 26462 72660 26514
rect 72492 26460 72660 26462
rect 74508 26852 74564 26862
rect 72492 26450 72548 26460
rect 72716 26404 72772 26414
rect 72716 26310 72772 26348
rect 73500 26404 73556 26414
rect 73500 26310 73556 26348
rect 73164 26292 73220 26302
rect 73164 26198 73220 26236
rect 74172 26292 74228 26302
rect 72604 26178 72660 26190
rect 72604 26126 72606 26178
rect 72658 26126 72660 26178
rect 69356 25620 69412 25630
rect 68908 25618 69412 25620
rect 68908 25566 69358 25618
rect 69410 25566 69412 25618
rect 68908 25564 69412 25566
rect 68908 25506 68964 25564
rect 69356 25554 69412 25564
rect 72044 25508 72100 25518
rect 68908 25454 68910 25506
rect 68962 25454 68964 25506
rect 68908 25442 68964 25454
rect 71820 25506 72100 25508
rect 71820 25454 72046 25506
rect 72098 25454 72100 25506
rect 71820 25452 72100 25454
rect 71820 25394 71876 25452
rect 72044 25442 72100 25452
rect 72604 25506 72660 26126
rect 72604 25454 72606 25506
rect 72658 25454 72660 25506
rect 72604 25442 72660 25454
rect 71820 25342 71822 25394
rect 71874 25342 71876 25394
rect 71820 25330 71876 25342
rect 68796 25282 68852 25294
rect 68796 25230 68798 25282
rect 68850 25230 68852 25282
rect 68796 24948 68852 25230
rect 71768 25116 72448 25126
rect 71824 25060 71872 25116
rect 71928 25114 71976 25116
rect 72032 25114 72080 25116
rect 71948 25062 71976 25114
rect 72072 25062 72080 25114
rect 71928 25060 71976 25062
rect 72032 25060 72080 25062
rect 72136 25114 72184 25116
rect 72240 25114 72288 25116
rect 72136 25062 72144 25114
rect 72240 25062 72268 25114
rect 72136 25060 72184 25062
rect 72240 25060 72288 25062
rect 72344 25060 72392 25116
rect 71768 25050 72448 25060
rect 68796 24882 68852 24892
rect 70252 24948 70308 24958
rect 70252 24854 70308 24892
rect 71148 24948 71204 24958
rect 69468 24834 69524 24846
rect 69468 24782 69470 24834
rect 69522 24782 69524 24834
rect 69468 23380 69524 24782
rect 71148 23938 71204 24892
rect 74172 24946 74228 26236
rect 74172 24894 74174 24946
rect 74226 24894 74228 24946
rect 74172 24882 74228 24894
rect 74508 26180 74564 26796
rect 74732 26516 74788 27020
rect 74732 26514 75124 26516
rect 74732 26462 74734 26514
rect 74786 26462 75124 26514
rect 74732 26460 75124 26462
rect 74732 26450 74788 26460
rect 75068 26290 75124 26460
rect 75068 26238 75070 26290
rect 75122 26238 75124 26290
rect 75068 26226 75124 26238
rect 74508 25284 74564 26124
rect 75068 25396 75124 25406
rect 74396 24836 74452 24846
rect 74396 24742 74452 24780
rect 74508 24834 74564 25228
rect 74956 25284 75012 25294
rect 74956 24948 75012 25228
rect 75068 25282 75124 25340
rect 75068 25230 75070 25282
rect 75122 25230 75124 25282
rect 75068 25218 75124 25230
rect 75068 24948 75124 24958
rect 74956 24946 75124 24948
rect 74956 24894 75070 24946
rect 75122 24894 75124 24946
rect 74956 24892 75124 24894
rect 75068 24882 75124 24892
rect 74508 24782 74510 24834
rect 74562 24782 74564 24834
rect 74508 24770 74564 24782
rect 71148 23886 71150 23938
rect 71202 23886 71204 23938
rect 71148 23874 71204 23886
rect 71484 23714 71540 23726
rect 71484 23662 71486 23714
rect 71538 23662 71540 23714
rect 69468 23314 69524 23324
rect 69804 23380 69860 23390
rect 69804 23286 69860 23324
rect 69356 22932 69412 22942
rect 68908 22372 68964 22382
rect 69132 22372 69188 22382
rect 68908 22370 69188 22372
rect 68908 22318 68910 22370
rect 68962 22318 69134 22370
rect 69186 22318 69188 22370
rect 68908 22316 69188 22318
rect 68908 22306 68964 22316
rect 69132 22306 69188 22316
rect 69356 22258 69412 22876
rect 70588 22932 70644 22942
rect 70644 22876 70756 22932
rect 70588 22838 70644 22876
rect 69916 22484 69972 22494
rect 69916 22390 69972 22428
rect 69356 22206 69358 22258
rect 69410 22206 69412 22258
rect 69356 22194 69412 22206
rect 69468 22258 69524 22270
rect 69468 22206 69470 22258
rect 69522 22206 69524 22258
rect 69468 21700 69524 22206
rect 69468 21634 69524 21644
rect 70364 22146 70420 22158
rect 70364 22094 70366 22146
rect 70418 22094 70420 22146
rect 70364 21700 70420 22094
rect 70364 21634 70420 21644
rect 68684 20850 68740 20860
rect 65884 20078 65886 20130
rect 65938 20078 65940 20130
rect 65884 20066 65940 20078
rect 66220 20130 66276 20142
rect 66220 20078 66222 20130
rect 66274 20078 66276 20130
rect 66220 16100 66276 20078
rect 67268 19628 67948 19638
rect 67324 19572 67372 19628
rect 67428 19626 67476 19628
rect 67532 19626 67580 19628
rect 67448 19574 67476 19626
rect 67572 19574 67580 19626
rect 67428 19572 67476 19574
rect 67532 19572 67580 19574
rect 67636 19626 67684 19628
rect 67740 19626 67788 19628
rect 67636 19574 67644 19626
rect 67740 19574 67768 19626
rect 67636 19572 67684 19574
rect 67740 19572 67788 19574
rect 67844 19572 67892 19628
rect 67268 19562 67948 19572
rect 67268 18060 67948 18070
rect 67324 18004 67372 18060
rect 67428 18058 67476 18060
rect 67532 18058 67580 18060
rect 67448 18006 67476 18058
rect 67572 18006 67580 18058
rect 67428 18004 67476 18006
rect 67532 18004 67580 18006
rect 67636 18058 67684 18060
rect 67740 18058 67788 18060
rect 67636 18006 67644 18058
rect 67740 18006 67768 18058
rect 67636 18004 67684 18006
rect 67740 18004 67788 18006
rect 67844 18004 67892 18060
rect 67268 17994 67948 18004
rect 67268 16492 67948 16502
rect 67324 16436 67372 16492
rect 67428 16490 67476 16492
rect 67532 16490 67580 16492
rect 67448 16438 67476 16490
rect 67572 16438 67580 16490
rect 67428 16436 67476 16438
rect 67532 16436 67580 16438
rect 67636 16490 67684 16492
rect 67740 16490 67788 16492
rect 67636 16438 67644 16490
rect 67740 16438 67768 16490
rect 67636 16436 67684 16438
rect 67740 16436 67788 16438
rect 67844 16436 67892 16492
rect 67268 16426 67948 16436
rect 66220 16034 66276 16044
rect 65324 15092 65492 15148
rect 62768 14140 63448 14150
rect 62824 14084 62872 14140
rect 62928 14138 62976 14140
rect 63032 14138 63080 14140
rect 62948 14086 62976 14138
rect 63072 14086 63080 14138
rect 62928 14084 62976 14086
rect 63032 14084 63080 14086
rect 63136 14138 63184 14140
rect 63240 14138 63288 14140
rect 63136 14086 63144 14138
rect 63240 14086 63268 14138
rect 63136 14084 63184 14086
rect 63240 14084 63288 14086
rect 63344 14084 63392 14140
rect 62768 14074 63448 14084
rect 61852 13860 61908 13870
rect 61292 11442 61348 11452
rect 61740 13858 62020 13860
rect 61740 13806 61854 13858
rect 61906 13806 62020 13858
rect 61740 13804 62020 13806
rect 61180 7074 61236 7084
rect 60284 4162 60340 4172
rect 60508 5964 60788 6020
rect 60060 3502 60062 3554
rect 60114 3502 60116 3554
rect 60060 3490 60116 3502
rect 60172 3892 60228 3902
rect 60172 3554 60228 3836
rect 60172 3502 60174 3554
rect 60226 3502 60228 3554
rect 46396 3278 46398 3330
rect 46450 3278 46452 3330
rect 46396 3266 46452 3278
rect 42700 3154 42756 3164
rect 44768 3164 45448 3174
rect 44824 3108 44872 3164
rect 44928 3162 44976 3164
rect 45032 3162 45080 3164
rect 44948 3110 44976 3162
rect 45072 3110 45080 3162
rect 44928 3108 44976 3110
rect 45032 3108 45080 3110
rect 45136 3162 45184 3164
rect 45240 3162 45288 3164
rect 45136 3110 45144 3162
rect 45240 3110 45268 3162
rect 45136 3108 45184 3110
rect 45240 3108 45288 3110
rect 45344 3108 45392 3164
rect 44768 3098 45448 3108
rect 50316 2212 50372 3388
rect 52668 3378 52724 3388
rect 59948 3442 60004 3454
rect 59948 3390 59950 3442
rect 60002 3390 60004 3442
rect 59948 3388 60004 3390
rect 60172 3388 60228 3502
rect 59948 3332 60228 3388
rect 60508 3442 60564 5964
rect 60732 5236 60788 5246
rect 60732 5142 60788 5180
rect 61740 3892 61796 13804
rect 61852 13794 61908 13804
rect 61964 13746 62020 13804
rect 61964 13694 61966 13746
rect 62018 13694 62020 13746
rect 61964 13682 62020 13694
rect 62768 12572 63448 12582
rect 62824 12516 62872 12572
rect 62928 12570 62976 12572
rect 63032 12570 63080 12572
rect 62948 12518 62976 12570
rect 63072 12518 63080 12570
rect 62928 12516 62976 12518
rect 63032 12516 63080 12518
rect 63136 12570 63184 12572
rect 63240 12570 63288 12572
rect 63136 12518 63144 12570
rect 63240 12518 63268 12570
rect 63136 12516 63184 12518
rect 63240 12516 63288 12518
rect 63344 12516 63392 12572
rect 62768 12506 63448 12516
rect 63756 12178 63812 12190
rect 63756 12126 63758 12178
rect 63810 12126 63812 12178
rect 62188 11508 62244 11518
rect 62188 11414 62244 11452
rect 63644 11508 63700 11518
rect 63644 11394 63700 11452
rect 63644 11342 63646 11394
rect 63698 11342 63700 11394
rect 62768 11004 63448 11014
rect 62824 10948 62872 11004
rect 62928 11002 62976 11004
rect 63032 11002 63080 11004
rect 62948 10950 62976 11002
rect 63072 10950 63080 11002
rect 62928 10948 62976 10950
rect 63032 10948 63080 10950
rect 63136 11002 63184 11004
rect 63240 11002 63288 11004
rect 63136 10950 63144 11002
rect 63240 10950 63268 11002
rect 63136 10948 63184 10950
rect 63240 10948 63288 10950
rect 63344 10948 63392 11004
rect 62768 10938 63448 10948
rect 63532 10498 63588 10510
rect 63532 10446 63534 10498
rect 63586 10446 63588 10498
rect 62412 9714 62468 9726
rect 62412 9662 62414 9714
rect 62466 9662 62468 9714
rect 62412 8372 62468 9662
rect 62768 9436 63448 9446
rect 62824 9380 62872 9436
rect 62928 9434 62976 9436
rect 63032 9434 63080 9436
rect 62948 9382 62976 9434
rect 63072 9382 63080 9434
rect 62928 9380 62976 9382
rect 63032 9380 63080 9382
rect 63136 9434 63184 9436
rect 63240 9434 63288 9436
rect 63136 9382 63144 9434
rect 63240 9382 63268 9434
rect 63136 9380 63184 9382
rect 63240 9380 63288 9382
rect 63344 9380 63392 9436
rect 62768 9370 63448 9380
rect 62412 8306 62468 8316
rect 63084 9044 63140 9054
rect 63532 9044 63588 10446
rect 63644 10164 63700 11342
rect 63644 10098 63700 10108
rect 63756 9828 63812 12126
rect 64316 9828 64372 9838
rect 63756 9826 64372 9828
rect 63756 9774 64318 9826
rect 64370 9774 64372 9826
rect 63756 9772 64372 9774
rect 63084 9042 63588 9044
rect 63084 8990 63086 9042
rect 63138 8990 63588 9042
rect 63084 8988 63588 8990
rect 61964 8260 62020 8270
rect 61964 8166 62020 8204
rect 63084 8036 63140 8988
rect 63084 7970 63140 7980
rect 63868 8146 63924 8158
rect 63868 8094 63870 8146
rect 63922 8094 63924 8146
rect 62768 7868 63448 7878
rect 62824 7812 62872 7868
rect 62928 7866 62976 7868
rect 63032 7866 63080 7868
rect 62948 7814 62976 7866
rect 63072 7814 63080 7866
rect 62928 7812 62976 7814
rect 63032 7812 63080 7814
rect 63136 7866 63184 7868
rect 63240 7866 63288 7868
rect 63136 7814 63144 7866
rect 63240 7814 63268 7866
rect 63136 7812 63184 7814
rect 63240 7812 63288 7814
rect 63344 7812 63392 7868
rect 62768 7802 63448 7812
rect 62188 7586 62244 7598
rect 62188 7534 62190 7586
rect 62242 7534 62244 7586
rect 62188 6356 62244 7534
rect 62188 6290 62244 6300
rect 62412 6692 62468 6702
rect 62636 6692 62692 6702
rect 62076 5908 62132 5918
rect 61852 5906 62132 5908
rect 61852 5854 62078 5906
rect 62130 5854 62132 5906
rect 61852 5852 62132 5854
rect 61852 4338 61908 5852
rect 62076 5842 62132 5852
rect 62412 5794 62468 6636
rect 62524 6636 62636 6692
rect 62524 5906 62580 6636
rect 62636 6626 62692 6636
rect 62768 6300 63448 6310
rect 62824 6244 62872 6300
rect 62928 6298 62976 6300
rect 63032 6298 63080 6300
rect 62948 6246 62976 6298
rect 63072 6246 63080 6298
rect 62928 6244 62976 6246
rect 63032 6244 63080 6246
rect 63136 6298 63184 6300
rect 63240 6298 63288 6300
rect 63136 6246 63144 6298
rect 63240 6246 63268 6298
rect 63136 6244 63184 6246
rect 63240 6244 63288 6246
rect 63344 6244 63392 6300
rect 62768 6234 63448 6244
rect 63756 6020 63812 6030
rect 62524 5854 62526 5906
rect 62578 5854 62580 5906
rect 62524 5842 62580 5854
rect 62860 6018 63812 6020
rect 62860 5966 63758 6018
rect 63810 5966 63812 6018
rect 62860 5964 63812 5966
rect 62860 5906 62916 5964
rect 63756 5954 63812 5964
rect 63868 6018 63924 8094
rect 64316 6802 64372 9772
rect 64652 7474 64708 7486
rect 64652 7422 64654 7474
rect 64706 7422 64708 7474
rect 64316 6750 64318 6802
rect 64370 6750 64372 6802
rect 64316 6738 64372 6750
rect 64428 7140 64484 7150
rect 63868 5966 63870 6018
rect 63922 5966 63924 6018
rect 63868 5954 63924 5966
rect 62860 5854 62862 5906
rect 62914 5854 62916 5906
rect 62860 5842 62916 5854
rect 64428 5906 64484 7084
rect 64428 5854 64430 5906
rect 64482 5854 64484 5906
rect 64428 5842 64484 5854
rect 62412 5742 62414 5794
rect 62466 5742 62468 5794
rect 62412 5730 62468 5742
rect 64652 5348 64708 7422
rect 64652 5282 64708 5292
rect 62768 4732 63448 4742
rect 62824 4676 62872 4732
rect 62928 4730 62976 4732
rect 63032 4730 63080 4732
rect 62948 4678 62976 4730
rect 63072 4678 63080 4730
rect 62928 4676 62976 4678
rect 63032 4676 63080 4678
rect 63136 4730 63184 4732
rect 63240 4730 63288 4732
rect 63136 4678 63144 4730
rect 63240 4678 63268 4730
rect 63136 4676 63184 4678
rect 63240 4676 63288 4678
rect 63344 4676 63392 4732
rect 62768 4666 63448 4676
rect 63196 4564 63252 4574
rect 62860 4508 63196 4564
rect 62748 4452 62804 4462
rect 62748 4358 62804 4396
rect 61852 4286 61854 4338
rect 61906 4286 61908 4338
rect 61852 4274 61908 4286
rect 62188 4228 62244 4238
rect 62188 4134 62244 4172
rect 60844 3780 60900 3790
rect 60844 3686 60900 3724
rect 60732 3668 60788 3678
rect 60732 3574 60788 3612
rect 61740 3666 61796 3836
rect 61740 3614 61742 3666
rect 61794 3614 61796 3666
rect 61740 3602 61796 3614
rect 62748 3668 62804 3678
rect 62860 3668 62916 4508
rect 63196 4470 63252 4508
rect 65324 4564 65380 15092
rect 67268 14924 67948 14934
rect 67324 14868 67372 14924
rect 67428 14922 67476 14924
rect 67532 14922 67580 14924
rect 67448 14870 67476 14922
rect 67572 14870 67580 14922
rect 67428 14868 67476 14870
rect 67532 14868 67580 14870
rect 67636 14922 67684 14924
rect 67740 14922 67788 14924
rect 67636 14870 67644 14922
rect 67740 14870 67768 14922
rect 67636 14868 67684 14870
rect 67740 14868 67788 14870
rect 67844 14868 67892 14924
rect 67268 14858 67948 14868
rect 68348 14532 68404 14542
rect 68236 14476 68348 14532
rect 65548 13748 65604 13758
rect 65548 10834 65604 13692
rect 67268 13356 67948 13366
rect 67324 13300 67372 13356
rect 67428 13354 67476 13356
rect 67532 13354 67580 13356
rect 67448 13302 67476 13354
rect 67572 13302 67580 13354
rect 67428 13300 67476 13302
rect 67532 13300 67580 13302
rect 67636 13354 67684 13356
rect 67740 13354 67788 13356
rect 67636 13302 67644 13354
rect 67740 13302 67768 13354
rect 67636 13300 67684 13302
rect 67740 13300 67788 13302
rect 67844 13300 67892 13356
rect 67268 13290 67948 13300
rect 66108 12964 66164 12974
rect 66108 12962 66612 12964
rect 66108 12910 66110 12962
rect 66162 12910 66612 12962
rect 66108 12908 66612 12910
rect 66108 12898 66164 12908
rect 66556 12738 66612 12908
rect 66556 12686 66558 12738
rect 66610 12686 66612 12738
rect 65548 10782 65550 10834
rect 65602 10782 65604 10834
rect 65548 10770 65604 10782
rect 65772 11396 65828 11406
rect 65548 8930 65604 8942
rect 65548 8878 65550 8930
rect 65602 8878 65604 8930
rect 65548 6692 65604 8878
rect 65548 6626 65604 6636
rect 65436 6580 65492 6590
rect 65436 5122 65492 6524
rect 65436 5070 65438 5122
rect 65490 5070 65492 5122
rect 65436 5058 65492 5070
rect 65324 4498 65380 4508
rect 63532 4450 63588 4462
rect 63532 4398 63534 4450
rect 63586 4398 63588 4450
rect 63532 3780 63588 4398
rect 65772 4450 65828 11340
rect 65772 4398 65774 4450
rect 65826 4398 65828 4450
rect 65772 4386 65828 4398
rect 65996 10164 66052 10174
rect 63532 3714 63588 3724
rect 62804 3612 62916 3668
rect 62748 3574 62804 3612
rect 60508 3390 60510 3442
rect 60562 3390 60564 3442
rect 60508 3378 60564 3390
rect 61292 3556 61348 3566
rect 61292 3388 61348 3500
rect 63196 3556 63252 3566
rect 63196 3462 63252 3500
rect 65996 3556 66052 10108
rect 66220 8260 66276 8270
rect 66556 8260 66612 12686
rect 67900 12180 67956 12190
rect 67900 12178 68180 12180
rect 67900 12126 67902 12178
rect 67954 12126 68180 12178
rect 67900 12124 68180 12126
rect 67900 12114 67956 12124
rect 67268 11788 67948 11798
rect 67324 11732 67372 11788
rect 67428 11786 67476 11788
rect 67532 11786 67580 11788
rect 67448 11734 67476 11786
rect 67572 11734 67580 11786
rect 67428 11732 67476 11734
rect 67532 11732 67580 11734
rect 67636 11786 67684 11788
rect 67740 11786 67788 11788
rect 67636 11734 67644 11786
rect 67740 11734 67768 11786
rect 67636 11732 67684 11734
rect 67740 11732 67788 11734
rect 67844 11732 67892 11788
rect 67268 11722 67948 11732
rect 67564 11620 67620 11630
rect 67564 11526 67620 11564
rect 67268 10220 67948 10230
rect 67324 10164 67372 10220
rect 67428 10218 67476 10220
rect 67532 10218 67580 10220
rect 67448 10166 67476 10218
rect 67572 10166 67580 10218
rect 67428 10164 67476 10166
rect 67532 10164 67580 10166
rect 67636 10218 67684 10220
rect 67740 10218 67788 10220
rect 67636 10166 67644 10218
rect 67740 10166 67768 10218
rect 67636 10164 67684 10166
rect 67740 10164 67788 10166
rect 67844 10164 67892 10220
rect 67268 10154 67948 10164
rect 67268 8652 67948 8662
rect 67324 8596 67372 8652
rect 67428 8650 67476 8652
rect 67532 8650 67580 8652
rect 67448 8598 67476 8650
rect 67572 8598 67580 8650
rect 67428 8596 67476 8598
rect 67532 8596 67580 8598
rect 67636 8650 67684 8652
rect 67740 8650 67788 8652
rect 67636 8598 67644 8650
rect 67740 8598 67768 8650
rect 67636 8596 67684 8598
rect 67740 8596 67788 8598
rect 67844 8596 67892 8652
rect 67268 8586 67948 8596
rect 66276 8204 66612 8260
rect 66220 8034 66276 8204
rect 66220 7982 66222 8034
rect 66274 7982 66276 8034
rect 66220 7924 66276 7982
rect 66220 7858 66276 7868
rect 66444 7588 66500 7598
rect 66444 7494 66500 7532
rect 68124 7140 68180 12124
rect 67268 7084 67948 7094
rect 67324 7028 67372 7084
rect 67428 7082 67476 7084
rect 67532 7082 67580 7084
rect 67448 7030 67476 7082
rect 67572 7030 67580 7082
rect 67428 7028 67476 7030
rect 67532 7028 67580 7030
rect 67636 7082 67684 7084
rect 67740 7082 67788 7084
rect 67636 7030 67644 7082
rect 67740 7030 67768 7082
rect 67636 7028 67684 7030
rect 67740 7028 67788 7030
rect 67844 7028 67892 7084
rect 68124 7074 68180 7084
rect 67268 7018 67948 7028
rect 67268 5516 67948 5526
rect 67324 5460 67372 5516
rect 67428 5514 67476 5516
rect 67532 5514 67580 5516
rect 67448 5462 67476 5514
rect 67572 5462 67580 5514
rect 67428 5460 67476 5462
rect 67532 5460 67580 5462
rect 67636 5514 67684 5516
rect 67740 5514 67788 5516
rect 67636 5462 67644 5514
rect 67740 5462 67768 5514
rect 67636 5460 67684 5462
rect 67740 5460 67788 5462
rect 67844 5460 67892 5516
rect 68236 5460 68292 14476
rect 68348 14466 68404 14476
rect 70028 14532 70084 14542
rect 70028 14438 70084 14476
rect 70588 14418 70644 14430
rect 70588 14366 70590 14418
rect 70642 14366 70644 14418
rect 67268 5450 67948 5460
rect 68124 5404 68292 5460
rect 68348 13748 68404 13758
rect 68348 11620 68404 13692
rect 69692 12850 69748 12862
rect 69692 12798 69694 12850
rect 69746 12798 69748 12850
rect 67788 5348 67844 5358
rect 68124 5348 68180 5404
rect 68348 5348 68404 11564
rect 67788 5346 68180 5348
rect 67788 5294 67790 5346
rect 67842 5294 68180 5346
rect 67788 5292 68180 5294
rect 68236 5292 68404 5348
rect 68460 12290 68516 12302
rect 68460 12238 68462 12290
rect 68514 12238 68516 12290
rect 67788 5282 67844 5292
rect 67340 5122 67396 5134
rect 67340 5070 67342 5122
rect 67394 5070 67396 5122
rect 67340 5012 67396 5070
rect 67340 4946 67396 4956
rect 68236 5012 68292 5292
rect 68348 5124 68404 5134
rect 68348 5030 68404 5068
rect 68236 4946 68292 4956
rect 67268 3948 67948 3958
rect 67324 3892 67372 3948
rect 67428 3946 67476 3948
rect 67532 3946 67580 3948
rect 67448 3894 67476 3946
rect 67572 3894 67580 3946
rect 67428 3892 67476 3894
rect 67532 3892 67580 3894
rect 67636 3946 67684 3948
rect 67740 3946 67788 3948
rect 67636 3894 67644 3946
rect 67740 3894 67768 3946
rect 67636 3892 67684 3894
rect 67740 3892 67788 3894
rect 67844 3892 67892 3948
rect 67268 3882 67948 3892
rect 68460 3780 68516 12238
rect 69692 12178 69748 12798
rect 69692 12126 69694 12178
rect 69746 12126 69748 12178
rect 69692 12114 69748 12126
rect 70140 12066 70196 12078
rect 70140 12014 70142 12066
rect 70194 12014 70196 12066
rect 69692 10610 69748 10622
rect 69692 10558 69694 10610
rect 69746 10558 69748 10610
rect 68908 9042 68964 9054
rect 68908 8990 68910 9042
rect 68962 8990 68964 9042
rect 68796 6020 68852 6030
rect 68908 6020 68964 8990
rect 69020 8258 69076 8270
rect 69020 8206 69022 8258
rect 69074 8206 69076 8258
rect 69020 6580 69076 8206
rect 69020 6486 69076 6524
rect 68796 6018 68964 6020
rect 68796 5966 68798 6018
rect 68850 5966 68964 6018
rect 68796 5964 68964 5966
rect 68796 5954 68852 5964
rect 68908 4338 68964 5964
rect 69692 6020 69748 10558
rect 70140 7028 70196 12014
rect 70140 6962 70196 6972
rect 70364 7362 70420 7374
rect 70364 7310 70366 7362
rect 70418 7310 70420 7362
rect 70364 6804 70420 7310
rect 69692 5954 69748 5964
rect 69916 6748 70420 6804
rect 68908 4286 68910 4338
rect 68962 4286 68964 4338
rect 68908 4274 68964 4286
rect 68460 3714 68516 3724
rect 69580 3780 69636 3790
rect 69580 3686 69636 3724
rect 67452 3666 67508 3678
rect 67452 3614 67454 3666
rect 67506 3614 67508 3666
rect 66444 3556 66500 3566
rect 65996 3554 66500 3556
rect 65996 3502 65998 3554
rect 66050 3502 66446 3554
rect 66498 3502 66500 3554
rect 65996 3500 66500 3502
rect 65996 3490 66052 3500
rect 66444 3490 66500 3500
rect 60956 3332 61348 3388
rect 67452 3444 67508 3614
rect 67452 3378 67508 3388
rect 69692 3444 69748 3482
rect 69916 3444 69972 6748
rect 70588 6692 70644 14366
rect 70700 13860 70756 22876
rect 71372 20580 71428 20590
rect 71036 20130 71092 20142
rect 71036 20078 71038 20130
rect 71090 20078 71092 20130
rect 70924 19236 70980 19246
rect 71036 19236 71092 20078
rect 70924 19234 71092 19236
rect 70924 19182 70926 19234
rect 70978 19182 71092 19234
rect 70924 19180 71092 19182
rect 71372 19234 71428 20524
rect 71372 19182 71374 19234
rect 71426 19182 71428 19234
rect 70924 19170 70980 19180
rect 71372 19170 71428 19182
rect 71484 19124 71540 23662
rect 73500 23716 73556 23726
rect 71768 23548 72448 23558
rect 71824 23492 71872 23548
rect 71928 23546 71976 23548
rect 72032 23546 72080 23548
rect 71948 23494 71976 23546
rect 72072 23494 72080 23546
rect 71928 23492 71976 23494
rect 72032 23492 72080 23494
rect 72136 23546 72184 23548
rect 72240 23546 72288 23548
rect 72136 23494 72144 23546
rect 72240 23494 72268 23546
rect 72136 23492 72184 23494
rect 72240 23492 72288 23494
rect 72344 23492 72392 23548
rect 71768 23482 72448 23492
rect 73500 23378 73556 23660
rect 73500 23326 73502 23378
rect 73554 23326 73556 23378
rect 73500 23314 73556 23326
rect 72156 23268 72212 23278
rect 72156 22370 72212 23212
rect 72940 23268 72996 23278
rect 72940 23174 72996 23212
rect 73724 23268 73780 23278
rect 73612 23042 73668 23054
rect 73612 22990 73614 23042
rect 73666 22990 73668 23042
rect 73612 22708 73668 22990
rect 72156 22318 72158 22370
rect 72210 22318 72212 22370
rect 72156 22306 72212 22318
rect 72716 22652 73668 22708
rect 72716 22370 72772 22652
rect 73724 22484 73780 23212
rect 74508 23268 74564 23278
rect 74508 23174 74564 23212
rect 74172 23156 74228 23166
rect 74172 23154 74452 23156
rect 74172 23102 74174 23154
rect 74226 23102 74452 23154
rect 74172 23100 74452 23102
rect 74172 23090 74228 23100
rect 73724 22418 73780 22428
rect 72716 22318 72718 22370
rect 72770 22318 72772 22370
rect 72716 22306 72772 22318
rect 74396 22372 74452 23100
rect 75068 22484 75124 22494
rect 74396 22316 75012 22372
rect 74844 22036 74900 22046
rect 71768 21980 72448 21990
rect 71824 21924 71872 21980
rect 71928 21978 71976 21980
rect 72032 21978 72080 21980
rect 71948 21926 71976 21978
rect 72072 21926 72080 21978
rect 71928 21924 71976 21926
rect 72032 21924 72080 21926
rect 72136 21978 72184 21980
rect 72240 21978 72288 21980
rect 72136 21926 72144 21978
rect 72240 21926 72268 21978
rect 72136 21924 72184 21926
rect 72240 21924 72288 21926
rect 72344 21924 72392 21980
rect 71768 21914 72448 21924
rect 73500 21588 73556 21598
rect 72044 20804 72100 20814
rect 72044 20710 72100 20748
rect 72716 20804 72772 20814
rect 72716 20802 73220 20804
rect 72716 20750 72718 20802
rect 72770 20750 73220 20802
rect 72716 20748 73220 20750
rect 72716 20738 72772 20748
rect 72156 20580 72212 20618
rect 72156 20514 72212 20524
rect 72268 20580 72324 20590
rect 72492 20580 72548 20590
rect 72268 20578 72492 20580
rect 72268 20526 72270 20578
rect 72322 20526 72492 20578
rect 72268 20524 72492 20526
rect 72268 20514 72324 20524
rect 72492 20514 72548 20524
rect 73052 20580 73108 20590
rect 73052 20486 73108 20524
rect 71768 20412 72448 20422
rect 71824 20356 71872 20412
rect 71928 20410 71976 20412
rect 72032 20410 72080 20412
rect 71948 20358 71976 20410
rect 72072 20358 72080 20410
rect 71928 20356 71976 20358
rect 72032 20356 72080 20358
rect 72136 20410 72184 20412
rect 72240 20410 72288 20412
rect 72136 20358 72144 20410
rect 72240 20358 72268 20410
rect 72136 20356 72184 20358
rect 72240 20356 72288 20358
rect 72344 20356 72392 20412
rect 71768 20346 72448 20356
rect 73164 20242 73220 20748
rect 73164 20190 73166 20242
rect 73218 20190 73220 20242
rect 73164 20178 73220 20190
rect 73388 20132 73444 20142
rect 73388 20038 73444 20076
rect 73500 20130 73556 21532
rect 74844 21026 74900 21980
rect 74956 21810 75012 22316
rect 75068 22146 75124 22428
rect 75068 22094 75070 22146
rect 75122 22094 75124 22146
rect 75068 22082 75124 22094
rect 75180 21924 75236 27692
rect 74956 21758 74958 21810
rect 75010 21758 75012 21810
rect 74956 21746 75012 21758
rect 75068 21868 75236 21924
rect 75292 26962 75348 26974
rect 75292 26910 75294 26962
rect 75346 26910 75348 26962
rect 75068 21588 75124 21868
rect 75180 21700 75236 21710
rect 75180 21606 75236 21644
rect 74844 20974 74846 21026
rect 74898 20974 74900 21026
rect 74844 20962 74900 20974
rect 74956 21532 75124 21588
rect 75292 21588 75348 26910
rect 75404 22372 75460 28588
rect 75740 28082 75796 32172
rect 76324 32116 76372 32172
rect 76428 32170 76476 32172
rect 76532 32170 76580 32172
rect 76448 32118 76476 32170
rect 76572 32118 76580 32170
rect 76428 32116 76476 32118
rect 76532 32116 76580 32118
rect 76636 32170 76684 32172
rect 76740 32170 76788 32172
rect 76636 32118 76644 32170
rect 76740 32118 76768 32170
rect 76636 32116 76684 32118
rect 76740 32116 76788 32118
rect 76844 32116 76892 32172
rect 76268 32106 76948 32116
rect 80768 31388 81448 31398
rect 80824 31332 80872 31388
rect 80928 31386 80976 31388
rect 81032 31386 81080 31388
rect 80948 31334 80976 31386
rect 81072 31334 81080 31386
rect 80928 31332 80976 31334
rect 81032 31332 81080 31334
rect 81136 31386 81184 31388
rect 81240 31386 81288 31388
rect 81136 31334 81144 31386
rect 81240 31334 81268 31386
rect 81136 31332 81184 31334
rect 81240 31332 81288 31334
rect 81344 31332 81392 31388
rect 80768 31322 81448 31332
rect 76268 30604 76948 30614
rect 76324 30548 76372 30604
rect 76428 30602 76476 30604
rect 76532 30602 76580 30604
rect 76448 30550 76476 30602
rect 76572 30550 76580 30602
rect 76428 30548 76476 30550
rect 76532 30548 76580 30550
rect 76636 30602 76684 30604
rect 76740 30602 76788 30604
rect 76636 30550 76644 30602
rect 76740 30550 76768 30602
rect 76636 30548 76684 30550
rect 76740 30548 76788 30550
rect 76844 30548 76892 30604
rect 76268 30538 76948 30548
rect 85148 30322 85204 35308
rect 85268 35308 85948 35318
rect 85324 35252 85372 35308
rect 85428 35306 85476 35308
rect 85532 35306 85580 35308
rect 85448 35254 85476 35306
rect 85572 35254 85580 35306
rect 85428 35252 85476 35254
rect 85532 35252 85580 35254
rect 85636 35306 85684 35308
rect 85740 35306 85788 35308
rect 85636 35254 85644 35306
rect 85740 35254 85768 35306
rect 85636 35252 85684 35254
rect 85740 35252 85788 35254
rect 85844 35252 85892 35308
rect 85268 35242 85948 35252
rect 85372 35140 85428 35150
rect 85372 34354 85428 35084
rect 85372 34302 85374 34354
rect 85426 34302 85428 34354
rect 85372 34244 85428 34302
rect 85820 34804 85876 34814
rect 85820 34354 85876 34748
rect 85820 34302 85822 34354
rect 85874 34302 85876 34354
rect 85820 34290 85876 34302
rect 85372 34178 85428 34188
rect 85932 34244 85988 34254
rect 85932 34150 85988 34188
rect 85820 33908 85876 33918
rect 86156 33908 86212 35644
rect 89964 35700 90020 35710
rect 89068 35586 89124 35598
rect 89068 35534 89070 35586
rect 89122 35534 89124 35586
rect 89068 35476 89124 35534
rect 89516 35476 89572 35486
rect 89068 35474 89572 35476
rect 89068 35422 89518 35474
rect 89570 35422 89572 35474
rect 89068 35420 89572 35422
rect 89068 34916 89124 35420
rect 89516 35410 89572 35420
rect 89964 35026 90020 35644
rect 90300 35700 90356 35710
rect 90636 35700 90692 37324
rect 90860 36258 90916 36270
rect 90860 36206 90862 36258
rect 90914 36206 90916 36258
rect 90300 35698 90692 35700
rect 90300 35646 90302 35698
rect 90354 35646 90692 35698
rect 90300 35644 90692 35646
rect 90748 35700 90804 35710
rect 90860 35700 90916 36206
rect 90748 35698 90916 35700
rect 90748 35646 90750 35698
rect 90802 35646 90916 35698
rect 90748 35644 90916 35646
rect 91308 36260 91364 38892
rect 91644 38834 91700 40124
rect 91756 39396 91812 40348
rect 91868 40402 91924 40414
rect 91868 40350 91870 40402
rect 91922 40350 91924 40402
rect 91868 39508 91924 40350
rect 92204 40402 92260 40572
rect 94780 40626 94836 41020
rect 94780 40574 94782 40626
rect 94834 40574 94836 40626
rect 94780 40516 94836 40574
rect 94780 40450 94836 40460
rect 92204 40350 92206 40402
rect 92258 40350 92260 40402
rect 92204 40338 92260 40350
rect 95340 40404 95396 40414
rect 95340 40310 95396 40348
rect 96124 40404 96180 42588
rect 96236 42578 96292 42588
rect 96236 41074 96292 41086
rect 96236 41022 96238 41074
rect 96290 41022 96292 41074
rect 96236 40628 96292 41022
rect 96236 40562 96292 40572
rect 96124 40338 96180 40348
rect 96236 40402 96292 40414
rect 96236 40350 96238 40402
rect 96290 40350 96292 40402
rect 94268 40012 94948 40022
rect 94324 39956 94372 40012
rect 94428 40010 94476 40012
rect 94532 40010 94580 40012
rect 94448 39958 94476 40010
rect 94572 39958 94580 40010
rect 94428 39956 94476 39958
rect 94532 39956 94580 39958
rect 94636 40010 94684 40012
rect 94740 40010 94788 40012
rect 94636 39958 94644 40010
rect 94740 39958 94768 40010
rect 94636 39956 94684 39958
rect 94740 39956 94788 39958
rect 94844 39956 94892 40012
rect 94268 39946 94948 39956
rect 92092 39508 92148 39518
rect 91868 39506 92148 39508
rect 91868 39454 92094 39506
rect 92146 39454 92148 39506
rect 91868 39452 92148 39454
rect 92092 39442 92148 39452
rect 96236 39396 96292 40350
rect 91756 39340 92036 39396
rect 91980 39058 92036 39340
rect 96236 39330 96292 39340
rect 91980 39006 91982 39058
rect 92034 39006 92036 39058
rect 91980 38994 92036 39006
rect 91644 38782 91646 38834
rect 91698 38782 91700 38834
rect 91644 38770 91700 38782
rect 94268 38444 94948 38454
rect 94324 38388 94372 38444
rect 94428 38442 94476 38444
rect 94532 38442 94580 38444
rect 94448 38390 94476 38442
rect 94572 38390 94580 38442
rect 94428 38388 94476 38390
rect 94532 38388 94580 38390
rect 94636 38442 94684 38444
rect 94740 38442 94788 38444
rect 94636 38390 94644 38442
rect 94740 38390 94768 38442
rect 94636 38388 94684 38390
rect 94740 38388 94788 38390
rect 94844 38388 94892 38444
rect 94268 38378 94948 38388
rect 96236 37938 96292 37950
rect 96236 37886 96238 37938
rect 96290 37886 96292 37938
rect 96124 37266 96180 37278
rect 96124 37214 96126 37266
rect 96178 37214 96180 37266
rect 94268 36876 94948 36886
rect 94324 36820 94372 36876
rect 94428 36874 94476 36876
rect 94532 36874 94580 36876
rect 94448 36822 94476 36874
rect 94572 36822 94580 36874
rect 94428 36820 94476 36822
rect 94532 36820 94580 36822
rect 94636 36874 94684 36876
rect 94740 36874 94788 36876
rect 94636 36822 94644 36874
rect 94740 36822 94768 36874
rect 94636 36820 94684 36822
rect 94740 36820 94788 36822
rect 94844 36820 94892 36876
rect 94268 36810 94948 36820
rect 92204 36484 92260 36494
rect 91756 36482 92260 36484
rect 91756 36430 92206 36482
rect 92258 36430 92260 36482
rect 91756 36428 92260 36430
rect 91756 36260 91812 36428
rect 92204 36418 92260 36428
rect 92428 36482 92484 36494
rect 92428 36430 92430 36482
rect 92482 36430 92484 36482
rect 91308 36258 91812 36260
rect 91308 36206 91310 36258
rect 91362 36206 91812 36258
rect 91308 36204 91812 36206
rect 91868 36260 91924 36270
rect 90300 35634 90356 35644
rect 90748 35634 90804 35644
rect 89964 34974 89966 35026
rect 90018 34974 90020 35026
rect 89964 34962 90020 34974
rect 89068 34850 89124 34860
rect 88172 34804 88228 34814
rect 88172 34710 88228 34748
rect 87388 34690 87444 34702
rect 87388 34638 87390 34690
rect 87442 34638 87444 34690
rect 87388 34356 87444 34638
rect 89768 34524 90448 34534
rect 89824 34468 89872 34524
rect 89928 34522 89976 34524
rect 90032 34522 90080 34524
rect 89948 34470 89976 34522
rect 90072 34470 90080 34522
rect 89928 34468 89976 34470
rect 90032 34468 90080 34470
rect 90136 34522 90184 34524
rect 90240 34522 90288 34524
rect 90136 34470 90144 34522
rect 90240 34470 90268 34522
rect 90136 34468 90184 34470
rect 90240 34468 90288 34470
rect 90344 34468 90392 34524
rect 89768 34458 90448 34468
rect 87388 34290 87444 34300
rect 85820 33906 86212 33908
rect 85820 33854 85822 33906
rect 85874 33854 86212 33906
rect 85820 33852 86212 33854
rect 85820 33842 85876 33852
rect 85268 33740 85948 33750
rect 85324 33684 85372 33740
rect 85428 33738 85476 33740
rect 85532 33738 85580 33740
rect 85448 33686 85476 33738
rect 85572 33686 85580 33738
rect 85428 33684 85476 33686
rect 85532 33684 85580 33686
rect 85636 33738 85684 33740
rect 85740 33738 85788 33740
rect 85636 33686 85644 33738
rect 85740 33686 85768 33738
rect 85636 33684 85684 33686
rect 85740 33684 85788 33686
rect 85844 33684 85892 33740
rect 85268 33674 85948 33684
rect 89768 32956 90448 32966
rect 89824 32900 89872 32956
rect 89928 32954 89976 32956
rect 90032 32954 90080 32956
rect 89948 32902 89976 32954
rect 90072 32902 90080 32954
rect 89928 32900 89976 32902
rect 90032 32900 90080 32902
rect 90136 32954 90184 32956
rect 90240 32954 90288 32956
rect 90136 32902 90144 32954
rect 90240 32902 90268 32954
rect 90136 32900 90184 32902
rect 90240 32900 90288 32902
rect 90344 32900 90392 32956
rect 89768 32890 90448 32900
rect 85268 32172 85948 32182
rect 85324 32116 85372 32172
rect 85428 32170 85476 32172
rect 85532 32170 85580 32172
rect 85448 32118 85476 32170
rect 85572 32118 85580 32170
rect 85428 32116 85476 32118
rect 85532 32116 85580 32118
rect 85636 32170 85684 32172
rect 85740 32170 85788 32172
rect 85636 32118 85644 32170
rect 85740 32118 85768 32170
rect 85636 32116 85684 32118
rect 85740 32116 85788 32118
rect 85844 32116 85892 32172
rect 85268 32106 85948 32116
rect 89768 31388 90448 31398
rect 89824 31332 89872 31388
rect 89928 31386 89976 31388
rect 90032 31386 90080 31388
rect 89948 31334 89976 31386
rect 90072 31334 90080 31386
rect 89928 31332 89976 31334
rect 90032 31332 90080 31334
rect 90136 31386 90184 31388
rect 90240 31386 90288 31388
rect 90136 31334 90144 31386
rect 90240 31334 90268 31386
rect 90136 31332 90184 31334
rect 90240 31332 90288 31334
rect 90344 31332 90392 31388
rect 89768 31322 90448 31332
rect 85268 30604 85948 30614
rect 85324 30548 85372 30604
rect 85428 30602 85476 30604
rect 85532 30602 85580 30604
rect 85448 30550 85476 30602
rect 85572 30550 85580 30602
rect 85428 30548 85476 30550
rect 85532 30548 85580 30550
rect 85636 30602 85684 30604
rect 85740 30602 85788 30604
rect 85636 30550 85644 30602
rect 85740 30550 85768 30602
rect 85636 30548 85684 30550
rect 85740 30548 85788 30550
rect 85844 30548 85892 30604
rect 85268 30538 85948 30548
rect 85148 30270 85150 30322
rect 85202 30270 85204 30322
rect 85148 30258 85204 30270
rect 77420 30212 77476 30222
rect 75852 29428 75908 29438
rect 75852 29334 75908 29372
rect 77420 29428 77476 30156
rect 83468 30212 83524 30222
rect 83468 30118 83524 30156
rect 84476 30212 84532 30222
rect 84476 30118 84532 30156
rect 91308 30212 91364 36204
rect 91868 36166 91924 36204
rect 92428 36036 92484 36430
rect 92428 35970 92484 35980
rect 92988 35924 93044 35934
rect 92988 35830 93044 35868
rect 93772 35924 93828 35934
rect 93772 35830 93828 35868
rect 96124 35924 96180 37214
rect 96236 37044 96292 37886
rect 96236 36978 96292 36988
rect 96236 36372 96292 36382
rect 96236 36278 96292 36316
rect 96124 35858 96180 35868
rect 94268 35308 94948 35318
rect 94324 35252 94372 35308
rect 94428 35306 94476 35308
rect 94532 35306 94580 35308
rect 94448 35254 94476 35306
rect 94572 35254 94580 35306
rect 94428 35252 94476 35254
rect 94532 35252 94580 35254
rect 94636 35306 94684 35308
rect 94740 35306 94788 35308
rect 94636 35254 94644 35306
rect 94740 35254 94768 35306
rect 94636 35252 94684 35254
rect 94740 35252 94788 35254
rect 94844 35252 94892 35308
rect 94268 35242 94948 35252
rect 96236 34804 96292 34814
rect 96236 34710 96292 34748
rect 94268 33740 94948 33750
rect 94324 33684 94372 33740
rect 94428 33738 94476 33740
rect 94532 33738 94580 33740
rect 94448 33686 94476 33738
rect 94572 33686 94580 33738
rect 94428 33684 94476 33686
rect 94532 33684 94580 33686
rect 94636 33738 94684 33740
rect 94740 33738 94788 33740
rect 94636 33686 94644 33738
rect 94740 33686 94768 33738
rect 94636 33684 94684 33686
rect 94740 33684 94788 33686
rect 94844 33684 94892 33740
rect 94268 33674 94948 33684
rect 94268 32172 94948 32182
rect 94324 32116 94372 32172
rect 94428 32170 94476 32172
rect 94532 32170 94580 32172
rect 94448 32118 94476 32170
rect 94572 32118 94580 32170
rect 94428 32116 94476 32118
rect 94532 32116 94580 32118
rect 94636 32170 94684 32172
rect 94740 32170 94788 32172
rect 94636 32118 94644 32170
rect 94740 32118 94768 32170
rect 94636 32116 94684 32118
rect 94740 32116 94788 32118
rect 94844 32116 94892 32172
rect 94268 32106 94948 32116
rect 94268 30604 94948 30614
rect 94324 30548 94372 30604
rect 94428 30602 94476 30604
rect 94532 30602 94580 30604
rect 94448 30550 94476 30602
rect 94572 30550 94580 30602
rect 94428 30548 94476 30550
rect 94532 30548 94580 30550
rect 94636 30602 94684 30604
rect 94740 30602 94788 30604
rect 94636 30550 94644 30602
rect 94740 30550 94768 30602
rect 94636 30548 94684 30550
rect 94740 30548 94788 30550
rect 94844 30548 94892 30604
rect 94268 30538 94948 30548
rect 91308 30146 91364 30156
rect 80768 29820 81448 29830
rect 80824 29764 80872 29820
rect 80928 29818 80976 29820
rect 81032 29818 81080 29820
rect 80948 29766 80976 29818
rect 81072 29766 81080 29818
rect 80928 29764 80976 29766
rect 81032 29764 81080 29766
rect 81136 29818 81184 29820
rect 81240 29818 81288 29820
rect 81136 29766 81144 29818
rect 81240 29766 81268 29818
rect 81136 29764 81184 29766
rect 81240 29764 81288 29766
rect 81344 29764 81392 29820
rect 80768 29754 81448 29764
rect 89768 29820 90448 29830
rect 89824 29764 89872 29820
rect 89928 29818 89976 29820
rect 90032 29818 90080 29820
rect 89948 29766 89976 29818
rect 90072 29766 90080 29818
rect 89928 29764 89976 29766
rect 90032 29764 90080 29766
rect 90136 29818 90184 29820
rect 90240 29818 90288 29820
rect 90136 29766 90144 29818
rect 90240 29766 90268 29818
rect 90136 29764 90184 29766
rect 90240 29764 90288 29766
rect 90344 29764 90392 29820
rect 89768 29754 90448 29764
rect 76268 29036 76948 29046
rect 76324 28980 76372 29036
rect 76428 29034 76476 29036
rect 76532 29034 76580 29036
rect 76448 28982 76476 29034
rect 76572 28982 76580 29034
rect 76428 28980 76476 28982
rect 76532 28980 76580 28982
rect 76636 29034 76684 29036
rect 76740 29034 76788 29036
rect 76636 28982 76644 29034
rect 76740 28982 76768 29034
rect 76636 28980 76684 28982
rect 76740 28980 76788 28982
rect 76844 28980 76892 29036
rect 76268 28970 76948 28980
rect 75740 28030 75742 28082
rect 75794 28030 75796 28082
rect 75740 26908 75796 28030
rect 76076 28868 76132 28878
rect 75964 27860 76020 27870
rect 75964 27188 76020 27804
rect 75964 27122 76020 27132
rect 76076 27076 76132 28812
rect 76748 28756 76804 28766
rect 76748 28754 77140 28756
rect 76748 28702 76750 28754
rect 76802 28702 77140 28754
rect 76748 28700 77140 28702
rect 76748 28690 76804 28700
rect 76188 28420 76244 28430
rect 76188 27858 76244 28364
rect 76188 27806 76190 27858
rect 76242 27806 76244 27858
rect 76188 27794 76244 27806
rect 76524 27860 76580 27870
rect 76524 27766 76580 27804
rect 76268 27468 76948 27478
rect 76324 27412 76372 27468
rect 76428 27466 76476 27468
rect 76532 27466 76580 27468
rect 76448 27414 76476 27466
rect 76572 27414 76580 27466
rect 76428 27412 76476 27414
rect 76532 27412 76580 27414
rect 76636 27466 76684 27468
rect 76740 27466 76788 27468
rect 76636 27414 76644 27466
rect 76740 27414 76768 27466
rect 76636 27412 76684 27414
rect 76740 27412 76788 27414
rect 76844 27412 76892 27468
rect 76268 27402 76948 27412
rect 77084 27300 77140 28700
rect 77420 28642 77476 29372
rect 85268 29036 85948 29046
rect 85324 28980 85372 29036
rect 85428 29034 85476 29036
rect 85532 29034 85580 29036
rect 85448 28982 85476 29034
rect 85572 28982 85580 29034
rect 85428 28980 85476 28982
rect 85532 28980 85580 28982
rect 85636 29034 85684 29036
rect 85740 29034 85788 29036
rect 85636 28982 85644 29034
rect 85740 28982 85768 29034
rect 85636 28980 85684 28982
rect 85740 28980 85788 28982
rect 85844 28980 85892 29036
rect 85268 28970 85948 28980
rect 94268 29036 94948 29046
rect 94324 28980 94372 29036
rect 94428 29034 94476 29036
rect 94532 29034 94580 29036
rect 94448 28982 94476 29034
rect 94572 28982 94580 29034
rect 94428 28980 94476 28982
rect 94532 28980 94580 28982
rect 94636 29034 94684 29036
rect 94740 29034 94788 29036
rect 94636 28982 94644 29034
rect 94740 28982 94768 29034
rect 94636 28980 94684 28982
rect 94740 28980 94788 28982
rect 94844 28980 94892 29036
rect 94268 28970 94948 28980
rect 77420 28590 77422 28642
rect 77474 28590 77476 28642
rect 77420 28578 77476 28590
rect 77756 28420 77812 28430
rect 77756 28326 77812 28364
rect 80768 28252 81448 28262
rect 80824 28196 80872 28252
rect 80928 28250 80976 28252
rect 81032 28250 81080 28252
rect 80948 28198 80976 28250
rect 81072 28198 81080 28250
rect 80928 28196 80976 28198
rect 81032 28196 81080 28198
rect 81136 28250 81184 28252
rect 81240 28250 81288 28252
rect 81136 28198 81144 28250
rect 81240 28198 81268 28250
rect 81136 28196 81184 28198
rect 81240 28196 81288 28198
rect 81344 28196 81392 28252
rect 80768 28186 81448 28196
rect 89768 28252 90448 28262
rect 89824 28196 89872 28252
rect 89928 28250 89976 28252
rect 90032 28250 90080 28252
rect 89948 28198 89976 28250
rect 90072 28198 90080 28250
rect 89928 28196 89976 28198
rect 90032 28196 90080 28198
rect 90136 28250 90184 28252
rect 90240 28250 90288 28252
rect 90136 28198 90144 28250
rect 90240 28198 90268 28250
rect 90136 28196 90184 28198
rect 90240 28196 90288 28198
rect 90344 28196 90392 28252
rect 89768 28186 90448 28196
rect 96348 28084 96404 43652
rect 96572 42642 96628 43652
rect 96908 42756 96964 42766
rect 96572 42590 96574 42642
rect 96626 42590 96628 42642
rect 96572 42578 96628 42590
rect 96684 42754 96964 42756
rect 96684 42702 96910 42754
rect 96962 42702 96964 42754
rect 96684 42700 96964 42702
rect 96684 41860 96740 42700
rect 96908 42690 96964 42700
rect 96572 41804 96740 41860
rect 96572 41074 96628 41804
rect 96908 41188 96964 41198
rect 96572 41022 96574 41074
rect 96626 41022 96628 41074
rect 96572 41010 96628 41022
rect 96684 41186 96964 41188
rect 96684 41134 96910 41186
rect 96962 41134 96964 41186
rect 96684 41132 96964 41134
rect 96572 40628 96628 40638
rect 96684 40628 96740 41132
rect 96908 41122 96964 41132
rect 96572 40626 96740 40628
rect 96572 40574 96574 40626
rect 96626 40574 96740 40626
rect 96572 40572 96740 40574
rect 96572 40562 96628 40572
rect 97020 40404 97076 43652
rect 98028 42642 98084 42654
rect 98028 42590 98030 42642
rect 98082 42590 98084 42642
rect 98028 42420 98084 42590
rect 98028 42354 98084 42364
rect 98028 41074 98084 41086
rect 98028 41022 98030 41074
rect 98082 41022 98084 41074
rect 98028 40628 98084 41022
rect 98028 40562 98084 40572
rect 96460 40348 97076 40404
rect 96460 37490 96516 40348
rect 96908 39620 96964 39630
rect 96572 39618 96964 39620
rect 96572 39566 96910 39618
rect 96962 39566 96964 39618
rect 96572 39564 96964 39566
rect 96572 37938 96628 39564
rect 96908 39554 96964 39564
rect 98028 39506 98084 39518
rect 98028 39454 98030 39506
rect 98082 39454 98084 39506
rect 98028 38836 98084 39454
rect 98028 38770 98084 38780
rect 96572 37886 96574 37938
rect 96626 37886 96628 37938
rect 96572 37874 96628 37886
rect 96460 37438 96462 37490
rect 96514 37438 96516 37490
rect 96460 37426 96516 37438
rect 96908 37268 96964 37278
rect 96572 37266 96964 37268
rect 96572 37214 96910 37266
rect 96962 37214 96964 37266
rect 96572 37212 96964 37214
rect 96572 36370 96628 37212
rect 96908 37202 96964 37212
rect 98028 37154 98084 37166
rect 98028 37102 98030 37154
rect 98082 37102 98084 37154
rect 98028 37044 98084 37102
rect 98028 36978 98084 36988
rect 96572 36318 96574 36370
rect 96626 36318 96628 36370
rect 96572 36306 96628 36318
rect 96908 35700 96964 35710
rect 96572 35698 96964 35700
rect 96572 35646 96910 35698
rect 96962 35646 96964 35698
rect 96572 35644 96964 35646
rect 96572 34802 96628 35644
rect 96908 35634 96964 35644
rect 97692 35474 97748 35486
rect 97692 35422 97694 35474
rect 97746 35422 97748 35474
rect 97692 35252 97748 35422
rect 97692 35186 97748 35196
rect 96572 34750 96574 34802
rect 96626 34750 96628 34802
rect 96572 34738 96628 34750
rect 96572 34132 96628 34142
rect 96572 34038 96628 34076
rect 97020 34132 97076 34142
rect 97020 34038 97076 34076
rect 97692 33906 97748 33918
rect 97692 33854 97694 33906
rect 97746 33854 97748 33906
rect 97692 33460 97748 33854
rect 97692 33394 97748 33404
rect 96908 31778 96964 31790
rect 96908 31726 96910 31778
rect 96962 31726 96964 31778
rect 96684 31556 96740 31566
rect 96908 31556 96964 31726
rect 98028 31668 98084 31678
rect 98028 31574 98084 31612
rect 96740 31500 96964 31556
rect 96684 31462 96740 31500
rect 96908 30210 96964 30222
rect 96908 30158 96910 30210
rect 96962 30158 96964 30210
rect 96684 30100 96740 30110
rect 96908 30100 96964 30158
rect 96740 30044 96964 30100
rect 98028 30098 98084 30110
rect 98028 30046 98030 30098
rect 98082 30046 98084 30098
rect 96684 30006 96740 30044
rect 98028 29876 98084 30046
rect 98028 29810 98084 29820
rect 96572 28644 96628 28654
rect 96572 28550 96628 28588
rect 97020 28644 97076 28654
rect 97020 28550 97076 28588
rect 97692 28642 97748 28654
rect 97692 28590 97694 28642
rect 97746 28590 97748 28642
rect 96348 28018 96404 28028
rect 97692 28084 97748 28590
rect 97692 28018 97748 28028
rect 78876 27970 78932 27982
rect 78876 27918 78878 27970
rect 78930 27918 78932 27970
rect 76524 27244 77140 27300
rect 77532 27636 77588 27646
rect 76412 27188 76468 27198
rect 76412 27094 76468 27132
rect 76300 27076 76356 27086
rect 76076 27074 76356 27076
rect 76076 27022 76302 27074
rect 76354 27022 76356 27074
rect 76076 27020 76356 27022
rect 76300 27010 76356 27020
rect 75740 26852 76020 26908
rect 75740 26180 75796 26190
rect 75740 26086 75796 26124
rect 75964 26180 76020 26852
rect 76524 26850 76580 27244
rect 76972 27076 77028 27086
rect 77308 27076 77364 27086
rect 76972 27074 77364 27076
rect 76972 27022 76974 27074
rect 77026 27022 77310 27074
rect 77362 27022 77364 27074
rect 76972 27020 77364 27022
rect 76972 27010 77028 27020
rect 77308 27010 77364 27020
rect 77532 26962 77588 27580
rect 77532 26910 77534 26962
rect 77586 26910 77588 26962
rect 77532 26898 77588 26910
rect 77644 26962 77700 26974
rect 77644 26910 77646 26962
rect 77698 26910 77700 26962
rect 77644 26908 77700 26910
rect 78092 26962 78148 26974
rect 78092 26910 78094 26962
rect 78146 26910 78148 26962
rect 78092 26908 78148 26910
rect 76524 26798 76526 26850
rect 76578 26798 76580 26850
rect 76524 26404 76580 26798
rect 77644 26852 78148 26908
rect 76524 26338 76580 26348
rect 77084 26404 77140 26414
rect 77140 26348 77588 26404
rect 77084 26310 77140 26348
rect 75964 25508 76020 26124
rect 76076 26068 76132 26078
rect 76076 25730 76132 26012
rect 76268 25900 76948 25910
rect 76324 25844 76372 25900
rect 76428 25898 76476 25900
rect 76532 25898 76580 25900
rect 76448 25846 76476 25898
rect 76572 25846 76580 25898
rect 76428 25844 76476 25846
rect 76532 25844 76580 25846
rect 76636 25898 76684 25900
rect 76740 25898 76788 25900
rect 76636 25846 76644 25898
rect 76740 25846 76768 25898
rect 76636 25844 76684 25846
rect 76740 25844 76788 25846
rect 76844 25844 76892 25900
rect 76268 25834 76948 25844
rect 76076 25678 76078 25730
rect 76130 25678 76132 25730
rect 76076 25666 76132 25678
rect 76748 25730 76804 25742
rect 76748 25678 76750 25730
rect 76802 25678 76804 25730
rect 76748 25618 76804 25678
rect 77084 25732 77140 25742
rect 77084 25730 77364 25732
rect 77084 25678 77086 25730
rect 77138 25678 77364 25730
rect 77084 25676 77364 25678
rect 77084 25666 77140 25676
rect 76748 25566 76750 25618
rect 76802 25566 76804 25618
rect 76748 25554 76804 25566
rect 76300 25508 76356 25518
rect 75964 25506 76356 25508
rect 75964 25454 76302 25506
rect 76354 25454 76356 25506
rect 75964 25452 76356 25454
rect 75964 25396 76020 25452
rect 76300 25442 76356 25452
rect 77308 25506 77364 25676
rect 77308 25454 77310 25506
rect 77362 25454 77364 25506
rect 77308 25442 77364 25454
rect 77420 25508 77476 25518
rect 77420 25414 77476 25452
rect 77532 25506 77588 26348
rect 77644 26292 77700 26852
rect 77700 26236 77812 26292
rect 77644 26226 77700 26236
rect 77532 25454 77534 25506
rect 77586 25454 77588 25506
rect 75740 25282 75796 25294
rect 75740 25230 75742 25282
rect 75794 25230 75796 25282
rect 75740 24836 75796 25230
rect 75740 23940 75796 24780
rect 75740 23874 75796 23884
rect 75964 22596 76020 25340
rect 77532 25284 77588 25454
rect 76972 25228 77588 25284
rect 76972 24946 77028 25228
rect 76972 24894 76974 24946
rect 77026 24894 77028 24946
rect 76972 24882 77028 24894
rect 76268 24332 76948 24342
rect 76324 24276 76372 24332
rect 76428 24330 76476 24332
rect 76532 24330 76580 24332
rect 76448 24278 76476 24330
rect 76572 24278 76580 24330
rect 76428 24276 76476 24278
rect 76532 24276 76580 24278
rect 76636 24330 76684 24332
rect 76740 24330 76788 24332
rect 76636 24278 76644 24330
rect 76740 24278 76768 24330
rect 76636 24276 76684 24278
rect 76740 24276 76788 24278
rect 76844 24276 76892 24332
rect 76268 24266 76948 24276
rect 76300 23940 76356 23950
rect 76300 23846 76356 23884
rect 76636 23714 76692 23726
rect 76636 23662 76638 23714
rect 76690 23662 76692 23714
rect 76636 23380 76692 23662
rect 76636 23314 76692 23324
rect 77420 23492 77476 25228
rect 77756 24946 77812 26236
rect 77980 26180 78036 26190
rect 77980 26086 78036 26124
rect 78876 26180 78932 27918
rect 79660 27636 79716 27646
rect 79660 27542 79716 27580
rect 84028 27636 84084 27646
rect 80768 26684 81448 26694
rect 80824 26628 80872 26684
rect 80928 26682 80976 26684
rect 81032 26682 81080 26684
rect 80948 26630 80976 26682
rect 81072 26630 81080 26682
rect 80928 26628 80976 26630
rect 81032 26628 81080 26630
rect 81136 26682 81184 26684
rect 81240 26682 81288 26684
rect 81136 26630 81144 26682
rect 81240 26630 81268 26682
rect 81136 26628 81184 26630
rect 81240 26628 81288 26630
rect 81344 26628 81392 26684
rect 80768 26618 81448 26628
rect 84028 26290 84084 27580
rect 85268 27468 85948 27478
rect 85324 27412 85372 27468
rect 85428 27466 85476 27468
rect 85532 27466 85580 27468
rect 85448 27414 85476 27466
rect 85572 27414 85580 27466
rect 85428 27412 85476 27414
rect 85532 27412 85580 27414
rect 85636 27466 85684 27468
rect 85740 27466 85788 27468
rect 85636 27414 85644 27466
rect 85740 27414 85768 27466
rect 85636 27412 85684 27414
rect 85740 27412 85788 27414
rect 85844 27412 85892 27468
rect 85268 27402 85948 27412
rect 94268 27468 94948 27478
rect 94324 27412 94372 27468
rect 94428 27466 94476 27468
rect 94532 27466 94580 27468
rect 94448 27414 94476 27466
rect 94572 27414 94580 27466
rect 94428 27412 94476 27414
rect 94532 27412 94580 27414
rect 94636 27466 94684 27468
rect 94740 27466 94788 27468
rect 94636 27414 94644 27466
rect 94740 27414 94768 27466
rect 94636 27412 94684 27414
rect 94740 27412 94788 27414
rect 94844 27412 94892 27468
rect 94268 27402 94948 27412
rect 96572 27300 96628 27310
rect 96572 27188 96628 27244
rect 96572 27186 96964 27188
rect 96572 27134 96574 27186
rect 96626 27134 96964 27186
rect 96572 27132 96964 27134
rect 96572 27122 96628 27132
rect 96908 27074 96964 27132
rect 96908 27022 96910 27074
rect 96962 27022 96964 27074
rect 96908 27010 96964 27022
rect 97692 26962 97748 26974
rect 97692 26910 97694 26962
rect 97746 26910 97748 26962
rect 89768 26684 90448 26694
rect 89824 26628 89872 26684
rect 89928 26682 89976 26684
rect 90032 26682 90080 26684
rect 89948 26630 89976 26682
rect 90072 26630 90080 26682
rect 89928 26628 89976 26630
rect 90032 26628 90080 26630
rect 90136 26682 90184 26684
rect 90240 26682 90288 26684
rect 90136 26630 90144 26682
rect 90240 26630 90268 26682
rect 90136 26628 90184 26630
rect 90240 26628 90288 26630
rect 90344 26628 90392 26684
rect 89768 26618 90448 26628
rect 84252 26404 84308 26414
rect 84252 26310 84308 26348
rect 96908 26404 96964 26414
rect 84028 26238 84030 26290
rect 84082 26238 84084 26290
rect 84028 26226 84084 26238
rect 78876 25620 78932 26124
rect 85268 25900 85948 25910
rect 85324 25844 85372 25900
rect 85428 25898 85476 25900
rect 85532 25898 85580 25900
rect 85448 25846 85476 25898
rect 85572 25846 85580 25898
rect 85428 25844 85476 25846
rect 85532 25844 85580 25846
rect 85636 25898 85684 25900
rect 85740 25898 85788 25900
rect 85636 25846 85644 25898
rect 85740 25846 85768 25898
rect 85636 25844 85684 25846
rect 85740 25844 85788 25846
rect 85844 25844 85892 25900
rect 85268 25834 85948 25844
rect 94268 25900 94948 25910
rect 94324 25844 94372 25900
rect 94428 25898 94476 25900
rect 94532 25898 94580 25900
rect 94448 25846 94476 25898
rect 94572 25846 94580 25898
rect 94428 25844 94476 25846
rect 94532 25844 94580 25846
rect 94636 25898 94684 25900
rect 94740 25898 94788 25900
rect 94636 25846 94644 25898
rect 94740 25846 94768 25898
rect 94636 25844 94684 25846
rect 94740 25844 94788 25846
rect 94844 25844 94892 25900
rect 94268 25834 94948 25844
rect 78876 25554 78932 25564
rect 77756 24894 77758 24946
rect 77810 24894 77812 24946
rect 77756 24724 77812 24894
rect 77868 25506 77924 25518
rect 77868 25454 77870 25506
rect 77922 25454 77924 25506
rect 77868 24946 77924 25454
rect 78428 25508 78484 25518
rect 78764 25508 78820 25518
rect 78428 25506 78596 25508
rect 78428 25454 78430 25506
rect 78482 25454 78596 25506
rect 78428 25452 78596 25454
rect 78428 25442 78484 25452
rect 77868 24894 77870 24946
rect 77922 24894 77924 24946
rect 77868 24882 77924 24894
rect 78092 24948 78148 24958
rect 78092 24854 78148 24892
rect 78540 24946 78596 25452
rect 78764 25414 78820 25452
rect 81116 25396 81172 25406
rect 81116 25302 81172 25340
rect 81900 25282 81956 25294
rect 81900 25230 81902 25282
rect 81954 25230 81956 25282
rect 80768 25116 81448 25126
rect 80824 25060 80872 25116
rect 80928 25114 80976 25116
rect 81032 25114 81080 25116
rect 80948 25062 80976 25114
rect 81072 25062 81080 25114
rect 80928 25060 80976 25062
rect 81032 25060 81080 25062
rect 81136 25114 81184 25116
rect 81240 25114 81288 25116
rect 81136 25062 81144 25114
rect 81240 25062 81268 25114
rect 81136 25060 81184 25062
rect 81240 25060 81288 25062
rect 81344 25060 81392 25116
rect 80768 25050 81448 25060
rect 78540 24894 78542 24946
rect 78594 24894 78596 24946
rect 78540 24882 78596 24894
rect 81900 24948 81956 25230
rect 89768 25116 90448 25126
rect 89824 25060 89872 25116
rect 89928 25114 89976 25116
rect 90032 25114 90080 25116
rect 89948 25062 89976 25114
rect 90072 25062 90080 25114
rect 89928 25060 89976 25062
rect 90032 25060 90080 25062
rect 90136 25114 90184 25116
rect 90240 25114 90288 25116
rect 90136 25062 90144 25114
rect 90240 25062 90268 25114
rect 90136 25060 90184 25062
rect 90240 25060 90288 25062
rect 90344 25060 90392 25116
rect 89768 25050 90448 25060
rect 81900 24882 81956 24892
rect 83132 24948 83188 24958
rect 83132 24834 83188 24892
rect 83132 24782 83134 24834
rect 83186 24782 83188 24834
rect 83132 24770 83188 24782
rect 83468 24834 83524 24846
rect 83468 24782 83470 24834
rect 83522 24782 83524 24834
rect 78204 24724 78260 24734
rect 77756 24722 78260 24724
rect 77756 24670 78206 24722
rect 78258 24670 78260 24722
rect 77756 24668 78260 24670
rect 78204 24658 78260 24668
rect 80768 23548 81448 23558
rect 80824 23492 80872 23548
rect 80928 23546 80976 23548
rect 81032 23546 81080 23548
rect 80948 23494 80976 23546
rect 81072 23494 81080 23546
rect 80928 23492 80976 23494
rect 81032 23492 81080 23494
rect 81136 23546 81184 23548
rect 81240 23546 81288 23548
rect 81136 23494 81144 23546
rect 81240 23494 81268 23546
rect 81136 23492 81184 23494
rect 81240 23492 81288 23494
rect 81344 23492 81392 23548
rect 77420 23436 78036 23492
rect 80768 23482 81448 23492
rect 77420 23378 77476 23436
rect 77420 23326 77422 23378
rect 77474 23326 77476 23378
rect 77420 23314 77476 23326
rect 77980 23378 78036 23436
rect 81004 23380 81060 23390
rect 82236 23380 82292 23390
rect 77980 23326 77982 23378
rect 78034 23326 78036 23378
rect 77980 23314 78036 23326
rect 80668 23378 82292 23380
rect 80668 23326 81006 23378
rect 81058 23326 82238 23378
rect 82290 23326 82292 23378
rect 80668 23324 82292 23326
rect 77756 23268 77812 23278
rect 77756 23174 77812 23212
rect 78652 23266 78708 23278
rect 78652 23214 78654 23266
rect 78706 23214 78708 23266
rect 78428 23156 78484 23166
rect 78428 23062 78484 23100
rect 77868 23042 77924 23054
rect 77868 22990 77870 23042
rect 77922 22990 77924 23042
rect 76268 22764 76948 22774
rect 76324 22708 76372 22764
rect 76428 22762 76476 22764
rect 76532 22762 76580 22764
rect 76448 22710 76476 22762
rect 76572 22710 76580 22762
rect 76428 22708 76476 22710
rect 76532 22708 76580 22710
rect 76636 22762 76684 22764
rect 76740 22762 76788 22764
rect 76636 22710 76644 22762
rect 76740 22710 76768 22762
rect 76636 22708 76684 22710
rect 76740 22708 76788 22710
rect 76844 22708 76892 22764
rect 76268 22698 76948 22708
rect 77868 22708 77924 22990
rect 77868 22652 78596 22708
rect 75964 22540 76356 22596
rect 75404 22036 75460 22316
rect 75628 22484 75684 22494
rect 75460 21980 75572 22036
rect 75404 21970 75460 21980
rect 73724 20916 73780 20926
rect 73724 20822 73780 20860
rect 74172 20916 74228 20926
rect 74172 20802 74228 20860
rect 74172 20750 74174 20802
rect 74226 20750 74228 20802
rect 74172 20738 74228 20750
rect 74956 20580 75012 21532
rect 75292 21494 75348 21532
rect 73500 20078 73502 20130
rect 73554 20078 73556 20130
rect 73052 19908 73108 19918
rect 73500 19908 73556 20078
rect 73052 19906 73556 19908
rect 73052 19854 73054 19906
rect 73106 19854 73556 19906
rect 73052 19852 73556 19854
rect 74396 20132 74452 20142
rect 73052 19842 73108 19852
rect 74396 19460 74452 20076
rect 74956 19908 75012 20524
rect 75516 20244 75572 21980
rect 75068 20242 75572 20244
rect 75068 20190 75518 20242
rect 75570 20190 75572 20242
rect 75068 20188 75572 20190
rect 75068 20130 75124 20188
rect 75516 20178 75572 20188
rect 75068 20078 75070 20130
rect 75122 20078 75124 20130
rect 75068 20066 75124 20078
rect 74956 19842 75012 19852
rect 74396 19366 74452 19404
rect 74508 19794 74564 19806
rect 74508 19742 74510 19794
rect 74562 19742 74564 19794
rect 71484 19058 71540 19068
rect 73836 19348 73892 19358
rect 74508 19348 74564 19742
rect 75180 19460 75236 19470
rect 74732 19348 74788 19358
rect 74508 19292 74732 19348
rect 73836 19010 73892 19292
rect 74732 19254 74788 19292
rect 73836 18958 73838 19010
rect 73890 18958 73892 19010
rect 73836 18946 73892 18958
rect 71768 18844 72448 18854
rect 71824 18788 71872 18844
rect 71928 18842 71976 18844
rect 72032 18842 72080 18844
rect 71948 18790 71976 18842
rect 72072 18790 72080 18842
rect 71928 18788 71976 18790
rect 72032 18788 72080 18790
rect 72136 18842 72184 18844
rect 72240 18842 72288 18844
rect 72136 18790 72144 18842
rect 72240 18790 72268 18842
rect 72136 18788 72184 18790
rect 72240 18788 72288 18790
rect 72344 18788 72392 18844
rect 71768 18778 72448 18788
rect 75180 18562 75236 19404
rect 75628 19348 75684 22428
rect 76300 22484 76356 22540
rect 76300 22390 76356 22428
rect 77756 22484 77812 22494
rect 75740 22146 75796 22158
rect 75740 22094 75742 22146
rect 75794 22094 75796 22146
rect 75740 21700 75796 22094
rect 77756 22148 77812 22428
rect 78204 22370 78260 22382
rect 78204 22318 78206 22370
rect 78258 22318 78260 22370
rect 78204 22148 78260 22318
rect 78540 22370 78596 22652
rect 78540 22318 78542 22370
rect 78594 22318 78596 22370
rect 78540 22306 78596 22318
rect 78652 22148 78708 23214
rect 78204 22092 78708 22148
rect 80220 23156 80276 23166
rect 77756 22082 77812 22092
rect 80220 21810 80276 23100
rect 80668 22148 80724 23324
rect 81004 23314 81060 23324
rect 82236 23314 82292 23324
rect 82572 23268 82628 23278
rect 82012 23154 82068 23166
rect 82012 23102 82014 23154
rect 82066 23102 82068 23154
rect 81452 23044 81508 23054
rect 82012 23044 82068 23102
rect 82124 23156 82180 23166
rect 82124 23062 82180 23100
rect 81452 23042 82068 23044
rect 81452 22990 81454 23042
rect 81506 22990 82068 23042
rect 81452 22988 82068 22990
rect 81452 22596 81508 22988
rect 81452 22530 81508 22540
rect 82572 22372 82628 23212
rect 82572 22278 82628 22316
rect 82684 23154 82740 23166
rect 82684 23102 82686 23154
rect 82738 23102 82740 23154
rect 82684 22260 82740 23102
rect 83020 23154 83076 23166
rect 83020 23102 83022 23154
rect 83074 23102 83076 23154
rect 83020 22260 83076 23102
rect 83356 23156 83412 23166
rect 83356 23062 83412 23100
rect 83132 22260 83188 22270
rect 83020 22258 83188 22260
rect 83020 22206 83134 22258
rect 83186 22206 83188 22258
rect 83020 22204 83188 22206
rect 82684 22194 82740 22204
rect 83132 22194 83188 22204
rect 80220 21758 80222 21810
rect 80274 21758 80276 21810
rect 80220 21746 80276 21758
rect 80556 22092 80724 22148
rect 80892 22148 80948 22186
rect 80556 21812 80612 22092
rect 80892 22082 80948 22092
rect 81676 22146 81732 22158
rect 81676 22094 81678 22146
rect 81730 22094 81732 22146
rect 80768 21980 81448 21990
rect 80824 21924 80872 21980
rect 80928 21978 80976 21980
rect 81032 21978 81080 21980
rect 80948 21926 80976 21978
rect 81072 21926 81080 21978
rect 80928 21924 80976 21926
rect 81032 21924 81080 21926
rect 81136 21978 81184 21980
rect 81240 21978 81288 21980
rect 81136 21926 81144 21978
rect 81240 21926 81268 21978
rect 81136 21924 81184 21926
rect 81240 21924 81288 21926
rect 81344 21924 81392 21980
rect 80768 21914 81448 21924
rect 80556 21756 80724 21812
rect 75740 21634 75796 21644
rect 77756 21700 77812 21710
rect 75852 21588 75908 21598
rect 75740 21476 75796 21486
rect 75852 21476 75908 21532
rect 75740 21474 75908 21476
rect 75740 21422 75742 21474
rect 75794 21422 75908 21474
rect 75740 21420 75908 21422
rect 75740 21410 75796 21420
rect 76268 21196 76948 21206
rect 76324 21140 76372 21196
rect 76428 21194 76476 21196
rect 76532 21194 76580 21196
rect 76448 21142 76476 21194
rect 76572 21142 76580 21194
rect 76428 21140 76476 21142
rect 76532 21140 76580 21142
rect 76636 21194 76684 21196
rect 76740 21194 76788 21196
rect 76636 21142 76644 21194
rect 76740 21142 76768 21194
rect 76636 21140 76684 21142
rect 76740 21140 76788 21142
rect 76844 21140 76892 21196
rect 76268 21130 76948 21140
rect 76300 20578 76356 20590
rect 76300 20526 76302 20578
rect 76354 20526 76356 20578
rect 76300 20244 76356 20526
rect 76300 20178 76356 20188
rect 77756 20188 77812 21644
rect 80444 21698 80500 21710
rect 80444 21646 80446 21698
rect 80498 21646 80500 21698
rect 78764 21588 78820 21598
rect 75628 19254 75684 19292
rect 75964 20130 76020 20142
rect 77756 20132 77924 20188
rect 75964 20078 75966 20130
rect 76018 20078 76020 20130
rect 75964 19236 76020 20078
rect 76524 20018 76580 20030
rect 76524 19966 76526 20018
rect 76578 19966 76580 20018
rect 76412 19908 76468 19918
rect 76076 19906 76468 19908
rect 76076 19854 76414 19906
rect 76466 19854 76468 19906
rect 76076 19852 76468 19854
rect 76076 19460 76132 19852
rect 76412 19842 76468 19852
rect 76524 19908 76580 19966
rect 76972 20020 77028 20030
rect 76972 19926 77028 19964
rect 76524 19842 76580 19852
rect 77420 19908 77476 19918
rect 77420 19814 77476 19852
rect 76268 19628 76948 19638
rect 76324 19572 76372 19628
rect 76428 19626 76476 19628
rect 76532 19626 76580 19628
rect 76448 19574 76476 19626
rect 76572 19574 76580 19626
rect 76428 19572 76476 19574
rect 76532 19572 76580 19574
rect 76636 19626 76684 19628
rect 76740 19626 76788 19628
rect 76636 19574 76644 19626
rect 76740 19574 76768 19626
rect 76636 19572 76684 19574
rect 76740 19572 76788 19574
rect 76844 19572 76892 19628
rect 76268 19562 76948 19572
rect 76076 19404 76692 19460
rect 76076 19236 76132 19246
rect 75964 19234 76132 19236
rect 75964 19182 76078 19234
rect 76130 19182 76132 19234
rect 75964 19180 76132 19182
rect 76076 19170 76132 19180
rect 76636 19234 76692 19404
rect 76636 19182 76638 19234
rect 76690 19182 76692 19234
rect 76636 19170 76692 19182
rect 75180 18510 75182 18562
rect 75234 18510 75236 18562
rect 75180 18498 75236 18510
rect 75516 18562 75572 18574
rect 75516 18510 75518 18562
rect 75570 18510 75572 18562
rect 71768 17276 72448 17286
rect 71824 17220 71872 17276
rect 71928 17274 71976 17276
rect 72032 17274 72080 17276
rect 71948 17222 71976 17274
rect 72072 17222 72080 17274
rect 71928 17220 71976 17222
rect 72032 17220 72080 17222
rect 72136 17274 72184 17276
rect 72240 17274 72288 17276
rect 72136 17222 72144 17274
rect 72240 17222 72268 17274
rect 72136 17220 72184 17222
rect 72240 17220 72288 17222
rect 72344 17220 72392 17276
rect 71768 17210 72448 17220
rect 71768 15708 72448 15718
rect 71824 15652 71872 15708
rect 71928 15706 71976 15708
rect 72032 15706 72080 15708
rect 71948 15654 71976 15706
rect 72072 15654 72080 15706
rect 71928 15652 71976 15654
rect 72032 15652 72080 15654
rect 72136 15706 72184 15708
rect 72240 15706 72288 15708
rect 72136 15654 72144 15706
rect 72240 15654 72268 15706
rect 72136 15652 72184 15654
rect 72240 15652 72288 15654
rect 72344 15652 72392 15708
rect 71768 15642 72448 15652
rect 71708 14532 71764 14542
rect 71148 14530 71764 14532
rect 71148 14478 71710 14530
rect 71762 14478 71764 14530
rect 71148 14476 71764 14478
rect 70812 13860 70868 13870
rect 70700 13804 70812 13860
rect 70812 13794 70868 13804
rect 71148 11506 71204 14476
rect 71708 14466 71764 14476
rect 74172 14530 74228 14542
rect 74172 14478 74174 14530
rect 74226 14478 74228 14530
rect 74172 14418 74228 14478
rect 74172 14366 74174 14418
rect 74226 14366 74228 14418
rect 73948 14308 74004 14318
rect 73724 14306 74004 14308
rect 73724 14254 73950 14306
rect 74002 14254 74004 14306
rect 73724 14252 74004 14254
rect 74172 14308 74228 14366
rect 74620 14308 74676 14318
rect 75068 14308 75124 14318
rect 74172 14306 75124 14308
rect 74172 14254 74622 14306
rect 74674 14254 75070 14306
rect 75122 14254 75124 14306
rect 74172 14252 75124 14254
rect 71768 14140 72448 14150
rect 71824 14084 71872 14140
rect 71928 14138 71976 14140
rect 72032 14138 72080 14140
rect 71948 14086 71976 14138
rect 72072 14086 72080 14138
rect 71928 14084 71976 14086
rect 72032 14084 72080 14086
rect 72136 14138 72184 14140
rect 72240 14138 72288 14140
rect 72136 14086 72144 14138
rect 72240 14086 72268 14138
rect 72136 14084 72184 14086
rect 72240 14084 72288 14086
rect 72344 14084 72392 14140
rect 71768 14074 72448 14084
rect 72268 13860 72324 13870
rect 72268 13766 72324 13804
rect 72604 13860 72660 13870
rect 72604 13858 72884 13860
rect 72604 13806 72606 13858
rect 72658 13806 72884 13858
rect 72604 13804 72884 13806
rect 72604 13794 72660 13804
rect 71768 12572 72448 12582
rect 71824 12516 71872 12572
rect 71928 12570 71976 12572
rect 72032 12570 72080 12572
rect 71948 12518 71976 12570
rect 72072 12518 72080 12570
rect 71928 12516 71976 12518
rect 72032 12516 72080 12518
rect 72136 12570 72184 12572
rect 72240 12570 72288 12572
rect 72136 12518 72144 12570
rect 72240 12518 72268 12570
rect 72136 12516 72184 12518
rect 72240 12516 72288 12518
rect 72344 12516 72392 12572
rect 71768 12506 72448 12516
rect 71708 12292 71764 12302
rect 71484 12290 71764 12292
rect 71484 12238 71710 12290
rect 71762 12238 71764 12290
rect 71484 12236 71764 12238
rect 71484 12178 71540 12236
rect 71708 12226 71764 12236
rect 72828 12292 72884 13804
rect 72828 12226 72884 12236
rect 71484 12126 71486 12178
rect 71538 12126 71540 12178
rect 71372 12068 71428 12078
rect 71148 11454 71150 11506
rect 71202 11454 71204 11506
rect 71148 11442 71204 11454
rect 71260 12012 71372 12068
rect 70140 6636 70644 6692
rect 70700 9714 70756 9726
rect 70700 9662 70702 9714
rect 70754 9662 70756 9714
rect 70028 5012 70084 5022
rect 70028 4338 70084 4956
rect 70140 4562 70196 6636
rect 70700 6580 70756 9662
rect 70924 8932 70980 8942
rect 70252 6524 70756 6580
rect 70812 7924 70868 7934
rect 70252 6018 70308 6524
rect 70812 6468 70868 7868
rect 70252 5966 70254 6018
rect 70306 5966 70308 6018
rect 70252 5954 70308 5966
rect 70700 6412 70868 6468
rect 70140 4510 70142 4562
rect 70194 4510 70196 4562
rect 70140 4498 70196 4510
rect 70364 5682 70420 5694
rect 70364 5630 70366 5682
rect 70418 5630 70420 5682
rect 70028 4286 70030 4338
rect 70082 4286 70084 4338
rect 70028 4116 70084 4286
rect 70028 4050 70084 4060
rect 70364 3668 70420 5630
rect 70700 5234 70756 6412
rect 70812 6244 70868 6254
rect 70812 6020 70868 6188
rect 70924 6132 70980 8876
rect 71036 8148 71092 8158
rect 71036 7474 71092 8092
rect 71036 7422 71038 7474
rect 71090 7422 71092 7474
rect 71036 7410 71092 7422
rect 71148 7250 71204 7262
rect 71148 7198 71150 7250
rect 71202 7198 71204 7250
rect 71148 6692 71204 7198
rect 71148 6626 71204 6636
rect 70924 6076 71204 6132
rect 70812 6018 71092 6020
rect 70812 5966 70814 6018
rect 70866 5966 71092 6018
rect 70812 5964 71092 5966
rect 70812 5954 70868 5964
rect 71036 5906 71092 5964
rect 71036 5854 71038 5906
rect 71090 5854 71092 5906
rect 71036 5842 71092 5854
rect 70812 5796 70868 5806
rect 70812 5702 70868 5740
rect 70700 5182 70702 5234
rect 70754 5182 70756 5234
rect 70700 5170 70756 5182
rect 70924 5684 70980 5694
rect 70700 4900 70756 4910
rect 70700 4340 70756 4844
rect 70924 4562 70980 5628
rect 70924 4510 70926 4562
rect 70978 4510 70980 4562
rect 70924 4498 70980 4510
rect 71036 4340 71092 4350
rect 70700 4338 71092 4340
rect 70700 4286 70702 4338
rect 70754 4286 71038 4338
rect 71090 4286 71092 4338
rect 70700 4284 71092 4286
rect 70700 4274 70756 4284
rect 71036 4274 71092 4284
rect 70364 3602 70420 3612
rect 71036 3668 71092 3678
rect 71036 3574 71092 3612
rect 71148 3556 71204 6076
rect 71260 6130 71316 12012
rect 71372 12002 71428 12012
rect 71484 9380 71540 12126
rect 72492 12068 72548 12078
rect 72492 11974 72548 12012
rect 73612 11394 73668 11406
rect 73612 11342 73614 11394
rect 73666 11342 73668 11394
rect 71768 11004 72448 11014
rect 71824 10948 71872 11004
rect 71928 11002 71976 11004
rect 72032 11002 72080 11004
rect 71948 10950 71976 11002
rect 72072 10950 72080 11002
rect 71928 10948 71976 10950
rect 72032 10948 72080 10950
rect 72136 11002 72184 11004
rect 72240 11002 72288 11004
rect 72136 10950 72144 11002
rect 72240 10950 72268 11002
rect 72136 10948 72184 10950
rect 72240 10948 72288 10950
rect 72344 10948 72392 11004
rect 71768 10938 72448 10948
rect 72604 10610 72660 10622
rect 72604 10558 72606 10610
rect 72658 10558 72660 10610
rect 71768 9436 72448 9446
rect 71824 9380 71872 9436
rect 71928 9434 71976 9436
rect 72032 9434 72080 9436
rect 71948 9382 71976 9434
rect 72072 9382 72080 9434
rect 71928 9380 71976 9382
rect 72032 9380 72080 9382
rect 72136 9434 72184 9436
rect 72240 9434 72288 9436
rect 72136 9382 72144 9434
rect 72240 9382 72268 9434
rect 72136 9380 72184 9382
rect 72240 9380 72288 9382
rect 72344 9380 72392 9436
rect 71484 9324 71652 9380
rect 71768 9370 72448 9380
rect 71372 8146 71428 8158
rect 71372 8094 71374 8146
rect 71426 8094 71428 8146
rect 71372 7474 71428 8094
rect 71372 7422 71374 7474
rect 71426 7422 71428 7474
rect 71372 7410 71428 7422
rect 71260 6078 71262 6130
rect 71314 6078 71316 6130
rect 71260 6066 71316 6078
rect 71484 7250 71540 7262
rect 71484 7198 71486 7250
rect 71538 7198 71540 7250
rect 71372 5348 71428 5358
rect 71372 4450 71428 5292
rect 71372 4398 71374 4450
rect 71426 4398 71428 4450
rect 71372 4386 71428 4398
rect 71484 3892 71540 7198
rect 71596 6468 71652 9324
rect 72492 8932 72548 8942
rect 72492 8838 72548 8876
rect 71768 7868 72448 7878
rect 71824 7812 71872 7868
rect 71928 7866 71976 7868
rect 72032 7866 72080 7868
rect 71948 7814 71976 7866
rect 72072 7814 72080 7866
rect 71928 7812 71976 7814
rect 72032 7812 72080 7814
rect 72136 7866 72184 7868
rect 72240 7866 72288 7868
rect 72136 7814 72144 7866
rect 72240 7814 72268 7866
rect 72136 7812 72184 7814
rect 72240 7812 72288 7814
rect 72344 7812 72392 7868
rect 71768 7802 72448 7812
rect 71596 6402 71652 6412
rect 71768 6300 72448 6310
rect 71824 6244 71872 6300
rect 71928 6298 71976 6300
rect 72032 6298 72080 6300
rect 71948 6246 71976 6298
rect 72072 6246 72080 6298
rect 71928 6244 71976 6246
rect 72032 6244 72080 6246
rect 72136 6298 72184 6300
rect 72240 6298 72288 6300
rect 72136 6246 72144 6298
rect 72240 6246 72268 6298
rect 72136 6244 72184 6246
rect 72240 6244 72288 6246
rect 72344 6244 72392 6300
rect 71768 6234 72448 6244
rect 71708 6132 71764 6142
rect 71708 5906 71764 6076
rect 72492 6020 72548 6030
rect 72492 5926 72548 5964
rect 71708 5854 71710 5906
rect 71762 5854 71764 5906
rect 71708 5842 71764 5854
rect 71596 5682 71652 5694
rect 71596 5630 71598 5682
rect 71650 5630 71652 5682
rect 71596 4564 71652 5630
rect 72604 5684 72660 10558
rect 73612 9044 73668 11342
rect 73612 8978 73668 8988
rect 72828 8036 72884 8046
rect 72604 5618 72660 5628
rect 72716 6690 72772 6702
rect 72716 6638 72718 6690
rect 72770 6638 72772 6690
rect 71768 4732 72448 4742
rect 71824 4676 71872 4732
rect 71928 4730 71976 4732
rect 72032 4730 72080 4732
rect 71948 4678 71976 4730
rect 72072 4678 72080 4730
rect 71928 4676 71976 4678
rect 72032 4676 72080 4678
rect 72136 4730 72184 4732
rect 72240 4730 72288 4732
rect 72136 4678 72144 4730
rect 72240 4678 72268 4730
rect 72136 4676 72184 4678
rect 72240 4676 72288 4678
rect 72344 4676 72392 4732
rect 71768 4666 72448 4676
rect 71596 4508 71988 4564
rect 71708 4228 71764 4238
rect 71708 4134 71764 4172
rect 71596 4116 71652 4126
rect 71596 4022 71652 4060
rect 71484 3836 71876 3892
rect 71260 3556 71316 3566
rect 71148 3554 71316 3556
rect 71148 3502 71262 3554
rect 71314 3502 71316 3554
rect 71148 3500 71316 3502
rect 71260 3490 71316 3500
rect 71596 3556 71652 3566
rect 69748 3388 69972 3444
rect 69692 3378 69748 3388
rect 53768 3164 54448 3174
rect 53824 3108 53872 3164
rect 53928 3162 53976 3164
rect 54032 3162 54080 3164
rect 53948 3110 53976 3162
rect 54072 3110 54080 3162
rect 53928 3108 53976 3110
rect 54032 3108 54080 3110
rect 54136 3162 54184 3164
rect 54240 3162 54288 3164
rect 54136 3110 54144 3162
rect 54240 3110 54268 3162
rect 54136 3108 54184 3110
rect 54240 3108 54288 3110
rect 54344 3108 54392 3164
rect 53768 3098 54448 3108
rect 49980 2156 50372 2212
rect 49980 800 50036 2156
rect 60956 800 61012 3332
rect 62768 3164 63448 3174
rect 62824 3108 62872 3164
rect 62928 3162 62976 3164
rect 63032 3162 63080 3164
rect 62948 3110 62976 3162
rect 63072 3110 63080 3162
rect 62928 3108 62976 3110
rect 63032 3108 63080 3110
rect 63136 3162 63184 3164
rect 63240 3162 63288 3164
rect 63136 3110 63144 3162
rect 63240 3110 63268 3162
rect 63136 3108 63184 3110
rect 63240 3108 63288 3110
rect 63344 3108 63392 3164
rect 62768 3098 63448 3108
rect 71596 2996 71652 3500
rect 71820 3442 71876 3836
rect 71820 3390 71822 3442
rect 71874 3390 71876 3442
rect 71820 3378 71876 3390
rect 71932 3444 71988 4508
rect 71932 3378 71988 3388
rect 72716 3330 72772 6638
rect 72828 4338 72884 7980
rect 73724 5124 73780 14252
rect 73948 14242 74004 14252
rect 74620 14242 74676 14252
rect 74060 13748 74116 13758
rect 74060 13654 74116 13692
rect 74844 13636 74900 14252
rect 75068 14242 75124 14252
rect 75516 13972 75572 18510
rect 76268 18060 76948 18070
rect 76324 18004 76372 18060
rect 76428 18058 76476 18060
rect 76532 18058 76580 18060
rect 76448 18006 76476 18058
rect 76572 18006 76580 18058
rect 76428 18004 76476 18006
rect 76532 18004 76580 18006
rect 76636 18058 76684 18060
rect 76740 18058 76788 18060
rect 76636 18006 76644 18058
rect 76740 18006 76768 18058
rect 76636 18004 76684 18006
rect 76740 18004 76788 18006
rect 76844 18004 76892 18060
rect 76268 17994 76948 18004
rect 76268 16492 76948 16502
rect 76324 16436 76372 16492
rect 76428 16490 76476 16492
rect 76532 16490 76580 16492
rect 76448 16438 76476 16490
rect 76572 16438 76580 16490
rect 76428 16436 76476 16438
rect 76532 16436 76580 16438
rect 76636 16490 76684 16492
rect 76740 16490 76788 16492
rect 76636 16438 76644 16490
rect 76740 16438 76768 16490
rect 76636 16436 76684 16438
rect 76740 16436 76788 16438
rect 76844 16436 76892 16492
rect 76268 16426 76948 16436
rect 76268 14924 76948 14934
rect 76324 14868 76372 14924
rect 76428 14922 76476 14924
rect 76532 14922 76580 14924
rect 76448 14870 76476 14922
rect 76572 14870 76580 14922
rect 76428 14868 76476 14870
rect 76532 14868 76580 14870
rect 76636 14922 76684 14924
rect 76740 14922 76788 14924
rect 76636 14870 76644 14922
rect 76740 14870 76768 14922
rect 76636 14868 76684 14870
rect 76740 14868 76788 14870
rect 76844 14868 76892 14924
rect 76268 14858 76948 14868
rect 77756 14084 77812 14094
rect 74844 13570 74900 13580
rect 74956 13916 75572 13972
rect 77644 14028 77756 14084
rect 73836 12962 73892 12974
rect 73836 12910 73838 12962
rect 73890 12910 73892 12962
rect 73836 12740 73892 12910
rect 73836 12674 73892 12684
rect 74284 12740 74340 12750
rect 74284 12646 74340 12684
rect 74060 7362 74116 7374
rect 74060 7310 74062 7362
rect 74114 7310 74116 7362
rect 73948 6692 74004 6702
rect 73948 6598 74004 6636
rect 74060 6690 74116 7310
rect 74620 6916 74676 6926
rect 74676 6860 74788 6916
rect 74620 6850 74676 6860
rect 74060 6638 74062 6690
rect 74114 6638 74116 6690
rect 74060 6626 74116 6638
rect 73948 6468 74004 6478
rect 73948 5234 74004 6412
rect 73948 5182 73950 5234
rect 74002 5182 74004 5234
rect 73948 5170 74004 5182
rect 74508 6468 74564 6478
rect 74508 5460 74564 6412
rect 74508 5236 74564 5404
rect 74732 5348 74788 6860
rect 74844 6466 74900 6478
rect 74844 6414 74846 6466
rect 74898 6414 74900 6466
rect 74844 6132 74900 6414
rect 74844 6066 74900 6076
rect 74844 5348 74900 5358
rect 74732 5346 74900 5348
rect 74732 5294 74846 5346
rect 74898 5294 74900 5346
rect 74732 5292 74900 5294
rect 74844 5282 74900 5292
rect 74508 5170 74564 5180
rect 73724 5058 73780 5068
rect 74396 5122 74452 5134
rect 74396 5070 74398 5122
rect 74450 5070 74452 5122
rect 72828 4286 72830 4338
rect 72882 4286 72884 4338
rect 72828 4274 72884 4286
rect 73276 4340 73332 4350
rect 73276 3444 73332 4284
rect 74396 4116 74452 5070
rect 74284 3668 74340 3678
rect 74284 3574 74340 3612
rect 73276 3378 73332 3388
rect 74396 3444 74452 4060
rect 74956 3780 75012 13916
rect 75516 13746 75572 13758
rect 75516 13694 75518 13746
rect 75570 13694 75572 13746
rect 75404 13636 75460 13646
rect 75516 13636 75572 13694
rect 76972 13748 77028 13758
rect 77308 13748 77364 13758
rect 76972 13746 77140 13748
rect 76972 13694 76974 13746
rect 77026 13694 77140 13746
rect 76972 13692 77140 13694
rect 76972 13682 77028 13692
rect 75404 13634 75516 13636
rect 75404 13582 75406 13634
rect 75458 13582 75516 13634
rect 75404 13580 75516 13582
rect 75404 13570 75460 13580
rect 75516 13570 75572 13580
rect 76268 13356 76948 13366
rect 76324 13300 76372 13356
rect 76428 13354 76476 13356
rect 76532 13354 76580 13356
rect 76448 13302 76476 13354
rect 76572 13302 76580 13354
rect 76428 13300 76476 13302
rect 76532 13300 76580 13302
rect 76636 13354 76684 13356
rect 76740 13354 76788 13356
rect 76636 13302 76644 13354
rect 76740 13302 76768 13354
rect 76636 13300 76684 13302
rect 76740 13300 76788 13302
rect 76844 13300 76892 13356
rect 76268 13290 76948 13300
rect 76076 12178 76132 12190
rect 76076 12126 76078 12178
rect 76130 12126 76132 12178
rect 75068 10724 75124 10734
rect 75068 9826 75124 10668
rect 76076 10724 76132 12126
rect 76268 11788 76948 11798
rect 76324 11732 76372 11788
rect 76428 11786 76476 11788
rect 76532 11786 76580 11788
rect 76448 11734 76476 11786
rect 76572 11734 76580 11786
rect 76428 11732 76476 11734
rect 76532 11732 76580 11734
rect 76636 11786 76684 11788
rect 76740 11786 76788 11788
rect 76636 11734 76644 11786
rect 76740 11734 76768 11786
rect 76636 11732 76684 11734
rect 76740 11732 76788 11734
rect 76844 11732 76892 11788
rect 76268 11722 76948 11732
rect 76076 10630 76132 10668
rect 76268 10220 76948 10230
rect 76324 10164 76372 10220
rect 76428 10218 76476 10220
rect 76532 10218 76580 10220
rect 76448 10166 76476 10218
rect 76572 10166 76580 10218
rect 76428 10164 76476 10166
rect 76532 10164 76580 10166
rect 76636 10218 76684 10220
rect 76740 10218 76788 10220
rect 76636 10166 76644 10218
rect 76740 10166 76768 10218
rect 76636 10164 76684 10166
rect 76740 10164 76788 10166
rect 76844 10164 76892 10220
rect 76268 10154 76948 10164
rect 75068 9774 75070 9826
rect 75122 9774 75124 9826
rect 75068 9762 75124 9774
rect 77084 9156 77140 13692
rect 77308 13654 77364 13692
rect 77308 9714 77364 9726
rect 77308 9662 77310 9714
rect 77362 9662 77364 9714
rect 77196 9156 77252 9166
rect 77084 9100 77196 9156
rect 77196 9090 77252 9100
rect 76076 9044 76132 9054
rect 76076 8950 76132 8988
rect 76268 8652 76948 8662
rect 76324 8596 76372 8652
rect 76428 8650 76476 8652
rect 76532 8650 76580 8652
rect 76448 8598 76476 8650
rect 76572 8598 76580 8650
rect 76428 8596 76476 8598
rect 76532 8596 76580 8598
rect 76636 8650 76684 8652
rect 76740 8650 76788 8652
rect 76636 8598 76644 8650
rect 76740 8598 76768 8650
rect 76636 8596 76684 8598
rect 76740 8596 76788 8598
rect 76844 8596 76892 8652
rect 76268 8586 76948 8596
rect 76412 8148 76468 8158
rect 76412 8054 76468 8092
rect 77196 7476 77252 7486
rect 77196 7382 77252 7420
rect 76268 7084 76948 7094
rect 76324 7028 76372 7084
rect 76428 7082 76476 7084
rect 76532 7082 76580 7084
rect 76448 7030 76476 7082
rect 76572 7030 76580 7082
rect 76428 7028 76476 7030
rect 76532 7028 76580 7030
rect 76636 7082 76684 7084
rect 76740 7082 76788 7084
rect 76636 7030 76644 7082
rect 76740 7030 76768 7082
rect 76636 7028 76684 7030
rect 76740 7028 76788 7030
rect 76844 7028 76892 7084
rect 76268 7018 76948 7028
rect 77084 6804 77140 6814
rect 76188 6690 76244 6702
rect 76188 6638 76190 6690
rect 76242 6638 76244 6690
rect 75516 6580 75572 6590
rect 75404 6468 75460 6478
rect 75404 6374 75460 6412
rect 75292 4898 75348 4910
rect 75292 4846 75294 4898
rect 75346 4846 75348 4898
rect 75292 4228 75348 4846
rect 75292 4162 75348 4172
rect 74956 3714 75012 3724
rect 75516 3666 75572 6524
rect 76188 6020 76244 6638
rect 76188 5954 76244 5964
rect 76076 5906 76132 5918
rect 76076 5854 76078 5906
rect 76130 5854 76132 5906
rect 75628 4452 75684 4462
rect 75628 4358 75684 4396
rect 75516 3614 75518 3666
rect 75570 3614 75572 3666
rect 75516 3602 75572 3614
rect 74396 3378 74452 3388
rect 75852 3444 75908 3454
rect 72716 3278 72718 3330
rect 72770 3278 72772 3330
rect 72716 3266 72772 3278
rect 75852 3330 75908 3388
rect 75852 3278 75854 3330
rect 75906 3278 75908 3330
rect 75852 3266 75908 3278
rect 76076 3332 76132 5854
rect 76268 5516 76948 5526
rect 76324 5460 76372 5516
rect 76428 5514 76476 5516
rect 76532 5514 76580 5516
rect 76448 5462 76476 5514
rect 76572 5462 76580 5514
rect 76428 5460 76476 5462
rect 76532 5460 76580 5462
rect 76636 5514 76684 5516
rect 76740 5514 76788 5516
rect 76636 5462 76644 5514
rect 76740 5462 76768 5514
rect 76636 5460 76684 5462
rect 76740 5460 76788 5462
rect 76844 5460 76892 5516
rect 76268 5450 76948 5460
rect 77084 5122 77140 6748
rect 77308 5908 77364 9662
rect 77084 5070 77086 5122
rect 77138 5070 77140 5122
rect 77084 5058 77140 5070
rect 77196 5852 77364 5908
rect 76268 3948 76948 3958
rect 76324 3892 76372 3948
rect 76428 3946 76476 3948
rect 76532 3946 76580 3948
rect 76448 3894 76476 3946
rect 76572 3894 76580 3946
rect 76428 3892 76476 3894
rect 76532 3892 76580 3894
rect 76636 3946 76684 3948
rect 76740 3946 76788 3948
rect 76636 3894 76644 3946
rect 76740 3894 76768 3946
rect 76636 3892 76684 3894
rect 76740 3892 76788 3894
rect 76844 3892 76892 3948
rect 76268 3882 76948 3892
rect 76748 3444 76804 3454
rect 77196 3444 77252 5852
rect 77308 5460 77364 5470
rect 77308 3554 77364 5404
rect 77644 4228 77700 14028
rect 77756 14018 77812 14028
rect 77644 4162 77700 4172
rect 77756 13860 77812 13870
rect 77756 3780 77812 13804
rect 77868 10722 77924 20132
rect 78092 20132 78148 20142
rect 78092 20038 78148 20076
rect 78204 20132 78260 20142
rect 78764 20132 78820 21532
rect 80444 21252 80500 21646
rect 80556 21588 80612 21598
rect 80556 21494 80612 21532
rect 80444 21186 80500 21196
rect 80668 20914 80724 21756
rect 81004 21588 81060 21598
rect 81004 21494 81060 21532
rect 81564 21588 81620 21598
rect 80668 20862 80670 20914
rect 80722 20862 80724 20914
rect 80668 20580 80724 20862
rect 80556 20524 80724 20580
rect 80108 20244 80164 20254
rect 80556 20244 80612 20524
rect 80768 20412 81448 20422
rect 80824 20356 80872 20412
rect 80928 20410 80976 20412
rect 81032 20410 81080 20412
rect 80948 20358 80976 20410
rect 81072 20358 81080 20410
rect 80928 20356 80976 20358
rect 81032 20356 81080 20358
rect 81136 20410 81184 20412
rect 81240 20410 81288 20412
rect 81136 20358 81144 20410
rect 81240 20358 81268 20410
rect 81136 20356 81184 20358
rect 81240 20356 81288 20358
rect 81344 20356 81392 20412
rect 80768 20346 81448 20356
rect 80556 20188 80724 20244
rect 81228 20242 81284 20254
rect 81228 20190 81230 20242
rect 81282 20190 81284 20242
rect 81228 20188 81284 20190
rect 78204 20130 78820 20132
rect 78204 20078 78206 20130
rect 78258 20078 78766 20130
rect 78818 20078 78820 20130
rect 78204 20076 78820 20078
rect 78204 20066 78260 20076
rect 78764 20038 78820 20076
rect 79772 20132 79828 20142
rect 77980 20020 78036 20030
rect 77980 19796 78036 19964
rect 78092 19796 78148 19806
rect 77980 19794 78148 19796
rect 77980 19742 78094 19794
rect 78146 19742 78148 19794
rect 77980 19740 78148 19742
rect 78092 19730 78148 19740
rect 79772 19460 79828 20076
rect 79772 19458 80052 19460
rect 79772 19406 79774 19458
rect 79826 19406 80052 19458
rect 79772 19404 80052 19406
rect 79772 19394 79828 19404
rect 79212 19348 79268 19358
rect 79212 19012 79268 19292
rect 79212 18918 79268 18956
rect 79660 19012 79716 19022
rect 79660 18674 79716 18956
rect 79660 18622 79662 18674
rect 79714 18622 79716 18674
rect 79660 18610 79716 18622
rect 79996 18564 80052 19404
rect 80108 19234 80164 20188
rect 80668 20132 81284 20188
rect 81564 20132 81620 21532
rect 81676 21252 81732 22094
rect 81676 21186 81732 21196
rect 82684 21252 82740 21262
rect 81900 20244 81956 20282
rect 81900 20178 81956 20188
rect 80444 19906 80500 19918
rect 80444 19854 80446 19906
rect 80498 19854 80500 19906
rect 80444 19796 80500 19854
rect 80668 19908 80724 20132
rect 81564 20066 81620 20076
rect 80668 19842 80724 19852
rect 81004 20018 81060 20030
rect 81004 19966 81006 20018
rect 81058 19966 81060 20018
rect 80444 19730 80500 19740
rect 81004 19796 81060 19966
rect 81676 20020 81732 20030
rect 81676 19926 81732 19964
rect 81004 19730 81060 19740
rect 81116 19906 81172 19918
rect 81116 19854 81118 19906
rect 81170 19854 81172 19906
rect 81116 19572 81172 19854
rect 80108 19182 80110 19234
rect 80162 19182 80164 19234
rect 80108 19170 80164 19182
rect 80556 19516 81172 19572
rect 80556 19234 80612 19516
rect 80556 19182 80558 19234
rect 80610 19182 80612 19234
rect 80556 19170 80612 19182
rect 80768 18844 81448 18854
rect 80824 18788 80872 18844
rect 80928 18842 80976 18844
rect 81032 18842 81080 18844
rect 80948 18790 80976 18842
rect 81072 18790 81080 18842
rect 80928 18788 80976 18790
rect 81032 18788 81080 18790
rect 81136 18842 81184 18844
rect 81240 18842 81288 18844
rect 81136 18790 81144 18842
rect 81240 18790 81268 18842
rect 81136 18788 81184 18790
rect 81240 18788 81288 18790
rect 81344 18788 81392 18844
rect 80768 18778 81448 18788
rect 80220 18564 80276 18574
rect 79996 18562 80276 18564
rect 79996 18510 80222 18562
rect 80274 18510 80276 18562
rect 79996 18508 80276 18510
rect 80220 18498 80276 18508
rect 80556 18562 80612 18574
rect 80556 18510 80558 18562
rect 80610 18510 80612 18562
rect 79660 15204 79716 15214
rect 80332 15204 80388 15214
rect 79660 15202 80388 15204
rect 79660 15150 79662 15202
rect 79714 15150 80334 15202
rect 80386 15150 80388 15202
rect 79660 15148 80388 15150
rect 78428 14530 78484 14542
rect 78428 14478 78430 14530
rect 78482 14478 78484 14530
rect 78316 14418 78372 14430
rect 78316 14366 78318 14418
rect 78370 14366 78372 14418
rect 77868 10670 77870 10722
rect 77922 10670 77924 10722
rect 77868 10658 77924 10670
rect 77980 13746 78036 13758
rect 77980 13694 77982 13746
rect 78034 13694 78036 13746
rect 77980 8428 78036 13694
rect 78316 11396 78372 14366
rect 78428 14084 78484 14478
rect 78428 14018 78484 14028
rect 78652 13748 78708 13758
rect 78316 11340 78484 11396
rect 78204 11172 78260 11182
rect 78204 11170 78372 11172
rect 78204 11118 78206 11170
rect 78258 11118 78372 11170
rect 78204 11116 78372 11118
rect 78204 11106 78260 11116
rect 78204 10724 78260 10734
rect 78204 10630 78260 10668
rect 77980 8372 78260 8428
rect 77980 7362 78036 7374
rect 77980 7310 77982 7362
rect 78034 7310 78036 7362
rect 77980 5460 78036 7310
rect 78204 6804 78260 8372
rect 78316 7474 78372 11116
rect 78316 7422 78318 7474
rect 78370 7422 78372 7474
rect 78316 7410 78372 7422
rect 78204 6748 78372 6804
rect 78204 6580 78260 6590
rect 78204 6486 78260 6524
rect 78092 6132 78148 6142
rect 78316 6132 78372 6748
rect 78092 6130 78372 6132
rect 78092 6078 78094 6130
rect 78146 6078 78372 6130
rect 78092 6076 78372 6078
rect 78092 6066 78148 6076
rect 77980 5394 78036 5404
rect 78428 4562 78484 11340
rect 78540 6132 78596 6142
rect 78540 6038 78596 6076
rect 78428 4510 78430 4562
rect 78482 4510 78484 4562
rect 78428 4498 78484 4510
rect 78316 4452 78372 4462
rect 78652 4452 78708 13692
rect 78876 13634 78932 13646
rect 78876 13582 78878 13634
rect 78930 13582 78932 13634
rect 78876 12628 78932 13582
rect 78876 12562 78932 12572
rect 79324 13636 79380 13646
rect 79660 13636 79716 15148
rect 80332 15138 80388 15148
rect 80556 14756 80612 18510
rect 80768 17276 81448 17286
rect 80824 17220 80872 17276
rect 80928 17274 80976 17276
rect 81032 17274 81080 17276
rect 80948 17222 80976 17274
rect 81072 17222 81080 17274
rect 80928 17220 80976 17222
rect 81032 17220 81080 17222
rect 81136 17274 81184 17276
rect 81240 17274 81288 17276
rect 81136 17222 81144 17274
rect 81240 17222 81268 17274
rect 81136 17220 81184 17222
rect 81240 17220 81288 17222
rect 81344 17220 81392 17276
rect 80768 17210 81448 17220
rect 80768 15708 81448 15718
rect 80824 15652 80872 15708
rect 80928 15706 80976 15708
rect 81032 15706 81080 15708
rect 80948 15654 80976 15706
rect 81072 15654 81080 15706
rect 80928 15652 80976 15654
rect 81032 15652 81080 15654
rect 81136 15706 81184 15708
rect 81240 15706 81288 15708
rect 81136 15654 81144 15706
rect 81240 15654 81268 15706
rect 81136 15652 81184 15654
rect 81240 15652 81288 15654
rect 81344 15652 81392 15708
rect 80768 15642 81448 15652
rect 80332 14700 80612 14756
rect 80220 13860 80276 13870
rect 80220 13766 80276 13804
rect 80108 13748 80164 13758
rect 80108 13654 80164 13692
rect 79380 13580 79716 13636
rect 78316 4358 78372 4396
rect 78540 4396 78708 4452
rect 78876 12068 78932 12078
rect 78876 6132 78932 12012
rect 79324 12066 79380 13580
rect 80108 12180 80164 12190
rect 80108 12086 80164 12124
rect 79324 12014 79326 12066
rect 79378 12014 79380 12066
rect 79100 9044 79156 9054
rect 78988 6132 79044 6142
rect 78876 6130 79044 6132
rect 78876 6078 78990 6130
rect 79042 6078 79044 6130
rect 78876 6076 79044 6078
rect 78876 4452 78932 6076
rect 78988 6066 79044 6076
rect 79100 5234 79156 8988
rect 79324 8428 79380 12014
rect 80332 8428 80388 14700
rect 80556 14532 80612 14542
rect 80556 14438 80612 14476
rect 81900 14530 81956 14542
rect 81900 14478 81902 14530
rect 81954 14478 81956 14530
rect 81676 14420 81732 14430
rect 81900 14420 81956 14478
rect 82684 14532 82740 21196
rect 83468 20188 83524 24782
rect 96908 24722 96964 26348
rect 97692 26292 97748 26910
rect 97692 26226 97748 26236
rect 96908 24670 96910 24722
rect 96962 24670 96964 24722
rect 96908 24658 96964 24670
rect 98028 24610 98084 24622
rect 98028 24558 98030 24610
rect 98082 24558 98084 24610
rect 98028 24500 98084 24558
rect 98028 24434 98084 24444
rect 85268 24332 85948 24342
rect 85324 24276 85372 24332
rect 85428 24330 85476 24332
rect 85532 24330 85580 24332
rect 85448 24278 85476 24330
rect 85572 24278 85580 24330
rect 85428 24276 85476 24278
rect 85532 24276 85580 24278
rect 85636 24330 85684 24332
rect 85740 24330 85788 24332
rect 85636 24278 85644 24330
rect 85740 24278 85768 24330
rect 85636 24276 85684 24278
rect 85740 24276 85788 24278
rect 85844 24276 85892 24332
rect 85268 24266 85948 24276
rect 94268 24332 94948 24342
rect 94324 24276 94372 24332
rect 94428 24330 94476 24332
rect 94532 24330 94580 24332
rect 94448 24278 94476 24330
rect 94572 24278 94580 24330
rect 94428 24276 94476 24278
rect 94532 24276 94580 24278
rect 94636 24330 94684 24332
rect 94740 24330 94788 24332
rect 94636 24278 94644 24330
rect 94740 24278 94768 24330
rect 94636 24276 94684 24278
rect 94740 24276 94788 24278
rect 94844 24276 94892 24332
rect 94268 24266 94948 24276
rect 89768 23548 90448 23558
rect 89824 23492 89872 23548
rect 89928 23546 89976 23548
rect 90032 23546 90080 23548
rect 89948 23494 89976 23546
rect 90072 23494 90080 23546
rect 89928 23492 89976 23494
rect 90032 23492 90080 23494
rect 90136 23546 90184 23548
rect 90240 23546 90288 23548
rect 90136 23494 90144 23546
rect 90240 23494 90268 23546
rect 90136 23492 90184 23494
rect 90240 23492 90288 23494
rect 90344 23492 90392 23548
rect 89768 23482 90448 23492
rect 96572 23380 96628 23390
rect 96628 23324 96964 23380
rect 96572 23286 96628 23324
rect 85036 23268 85092 23278
rect 84364 22428 84980 22484
rect 84364 22148 84420 22428
rect 84924 22370 84980 22428
rect 84924 22318 84926 22370
rect 84978 22318 84980 22370
rect 84924 22306 84980 22318
rect 84588 22260 84644 22270
rect 84588 22166 84644 22204
rect 84812 22260 84868 22270
rect 84812 22166 84868 22204
rect 84252 22146 84420 22148
rect 84252 22094 84366 22146
rect 84418 22094 84420 22146
rect 84252 22092 84420 22094
rect 82908 20132 82964 20142
rect 82908 20038 82964 20076
rect 83244 20130 83300 20142
rect 83244 20078 83246 20130
rect 83298 20078 83300 20130
rect 83020 20020 83076 20030
rect 83020 19926 83076 19964
rect 82796 19012 82852 19022
rect 83244 19012 83300 20078
rect 83356 20132 83412 20142
rect 83468 20132 83748 20188
rect 83356 20038 83412 20076
rect 83580 19012 83636 19022
rect 83244 19010 83636 19012
rect 83244 18958 83582 19010
rect 83634 18958 83636 19010
rect 83244 18956 83636 18958
rect 82796 18918 82852 18956
rect 83580 17668 83636 18956
rect 83580 17602 83636 17612
rect 83692 17444 83748 20132
rect 84252 20132 84308 22092
rect 84364 22082 84420 22092
rect 84364 21364 84420 21374
rect 84364 20916 84420 21308
rect 84364 20914 84980 20916
rect 84364 20862 84366 20914
rect 84418 20862 84980 20914
rect 84364 20860 84980 20862
rect 84364 20850 84420 20860
rect 84924 20802 84980 20860
rect 84924 20750 84926 20802
rect 84978 20750 84980 20802
rect 84924 20738 84980 20750
rect 85036 20804 85092 23212
rect 85708 23268 85764 23278
rect 85708 23174 85764 23212
rect 96908 23154 96964 23324
rect 96908 23102 96910 23154
rect 96962 23102 96964 23154
rect 96908 23090 96964 23102
rect 98028 23042 98084 23054
rect 98028 22990 98030 23042
rect 98082 22990 98084 23042
rect 86492 22930 86548 22942
rect 86492 22878 86494 22930
rect 86546 22878 86548 22930
rect 85268 22764 85948 22774
rect 85324 22708 85372 22764
rect 85428 22762 85476 22764
rect 85532 22762 85580 22764
rect 85448 22710 85476 22762
rect 85572 22710 85580 22762
rect 85428 22708 85476 22710
rect 85532 22708 85580 22710
rect 85636 22762 85684 22764
rect 85740 22762 85788 22764
rect 85636 22710 85644 22762
rect 85740 22710 85768 22762
rect 85636 22708 85684 22710
rect 85740 22708 85788 22710
rect 85844 22708 85892 22764
rect 85268 22698 85948 22708
rect 86492 22260 86548 22878
rect 94268 22764 94948 22774
rect 94324 22708 94372 22764
rect 94428 22762 94476 22764
rect 94532 22762 94580 22764
rect 94448 22710 94476 22762
rect 94572 22710 94580 22762
rect 94428 22708 94476 22710
rect 94532 22708 94580 22710
rect 94636 22762 94684 22764
rect 94740 22762 94788 22764
rect 94636 22710 94644 22762
rect 94740 22710 94768 22762
rect 94636 22708 94684 22710
rect 94740 22708 94788 22710
rect 94844 22708 94892 22764
rect 94268 22698 94948 22708
rect 98028 22708 98084 22990
rect 98028 22642 98084 22652
rect 86492 21700 86548 22204
rect 89768 21980 90448 21990
rect 89824 21924 89872 21980
rect 89928 21978 89976 21980
rect 90032 21978 90080 21980
rect 89948 21926 89976 21978
rect 90072 21926 90080 21978
rect 89928 21924 89976 21926
rect 90032 21924 90080 21926
rect 90136 21978 90184 21980
rect 90240 21978 90288 21980
rect 90136 21926 90144 21978
rect 90240 21926 90268 21978
rect 90136 21924 90184 21926
rect 90240 21924 90288 21926
rect 90344 21924 90392 21980
rect 89768 21914 90448 21924
rect 96572 21812 96628 21822
rect 96628 21756 96964 21812
rect 96572 21718 96628 21756
rect 87052 21700 87108 21710
rect 86492 21698 87108 21700
rect 86492 21646 87054 21698
rect 87106 21646 87108 21698
rect 86492 21644 87108 21646
rect 87052 21634 87108 21644
rect 87388 21698 87444 21710
rect 87388 21646 87390 21698
rect 87442 21646 87444 21698
rect 85268 21196 85948 21206
rect 85324 21140 85372 21196
rect 85428 21194 85476 21196
rect 85532 21194 85580 21196
rect 85448 21142 85476 21194
rect 85572 21142 85580 21194
rect 85428 21140 85476 21142
rect 85532 21140 85580 21142
rect 85636 21194 85684 21196
rect 85740 21194 85788 21196
rect 85636 21142 85644 21194
rect 85740 21142 85768 21194
rect 85636 21140 85684 21142
rect 85740 21140 85788 21142
rect 85844 21140 85892 21196
rect 85268 21130 85948 21140
rect 85596 20804 85652 20814
rect 85036 20748 85316 20804
rect 85036 20580 85092 20590
rect 85036 20486 85092 20524
rect 85148 20578 85204 20590
rect 85148 20526 85150 20578
rect 85202 20526 85204 20578
rect 85148 20244 85204 20526
rect 84252 20066 84308 20076
rect 85036 20188 85204 20244
rect 84700 19908 84756 19918
rect 84700 19814 84756 19852
rect 85036 19908 85092 20188
rect 85260 20132 85316 20748
rect 85596 20802 85876 20804
rect 85596 20750 85598 20802
rect 85650 20750 85876 20802
rect 85596 20748 85876 20750
rect 85596 20738 85652 20748
rect 85036 19842 85092 19852
rect 85148 20076 85316 20132
rect 85372 20132 85428 20142
rect 85148 19012 85204 20076
rect 85372 20020 85428 20076
rect 85596 20132 85652 20142
rect 85596 20038 85652 20076
rect 85820 20130 85876 20748
rect 86156 20580 86212 20590
rect 85820 20078 85822 20130
rect 85874 20078 85876 20130
rect 85820 20066 85876 20078
rect 86044 20242 86100 20254
rect 86044 20190 86046 20242
rect 86098 20190 86100 20242
rect 85484 20020 85540 20030
rect 85372 20018 85540 20020
rect 85372 19966 85486 20018
rect 85538 19966 85540 20018
rect 85372 19964 85540 19966
rect 85260 19908 85316 19918
rect 85372 19908 85428 19964
rect 85484 19954 85540 19964
rect 85260 19906 85428 19908
rect 85260 19854 85262 19906
rect 85314 19854 85428 19906
rect 85260 19852 85428 19854
rect 85260 19842 85316 19852
rect 85268 19628 85948 19638
rect 85324 19572 85372 19628
rect 85428 19626 85476 19628
rect 85532 19626 85580 19628
rect 85448 19574 85476 19626
rect 85572 19574 85580 19626
rect 85428 19572 85476 19574
rect 85532 19572 85580 19574
rect 85636 19626 85684 19628
rect 85740 19626 85788 19628
rect 85636 19574 85644 19626
rect 85740 19574 85768 19626
rect 85636 19572 85684 19574
rect 85740 19572 85788 19574
rect 85844 19572 85892 19628
rect 85268 19562 85948 19572
rect 86044 19460 86100 20190
rect 85596 19404 86100 19460
rect 85596 19234 85652 19404
rect 85596 19182 85598 19234
rect 85650 19182 85652 19234
rect 85596 19170 85652 19182
rect 86044 19236 86100 19246
rect 86156 19236 86212 20524
rect 86044 19234 86212 19236
rect 86044 19182 86046 19234
rect 86098 19182 86212 19234
rect 86044 19180 86212 19182
rect 86044 19170 86100 19180
rect 85148 18918 85204 18956
rect 85268 18060 85948 18070
rect 85324 18004 85372 18060
rect 85428 18058 85476 18060
rect 85532 18058 85580 18060
rect 85448 18006 85476 18058
rect 85572 18006 85580 18058
rect 85428 18004 85476 18006
rect 85532 18004 85580 18006
rect 85636 18058 85684 18060
rect 85740 18058 85788 18060
rect 85636 18006 85644 18058
rect 85740 18006 85768 18058
rect 85636 18004 85684 18006
rect 85740 18004 85788 18006
rect 85844 18004 85892 18060
rect 85268 17994 85948 18004
rect 85708 17668 85764 17678
rect 85708 17574 85764 17612
rect 83692 17378 83748 17388
rect 86044 17442 86100 17454
rect 86044 17390 86046 17442
rect 86098 17390 86100 17442
rect 85268 16492 85948 16502
rect 85324 16436 85372 16492
rect 85428 16490 85476 16492
rect 85532 16490 85580 16492
rect 85448 16438 85476 16490
rect 85572 16438 85580 16490
rect 85428 16436 85476 16438
rect 85532 16436 85580 16438
rect 85636 16490 85684 16492
rect 85740 16490 85788 16492
rect 85636 16438 85644 16490
rect 85740 16438 85768 16490
rect 85636 16436 85684 16438
rect 85740 16436 85788 16438
rect 85844 16436 85892 16492
rect 85268 16426 85948 16436
rect 82796 15204 82852 15214
rect 82796 15202 82964 15204
rect 82796 15150 82798 15202
rect 82850 15150 82964 15202
rect 82796 15148 82964 15150
rect 82796 15138 82852 15148
rect 82796 14532 82852 14542
rect 82684 14530 82852 14532
rect 82684 14478 82798 14530
rect 82850 14478 82852 14530
rect 82684 14476 82852 14478
rect 82908 14532 82964 15148
rect 86044 15148 86100 17390
rect 86044 15092 86324 15148
rect 85268 14924 85948 14934
rect 85324 14868 85372 14924
rect 85428 14922 85476 14924
rect 85532 14922 85580 14924
rect 85448 14870 85476 14922
rect 85572 14870 85580 14922
rect 85428 14868 85476 14870
rect 85532 14868 85580 14870
rect 85636 14922 85684 14924
rect 85740 14922 85788 14924
rect 85636 14870 85644 14922
rect 85740 14870 85768 14922
rect 85636 14868 85684 14870
rect 85740 14868 85788 14870
rect 85844 14868 85892 14924
rect 85268 14858 85948 14868
rect 83020 14532 83076 14542
rect 82908 14476 83020 14532
rect 82796 14466 82852 14476
rect 83020 14466 83076 14476
rect 81676 14418 81956 14420
rect 81676 14366 81678 14418
rect 81730 14366 81956 14418
rect 81676 14364 81956 14366
rect 81676 14354 81732 14364
rect 80768 14140 81448 14150
rect 80824 14084 80872 14140
rect 80928 14138 80976 14140
rect 81032 14138 81080 14140
rect 80948 14086 80976 14138
rect 81072 14086 81080 14138
rect 80928 14084 80976 14086
rect 81032 14084 81080 14086
rect 81136 14138 81184 14140
rect 81240 14138 81288 14140
rect 81136 14086 81144 14138
rect 81240 14086 81268 14138
rect 81136 14084 81184 14086
rect 81240 14084 81288 14086
rect 81344 14084 81392 14140
rect 80768 14074 81448 14084
rect 80444 13748 80500 13758
rect 80444 13074 80500 13692
rect 81788 13748 81844 13758
rect 81788 13654 81844 13692
rect 80444 13022 80446 13074
rect 80498 13022 80500 13074
rect 80444 13010 80500 13022
rect 81788 12740 81844 12750
rect 80768 12572 81448 12582
rect 80824 12516 80872 12572
rect 80928 12570 80976 12572
rect 81032 12570 81080 12572
rect 80948 12518 80976 12570
rect 81072 12518 81080 12570
rect 80928 12516 80976 12518
rect 81032 12516 81080 12518
rect 81136 12570 81184 12572
rect 81240 12570 81288 12572
rect 81136 12518 81144 12570
rect 81240 12518 81268 12570
rect 81136 12516 81184 12518
rect 81240 12516 81288 12518
rect 81344 12516 81392 12572
rect 80768 12506 81448 12516
rect 81564 12292 81620 12302
rect 81340 12180 81396 12190
rect 81340 12178 81508 12180
rect 81340 12126 81342 12178
rect 81394 12126 81508 12178
rect 81340 12124 81508 12126
rect 81340 12114 81396 12124
rect 81452 11172 81508 12124
rect 81452 11106 81508 11116
rect 80768 11004 81448 11014
rect 80824 10948 80872 11004
rect 80928 11002 80976 11004
rect 81032 11002 81080 11004
rect 80948 10950 80976 11002
rect 81072 10950 81080 11002
rect 80928 10948 80976 10950
rect 81032 10948 81080 10950
rect 81136 11002 81184 11004
rect 81240 11002 81288 11004
rect 81136 10950 81144 11002
rect 81240 10950 81268 11002
rect 81136 10948 81184 10950
rect 81240 10948 81288 10950
rect 81344 10948 81392 11004
rect 80768 10938 81448 10948
rect 81564 10610 81620 12236
rect 81564 10558 81566 10610
rect 81618 10558 81620 10610
rect 81564 10546 81620 10558
rect 81452 9828 81508 9838
rect 81452 9826 81620 9828
rect 81452 9774 81454 9826
rect 81506 9774 81620 9826
rect 81452 9772 81620 9774
rect 81452 9762 81508 9772
rect 80768 9436 81448 9446
rect 80824 9380 80872 9436
rect 80928 9434 80976 9436
rect 81032 9434 81080 9436
rect 80948 9382 80976 9434
rect 81072 9382 81080 9434
rect 80928 9380 80976 9382
rect 81032 9380 81080 9382
rect 81136 9434 81184 9436
rect 81240 9434 81288 9436
rect 81136 9382 81144 9434
rect 81240 9382 81268 9434
rect 81136 9380 81184 9382
rect 81240 9380 81288 9382
rect 81344 9380 81392 9436
rect 80768 9370 81448 9380
rect 80668 9156 80724 9166
rect 80668 9062 80724 9100
rect 81564 8428 81620 9772
rect 81788 8428 81844 12684
rect 81900 12068 81956 14364
rect 83132 14420 83188 14430
rect 83132 14326 83188 14364
rect 82236 14308 82292 14318
rect 82236 14214 82292 14252
rect 82796 13746 82852 13758
rect 82796 13694 82798 13746
rect 82850 13694 82852 13746
rect 82684 13634 82740 13646
rect 82684 13582 82686 13634
rect 82738 13582 82740 13634
rect 81900 12002 81956 12012
rect 82236 12962 82292 12974
rect 82236 12910 82238 12962
rect 82290 12910 82292 12962
rect 81900 11394 81956 11406
rect 81900 11342 81902 11394
rect 81954 11342 81956 11394
rect 81900 9044 81956 11342
rect 81900 8978 81956 8988
rect 82124 11172 82180 11182
rect 79324 8372 80052 8428
rect 80332 8372 80500 8428
rect 79100 5182 79102 5234
rect 79154 5182 79156 5234
rect 79100 5170 79156 5182
rect 79436 5794 79492 5806
rect 79436 5742 79438 5794
rect 79490 5742 79492 5794
rect 77868 4340 77924 4350
rect 77868 4004 77924 4284
rect 77980 4228 78036 4238
rect 78540 4228 78596 4396
rect 78876 4386 78932 4396
rect 79436 4340 79492 5742
rect 79436 4274 79492 4284
rect 79996 4564 80052 8372
rect 80108 5908 80164 5918
rect 80108 5814 80164 5852
rect 80444 5460 80500 8372
rect 81452 8370 81508 8382
rect 81564 8372 81732 8428
rect 81452 8318 81454 8370
rect 81506 8318 81508 8370
rect 81452 8258 81508 8318
rect 81452 8206 81454 8258
rect 81506 8206 81508 8258
rect 81452 8194 81508 8206
rect 80768 7868 81448 7878
rect 80824 7812 80872 7868
rect 80928 7866 80976 7868
rect 81032 7866 81080 7868
rect 80948 7814 80976 7866
rect 81072 7814 81080 7866
rect 80928 7812 80976 7814
rect 81032 7812 81080 7814
rect 81136 7866 81184 7868
rect 81240 7866 81288 7868
rect 81136 7814 81144 7866
rect 81240 7814 81268 7866
rect 81136 7812 81184 7814
rect 81240 7812 81288 7814
rect 81344 7812 81392 7868
rect 80768 7802 81448 7812
rect 81564 7362 81620 7374
rect 81564 7310 81566 7362
rect 81618 7310 81620 7362
rect 80768 6300 81448 6310
rect 80824 6244 80872 6300
rect 80928 6298 80976 6300
rect 81032 6298 81080 6300
rect 80948 6246 80976 6298
rect 81072 6246 81080 6298
rect 80928 6244 80976 6246
rect 81032 6244 81080 6246
rect 81136 6298 81184 6300
rect 81240 6298 81288 6300
rect 81136 6246 81144 6298
rect 81240 6246 81268 6298
rect 81136 6244 81184 6246
rect 81240 6244 81288 6246
rect 81344 6244 81392 6300
rect 80768 6234 81448 6244
rect 80444 5394 80500 5404
rect 81564 5348 81620 7310
rect 81676 6804 81732 8372
rect 81788 8372 81956 8428
rect 81788 8370 81844 8372
rect 81788 8318 81790 8370
rect 81842 8318 81844 8370
rect 81788 8306 81844 8318
rect 81900 8036 81956 8372
rect 81900 8034 82068 8036
rect 81900 7982 81902 8034
rect 81954 7982 82068 8034
rect 81900 7980 82068 7982
rect 81900 7970 81956 7980
rect 81676 6738 81732 6748
rect 81788 6580 81844 6590
rect 81788 6486 81844 6524
rect 81564 5282 81620 5292
rect 81676 6468 81732 6478
rect 80668 5236 80724 5246
rect 80668 4900 80724 5180
rect 80556 4844 80724 4900
rect 81676 5124 81732 6412
rect 80556 4564 80612 4844
rect 80768 4732 81448 4742
rect 80824 4676 80872 4732
rect 80928 4730 80976 4732
rect 81032 4730 81080 4732
rect 80948 4678 80976 4730
rect 81072 4678 81080 4730
rect 80928 4676 80976 4678
rect 81032 4676 81080 4678
rect 81136 4730 81184 4732
rect 81240 4730 81288 4732
rect 81136 4678 81144 4730
rect 81240 4678 81268 4730
rect 81136 4676 81184 4678
rect 81240 4676 81288 4678
rect 81344 4676 81392 4732
rect 80768 4666 81448 4676
rect 80556 4508 80724 4564
rect 77980 4226 78596 4228
rect 77980 4174 77982 4226
rect 78034 4174 78596 4226
rect 77980 4172 78596 4174
rect 78876 4226 78932 4238
rect 78876 4174 78878 4226
rect 78930 4174 78932 4226
rect 77980 4162 78036 4172
rect 78876 4116 78932 4174
rect 79212 4228 79268 4238
rect 79268 4172 79380 4228
rect 79212 4162 79268 4172
rect 79324 4116 79380 4172
rect 79436 4116 79492 4126
rect 79324 4114 79492 4116
rect 79324 4062 79438 4114
rect 79490 4062 79492 4114
rect 79324 4060 79492 4062
rect 78876 4050 78932 4060
rect 79436 4050 79492 4060
rect 77868 3948 78148 4004
rect 77980 3780 78036 3790
rect 77756 3778 78036 3780
rect 77756 3726 77982 3778
rect 78034 3726 78036 3778
rect 77756 3724 78036 3726
rect 77980 3714 78036 3724
rect 77308 3502 77310 3554
rect 77362 3502 77364 3554
rect 77308 3490 77364 3502
rect 78092 3668 78148 3948
rect 78092 3554 78148 3612
rect 79996 3666 80052 4508
rect 79996 3614 79998 3666
rect 80050 3614 80052 3666
rect 79996 3602 80052 3614
rect 78092 3502 78094 3554
rect 78146 3502 78148 3554
rect 78092 3490 78148 3502
rect 80668 3554 80724 4508
rect 81564 4340 81620 4350
rect 81676 4340 81732 5068
rect 81900 6466 81956 6478
rect 81900 6414 81902 6466
rect 81954 6414 81956 6466
rect 81900 5124 81956 6414
rect 81900 5058 81956 5068
rect 82012 4452 82068 7980
rect 82124 6692 82180 11116
rect 82236 10388 82292 12910
rect 82572 12180 82628 12190
rect 82572 12086 82628 12124
rect 82236 10322 82292 10332
rect 82124 6626 82180 6636
rect 82684 6692 82740 13582
rect 82796 13636 82852 13694
rect 82796 13570 82852 13580
rect 83580 13746 83636 13758
rect 83580 13694 83582 13746
rect 83634 13694 83636 13746
rect 83580 13636 83636 13694
rect 83580 13570 83636 13580
rect 85268 13356 85948 13366
rect 85324 13300 85372 13356
rect 85428 13354 85476 13356
rect 85532 13354 85580 13356
rect 85448 13302 85476 13354
rect 85572 13302 85580 13354
rect 85428 13300 85476 13302
rect 85532 13300 85580 13302
rect 85636 13354 85684 13356
rect 85740 13354 85788 13356
rect 85636 13302 85644 13354
rect 85740 13302 85768 13354
rect 85636 13300 85684 13302
rect 85740 13300 85788 13302
rect 85844 13300 85892 13356
rect 85268 13290 85948 13300
rect 83468 12178 83524 12190
rect 83468 12126 83470 12178
rect 83522 12126 83524 12178
rect 83468 12068 83524 12126
rect 83804 12068 83860 12078
rect 83468 12012 83804 12068
rect 83804 11974 83860 12012
rect 86044 12068 86100 12078
rect 83916 11954 83972 11966
rect 83916 11902 83918 11954
rect 83970 11902 83972 11954
rect 83916 10052 83972 11902
rect 85268 11788 85948 11798
rect 85324 11732 85372 11788
rect 85428 11786 85476 11788
rect 85532 11786 85580 11788
rect 85448 11734 85476 11786
rect 85572 11734 85580 11786
rect 85428 11732 85476 11734
rect 85532 11732 85580 11734
rect 85636 11786 85684 11788
rect 85740 11786 85788 11788
rect 85636 11734 85644 11786
rect 85740 11734 85768 11786
rect 85636 11732 85684 11734
rect 85740 11732 85788 11734
rect 85844 11732 85892 11788
rect 85268 11722 85948 11732
rect 85148 10498 85204 10510
rect 85148 10446 85150 10498
rect 85202 10446 85204 10498
rect 85148 10052 85204 10446
rect 85268 10220 85948 10230
rect 85324 10164 85372 10220
rect 85428 10218 85476 10220
rect 85532 10218 85580 10220
rect 85448 10166 85476 10218
rect 85572 10166 85580 10218
rect 85428 10164 85476 10166
rect 85532 10164 85580 10166
rect 85636 10218 85684 10220
rect 85740 10218 85788 10220
rect 85636 10166 85644 10218
rect 85740 10166 85768 10218
rect 85636 10164 85684 10166
rect 85740 10164 85788 10166
rect 85844 10164 85892 10220
rect 85268 10154 85948 10164
rect 83916 9996 84308 10052
rect 82684 6626 82740 6636
rect 82796 9716 82852 9726
rect 82348 6468 82404 6478
rect 82348 6374 82404 6412
rect 82124 5236 82180 5246
rect 82124 5010 82180 5180
rect 82124 4958 82126 5010
rect 82178 4958 82180 5010
rect 82124 4946 82180 4958
rect 82460 5124 82516 5134
rect 82124 4452 82180 4462
rect 82012 4450 82180 4452
rect 82012 4398 82126 4450
rect 82178 4398 82180 4450
rect 82012 4396 82180 4398
rect 82124 4386 82180 4396
rect 81564 4338 81732 4340
rect 81564 4286 81566 4338
rect 81618 4286 81732 4338
rect 81564 4284 81732 4286
rect 81564 4274 81620 4284
rect 82460 3666 82516 5068
rect 82460 3614 82462 3666
rect 82514 3614 82516 3666
rect 82460 3602 82516 3614
rect 80668 3502 80670 3554
rect 80722 3502 80724 3554
rect 80668 3490 80724 3502
rect 82796 3554 82852 9660
rect 84028 9044 84084 9054
rect 84028 8950 84084 8988
rect 83916 7476 83972 7486
rect 84028 7476 84084 7486
rect 83972 7474 84084 7476
rect 83972 7422 84030 7474
rect 84082 7422 84084 7474
rect 83972 7420 84084 7422
rect 83916 6018 83972 7420
rect 84028 7410 84084 7420
rect 84028 6692 84084 6702
rect 84028 6598 84084 6636
rect 83916 5966 83918 6018
rect 83970 5966 83972 6018
rect 83916 5954 83972 5966
rect 83244 5122 83300 5134
rect 83244 5070 83246 5122
rect 83298 5070 83300 5122
rect 83244 3668 83300 5070
rect 84252 5122 84308 9996
rect 85148 9986 85204 9996
rect 84364 9716 84420 9726
rect 84364 9622 84420 9660
rect 85268 8652 85948 8662
rect 85324 8596 85372 8652
rect 85428 8650 85476 8652
rect 85532 8650 85580 8652
rect 85448 8598 85476 8650
rect 85572 8598 85580 8650
rect 85428 8596 85476 8598
rect 85532 8596 85580 8598
rect 85636 8650 85684 8652
rect 85740 8650 85788 8652
rect 85636 8598 85644 8650
rect 85740 8598 85768 8650
rect 85636 8596 85684 8598
rect 85740 8596 85788 8598
rect 85844 8596 85892 8652
rect 85268 8586 85948 8596
rect 85268 7084 85948 7094
rect 85324 7028 85372 7084
rect 85428 7082 85476 7084
rect 85532 7082 85580 7084
rect 85448 7030 85476 7082
rect 85572 7030 85580 7082
rect 85428 7028 85476 7030
rect 85532 7028 85580 7030
rect 85636 7082 85684 7084
rect 85740 7082 85788 7084
rect 85636 7030 85644 7082
rect 85740 7030 85768 7082
rect 85636 7028 85684 7030
rect 85740 7028 85788 7030
rect 85844 7028 85892 7084
rect 85268 7018 85948 7028
rect 85268 5516 85948 5526
rect 85324 5460 85372 5516
rect 85428 5514 85476 5516
rect 85532 5514 85580 5516
rect 85448 5462 85476 5514
rect 85572 5462 85580 5514
rect 85428 5460 85476 5462
rect 85532 5460 85580 5462
rect 85636 5514 85684 5516
rect 85740 5514 85788 5516
rect 85636 5462 85644 5514
rect 85740 5462 85768 5514
rect 85636 5460 85684 5462
rect 85740 5460 85788 5462
rect 85844 5460 85892 5516
rect 85268 5450 85948 5460
rect 84252 5070 84254 5122
rect 84306 5070 84308 5122
rect 84252 5058 84308 5070
rect 84700 5236 84756 5246
rect 83244 3602 83300 3612
rect 84700 3666 84756 5180
rect 85932 4228 85988 4238
rect 85932 4134 85988 4172
rect 85268 3948 85948 3958
rect 85324 3892 85372 3948
rect 85428 3946 85476 3948
rect 85532 3946 85580 3948
rect 85448 3894 85476 3946
rect 85572 3894 85580 3946
rect 85428 3892 85476 3894
rect 85532 3892 85580 3894
rect 85636 3946 85684 3948
rect 85740 3946 85788 3948
rect 85636 3894 85644 3946
rect 85740 3894 85768 3946
rect 85636 3892 85684 3894
rect 85740 3892 85788 3894
rect 85844 3892 85892 3948
rect 85268 3882 85948 3892
rect 84700 3614 84702 3666
rect 84754 3614 84756 3666
rect 84700 3602 84756 3614
rect 85708 3668 85764 3678
rect 86044 3668 86100 12012
rect 86156 8146 86212 8158
rect 86156 8094 86158 8146
rect 86210 8094 86212 8146
rect 86156 6580 86212 8094
rect 86156 6514 86212 6524
rect 86268 4564 86324 15092
rect 87388 9268 87444 21646
rect 96908 21586 96964 21756
rect 96908 21534 96910 21586
rect 96962 21534 96964 21586
rect 96908 21522 96964 21534
rect 98028 21474 98084 21486
rect 98028 21422 98030 21474
rect 98082 21422 98084 21474
rect 94268 21196 94948 21206
rect 94324 21140 94372 21196
rect 94428 21194 94476 21196
rect 94532 21194 94580 21196
rect 94448 21142 94476 21194
rect 94572 21142 94580 21194
rect 94428 21140 94476 21142
rect 94532 21140 94580 21142
rect 94636 21194 94684 21196
rect 94740 21194 94788 21196
rect 94636 21142 94644 21194
rect 94740 21142 94768 21194
rect 94636 21140 94684 21142
rect 94740 21140 94788 21142
rect 94844 21140 94892 21196
rect 94268 21130 94948 21140
rect 98028 20916 98084 21422
rect 98028 20850 98084 20860
rect 89768 20412 90448 20422
rect 89824 20356 89872 20412
rect 89928 20410 89976 20412
rect 90032 20410 90080 20412
rect 89948 20358 89976 20410
rect 90072 20358 90080 20410
rect 89928 20356 89976 20358
rect 90032 20356 90080 20358
rect 90136 20410 90184 20412
rect 90240 20410 90288 20412
rect 90136 20358 90144 20410
rect 90240 20358 90268 20410
rect 90136 20356 90184 20358
rect 90240 20356 90288 20358
rect 90344 20356 90392 20412
rect 89768 20346 90448 20356
rect 89068 20132 89124 20142
rect 89068 19458 89124 20076
rect 94268 19628 94948 19638
rect 94324 19572 94372 19628
rect 94428 19626 94476 19628
rect 94532 19626 94580 19628
rect 94448 19574 94476 19626
rect 94572 19574 94580 19626
rect 94428 19572 94476 19574
rect 94532 19572 94580 19574
rect 94636 19626 94684 19628
rect 94740 19626 94788 19628
rect 94636 19574 94644 19626
rect 94740 19574 94768 19626
rect 94636 19572 94684 19574
rect 94740 19572 94788 19574
rect 94844 19572 94892 19628
rect 94268 19562 94948 19572
rect 89068 19406 89070 19458
rect 89122 19406 89124 19458
rect 88284 19012 88340 19022
rect 88284 18918 88340 18956
rect 89068 18564 89124 19406
rect 96908 19234 96964 19246
rect 96908 19182 96910 19234
rect 96962 19182 96964 19234
rect 96684 19124 96740 19134
rect 96908 19124 96964 19182
rect 96740 19068 96964 19124
rect 98028 19124 98084 19134
rect 96684 19030 96740 19068
rect 98028 19030 98084 19068
rect 89768 18844 90448 18854
rect 89824 18788 89872 18844
rect 89928 18842 89976 18844
rect 90032 18842 90080 18844
rect 89948 18790 89976 18842
rect 90072 18790 90080 18842
rect 89928 18788 89976 18790
rect 90032 18788 90080 18790
rect 90136 18842 90184 18844
rect 90240 18842 90288 18844
rect 90136 18790 90144 18842
rect 90240 18790 90268 18842
rect 90136 18788 90184 18790
rect 90240 18788 90288 18790
rect 90344 18788 90392 18844
rect 89768 18778 90448 18788
rect 89068 18498 89124 18508
rect 89964 18564 90020 18574
rect 89964 18470 90020 18508
rect 90300 18562 90356 18574
rect 90300 18510 90302 18562
rect 90354 18510 90356 18562
rect 90300 17444 90356 18510
rect 94268 18060 94948 18070
rect 94324 18004 94372 18060
rect 94428 18058 94476 18060
rect 94532 18058 94580 18060
rect 94448 18006 94476 18058
rect 94572 18006 94580 18058
rect 94428 18004 94476 18006
rect 94532 18004 94580 18006
rect 94636 18058 94684 18060
rect 94740 18058 94788 18060
rect 94636 18006 94644 18058
rect 94740 18006 94768 18058
rect 94636 18004 94684 18006
rect 94740 18004 94788 18006
rect 94844 18004 94892 18060
rect 94268 17994 94948 18004
rect 96908 17666 96964 17678
rect 96908 17614 96910 17666
rect 96962 17614 96964 17666
rect 96684 17444 96740 17454
rect 96908 17444 96964 17614
rect 90300 17388 90580 17444
rect 89768 17276 90448 17286
rect 89824 17220 89872 17276
rect 89928 17274 89976 17276
rect 90032 17274 90080 17276
rect 89948 17222 89976 17274
rect 90072 17222 90080 17274
rect 89928 17220 89976 17222
rect 90032 17220 90080 17222
rect 90136 17274 90184 17276
rect 90240 17274 90288 17276
rect 90136 17222 90144 17274
rect 90240 17222 90268 17274
rect 90136 17220 90184 17222
rect 90240 17220 90288 17222
rect 90344 17220 90392 17276
rect 89768 17210 90448 17220
rect 89768 15708 90448 15718
rect 89824 15652 89872 15708
rect 89928 15706 89976 15708
rect 90032 15706 90080 15708
rect 89948 15654 89976 15706
rect 90072 15654 90080 15706
rect 89928 15652 89976 15654
rect 90032 15652 90080 15654
rect 90136 15706 90184 15708
rect 90240 15706 90288 15708
rect 90136 15654 90144 15706
rect 90240 15654 90268 15706
rect 90136 15652 90184 15654
rect 90240 15652 90288 15654
rect 90344 15652 90392 15708
rect 89768 15642 90448 15652
rect 88172 14308 88228 14318
rect 87388 9202 87444 9212
rect 88060 10052 88116 10062
rect 87500 9044 87556 9054
rect 87500 5234 87556 8988
rect 88060 8258 88116 9996
rect 88060 8206 88062 8258
rect 88114 8206 88116 8258
rect 87948 7474 88004 7486
rect 87948 7422 87950 7474
rect 88002 7422 88004 7474
rect 87948 6804 88004 7422
rect 87948 6710 88004 6748
rect 87500 5182 87502 5234
rect 87554 5182 87556 5234
rect 87500 5170 87556 5182
rect 86268 4498 86324 4508
rect 88060 4338 88116 8206
rect 88172 5906 88228 14252
rect 89768 14140 90448 14150
rect 89824 14084 89872 14140
rect 89928 14138 89976 14140
rect 90032 14138 90080 14140
rect 89948 14086 89976 14138
rect 90072 14086 90080 14138
rect 89928 14084 89976 14086
rect 90032 14084 90080 14086
rect 90136 14138 90184 14140
rect 90240 14138 90288 14140
rect 90136 14086 90144 14138
rect 90240 14086 90268 14138
rect 90136 14084 90184 14086
rect 90240 14084 90288 14086
rect 90344 14084 90392 14140
rect 89768 14074 90448 14084
rect 89768 12572 90448 12582
rect 89824 12516 89872 12572
rect 89928 12570 89976 12572
rect 90032 12570 90080 12572
rect 89948 12518 89976 12570
rect 90072 12518 90080 12570
rect 89928 12516 89976 12518
rect 90032 12516 90080 12518
rect 90136 12570 90184 12572
rect 90240 12570 90288 12572
rect 90136 12518 90144 12570
rect 90240 12518 90268 12570
rect 90136 12516 90184 12518
rect 90240 12516 90288 12518
rect 90344 12516 90392 12572
rect 89768 12506 90448 12516
rect 89768 11004 90448 11014
rect 89824 10948 89872 11004
rect 89928 11002 89976 11004
rect 90032 11002 90080 11004
rect 89948 10950 89976 11002
rect 90072 10950 90080 11002
rect 89928 10948 89976 10950
rect 90032 10948 90080 10950
rect 90136 11002 90184 11004
rect 90240 11002 90288 11004
rect 90136 10950 90144 11002
rect 90240 10950 90268 11002
rect 90136 10948 90184 10950
rect 90240 10948 90288 10950
rect 90344 10948 90392 11004
rect 89768 10938 90448 10948
rect 88956 10388 89012 10398
rect 88956 9826 89012 10332
rect 88956 9774 88958 9826
rect 89010 9774 89012 9826
rect 88956 8372 89012 9774
rect 89768 9436 90448 9446
rect 89824 9380 89872 9436
rect 89928 9434 89976 9436
rect 90032 9434 90080 9436
rect 89948 9382 89976 9434
rect 90072 9382 90080 9434
rect 89928 9380 89976 9382
rect 90032 9380 90080 9382
rect 90136 9434 90184 9436
rect 90240 9434 90288 9436
rect 90136 9382 90144 9434
rect 90240 9382 90268 9434
rect 90136 9380 90184 9382
rect 90240 9380 90288 9382
rect 90344 9380 90392 9436
rect 89768 9370 90448 9380
rect 88956 8306 89012 8316
rect 89768 7868 90448 7878
rect 89824 7812 89872 7868
rect 89928 7866 89976 7868
rect 90032 7866 90080 7868
rect 89948 7814 89976 7866
rect 90072 7814 90080 7866
rect 89928 7812 89976 7814
rect 90032 7812 90080 7814
rect 90136 7866 90184 7868
rect 90240 7866 90288 7868
rect 90136 7814 90144 7866
rect 90240 7814 90268 7866
rect 90136 7812 90184 7814
rect 90240 7812 90288 7814
rect 90344 7812 90392 7868
rect 89768 7802 90448 7812
rect 90524 6692 90580 17388
rect 96740 17388 96964 17444
rect 98028 17554 98084 17566
rect 98028 17502 98030 17554
rect 98082 17502 98084 17554
rect 96684 17350 96740 17388
rect 98028 17332 98084 17502
rect 98028 17266 98084 17276
rect 94268 16492 94948 16502
rect 94324 16436 94372 16492
rect 94428 16490 94476 16492
rect 94532 16490 94580 16492
rect 94448 16438 94476 16490
rect 94572 16438 94580 16490
rect 94428 16436 94476 16438
rect 94532 16436 94580 16438
rect 94636 16490 94684 16492
rect 94740 16490 94788 16492
rect 94636 16438 94644 16490
rect 94740 16438 94768 16490
rect 94636 16436 94684 16438
rect 94740 16436 94788 16438
rect 94844 16436 94892 16492
rect 94268 16426 94948 16436
rect 96684 16100 96740 16110
rect 96908 16100 96964 16110
rect 96740 16098 96964 16100
rect 96740 16046 96910 16098
rect 96962 16046 96964 16098
rect 96740 16044 96964 16046
rect 96684 16006 96740 16044
rect 96908 16034 96964 16044
rect 98028 15986 98084 15998
rect 98028 15934 98030 15986
rect 98082 15934 98084 15986
rect 98028 15540 98084 15934
rect 98028 15474 98084 15484
rect 94268 14924 94948 14934
rect 94324 14868 94372 14924
rect 94428 14922 94476 14924
rect 94532 14922 94580 14924
rect 94448 14870 94476 14922
rect 94572 14870 94580 14922
rect 94428 14868 94476 14870
rect 94532 14868 94580 14870
rect 94636 14922 94684 14924
rect 94740 14922 94788 14924
rect 94636 14870 94644 14922
rect 94740 14870 94768 14922
rect 94636 14868 94684 14870
rect 94740 14868 94788 14870
rect 94844 14868 94892 14924
rect 94268 14858 94948 14868
rect 90860 14532 90916 14542
rect 90524 6626 90580 6636
rect 90748 8372 90804 8382
rect 89768 6300 90448 6310
rect 89824 6244 89872 6300
rect 89928 6298 89976 6300
rect 90032 6298 90080 6300
rect 89948 6246 89976 6298
rect 90072 6246 90080 6298
rect 89928 6244 89976 6246
rect 90032 6244 90080 6246
rect 90136 6298 90184 6300
rect 90240 6298 90288 6300
rect 90136 6246 90144 6298
rect 90240 6246 90268 6298
rect 90136 6244 90184 6246
rect 90240 6244 90288 6246
rect 90344 6244 90392 6300
rect 89768 6234 90448 6244
rect 90748 6018 90804 8316
rect 90860 7586 90916 14476
rect 96908 14532 96964 14542
rect 96908 14438 96964 14476
rect 98028 14418 98084 14430
rect 98028 14366 98030 14418
rect 98082 14366 98084 14418
rect 98028 13748 98084 14366
rect 98028 13682 98084 13692
rect 94268 13356 94948 13366
rect 94324 13300 94372 13356
rect 94428 13354 94476 13356
rect 94532 13354 94580 13356
rect 94448 13302 94476 13354
rect 94572 13302 94580 13354
rect 94428 13300 94476 13302
rect 94532 13300 94580 13302
rect 94636 13354 94684 13356
rect 94740 13354 94788 13356
rect 94636 13302 94644 13354
rect 94740 13302 94768 13354
rect 94636 13300 94684 13302
rect 94740 13300 94788 13302
rect 94844 13300 94892 13356
rect 94268 13290 94948 13300
rect 96572 12292 96628 12302
rect 96628 12236 96964 12292
rect 96572 12198 96628 12236
rect 90860 7534 90862 7586
rect 90914 7534 90916 7586
rect 90860 7522 90916 7534
rect 91196 12180 91252 12190
rect 90748 5966 90750 6018
rect 90802 5966 90804 6018
rect 90748 5954 90804 5966
rect 88172 5854 88174 5906
rect 88226 5854 88228 5906
rect 88172 5842 88228 5854
rect 89768 4732 90448 4742
rect 89824 4676 89872 4732
rect 89928 4730 89976 4732
rect 90032 4730 90080 4732
rect 89948 4678 89976 4730
rect 90072 4678 90080 4730
rect 89928 4676 89976 4678
rect 90032 4676 90080 4678
rect 90136 4730 90184 4732
rect 90240 4730 90288 4732
rect 90136 4678 90144 4730
rect 90240 4678 90268 4730
rect 90136 4676 90184 4678
rect 90240 4676 90288 4678
rect 90344 4676 90392 4732
rect 89768 4666 90448 4676
rect 91196 4562 91252 12124
rect 96908 12178 96964 12236
rect 96908 12126 96910 12178
rect 96962 12126 96964 12178
rect 96908 12114 96964 12126
rect 98028 12066 98084 12078
rect 98028 12014 98030 12066
rect 98082 12014 98084 12066
rect 98028 11956 98084 12014
rect 98028 11890 98084 11900
rect 94268 11788 94948 11798
rect 94324 11732 94372 11788
rect 94428 11786 94476 11788
rect 94532 11786 94580 11788
rect 94448 11734 94476 11786
rect 94572 11734 94580 11786
rect 94428 11732 94476 11734
rect 94532 11732 94580 11734
rect 94636 11786 94684 11788
rect 94740 11786 94788 11788
rect 94636 11734 94644 11786
rect 94740 11734 94768 11786
rect 94636 11732 94684 11734
rect 94740 11732 94788 11734
rect 94844 11732 94892 11788
rect 94268 11722 94948 11732
rect 96684 10724 96740 10734
rect 96740 10668 96964 10724
rect 96684 10630 96740 10668
rect 96908 10610 96964 10668
rect 96908 10558 96910 10610
rect 96962 10558 96964 10610
rect 96908 10546 96964 10558
rect 98028 10498 98084 10510
rect 98028 10446 98030 10498
rect 98082 10446 98084 10498
rect 94268 10220 94948 10230
rect 94324 10164 94372 10220
rect 94428 10218 94476 10220
rect 94532 10218 94580 10220
rect 94448 10166 94476 10218
rect 94572 10166 94580 10218
rect 94428 10164 94476 10166
rect 94532 10164 94580 10166
rect 94636 10218 94684 10220
rect 94740 10218 94788 10220
rect 94636 10166 94644 10218
rect 94740 10166 94768 10218
rect 94636 10164 94684 10166
rect 94740 10164 94788 10166
rect 94844 10164 94892 10220
rect 94268 10154 94948 10164
rect 98028 10164 98084 10446
rect 98028 10098 98084 10108
rect 96684 9268 96740 9278
rect 96908 9268 96964 9278
rect 96740 9266 96964 9268
rect 96740 9214 96910 9266
rect 96962 9214 96964 9266
rect 96740 9212 96964 9214
rect 96684 9174 96740 9212
rect 96908 9202 96964 9212
rect 97692 8818 97748 8830
rect 97692 8766 97694 8818
rect 97746 8766 97748 8818
rect 94268 8652 94948 8662
rect 94324 8596 94372 8652
rect 94428 8650 94476 8652
rect 94532 8650 94580 8652
rect 94448 8598 94476 8650
rect 94572 8598 94580 8650
rect 94428 8596 94476 8598
rect 94532 8596 94580 8598
rect 94636 8650 94684 8652
rect 94740 8650 94788 8652
rect 94636 8598 94644 8650
rect 94740 8598 94768 8650
rect 94636 8596 94684 8598
rect 94740 8596 94788 8598
rect 94844 8596 94892 8652
rect 94268 8586 94948 8596
rect 97692 8372 97748 8766
rect 97692 8306 97748 8316
rect 94268 7084 94948 7094
rect 94324 7028 94372 7084
rect 94428 7082 94476 7084
rect 94532 7082 94580 7084
rect 94448 7030 94476 7082
rect 94572 7030 94580 7082
rect 94428 7028 94476 7030
rect 94532 7028 94580 7030
rect 94636 7082 94684 7084
rect 94740 7082 94788 7084
rect 94636 7030 94644 7082
rect 94740 7030 94768 7082
rect 94636 7028 94684 7030
rect 94740 7028 94788 7030
rect 94844 7028 94892 7084
rect 94268 7018 94948 7028
rect 96684 6692 96740 6702
rect 96908 6692 96964 6702
rect 96740 6690 96964 6692
rect 96740 6638 96910 6690
rect 96962 6638 96964 6690
rect 96740 6636 96964 6638
rect 96684 6598 96740 6636
rect 96908 6626 96964 6636
rect 98028 6580 98084 6590
rect 98028 6486 98084 6524
rect 94268 5516 94948 5526
rect 94324 5460 94372 5516
rect 94428 5514 94476 5516
rect 94532 5514 94580 5516
rect 94448 5462 94476 5514
rect 94572 5462 94580 5514
rect 94428 5460 94476 5462
rect 94532 5460 94580 5462
rect 94636 5514 94684 5516
rect 94740 5514 94788 5516
rect 94636 5462 94644 5514
rect 94740 5462 94768 5514
rect 94636 5460 94684 5462
rect 94740 5460 94788 5462
rect 94844 5460 94892 5516
rect 94268 5450 94948 5460
rect 96572 5348 96628 5358
rect 96572 5236 96628 5292
rect 96572 5234 96964 5236
rect 96572 5182 96574 5234
rect 96626 5182 96964 5234
rect 96572 5180 96964 5182
rect 96572 5170 96628 5180
rect 96908 5122 96964 5180
rect 96908 5070 96910 5122
rect 96962 5070 96964 5122
rect 96908 5058 96964 5070
rect 97692 5122 97748 5134
rect 97692 5070 97694 5122
rect 97746 5070 97748 5122
rect 97692 4788 97748 5070
rect 97692 4722 97748 4732
rect 91196 4510 91198 4562
rect 91250 4510 91252 4562
rect 91196 4498 91252 4510
rect 96684 4564 96740 4574
rect 96908 4564 96964 4574
rect 96740 4562 96964 4564
rect 96740 4510 96910 4562
rect 96962 4510 96964 4562
rect 96740 4508 96964 4510
rect 96684 4470 96740 4508
rect 96908 4498 96964 4508
rect 88060 4286 88062 4338
rect 88114 4286 88116 4338
rect 88060 4274 88116 4286
rect 85708 3666 86100 3668
rect 85708 3614 85710 3666
rect 85762 3614 86100 3666
rect 85708 3612 86100 3614
rect 86156 4228 86212 4238
rect 85708 3602 85764 3612
rect 82796 3502 82798 3554
rect 82850 3502 82852 3554
rect 82796 3490 82852 3502
rect 82908 3556 82964 3566
rect 76748 3442 77252 3444
rect 76748 3390 76750 3442
rect 76802 3390 77252 3442
rect 76748 3388 77252 3390
rect 76748 3378 76804 3388
rect 76188 3332 76244 3342
rect 76076 3276 76188 3332
rect 76188 3266 76244 3276
rect 81900 3332 81956 3342
rect 81900 3238 81956 3276
rect 71768 3164 72448 3174
rect 71824 3108 71872 3164
rect 71928 3162 71976 3164
rect 72032 3162 72080 3164
rect 71948 3110 71976 3162
rect 72072 3110 72080 3162
rect 71928 3108 71976 3110
rect 72032 3108 72080 3110
rect 72136 3162 72184 3164
rect 72240 3162 72288 3164
rect 72136 3110 72144 3162
rect 72240 3110 72268 3162
rect 72136 3108 72184 3110
rect 72240 3108 72288 3110
rect 72344 3108 72392 3164
rect 71768 3098 72448 3108
rect 80768 3164 81448 3174
rect 80824 3108 80872 3164
rect 80928 3162 80976 3164
rect 81032 3162 81080 3164
rect 80948 3110 80976 3162
rect 81072 3110 81080 3162
rect 80928 3108 80976 3110
rect 81032 3108 81080 3110
rect 81136 3162 81184 3164
rect 81240 3162 81288 3164
rect 81136 3110 81144 3162
rect 81240 3110 81268 3162
rect 81136 3108 81184 3110
rect 81240 3108 81288 3110
rect 81344 3108 81392 3164
rect 80768 3098 81448 3108
rect 71596 2940 71988 2996
rect 71932 800 71988 2940
rect 82908 800 82964 3500
rect 86156 3556 86212 4172
rect 97692 4116 97748 4126
rect 97692 4114 97860 4116
rect 97692 4062 97694 4114
rect 97746 4062 97860 4114
rect 97692 4060 97860 4062
rect 97692 4050 97748 4060
rect 94268 3948 94948 3958
rect 94324 3892 94372 3948
rect 94428 3946 94476 3948
rect 94532 3946 94580 3948
rect 94448 3894 94476 3946
rect 94572 3894 94580 3946
rect 94428 3892 94476 3894
rect 94532 3892 94580 3894
rect 94636 3946 94684 3948
rect 94740 3946 94788 3948
rect 94636 3894 94644 3946
rect 94740 3894 94768 3946
rect 94636 3892 94684 3894
rect 94740 3892 94788 3894
rect 94844 3892 94892 3948
rect 94268 3882 94948 3892
rect 96348 3780 96404 3790
rect 86156 3462 86212 3500
rect 93884 3612 94276 3668
rect 83244 3444 83300 3454
rect 83244 3350 83300 3388
rect 93884 3442 93940 3612
rect 94220 3556 94276 3612
rect 96348 3666 96404 3724
rect 96348 3614 96350 3666
rect 96402 3614 96404 3666
rect 96348 3602 96404 3614
rect 96908 3780 96964 3790
rect 94332 3556 94388 3566
rect 94220 3554 94388 3556
rect 94220 3502 94334 3554
rect 94386 3502 94388 3554
rect 94220 3500 94388 3502
rect 94332 3490 94388 3500
rect 96908 3554 96964 3724
rect 96908 3502 96910 3554
rect 96962 3502 96964 3554
rect 96908 3490 96964 3502
rect 93884 3390 93886 3442
rect 93938 3390 93940 3442
rect 89768 3164 90448 3174
rect 89824 3108 89872 3164
rect 89928 3162 89976 3164
rect 90032 3162 90080 3164
rect 89948 3110 89976 3162
rect 90072 3110 90080 3162
rect 89928 3108 89976 3110
rect 90032 3108 90080 3110
rect 90136 3162 90184 3164
rect 90240 3162 90288 3164
rect 90136 3110 90144 3162
rect 90240 3110 90268 3162
rect 90136 3108 90184 3110
rect 90240 3108 90288 3110
rect 90344 3108 90392 3164
rect 89768 3098 90448 3108
rect 93884 800 93940 3390
rect 94108 3444 94164 3482
rect 94108 3378 94164 3388
rect 97692 3442 97748 3454
rect 97692 3390 97694 3442
rect 97746 3390 97748 3442
rect 97692 2996 97748 3390
rect 97692 2930 97748 2940
rect 97804 1204 97860 4060
rect 97804 1138 97860 1148
rect 6048 0 6160 800
rect 17024 0 17136 800
rect 28000 0 28112 800
rect 38976 0 39088 800
rect 49952 0 50064 800
rect 60928 0 61040 800
rect 71904 0 72016 800
rect 82880 0 82992 800
rect 93856 0 93968 800
<< via2 >>
rect 2044 56194 2100 56196
rect 2044 56142 2046 56194
rect 2046 56142 2098 56194
rect 2098 56142 2100 56194
rect 2044 56140 2100 56142
rect 8768 56420 8824 56476
rect 8872 56474 8928 56476
rect 8976 56474 9032 56476
rect 8872 56422 8896 56474
rect 8896 56422 8928 56474
rect 8976 56422 9020 56474
rect 9020 56422 9032 56474
rect 8872 56420 8928 56422
rect 8976 56420 9032 56422
rect 9080 56420 9136 56476
rect 9184 56474 9240 56476
rect 9288 56474 9344 56476
rect 9184 56422 9196 56474
rect 9196 56422 9240 56474
rect 9288 56422 9320 56474
rect 9320 56422 9344 56474
rect 9184 56420 9240 56422
rect 9288 56420 9344 56422
rect 9392 56420 9448 56476
rect 17768 56420 17824 56476
rect 17872 56474 17928 56476
rect 17976 56474 18032 56476
rect 17872 56422 17896 56474
rect 17896 56422 17928 56474
rect 17976 56422 18020 56474
rect 18020 56422 18032 56474
rect 17872 56420 17928 56422
rect 17976 56420 18032 56422
rect 18080 56420 18136 56476
rect 18184 56474 18240 56476
rect 18288 56474 18344 56476
rect 18184 56422 18196 56474
rect 18196 56422 18240 56474
rect 18288 56422 18320 56474
rect 18320 56422 18344 56474
rect 18184 56420 18240 56422
rect 18288 56420 18344 56422
rect 18392 56420 18448 56476
rect 12124 56140 12180 56196
rect 1708 55580 1764 55636
rect 8204 55916 8260 55972
rect 8764 55970 8820 55972
rect 8764 55918 8766 55970
rect 8766 55918 8818 55970
rect 8818 55918 8820 55970
rect 8764 55916 8820 55918
rect 2492 55580 2548 55636
rect 4268 55636 4324 55692
rect 4372 55690 4428 55692
rect 4476 55690 4532 55692
rect 4372 55638 4396 55690
rect 4396 55638 4428 55690
rect 4476 55638 4520 55690
rect 4520 55638 4532 55690
rect 4372 55636 4428 55638
rect 4476 55636 4532 55638
rect 4580 55636 4636 55692
rect 4684 55690 4740 55692
rect 4788 55690 4844 55692
rect 4684 55638 4696 55690
rect 4696 55638 4740 55690
rect 4788 55638 4820 55690
rect 4820 55638 4844 55690
rect 4684 55636 4740 55638
rect 4788 55636 4844 55638
rect 4892 55636 4948 55692
rect 1708 55020 1764 55076
rect 1708 54460 1764 54516
rect 2492 55074 2548 55076
rect 2492 55022 2494 55074
rect 2494 55022 2546 55074
rect 2546 55022 2548 55074
rect 2492 55020 2548 55022
rect 8768 54852 8824 54908
rect 8872 54906 8928 54908
rect 8976 54906 9032 54908
rect 8872 54854 8896 54906
rect 8896 54854 8928 54906
rect 8976 54854 9020 54906
rect 9020 54854 9032 54906
rect 8872 54852 8928 54854
rect 8976 54852 9032 54854
rect 9080 54852 9136 54908
rect 9184 54906 9240 54908
rect 9288 54906 9344 54908
rect 9184 54854 9196 54906
rect 9196 54854 9240 54906
rect 9288 54854 9320 54906
rect 9320 54854 9344 54906
rect 9184 54852 9240 54854
rect 9288 54852 9344 54854
rect 9392 54852 9448 54908
rect 4268 54068 4324 54124
rect 4372 54122 4428 54124
rect 4476 54122 4532 54124
rect 4372 54070 4396 54122
rect 4396 54070 4428 54122
rect 4476 54070 4520 54122
rect 4520 54070 4532 54122
rect 4372 54068 4428 54070
rect 4476 54068 4532 54070
rect 4580 54068 4636 54124
rect 4684 54122 4740 54124
rect 4788 54122 4844 54124
rect 4684 54070 4696 54122
rect 4696 54070 4740 54122
rect 4788 54070 4820 54122
rect 4820 54070 4844 54122
rect 4684 54068 4740 54070
rect 4788 54068 4844 54070
rect 4892 54068 4948 54124
rect 1708 53340 1764 53396
rect 1708 52780 1764 52836
rect 1708 52220 1764 52276
rect 1708 51100 1764 51156
rect 2492 53340 2548 53396
rect 8768 53284 8824 53340
rect 8872 53338 8928 53340
rect 8976 53338 9032 53340
rect 8872 53286 8896 53338
rect 8896 53286 8928 53338
rect 8976 53286 9020 53338
rect 9020 53286 9032 53338
rect 8872 53284 8928 53286
rect 8976 53284 9032 53286
rect 9080 53284 9136 53340
rect 9184 53338 9240 53340
rect 9288 53338 9344 53340
rect 9184 53286 9196 53338
rect 9196 53286 9240 53338
rect 9288 53286 9320 53338
rect 9320 53286 9344 53338
rect 9184 53284 9240 53286
rect 9288 53284 9344 53286
rect 9392 53284 9448 53340
rect 2492 52834 2548 52836
rect 2492 52782 2494 52834
rect 2494 52782 2546 52834
rect 2546 52782 2548 52834
rect 2492 52780 2548 52782
rect 4268 52500 4324 52556
rect 4372 52554 4428 52556
rect 4476 52554 4532 52556
rect 4372 52502 4396 52554
rect 4396 52502 4428 52554
rect 4476 52502 4520 52554
rect 4520 52502 4532 52554
rect 4372 52500 4428 52502
rect 4476 52500 4532 52502
rect 4580 52500 4636 52556
rect 4684 52554 4740 52556
rect 4788 52554 4844 52556
rect 4684 52502 4696 52554
rect 4696 52502 4740 52554
rect 4788 52502 4820 52554
rect 4820 52502 4844 52554
rect 4684 52500 4740 52502
rect 4788 52500 4844 52502
rect 4892 52500 4948 52556
rect 2044 51660 2100 51716
rect 5852 51660 5908 51716
rect 8768 51716 8824 51772
rect 8872 51770 8928 51772
rect 8976 51770 9032 51772
rect 8872 51718 8896 51770
rect 8896 51718 8928 51770
rect 8976 51718 9020 51770
rect 9020 51718 9032 51770
rect 8872 51716 8928 51718
rect 8976 51716 9032 51718
rect 9080 51716 9136 51772
rect 9184 51770 9240 51772
rect 9288 51770 9344 51772
rect 9184 51718 9196 51770
rect 9196 51718 9240 51770
rect 9288 51718 9320 51770
rect 9320 51718 9344 51770
rect 9184 51716 9240 51718
rect 9288 51716 9344 51718
rect 9392 51716 9448 51772
rect 1932 50428 1988 50484
rect 2044 50316 2100 50372
rect 1708 49980 1764 50036
rect 1708 48636 1764 48692
rect 1708 47740 1764 47796
rect 2492 51100 2548 51156
rect 4268 50932 4324 50988
rect 4372 50986 4428 50988
rect 4476 50986 4532 50988
rect 4372 50934 4396 50986
rect 4396 50934 4428 50986
rect 4476 50934 4520 50986
rect 4520 50934 4532 50986
rect 4372 50932 4428 50934
rect 4476 50932 4532 50934
rect 4580 50932 4636 50988
rect 4684 50986 4740 50988
rect 4788 50986 4844 50988
rect 4684 50934 4696 50986
rect 4696 50934 4740 50986
rect 4788 50934 4820 50986
rect 4820 50934 4844 50986
rect 4684 50932 4740 50934
rect 4788 50932 4844 50934
rect 4892 50932 4948 50988
rect 2492 49980 2548 50036
rect 2828 50316 2884 50372
rect 2268 48972 2324 49028
rect 2380 48914 2436 48916
rect 2380 48862 2382 48914
rect 2382 48862 2434 48914
rect 2434 48862 2436 48914
rect 2380 48860 2436 48862
rect 2492 48636 2548 48692
rect 2044 47346 2100 47348
rect 2044 47294 2046 47346
rect 2046 47294 2098 47346
rect 2098 47294 2100 47346
rect 2044 47292 2100 47294
rect 1820 46674 1876 46676
rect 1820 46622 1822 46674
rect 1822 46622 1874 46674
rect 1874 46622 1876 46674
rect 1820 46620 1876 46622
rect 1708 45500 1764 45556
rect 1708 44940 1764 44996
rect 1708 44380 1764 44436
rect 1820 43260 1876 43316
rect 1708 42140 1764 42196
rect 1708 39900 1764 39956
rect 2492 45500 2548 45556
rect 8768 50148 8824 50204
rect 8872 50202 8928 50204
rect 8976 50202 9032 50204
rect 8872 50150 8896 50202
rect 8896 50150 8928 50202
rect 8976 50150 9020 50202
rect 9020 50150 9032 50202
rect 8872 50148 8928 50150
rect 8976 50148 9032 50150
rect 9080 50148 9136 50204
rect 9184 50202 9240 50204
rect 9288 50202 9344 50204
rect 9184 50150 9196 50202
rect 9196 50150 9240 50202
rect 9288 50150 9320 50202
rect 9320 50150 9344 50202
rect 9184 50148 9240 50150
rect 9288 50148 9344 50150
rect 9392 50148 9448 50204
rect 8316 49644 8372 49700
rect 5852 49532 5908 49588
rect 4268 49364 4324 49420
rect 4372 49418 4428 49420
rect 4476 49418 4532 49420
rect 4372 49366 4396 49418
rect 4396 49366 4428 49418
rect 4476 49366 4520 49418
rect 4520 49366 4532 49418
rect 4372 49364 4428 49366
rect 4476 49364 4532 49366
rect 4580 49364 4636 49420
rect 4684 49418 4740 49420
rect 4788 49418 4844 49420
rect 4684 49366 4696 49418
rect 4696 49366 4740 49418
rect 4788 49366 4820 49418
rect 4820 49366 4844 49418
rect 4684 49364 4740 49366
rect 4788 49364 4844 49366
rect 4892 49364 4948 49420
rect 3164 48914 3220 48916
rect 3164 48862 3166 48914
rect 3166 48862 3218 48914
rect 3218 48862 3220 48914
rect 3164 48860 3220 48862
rect 4732 48076 4788 48132
rect 5628 48130 5684 48132
rect 5628 48078 5630 48130
rect 5630 48078 5682 48130
rect 5682 48078 5684 48130
rect 5628 48076 5684 48078
rect 5292 48018 5348 48020
rect 5292 47966 5294 48018
rect 5294 47966 5346 48018
rect 5346 47966 5348 48018
rect 5292 47964 5348 47966
rect 4268 47796 4324 47852
rect 4372 47850 4428 47852
rect 4476 47850 4532 47852
rect 4372 47798 4396 47850
rect 4396 47798 4428 47850
rect 4476 47798 4520 47850
rect 4520 47798 4532 47850
rect 4372 47796 4428 47798
rect 4476 47796 4532 47798
rect 4580 47796 4636 47852
rect 4684 47850 4740 47852
rect 4788 47850 4844 47852
rect 4684 47798 4696 47850
rect 4696 47798 4740 47850
rect 4788 47798 4820 47850
rect 4820 47798 4844 47850
rect 4684 47796 4740 47798
rect 4788 47796 4844 47798
rect 4892 47796 4948 47852
rect 4268 46228 4324 46284
rect 4372 46282 4428 46284
rect 4476 46282 4532 46284
rect 4372 46230 4396 46282
rect 4396 46230 4428 46282
rect 4476 46230 4520 46282
rect 4520 46230 4532 46282
rect 4372 46228 4428 46230
rect 4476 46228 4532 46230
rect 4580 46228 4636 46284
rect 4684 46282 4740 46284
rect 4788 46282 4844 46284
rect 4684 46230 4696 46282
rect 4696 46230 4740 46282
rect 4788 46230 4820 46282
rect 4820 46230 4844 46282
rect 4684 46228 4740 46230
rect 4788 46228 4844 46230
rect 4892 46228 4948 46284
rect 2716 45052 2772 45108
rect 3388 45106 3444 45108
rect 3388 45054 3390 45106
rect 3390 45054 3442 45106
rect 3442 45054 3444 45106
rect 3388 45052 3444 45054
rect 2492 44994 2548 44996
rect 2492 44942 2494 44994
rect 2494 44942 2546 44994
rect 2546 44942 2548 44994
rect 2492 44940 2548 44942
rect 4268 44660 4324 44716
rect 4372 44714 4428 44716
rect 4476 44714 4532 44716
rect 4372 44662 4396 44714
rect 4396 44662 4428 44714
rect 4476 44662 4520 44714
rect 4520 44662 4532 44714
rect 4372 44660 4428 44662
rect 4476 44660 4532 44662
rect 4580 44660 4636 44716
rect 4684 44714 4740 44716
rect 4788 44714 4844 44716
rect 4684 44662 4696 44714
rect 4696 44662 4740 44714
rect 4788 44662 4820 44714
rect 4820 44662 4844 44714
rect 4684 44660 4740 44662
rect 4788 44660 4844 44662
rect 4892 44660 4948 44716
rect 5740 43596 5796 43652
rect 4268 43092 4324 43148
rect 4372 43146 4428 43148
rect 4476 43146 4532 43148
rect 4372 43094 4396 43146
rect 4396 43094 4428 43146
rect 4476 43094 4520 43146
rect 4520 43094 4532 43146
rect 4372 43092 4428 43094
rect 4476 43092 4532 43094
rect 4580 43092 4636 43148
rect 4684 43146 4740 43148
rect 4788 43146 4844 43148
rect 4684 43094 4696 43146
rect 4696 43094 4740 43146
rect 4788 43094 4820 43146
rect 4820 43094 4844 43146
rect 4684 43092 4740 43094
rect 4788 43092 4844 43094
rect 4892 43092 4948 43148
rect 2492 42140 2548 42196
rect 2044 41356 2100 41412
rect 2380 41074 2436 41076
rect 2380 41022 2382 41074
rect 2382 41022 2434 41074
rect 2434 41022 2436 41074
rect 2380 41020 2436 41022
rect 2044 39394 2100 39396
rect 2044 39342 2046 39394
rect 2046 39342 2098 39394
rect 2098 39342 2100 39394
rect 2044 39340 2100 39342
rect 1820 38834 1876 38836
rect 1820 38782 1822 38834
rect 1822 38782 1874 38834
rect 1874 38782 1876 38834
rect 1820 38780 1876 38782
rect 1708 37660 1764 37716
rect 1708 36540 1764 36596
rect 1708 35420 1764 35476
rect 1708 34300 1764 34356
rect 1820 34412 1876 34468
rect 2044 35810 2100 35812
rect 2044 35758 2046 35810
rect 2046 35758 2098 35810
rect 2098 35758 2100 35810
rect 2044 35756 2100 35758
rect 2156 34860 2212 34916
rect 2044 34690 2100 34692
rect 2044 34638 2046 34690
rect 2046 34638 2098 34690
rect 2098 34638 2100 34690
rect 2044 34636 2100 34638
rect 2492 37660 2548 37716
rect 10108 49922 10164 49924
rect 10108 49870 10110 49922
rect 10110 49870 10162 49922
rect 10162 49870 10164 49922
rect 10108 49868 10164 49870
rect 11340 49922 11396 49924
rect 11340 49870 11342 49922
rect 11342 49870 11394 49922
rect 11394 49870 11396 49922
rect 11340 49868 11396 49870
rect 26768 56420 26824 56476
rect 26872 56474 26928 56476
rect 26976 56474 27032 56476
rect 26872 56422 26896 56474
rect 26896 56422 26928 56474
rect 26976 56422 27020 56474
rect 27020 56422 27032 56474
rect 26872 56420 26928 56422
rect 26976 56420 27032 56422
rect 27080 56420 27136 56476
rect 27184 56474 27240 56476
rect 27288 56474 27344 56476
rect 27184 56422 27196 56474
rect 27196 56422 27240 56474
rect 27288 56422 27320 56474
rect 27320 56422 27344 56474
rect 27184 56420 27240 56422
rect 27288 56420 27344 56422
rect 27392 56420 27448 56476
rect 35768 56420 35824 56476
rect 35872 56474 35928 56476
rect 35976 56474 36032 56476
rect 35872 56422 35896 56474
rect 35896 56422 35928 56474
rect 35976 56422 36020 56474
rect 36020 56422 36032 56474
rect 35872 56420 35928 56422
rect 35976 56420 36032 56422
rect 36080 56420 36136 56476
rect 36184 56474 36240 56476
rect 36288 56474 36344 56476
rect 36184 56422 36196 56474
rect 36196 56422 36240 56474
rect 36288 56422 36320 56474
rect 36320 56422 36344 56474
rect 36184 56420 36240 56422
rect 36288 56420 36344 56422
rect 36392 56420 36448 56476
rect 31388 56252 31444 56308
rect 32172 56306 32228 56308
rect 32172 56254 32174 56306
rect 32174 56254 32226 56306
rect 32226 56254 32228 56306
rect 32172 56252 32228 56254
rect 20076 56082 20132 56084
rect 20076 56030 20078 56082
rect 20078 56030 20130 56082
rect 20130 56030 20132 56082
rect 20076 56028 20132 56030
rect 25452 56028 25508 56084
rect 13268 55636 13324 55692
rect 13372 55690 13428 55692
rect 13476 55690 13532 55692
rect 13372 55638 13396 55690
rect 13396 55638 13428 55690
rect 13476 55638 13520 55690
rect 13520 55638 13532 55690
rect 13372 55636 13428 55638
rect 13476 55636 13532 55638
rect 13580 55636 13636 55692
rect 13684 55690 13740 55692
rect 13788 55690 13844 55692
rect 13684 55638 13696 55690
rect 13696 55638 13740 55690
rect 13788 55638 13820 55690
rect 13820 55638 13844 55690
rect 13684 55636 13740 55638
rect 13788 55636 13844 55638
rect 13892 55636 13948 55692
rect 22268 55636 22324 55692
rect 22372 55690 22428 55692
rect 22476 55690 22532 55692
rect 22372 55638 22396 55690
rect 22396 55638 22428 55690
rect 22476 55638 22520 55690
rect 22520 55638 22532 55690
rect 22372 55636 22428 55638
rect 22476 55636 22532 55638
rect 22580 55636 22636 55692
rect 22684 55690 22740 55692
rect 22788 55690 22844 55692
rect 22684 55638 22696 55690
rect 22696 55638 22740 55690
rect 22788 55638 22820 55690
rect 22820 55638 22844 55690
rect 22684 55636 22740 55638
rect 22788 55636 22844 55638
rect 22892 55636 22948 55692
rect 26124 55916 26180 55972
rect 17768 54852 17824 54908
rect 17872 54906 17928 54908
rect 17976 54906 18032 54908
rect 17872 54854 17896 54906
rect 17896 54854 17928 54906
rect 17976 54854 18020 54906
rect 18020 54854 18032 54906
rect 17872 54852 17928 54854
rect 17976 54852 18032 54854
rect 18080 54852 18136 54908
rect 18184 54906 18240 54908
rect 18288 54906 18344 54908
rect 18184 54854 18196 54906
rect 18196 54854 18240 54906
rect 18288 54854 18320 54906
rect 18320 54854 18344 54906
rect 18184 54852 18240 54854
rect 18288 54852 18344 54854
rect 18392 54852 18448 54908
rect 13268 54068 13324 54124
rect 13372 54122 13428 54124
rect 13476 54122 13532 54124
rect 13372 54070 13396 54122
rect 13396 54070 13428 54122
rect 13476 54070 13520 54122
rect 13520 54070 13532 54122
rect 13372 54068 13428 54070
rect 13476 54068 13532 54070
rect 13580 54068 13636 54124
rect 13684 54122 13740 54124
rect 13788 54122 13844 54124
rect 13684 54070 13696 54122
rect 13696 54070 13740 54122
rect 13788 54070 13820 54122
rect 13820 54070 13844 54122
rect 13684 54068 13740 54070
rect 13788 54068 13844 54070
rect 13892 54068 13948 54124
rect 22268 54068 22324 54124
rect 22372 54122 22428 54124
rect 22476 54122 22532 54124
rect 22372 54070 22396 54122
rect 22396 54070 22428 54122
rect 22476 54070 22520 54122
rect 22520 54070 22532 54122
rect 22372 54068 22428 54070
rect 22476 54068 22532 54070
rect 22580 54068 22636 54124
rect 22684 54122 22740 54124
rect 22788 54122 22844 54124
rect 22684 54070 22696 54122
rect 22696 54070 22740 54122
rect 22788 54070 22820 54122
rect 22820 54070 22844 54122
rect 22684 54068 22740 54070
rect 22788 54068 22844 54070
rect 22892 54068 22948 54124
rect 17768 53284 17824 53340
rect 17872 53338 17928 53340
rect 17976 53338 18032 53340
rect 17872 53286 17896 53338
rect 17896 53286 17928 53338
rect 17976 53286 18020 53338
rect 18020 53286 18032 53338
rect 17872 53284 17928 53286
rect 17976 53284 18032 53286
rect 18080 53284 18136 53340
rect 18184 53338 18240 53340
rect 18288 53338 18344 53340
rect 18184 53286 18196 53338
rect 18196 53286 18240 53338
rect 18288 53286 18320 53338
rect 18320 53286 18344 53338
rect 18184 53284 18240 53286
rect 18288 53284 18344 53286
rect 18392 53284 18448 53340
rect 31268 55636 31324 55692
rect 31372 55690 31428 55692
rect 31476 55690 31532 55692
rect 31372 55638 31396 55690
rect 31396 55638 31428 55690
rect 31476 55638 31520 55690
rect 31520 55638 31532 55690
rect 31372 55636 31428 55638
rect 31476 55636 31532 55638
rect 31580 55636 31636 55692
rect 31684 55690 31740 55692
rect 31788 55690 31844 55692
rect 31684 55638 31696 55690
rect 31696 55638 31740 55690
rect 31788 55638 31820 55690
rect 31820 55638 31844 55690
rect 31684 55636 31740 55638
rect 31788 55636 31844 55638
rect 31892 55636 31948 55692
rect 29260 55298 29316 55300
rect 29260 55246 29262 55298
rect 29262 55246 29314 55298
rect 29314 55246 29316 55298
rect 29260 55244 29316 55246
rect 26768 54852 26824 54908
rect 26872 54906 26928 54908
rect 26976 54906 27032 54908
rect 26872 54854 26896 54906
rect 26896 54854 26928 54906
rect 26976 54854 27020 54906
rect 27020 54854 27032 54906
rect 26872 54852 26928 54854
rect 26976 54852 27032 54854
rect 27080 54852 27136 54908
rect 27184 54906 27240 54908
rect 27288 54906 27344 54908
rect 27184 54854 27196 54906
rect 27196 54854 27240 54906
rect 27288 54854 27320 54906
rect 27320 54854 27344 54906
rect 27184 54852 27240 54854
rect 27288 54852 27344 54854
rect 27392 54852 27448 54908
rect 28476 53900 28532 53956
rect 31268 54068 31324 54124
rect 31372 54122 31428 54124
rect 31476 54122 31532 54124
rect 31372 54070 31396 54122
rect 31396 54070 31428 54122
rect 31476 54070 31520 54122
rect 31520 54070 31532 54122
rect 31372 54068 31428 54070
rect 31476 54068 31532 54070
rect 31580 54068 31636 54124
rect 31684 54122 31740 54124
rect 31788 54122 31844 54124
rect 31684 54070 31696 54122
rect 31696 54070 31740 54122
rect 31788 54070 31820 54122
rect 31820 54070 31844 54122
rect 31684 54068 31740 54070
rect 31788 54068 31844 54070
rect 31892 54068 31948 54124
rect 26768 53284 26824 53340
rect 26872 53338 26928 53340
rect 26976 53338 27032 53340
rect 26872 53286 26896 53338
rect 26896 53286 26928 53338
rect 26976 53286 27020 53338
rect 27020 53286 27032 53338
rect 26872 53284 26928 53286
rect 26976 53284 27032 53286
rect 27080 53284 27136 53340
rect 27184 53338 27240 53340
rect 27288 53338 27344 53340
rect 27184 53286 27196 53338
rect 27196 53286 27240 53338
rect 27288 53286 27320 53338
rect 27320 53286 27344 53338
rect 27184 53284 27240 53286
rect 27288 53284 27344 53286
rect 27392 53284 27448 53340
rect 25788 53004 25844 53060
rect 25116 52780 25172 52836
rect 13268 52500 13324 52556
rect 13372 52554 13428 52556
rect 13476 52554 13532 52556
rect 13372 52502 13396 52554
rect 13396 52502 13428 52554
rect 13476 52502 13520 52554
rect 13520 52502 13532 52554
rect 13372 52500 13428 52502
rect 13476 52500 13532 52502
rect 13580 52500 13636 52556
rect 13684 52554 13740 52556
rect 13788 52554 13844 52556
rect 13684 52502 13696 52554
rect 13696 52502 13740 52554
rect 13788 52502 13820 52554
rect 13820 52502 13844 52554
rect 13684 52500 13740 52502
rect 13788 52500 13844 52502
rect 13892 52500 13948 52556
rect 22268 52500 22324 52556
rect 22372 52554 22428 52556
rect 22476 52554 22532 52556
rect 22372 52502 22396 52554
rect 22396 52502 22428 52554
rect 22476 52502 22520 52554
rect 22520 52502 22532 52554
rect 22372 52500 22428 52502
rect 22476 52500 22532 52502
rect 22580 52500 22636 52556
rect 22684 52554 22740 52556
rect 22788 52554 22844 52556
rect 22684 52502 22696 52554
rect 22696 52502 22740 52554
rect 22788 52502 22820 52554
rect 22820 52502 22844 52554
rect 22684 52500 22740 52502
rect 22788 52500 22844 52502
rect 22892 52500 22948 52556
rect 22988 52274 23044 52276
rect 22988 52222 22990 52274
rect 22990 52222 23042 52274
rect 23042 52222 23044 52274
rect 22988 52220 23044 52222
rect 26236 51884 26292 51940
rect 17768 51716 17824 51772
rect 17872 51770 17928 51772
rect 17976 51770 18032 51772
rect 17872 51718 17896 51770
rect 17896 51718 17928 51770
rect 17976 51718 18020 51770
rect 18020 51718 18032 51770
rect 17872 51716 17928 51718
rect 17976 51716 18032 51718
rect 18080 51716 18136 51772
rect 18184 51770 18240 51772
rect 18288 51770 18344 51772
rect 18184 51718 18196 51770
rect 18196 51718 18240 51770
rect 18288 51718 18320 51770
rect 18320 51718 18344 51770
rect 18184 51716 18240 51718
rect 18288 51716 18344 51718
rect 18392 51716 18448 51772
rect 13268 50932 13324 50988
rect 13372 50986 13428 50988
rect 13476 50986 13532 50988
rect 13372 50934 13396 50986
rect 13396 50934 13428 50986
rect 13476 50934 13520 50986
rect 13520 50934 13532 50986
rect 13372 50932 13428 50934
rect 13476 50932 13532 50934
rect 13580 50932 13636 50988
rect 13684 50986 13740 50988
rect 13788 50986 13844 50988
rect 13684 50934 13696 50986
rect 13696 50934 13740 50986
rect 13788 50934 13820 50986
rect 13820 50934 13844 50986
rect 13684 50932 13740 50934
rect 13788 50932 13844 50934
rect 13892 50932 13948 50988
rect 22268 50932 22324 50988
rect 22372 50986 22428 50988
rect 22476 50986 22532 50988
rect 22372 50934 22396 50986
rect 22396 50934 22428 50986
rect 22476 50934 22520 50986
rect 22520 50934 22532 50986
rect 22372 50932 22428 50934
rect 22476 50932 22532 50934
rect 22580 50932 22636 50988
rect 22684 50986 22740 50988
rect 22788 50986 22844 50988
rect 22684 50934 22696 50986
rect 22696 50934 22740 50986
rect 22788 50934 22820 50986
rect 22820 50934 22844 50986
rect 22684 50932 22740 50934
rect 22788 50932 22844 50934
rect 22892 50932 22948 50988
rect 16156 50482 16212 50484
rect 16156 50430 16158 50482
rect 16158 50430 16210 50482
rect 16210 50430 16212 50482
rect 16156 50428 16212 50430
rect 17276 50428 17332 50484
rect 19628 50482 19684 50484
rect 19628 50430 19630 50482
rect 19630 50430 19682 50482
rect 19682 50430 19684 50482
rect 19628 50428 19684 50430
rect 20524 50428 20580 50484
rect 17768 50148 17824 50204
rect 17872 50202 17928 50204
rect 17976 50202 18032 50204
rect 17872 50150 17896 50202
rect 17896 50150 17928 50202
rect 17976 50150 18020 50202
rect 18020 50150 18032 50202
rect 17872 50148 17928 50150
rect 17976 50148 18032 50150
rect 18080 50148 18136 50204
rect 18184 50202 18240 50204
rect 18288 50202 18344 50204
rect 18184 50150 18196 50202
rect 18196 50150 18240 50202
rect 18288 50150 18320 50202
rect 18320 50150 18344 50202
rect 18184 50148 18240 50150
rect 18288 50148 18344 50150
rect 18392 50148 18448 50204
rect 14476 49922 14532 49924
rect 14476 49870 14478 49922
rect 14478 49870 14530 49922
rect 14530 49870 14532 49922
rect 14476 49868 14532 49870
rect 13268 49364 13324 49420
rect 13372 49418 13428 49420
rect 13476 49418 13532 49420
rect 13372 49366 13396 49418
rect 13396 49366 13428 49418
rect 13476 49366 13520 49418
rect 13520 49366 13532 49418
rect 13372 49364 13428 49366
rect 13476 49364 13532 49366
rect 13580 49364 13636 49420
rect 13684 49418 13740 49420
rect 13788 49418 13844 49420
rect 13684 49366 13696 49418
rect 13696 49366 13740 49418
rect 13788 49366 13820 49418
rect 13820 49366 13844 49418
rect 13684 49364 13740 49366
rect 13788 49364 13844 49366
rect 13892 49364 13948 49420
rect 9324 49026 9380 49028
rect 9324 48974 9326 49026
rect 9326 48974 9378 49026
rect 9378 48974 9380 49026
rect 9324 48972 9380 48974
rect 8768 48580 8824 48636
rect 8872 48634 8928 48636
rect 8976 48634 9032 48636
rect 8872 48582 8896 48634
rect 8896 48582 8928 48634
rect 8976 48582 9020 48634
rect 9020 48582 9032 48634
rect 8872 48580 8928 48582
rect 8976 48580 9032 48582
rect 9080 48580 9136 48636
rect 9184 48634 9240 48636
rect 9288 48634 9344 48636
rect 9184 48582 9196 48634
rect 9196 48582 9240 48634
rect 9288 48582 9320 48634
rect 9320 48582 9344 48634
rect 9184 48580 9240 48582
rect 9288 48580 9344 48582
rect 9392 48580 9448 48636
rect 9660 47964 9716 48020
rect 10108 47404 10164 47460
rect 8540 46844 8596 46900
rect 8764 47180 8820 47236
rect 8768 47012 8824 47068
rect 8872 47066 8928 47068
rect 8976 47066 9032 47068
rect 8872 47014 8896 47066
rect 8896 47014 8928 47066
rect 8976 47014 9020 47066
rect 9020 47014 9032 47066
rect 8872 47012 8928 47014
rect 8976 47012 9032 47014
rect 9080 47012 9136 47068
rect 9184 47066 9240 47068
rect 9288 47066 9344 47068
rect 9184 47014 9196 47066
rect 9196 47014 9240 47066
rect 9288 47014 9320 47066
rect 9320 47014 9344 47066
rect 9184 47012 9240 47014
rect 9288 47012 9344 47014
rect 9392 47012 9448 47068
rect 8988 46620 9044 46676
rect 9996 46674 10052 46676
rect 9996 46622 9998 46674
rect 9998 46622 10050 46674
rect 10050 46622 10052 46674
rect 9996 46620 10052 46622
rect 8768 45444 8824 45500
rect 8872 45498 8928 45500
rect 8976 45498 9032 45500
rect 8872 45446 8896 45498
rect 8896 45446 8928 45498
rect 8976 45446 9020 45498
rect 9020 45446 9032 45498
rect 8872 45444 8928 45446
rect 8976 45444 9032 45446
rect 9080 45444 9136 45500
rect 9184 45498 9240 45500
rect 9288 45498 9344 45500
rect 9184 45446 9196 45498
rect 9196 45446 9240 45498
rect 9288 45446 9320 45498
rect 9320 45446 9344 45498
rect 9184 45444 9240 45446
rect 9288 45444 9344 45446
rect 9392 45444 9448 45500
rect 5964 45164 6020 45220
rect 6524 44492 6580 44548
rect 10444 47458 10500 47460
rect 10444 47406 10446 47458
rect 10446 47406 10498 47458
rect 10498 47406 10500 47458
rect 10444 47404 10500 47406
rect 9772 44322 9828 44324
rect 9772 44270 9774 44322
rect 9774 44270 9826 44322
rect 9826 44270 9828 44322
rect 9772 44268 9828 44270
rect 10220 47346 10276 47348
rect 10220 47294 10222 47346
rect 10222 47294 10274 47346
rect 10274 47294 10276 47346
rect 10220 47292 10276 47294
rect 11340 47346 11396 47348
rect 11340 47294 11342 47346
rect 11342 47294 11394 47346
rect 11394 47294 11396 47346
rect 11340 47292 11396 47294
rect 10780 47234 10836 47236
rect 10780 47182 10782 47234
rect 10782 47182 10834 47234
rect 10834 47182 10836 47234
rect 10780 47180 10836 47182
rect 7196 44156 7252 44212
rect 6300 43596 6356 43652
rect 8988 44098 9044 44100
rect 8988 44046 8990 44098
rect 8990 44046 9042 44098
rect 9042 44046 9044 44098
rect 8988 44044 9044 44046
rect 9772 44044 9828 44100
rect 8768 43876 8824 43932
rect 8872 43930 8928 43932
rect 8976 43930 9032 43932
rect 8872 43878 8896 43930
rect 8896 43878 8928 43930
rect 8976 43878 9020 43930
rect 9020 43878 9032 43930
rect 8872 43876 8928 43878
rect 8976 43876 9032 43878
rect 9080 43876 9136 43932
rect 9184 43930 9240 43932
rect 9288 43930 9344 43932
rect 9184 43878 9196 43930
rect 9196 43878 9240 43930
rect 9288 43878 9320 43930
rect 9320 43878 9344 43930
rect 9184 43876 9240 43878
rect 9288 43876 9344 43878
rect 9392 43876 9448 43932
rect 8316 43708 8372 43764
rect 9436 43708 9492 43764
rect 5964 43314 6020 43316
rect 5964 43262 5966 43314
rect 5966 43262 6018 43314
rect 6018 43262 6020 43314
rect 5964 43260 6020 43262
rect 6188 42140 6244 42196
rect 4268 41524 4324 41580
rect 4372 41578 4428 41580
rect 4476 41578 4532 41580
rect 4372 41526 4396 41578
rect 4396 41526 4428 41578
rect 4476 41526 4520 41578
rect 4520 41526 4532 41578
rect 4372 41524 4428 41526
rect 4476 41524 4532 41526
rect 4580 41524 4636 41580
rect 4684 41578 4740 41580
rect 4788 41578 4844 41580
rect 4684 41526 4696 41578
rect 4696 41526 4740 41578
rect 4788 41526 4820 41578
rect 4820 41526 4844 41578
rect 4684 41524 4740 41526
rect 4788 41524 4844 41526
rect 4892 41524 4948 41580
rect 2380 35756 2436 35812
rect 2380 34412 2436 34468
rect 1708 33234 1764 33236
rect 1708 33182 1710 33234
rect 1710 33182 1762 33234
rect 1762 33182 1764 33234
rect 1708 33180 1764 33182
rect 1708 32060 1764 32116
rect 2492 33234 2548 33236
rect 2492 33182 2494 33234
rect 2494 33182 2546 33234
rect 2546 33182 2548 33234
rect 2492 33180 2548 33182
rect 1820 31948 1876 32004
rect 1708 31500 1764 31556
rect 1708 30940 1764 30996
rect 1820 31164 1876 31220
rect 2492 32060 2548 32116
rect 5964 41356 6020 41412
rect 4732 40626 4788 40628
rect 4732 40574 4734 40626
rect 4734 40574 4786 40626
rect 4786 40574 4788 40626
rect 4732 40572 4788 40574
rect 5852 40572 5908 40628
rect 3164 39900 3220 39956
rect 4268 39956 4324 40012
rect 4372 40010 4428 40012
rect 4476 40010 4532 40012
rect 4372 39958 4396 40010
rect 4396 39958 4428 40010
rect 4476 39958 4520 40010
rect 4520 39958 4532 40010
rect 4372 39956 4428 39958
rect 4476 39956 4532 39958
rect 4580 39956 4636 40012
rect 4684 40010 4740 40012
rect 4788 40010 4844 40012
rect 4684 39958 4696 40010
rect 4696 39958 4740 40010
rect 4788 39958 4820 40010
rect 4820 39958 4844 40010
rect 4684 39956 4740 39958
rect 4788 39956 4844 39958
rect 4892 39956 4948 40012
rect 4268 38388 4324 38444
rect 4372 38442 4428 38444
rect 4476 38442 4532 38444
rect 4372 38390 4396 38442
rect 4396 38390 4428 38442
rect 4476 38390 4520 38442
rect 4520 38390 4532 38442
rect 4372 38388 4428 38390
rect 4476 38388 4532 38390
rect 4580 38388 4636 38444
rect 4684 38442 4740 38444
rect 4788 38442 4844 38444
rect 4684 38390 4696 38442
rect 4696 38390 4740 38442
rect 4788 38390 4820 38442
rect 4820 38390 4844 38442
rect 4684 38388 4740 38390
rect 4788 38388 4844 38390
rect 4892 38388 4948 38444
rect 5292 37772 5348 37828
rect 4268 36820 4324 36876
rect 4372 36874 4428 36876
rect 4476 36874 4532 36876
rect 4372 36822 4396 36874
rect 4396 36822 4428 36874
rect 4476 36822 4520 36874
rect 4520 36822 4532 36874
rect 4372 36820 4428 36822
rect 4476 36820 4532 36822
rect 4580 36820 4636 36876
rect 4684 36874 4740 36876
rect 4788 36874 4844 36876
rect 4684 36822 4696 36874
rect 4696 36822 4740 36874
rect 4788 36822 4820 36874
rect 4820 36822 4844 36874
rect 4684 36820 4740 36822
rect 4788 36820 4844 36822
rect 4892 36820 4948 36876
rect 3276 36594 3332 36596
rect 3276 36542 3278 36594
rect 3278 36542 3330 36594
rect 3330 36542 3332 36594
rect 3276 36540 3332 36542
rect 5852 37378 5908 37380
rect 5852 37326 5854 37378
rect 5854 37326 5906 37378
rect 5906 37326 5908 37378
rect 5852 37324 5908 37326
rect 5068 36204 5124 36260
rect 5628 36204 5684 36260
rect 10332 46844 10388 46900
rect 12460 48802 12516 48804
rect 12460 48750 12462 48802
rect 12462 48750 12514 48802
rect 12514 48750 12516 48802
rect 12460 48748 12516 48750
rect 13580 48354 13636 48356
rect 13580 48302 13582 48354
rect 13582 48302 13634 48354
rect 13634 48302 13636 48354
rect 13580 48300 13636 48302
rect 14028 48242 14084 48244
rect 14028 48190 14030 48242
rect 14030 48190 14082 48242
rect 14082 48190 14084 48242
rect 14028 48188 14084 48190
rect 13268 47796 13324 47852
rect 13372 47850 13428 47852
rect 13476 47850 13532 47852
rect 13372 47798 13396 47850
rect 13396 47798 13428 47850
rect 13476 47798 13520 47850
rect 13520 47798 13532 47850
rect 13372 47796 13428 47798
rect 13476 47796 13532 47798
rect 13580 47796 13636 47852
rect 13684 47850 13740 47852
rect 13788 47850 13844 47852
rect 13684 47798 13696 47850
rect 13696 47798 13740 47850
rect 13788 47798 13820 47850
rect 13820 47798 13844 47850
rect 13684 47796 13740 47798
rect 13788 47796 13844 47798
rect 13892 47796 13948 47852
rect 14924 48748 14980 48804
rect 15036 48300 15092 48356
rect 11788 47234 11844 47236
rect 11788 47182 11790 47234
rect 11790 47182 11842 47234
rect 11842 47182 11844 47234
rect 11788 47180 11844 47182
rect 13132 47180 13188 47236
rect 11564 44322 11620 44324
rect 11564 44270 11566 44322
rect 11566 44270 11618 44322
rect 11618 44270 11620 44322
rect 11564 44268 11620 44270
rect 8768 42308 8824 42364
rect 8872 42362 8928 42364
rect 8976 42362 9032 42364
rect 8872 42310 8896 42362
rect 8896 42310 8928 42362
rect 8976 42310 9020 42362
rect 9020 42310 9032 42362
rect 8872 42308 8928 42310
rect 8976 42308 9032 42310
rect 9080 42308 9136 42364
rect 9184 42362 9240 42364
rect 9288 42362 9344 42364
rect 9184 42310 9196 42362
rect 9196 42310 9240 42362
rect 9288 42310 9320 42362
rect 9320 42310 9344 42362
rect 9184 42308 9240 42310
rect 9288 42308 9344 42310
rect 9392 42308 9448 42364
rect 6748 42140 6804 42196
rect 6300 41746 6356 41748
rect 6300 41694 6302 41746
rect 6302 41694 6354 41746
rect 6354 41694 6356 41746
rect 6300 41692 6356 41694
rect 9324 40962 9380 40964
rect 9324 40910 9326 40962
rect 9326 40910 9378 40962
rect 9378 40910 9380 40962
rect 9324 40908 9380 40910
rect 8768 40740 8824 40796
rect 8872 40794 8928 40796
rect 8976 40794 9032 40796
rect 8872 40742 8896 40794
rect 8896 40742 8928 40794
rect 8976 40742 9020 40794
rect 9020 40742 9032 40794
rect 8872 40740 8928 40742
rect 8976 40740 9032 40742
rect 9080 40740 9136 40796
rect 9184 40794 9240 40796
rect 9288 40794 9344 40796
rect 9184 40742 9196 40794
rect 9196 40742 9240 40794
rect 9288 40742 9320 40794
rect 9320 40742 9344 40794
rect 9184 40740 9240 40742
rect 9288 40740 9344 40742
rect 9392 40740 9448 40796
rect 6636 40572 6692 40628
rect 8316 40626 8372 40628
rect 8316 40574 8318 40626
rect 8318 40574 8370 40626
rect 8370 40574 8372 40626
rect 8316 40572 8372 40574
rect 9660 40908 9716 40964
rect 13268 46228 13324 46284
rect 13372 46282 13428 46284
rect 13476 46282 13532 46284
rect 13372 46230 13396 46282
rect 13396 46230 13428 46282
rect 13476 46230 13520 46282
rect 13520 46230 13532 46282
rect 13372 46228 13428 46230
rect 13476 46228 13532 46230
rect 13580 46228 13636 46284
rect 13684 46282 13740 46284
rect 13788 46282 13844 46284
rect 13684 46230 13696 46282
rect 13696 46230 13740 46282
rect 13788 46230 13820 46282
rect 13820 46230 13844 46282
rect 13684 46228 13740 46230
rect 13788 46228 13844 46230
rect 13892 46228 13948 46284
rect 13244 45948 13300 46004
rect 15484 48018 15540 48020
rect 15484 47966 15486 48018
rect 15486 47966 15538 48018
rect 15538 47966 15540 48018
rect 15484 47964 15540 47966
rect 13268 44660 13324 44716
rect 13372 44714 13428 44716
rect 13476 44714 13532 44716
rect 13372 44662 13396 44714
rect 13396 44662 13428 44714
rect 13476 44662 13520 44714
rect 13520 44662 13532 44714
rect 13372 44660 13428 44662
rect 13476 44660 13532 44662
rect 13580 44660 13636 44716
rect 13684 44714 13740 44716
rect 13788 44714 13844 44716
rect 13684 44662 13696 44714
rect 13696 44662 13740 44714
rect 13788 44662 13820 44714
rect 13820 44662 13844 44714
rect 13684 44660 13740 44662
rect 13788 44660 13844 44662
rect 13892 44660 13948 44716
rect 12348 43650 12404 43652
rect 12348 43598 12350 43650
rect 12350 43598 12402 43650
rect 12402 43598 12404 43650
rect 12348 43596 12404 43598
rect 13132 44268 13188 44324
rect 14924 45106 14980 45108
rect 14924 45054 14926 45106
rect 14926 45054 14978 45106
rect 14978 45054 14980 45106
rect 14924 45052 14980 45054
rect 15484 45218 15540 45220
rect 15484 45166 15486 45218
rect 15486 45166 15538 45218
rect 15538 45166 15540 45218
rect 15484 45164 15540 45166
rect 14028 44210 14084 44212
rect 14028 44158 14030 44210
rect 14030 44158 14082 44210
rect 14082 44158 14084 44210
rect 14028 44156 14084 44158
rect 12684 42588 12740 42644
rect 10332 42476 10388 42532
rect 9100 39564 9156 39620
rect 8768 39172 8824 39228
rect 8872 39226 8928 39228
rect 8976 39226 9032 39228
rect 8872 39174 8896 39226
rect 8896 39174 8928 39226
rect 8976 39174 9020 39226
rect 9020 39174 9032 39226
rect 8872 39172 8928 39174
rect 8976 39172 9032 39174
rect 9080 39172 9136 39228
rect 9184 39226 9240 39228
rect 9288 39226 9344 39228
rect 9184 39174 9196 39226
rect 9196 39174 9240 39226
rect 9288 39174 9320 39226
rect 9320 39174 9344 39226
rect 9184 39172 9240 39174
rect 9288 39172 9344 39174
rect 9392 39172 9448 39228
rect 8768 37604 8824 37660
rect 8872 37658 8928 37660
rect 8976 37658 9032 37660
rect 8872 37606 8896 37658
rect 8896 37606 8928 37658
rect 8976 37606 9020 37658
rect 9020 37606 9032 37658
rect 8872 37604 8928 37606
rect 8976 37604 9032 37606
rect 9080 37604 9136 37660
rect 9184 37658 9240 37660
rect 9288 37658 9344 37660
rect 9184 37606 9196 37658
rect 9196 37606 9240 37658
rect 9288 37606 9320 37658
rect 9320 37606 9344 37658
rect 9184 37604 9240 37606
rect 9288 37604 9344 37606
rect 9392 37604 9448 37660
rect 7308 37436 7364 37492
rect 6076 36988 6132 37044
rect 5964 36204 6020 36260
rect 6300 36258 6356 36260
rect 6300 36206 6302 36258
rect 6302 36206 6354 36258
rect 6354 36206 6356 36258
rect 6300 36204 6356 36206
rect 6188 35698 6244 35700
rect 6188 35646 6190 35698
rect 6190 35646 6242 35698
rect 6242 35646 6244 35698
rect 6188 35644 6244 35646
rect 4268 35252 4324 35308
rect 4372 35306 4428 35308
rect 4476 35306 4532 35308
rect 4372 35254 4396 35306
rect 4396 35254 4428 35306
rect 4476 35254 4520 35306
rect 4520 35254 4532 35306
rect 4372 35252 4428 35254
rect 4476 35252 4532 35254
rect 4580 35252 4636 35308
rect 4684 35306 4740 35308
rect 4788 35306 4844 35308
rect 4684 35254 4696 35306
rect 4696 35254 4740 35306
rect 4788 35254 4820 35306
rect 4820 35254 4844 35306
rect 4684 35252 4740 35254
rect 4788 35252 4844 35254
rect 4892 35252 4948 35308
rect 6076 34914 6132 34916
rect 6076 34862 6078 34914
rect 6078 34862 6130 34914
rect 6130 34862 6132 34914
rect 6076 34860 6132 34862
rect 1708 29820 1764 29876
rect 2380 31164 2436 31220
rect 2604 31724 2660 31780
rect 2716 34636 2772 34692
rect 2604 30156 2660 30212
rect 2492 29820 2548 29876
rect 1708 28700 1764 28756
rect 2044 28588 2100 28644
rect 2380 29372 2436 29428
rect 2940 34300 2996 34356
rect 4732 34188 4788 34244
rect 5628 34188 5684 34244
rect 5292 34018 5348 34020
rect 5292 33966 5294 34018
rect 5294 33966 5346 34018
rect 5346 33966 5348 34018
rect 5292 33964 5348 33966
rect 4268 33684 4324 33740
rect 4372 33738 4428 33740
rect 4476 33738 4532 33740
rect 4372 33686 4396 33738
rect 4396 33686 4428 33738
rect 4476 33686 4520 33738
rect 4520 33686 4532 33738
rect 4372 33684 4428 33686
rect 4476 33684 4532 33686
rect 4580 33684 4636 33740
rect 4684 33738 4740 33740
rect 4788 33738 4844 33740
rect 4684 33686 4696 33738
rect 4696 33686 4740 33738
rect 4788 33686 4820 33738
rect 4820 33686 4844 33738
rect 4684 33684 4740 33686
rect 4788 33684 4844 33686
rect 4892 33684 4948 33740
rect 5628 32508 5684 32564
rect 4268 32116 4324 32172
rect 4372 32170 4428 32172
rect 4476 32170 4532 32172
rect 4372 32118 4396 32170
rect 4396 32118 4428 32170
rect 4476 32118 4520 32170
rect 4520 32118 4532 32170
rect 4372 32116 4428 32118
rect 4476 32116 4532 32118
rect 4580 32116 4636 32172
rect 4684 32170 4740 32172
rect 4788 32170 4844 32172
rect 4684 32118 4696 32170
rect 4696 32118 4740 32170
rect 4788 32118 4820 32170
rect 4820 32118 4844 32170
rect 4684 32116 4740 32118
rect 4788 32116 4844 32118
rect 4892 32116 4948 32172
rect 6748 36876 6804 36932
rect 8652 37378 8708 37380
rect 8652 37326 8654 37378
rect 8654 37326 8706 37378
rect 8706 37326 8708 37378
rect 8652 37324 8708 37326
rect 9660 37378 9716 37380
rect 9660 37326 9662 37378
rect 9662 37326 9714 37378
rect 9714 37326 9716 37378
rect 9660 37324 9716 37326
rect 9996 37042 10052 37044
rect 9996 36990 9998 37042
rect 9998 36990 10050 37042
rect 10050 36990 10052 37042
rect 9996 36988 10052 36990
rect 10108 36876 10164 36932
rect 6636 36204 6692 36260
rect 8428 36258 8484 36260
rect 8428 36206 8430 36258
rect 8430 36206 8482 36258
rect 8482 36206 8484 36258
rect 8428 36204 8484 36206
rect 8768 36036 8824 36092
rect 8872 36090 8928 36092
rect 8976 36090 9032 36092
rect 8872 36038 8896 36090
rect 8896 36038 8928 36090
rect 8976 36038 9020 36090
rect 9020 36038 9032 36090
rect 8872 36036 8928 36038
rect 8976 36036 9032 36038
rect 9080 36036 9136 36092
rect 9184 36090 9240 36092
rect 9288 36090 9344 36092
rect 9184 36038 9196 36090
rect 9196 36038 9240 36090
rect 9288 36038 9320 36090
rect 9320 36038 9344 36090
rect 9184 36036 9240 36038
rect 9288 36036 9344 36038
rect 9392 36036 9448 36092
rect 8768 34468 8824 34524
rect 8872 34522 8928 34524
rect 8976 34522 9032 34524
rect 8872 34470 8896 34522
rect 8896 34470 8928 34522
rect 8976 34470 9020 34522
rect 9020 34470 9032 34522
rect 8872 34468 8928 34470
rect 8976 34468 9032 34470
rect 9080 34468 9136 34524
rect 9184 34522 9240 34524
rect 9288 34522 9344 34524
rect 9184 34470 9196 34522
rect 9196 34470 9240 34522
rect 9288 34470 9320 34522
rect 9320 34470 9344 34522
rect 9184 34468 9240 34470
rect 9288 34468 9344 34470
rect 9392 34468 9448 34524
rect 8652 33628 8708 33684
rect 8540 32674 8596 32676
rect 8540 32622 8542 32674
rect 8542 32622 8594 32674
rect 8594 32622 8596 32674
rect 8540 32620 8596 32622
rect 3276 31836 3332 31892
rect 2940 31554 2996 31556
rect 2940 31502 2942 31554
rect 2942 31502 2994 31554
rect 2994 31502 2996 31554
rect 2940 31500 2996 31502
rect 6076 31778 6132 31780
rect 6076 31726 6078 31778
rect 6078 31726 6130 31778
rect 6130 31726 6132 31778
rect 6076 31724 6132 31726
rect 3276 30828 3332 30884
rect 4268 30548 4324 30604
rect 4372 30602 4428 30604
rect 4476 30602 4532 30604
rect 4372 30550 4396 30602
rect 4396 30550 4428 30602
rect 4476 30550 4520 30602
rect 4520 30550 4532 30602
rect 4372 30548 4428 30550
rect 4476 30548 4532 30550
rect 4580 30548 4636 30604
rect 4684 30602 4740 30604
rect 4788 30602 4844 30604
rect 4684 30550 4696 30602
rect 4696 30550 4740 30602
rect 4788 30550 4820 30602
rect 4820 30550 4844 30602
rect 4684 30548 4740 30550
rect 4788 30548 4844 30550
rect 4892 30548 4948 30604
rect 4268 28980 4324 29036
rect 4372 29034 4428 29036
rect 4476 29034 4532 29036
rect 4372 28982 4396 29034
rect 4396 28982 4428 29034
rect 4476 28982 4520 29034
rect 4520 28982 4532 29034
rect 4372 28980 4428 28982
rect 4476 28980 4532 28982
rect 4580 28980 4636 29036
rect 4684 29034 4740 29036
rect 4788 29034 4844 29036
rect 4684 28982 4696 29034
rect 4696 28982 4740 29034
rect 4788 28982 4820 29034
rect 4820 28982 4844 29034
rect 4684 28980 4740 28982
rect 4788 28980 4844 28982
rect 4892 28980 4948 29036
rect 2492 28754 2548 28756
rect 2492 28702 2494 28754
rect 2494 28702 2546 28754
rect 2546 28702 2548 28754
rect 2492 28700 2548 28702
rect 5292 29596 5348 29652
rect 6076 29260 6132 29316
rect 5068 28082 5124 28084
rect 5068 28030 5070 28082
rect 5070 28030 5122 28082
rect 5122 28030 5124 28082
rect 5068 28028 5124 28030
rect 1708 27580 1764 27636
rect 4268 27412 4324 27468
rect 4372 27466 4428 27468
rect 4476 27466 4532 27468
rect 4372 27414 4396 27466
rect 4396 27414 4428 27466
rect 4476 27414 4520 27466
rect 4520 27414 4532 27466
rect 4372 27412 4428 27414
rect 4476 27412 4532 27414
rect 4580 27412 4636 27468
rect 4684 27466 4740 27468
rect 4788 27466 4844 27468
rect 4684 27414 4696 27466
rect 4696 27414 4740 27466
rect 4788 27414 4820 27466
rect 4820 27414 4844 27466
rect 4684 27412 4740 27414
rect 4788 27412 4844 27414
rect 4892 27412 4948 27468
rect 7644 28588 7700 28644
rect 5628 27244 5684 27300
rect 1708 27074 1764 27076
rect 1708 27022 1710 27074
rect 1710 27022 1762 27074
rect 1762 27022 1764 27074
rect 1708 27020 1764 27022
rect 2492 27020 2548 27076
rect 1708 25394 1764 25396
rect 1708 25342 1710 25394
rect 1710 25342 1762 25394
rect 1762 25342 1764 25394
rect 1708 25340 1764 25342
rect 2044 25676 2100 25732
rect 2156 25452 2212 25508
rect 6748 28028 6804 28084
rect 2604 26460 2660 26516
rect 4268 25844 4324 25900
rect 4372 25898 4428 25900
rect 4476 25898 4532 25900
rect 4372 25846 4396 25898
rect 4396 25846 4428 25898
rect 4476 25846 4520 25898
rect 4520 25846 4532 25898
rect 4372 25844 4428 25846
rect 4476 25844 4532 25846
rect 4580 25844 4636 25900
rect 4684 25898 4740 25900
rect 4788 25898 4844 25900
rect 4684 25846 4696 25898
rect 4696 25846 4740 25898
rect 4788 25846 4820 25898
rect 4820 25846 4844 25898
rect 4684 25844 4740 25846
rect 4788 25844 4844 25846
rect 4892 25844 4948 25900
rect 2492 25394 2548 25396
rect 2492 25342 2494 25394
rect 2494 25342 2546 25394
rect 2546 25342 2548 25394
rect 2492 25340 2548 25342
rect 5852 25564 5908 25620
rect 6076 25506 6132 25508
rect 6076 25454 6078 25506
rect 6078 25454 6130 25506
rect 6130 25454 6132 25506
rect 6076 25452 6132 25454
rect 5292 24946 5348 24948
rect 5292 24894 5294 24946
rect 5294 24894 5346 24946
rect 5346 24894 5348 24946
rect 5292 24892 5348 24894
rect 4732 24780 4788 24836
rect 5068 24780 5124 24836
rect 1708 24220 1764 24276
rect 3612 24220 3668 24276
rect 4268 24276 4324 24332
rect 4372 24330 4428 24332
rect 4476 24330 4532 24332
rect 4372 24278 4396 24330
rect 4396 24278 4428 24330
rect 4476 24278 4520 24330
rect 4520 24278 4532 24330
rect 4372 24276 4428 24278
rect 4476 24276 4532 24278
rect 4580 24276 4636 24332
rect 4684 24330 4740 24332
rect 4788 24330 4844 24332
rect 4684 24278 4696 24330
rect 4696 24278 4740 24330
rect 4788 24278 4820 24330
rect 4820 24278 4844 24330
rect 4684 24276 4740 24278
rect 4788 24276 4844 24278
rect 4892 24276 4948 24332
rect 2044 23324 2100 23380
rect 2380 23436 2436 23492
rect 2156 23100 2212 23156
rect 1708 21980 1764 22036
rect 1932 21532 1988 21588
rect 1708 21420 1764 21476
rect 1708 20860 1764 20916
rect 2044 20748 2100 20804
rect 1708 19740 1764 19796
rect 1708 19292 1764 19348
rect 1708 17554 1764 17556
rect 1708 17502 1710 17554
rect 1710 17502 1762 17554
rect 1762 17502 1764 17554
rect 1708 17500 1764 17502
rect 2044 19010 2100 19012
rect 2044 18958 2046 19010
rect 2046 18958 2098 19010
rect 2098 18958 2100 19010
rect 2044 18956 2100 18958
rect 2492 21474 2548 21476
rect 2492 21422 2494 21474
rect 2494 21422 2546 21474
rect 2546 21422 2548 21474
rect 2492 21420 2548 21422
rect 5740 24780 5796 24836
rect 9548 33292 9604 33348
rect 10108 33404 10164 33460
rect 8768 32900 8824 32956
rect 8872 32954 8928 32956
rect 8976 32954 9032 32956
rect 8872 32902 8896 32954
rect 8896 32902 8928 32954
rect 8976 32902 9020 32954
rect 9020 32902 9032 32954
rect 8872 32900 8928 32902
rect 8976 32900 9032 32902
rect 9080 32900 9136 32956
rect 9184 32954 9240 32956
rect 9288 32954 9344 32956
rect 9184 32902 9196 32954
rect 9196 32902 9240 32954
rect 9288 32902 9320 32954
rect 9320 32902 9344 32954
rect 9184 32900 9240 32902
rect 9288 32900 9344 32902
rect 9392 32900 9448 32956
rect 9100 32562 9156 32564
rect 9100 32510 9102 32562
rect 9102 32510 9154 32562
rect 9154 32510 9156 32562
rect 9100 32508 9156 32510
rect 9996 32562 10052 32564
rect 9996 32510 9998 32562
rect 9998 32510 10050 32562
rect 10050 32510 10052 32562
rect 9996 32508 10052 32510
rect 9212 31890 9268 31892
rect 9212 31838 9214 31890
rect 9214 31838 9266 31890
rect 9266 31838 9268 31890
rect 9212 31836 9268 31838
rect 8768 31332 8824 31388
rect 8872 31386 8928 31388
rect 8976 31386 9032 31388
rect 8872 31334 8896 31386
rect 8896 31334 8928 31386
rect 8976 31334 9020 31386
rect 9020 31334 9032 31386
rect 8872 31332 8928 31334
rect 8976 31332 9032 31334
rect 9080 31332 9136 31388
rect 9184 31386 9240 31388
rect 9288 31386 9344 31388
rect 9184 31334 9196 31386
rect 9196 31334 9240 31386
rect 9288 31334 9320 31386
rect 9320 31334 9344 31386
rect 9184 31332 9240 31334
rect 9288 31332 9344 31334
rect 9392 31332 9448 31388
rect 9436 30210 9492 30212
rect 9436 30158 9438 30210
rect 9438 30158 9490 30210
rect 9490 30158 9492 30210
rect 9436 30156 9492 30158
rect 8768 29764 8824 29820
rect 8872 29818 8928 29820
rect 8976 29818 9032 29820
rect 8872 29766 8896 29818
rect 8896 29766 8928 29818
rect 8976 29766 9020 29818
rect 9020 29766 9032 29818
rect 8872 29764 8928 29766
rect 8976 29764 9032 29766
rect 9080 29764 9136 29820
rect 9184 29818 9240 29820
rect 9288 29818 9344 29820
rect 9184 29766 9196 29818
rect 9196 29766 9240 29818
rect 9288 29766 9320 29818
rect 9320 29766 9344 29818
rect 9184 29764 9240 29766
rect 9288 29764 9344 29766
rect 9392 29764 9448 29820
rect 8768 28196 8824 28252
rect 8872 28250 8928 28252
rect 8976 28250 9032 28252
rect 8872 28198 8896 28250
rect 8896 28198 8928 28250
rect 8976 28198 9020 28250
rect 9020 28198 9032 28250
rect 8872 28196 8928 28198
rect 8976 28196 9032 28198
rect 9080 28196 9136 28252
rect 9184 28250 9240 28252
rect 9288 28250 9344 28252
rect 9184 28198 9196 28250
rect 9196 28198 9240 28250
rect 9288 28198 9320 28250
rect 9320 28198 9344 28250
rect 9184 28196 9240 28198
rect 9288 28196 9344 28198
rect 9392 28196 9448 28252
rect 8768 26628 8824 26684
rect 8872 26682 8928 26684
rect 8976 26682 9032 26684
rect 8872 26630 8896 26682
rect 8896 26630 8928 26682
rect 8976 26630 9020 26682
rect 9020 26630 9032 26682
rect 8872 26628 8928 26630
rect 8976 26628 9032 26630
rect 9080 26628 9136 26684
rect 9184 26682 9240 26684
rect 9288 26682 9344 26684
rect 9184 26630 9196 26682
rect 9196 26630 9240 26682
rect 9288 26630 9320 26682
rect 9320 26630 9344 26682
rect 9184 26628 9240 26630
rect 9288 26628 9344 26630
rect 9392 26628 9448 26684
rect 3164 23436 3220 23492
rect 6076 24780 6132 24836
rect 5292 23266 5348 23268
rect 5292 23214 5294 23266
rect 5294 23214 5346 23266
rect 5346 23214 5348 23266
rect 5292 23212 5348 23214
rect 4268 22708 4324 22764
rect 4372 22762 4428 22764
rect 4476 22762 4532 22764
rect 4372 22710 4396 22762
rect 4396 22710 4428 22762
rect 4476 22710 4520 22762
rect 4520 22710 4532 22762
rect 4372 22708 4428 22710
rect 4476 22708 4532 22710
rect 4580 22708 4636 22764
rect 4684 22762 4740 22764
rect 4788 22762 4844 22764
rect 4684 22710 4696 22762
rect 4696 22710 4740 22762
rect 4788 22710 4820 22762
rect 4820 22710 4844 22762
rect 4684 22708 4740 22710
rect 4788 22708 4844 22710
rect 4892 22708 4948 22764
rect 2716 21420 2772 21476
rect 2828 22316 2884 22372
rect 2380 19404 2436 19460
rect 2268 18620 2324 18676
rect 2940 21980 2996 22036
rect 4268 21140 4324 21196
rect 4372 21194 4428 21196
rect 4476 21194 4532 21196
rect 4372 21142 4396 21194
rect 4396 21142 4428 21194
rect 4476 21142 4520 21194
rect 4520 21142 4532 21194
rect 4372 21140 4428 21142
rect 4476 21140 4532 21142
rect 4580 21140 4636 21196
rect 4684 21194 4740 21196
rect 4788 21194 4844 21196
rect 4684 21142 4696 21194
rect 4696 21142 4740 21194
rect 4788 21142 4820 21194
rect 4820 21142 4844 21194
rect 4684 21140 4740 21142
rect 4788 21140 4844 21142
rect 4892 21140 4948 21196
rect 4620 20972 4676 21028
rect 4508 19964 4564 20020
rect 5292 20130 5348 20132
rect 5292 20078 5294 20130
rect 5294 20078 5346 20130
rect 5346 20078 5348 20130
rect 5292 20076 5348 20078
rect 5068 19852 5124 19908
rect 8768 25060 8824 25116
rect 8872 25114 8928 25116
rect 8976 25114 9032 25116
rect 8872 25062 8896 25114
rect 8896 25062 8928 25114
rect 8976 25062 9020 25114
rect 9020 25062 9032 25114
rect 8872 25060 8928 25062
rect 8976 25060 9032 25062
rect 9080 25060 9136 25116
rect 9184 25114 9240 25116
rect 9288 25114 9344 25116
rect 9184 25062 9196 25114
rect 9196 25062 9240 25114
rect 9288 25062 9320 25114
rect 9320 25062 9344 25114
rect 9184 25060 9240 25062
rect 9288 25060 9344 25062
rect 9392 25060 9448 25116
rect 8428 24780 8484 24836
rect 6076 22370 6132 22372
rect 6076 22318 6078 22370
rect 6078 22318 6130 22370
rect 6130 22318 6132 22370
rect 6076 22316 6132 22318
rect 5852 20972 5908 21028
rect 9660 23772 9716 23828
rect 8768 23492 8824 23548
rect 8872 23546 8928 23548
rect 8976 23546 9032 23548
rect 8872 23494 8896 23546
rect 8896 23494 8928 23546
rect 8976 23494 9020 23546
rect 9020 23494 9032 23546
rect 8872 23492 8928 23494
rect 8976 23492 9032 23494
rect 9080 23492 9136 23548
rect 9184 23546 9240 23548
rect 9288 23546 9344 23548
rect 9184 23494 9196 23546
rect 9196 23494 9240 23546
rect 9288 23494 9320 23546
rect 9320 23494 9344 23546
rect 9184 23492 9240 23494
rect 9288 23492 9344 23494
rect 9392 23492 9448 23548
rect 9996 29932 10052 29988
rect 9996 27916 10052 27972
rect 8428 22428 8484 22484
rect 9548 22482 9604 22484
rect 9548 22430 9550 22482
rect 9550 22430 9602 22482
rect 9602 22430 9604 22482
rect 9548 22428 9604 22430
rect 8768 21924 8824 21980
rect 8872 21978 8928 21980
rect 8976 21978 9032 21980
rect 8872 21926 8896 21978
rect 8896 21926 8928 21978
rect 8976 21926 9020 21978
rect 9020 21926 9032 21978
rect 8872 21924 8928 21926
rect 8976 21924 9032 21926
rect 9080 21924 9136 21980
rect 9184 21978 9240 21980
rect 9288 21978 9344 21980
rect 9184 21926 9196 21978
rect 9196 21926 9240 21978
rect 9288 21926 9320 21978
rect 9320 21926 9344 21978
rect 9184 21924 9240 21926
rect 9288 21924 9344 21926
rect 9392 21924 9448 21980
rect 9100 21756 9156 21812
rect 6748 20802 6804 20804
rect 6748 20750 6750 20802
rect 6750 20750 6802 20802
rect 6802 20750 6804 20802
rect 6748 20748 6804 20750
rect 8768 20356 8824 20412
rect 8872 20410 8928 20412
rect 8976 20410 9032 20412
rect 8872 20358 8896 20410
rect 8896 20358 8928 20410
rect 8976 20358 9020 20410
rect 9020 20358 9032 20410
rect 8872 20356 8928 20358
rect 8976 20356 9032 20358
rect 9080 20356 9136 20412
rect 9184 20410 9240 20412
rect 9288 20410 9344 20412
rect 9184 20358 9196 20410
rect 9196 20358 9240 20410
rect 9288 20358 9320 20410
rect 9320 20358 9344 20410
rect 9184 20356 9240 20358
rect 9288 20356 9344 20358
rect 9392 20356 9448 20412
rect 5740 19852 5796 19908
rect 6076 19964 6132 20020
rect 4268 19572 4324 19628
rect 4372 19626 4428 19628
rect 4476 19626 4532 19628
rect 4372 19574 4396 19626
rect 4396 19574 4428 19626
rect 4476 19574 4520 19626
rect 4520 19574 4532 19626
rect 4372 19572 4428 19574
rect 4476 19572 4532 19574
rect 4580 19572 4636 19628
rect 4684 19626 4740 19628
rect 4788 19626 4844 19628
rect 4684 19574 4696 19626
rect 4696 19574 4740 19626
rect 4788 19574 4820 19626
rect 4820 19574 4844 19626
rect 4684 19572 4740 19574
rect 4788 19572 4844 19574
rect 4892 19572 4948 19628
rect 3164 19346 3220 19348
rect 3164 19294 3166 19346
rect 3166 19294 3218 19346
rect 3218 19294 3220 19346
rect 3164 19292 3220 19294
rect 2828 18956 2884 19012
rect 2716 18620 2772 18676
rect 4268 18004 4324 18060
rect 4372 18058 4428 18060
rect 4476 18058 4532 18060
rect 4372 18006 4396 18058
rect 4396 18006 4428 18058
rect 4476 18006 4520 18058
rect 4520 18006 4532 18058
rect 4372 18004 4428 18006
rect 4476 18004 4532 18006
rect 4580 18004 4636 18060
rect 4684 18058 4740 18060
rect 4788 18058 4844 18060
rect 4684 18006 4696 18058
rect 4696 18006 4740 18058
rect 4788 18006 4820 18058
rect 4820 18006 4844 18058
rect 4684 18004 4740 18006
rect 4788 18004 4844 18006
rect 4892 18004 4948 18060
rect 2492 17554 2548 17556
rect 2492 17502 2494 17554
rect 2494 17502 2546 17554
rect 2546 17502 2548 17554
rect 2492 17500 2548 17502
rect 1708 16380 1764 16436
rect 2492 16380 2548 16436
rect 4268 16436 4324 16492
rect 4372 16490 4428 16492
rect 4476 16490 4532 16492
rect 4372 16438 4396 16490
rect 4396 16438 4428 16490
rect 4476 16438 4520 16490
rect 4520 16438 4532 16490
rect 4372 16436 4428 16438
rect 4476 16436 4532 16438
rect 4580 16436 4636 16492
rect 4684 16490 4740 16492
rect 4788 16490 4844 16492
rect 4684 16438 4696 16490
rect 4696 16438 4740 16490
rect 4788 16438 4820 16490
rect 4820 16438 4844 16490
rect 4684 16436 4740 16438
rect 4788 16436 4844 16438
rect 4892 16436 4948 16492
rect 4268 14868 4324 14924
rect 4372 14922 4428 14924
rect 4476 14922 4532 14924
rect 4372 14870 4396 14922
rect 4396 14870 4428 14922
rect 4476 14870 4520 14922
rect 4520 14870 4532 14922
rect 4372 14868 4428 14870
rect 4476 14868 4532 14870
rect 4580 14868 4636 14924
rect 4684 14922 4740 14924
rect 4788 14922 4844 14924
rect 4684 14870 4696 14922
rect 4696 14870 4740 14922
rect 4788 14870 4820 14922
rect 4820 14870 4844 14922
rect 4684 14868 4740 14870
rect 4788 14868 4844 14870
rect 4892 14868 4948 14924
rect 2044 13970 2100 13972
rect 2044 13918 2046 13970
rect 2046 13918 2098 13970
rect 2098 13918 2100 13970
rect 2044 13916 2100 13918
rect 1708 13020 1764 13076
rect 4268 13300 4324 13356
rect 4372 13354 4428 13356
rect 4476 13354 4532 13356
rect 4372 13302 4396 13354
rect 4396 13302 4428 13354
rect 4476 13302 4520 13354
rect 4520 13302 4532 13354
rect 4372 13300 4428 13302
rect 4476 13300 4532 13302
rect 4580 13300 4636 13356
rect 4684 13354 4740 13356
rect 4788 13354 4844 13356
rect 4684 13302 4696 13354
rect 4696 13302 4740 13354
rect 4788 13302 4820 13354
rect 4820 13302 4844 13354
rect 4684 13300 4740 13302
rect 4788 13300 4844 13302
rect 4892 13300 4948 13356
rect 2492 13020 2548 13076
rect 2044 12290 2100 12292
rect 2044 12238 2046 12290
rect 2046 12238 2098 12290
rect 2098 12238 2100 12290
rect 2044 12236 2100 12238
rect 1708 11900 1764 11956
rect 2492 11900 2548 11956
rect 4268 11732 4324 11788
rect 4372 11786 4428 11788
rect 4476 11786 4532 11788
rect 4372 11734 4396 11786
rect 4396 11734 4428 11786
rect 4476 11734 4520 11786
rect 4520 11734 4532 11786
rect 4372 11732 4428 11734
rect 4476 11732 4532 11734
rect 4580 11732 4636 11788
rect 4684 11786 4740 11788
rect 4788 11786 4844 11788
rect 4684 11734 4696 11786
rect 4696 11734 4740 11786
rect 4788 11734 4820 11786
rect 4820 11734 4844 11786
rect 4684 11732 4740 11734
rect 4788 11732 4844 11734
rect 4892 11732 4948 11788
rect 2044 11170 2100 11172
rect 2044 11118 2046 11170
rect 2046 11118 2098 11170
rect 2098 11118 2100 11170
rect 2044 11116 2100 11118
rect 1708 10780 1764 10836
rect 2492 10780 2548 10836
rect 4268 10164 4324 10220
rect 4372 10218 4428 10220
rect 4476 10218 4532 10220
rect 4372 10166 4396 10218
rect 4396 10166 4428 10218
rect 4476 10166 4520 10218
rect 4520 10166 4532 10218
rect 4372 10164 4428 10166
rect 4476 10164 4532 10166
rect 4580 10164 4636 10220
rect 4684 10218 4740 10220
rect 4788 10218 4844 10220
rect 4684 10166 4696 10218
rect 4696 10166 4740 10218
rect 4788 10166 4820 10218
rect 4820 10166 4844 10218
rect 4684 10164 4740 10166
rect 4788 10164 4844 10166
rect 4892 10164 4948 10220
rect 1708 9714 1764 9716
rect 1708 9662 1710 9714
rect 1710 9662 1762 9714
rect 1762 9662 1764 9714
rect 1708 9660 1764 9662
rect 2492 9714 2548 9716
rect 2492 9662 2494 9714
rect 2494 9662 2546 9714
rect 2546 9662 2548 9714
rect 2492 9660 2548 9662
rect 2044 9602 2100 9604
rect 2044 9550 2046 9602
rect 2046 9550 2098 9602
rect 2098 9550 2100 9602
rect 2044 9548 2100 9550
rect 4268 8596 4324 8652
rect 4372 8650 4428 8652
rect 4476 8650 4532 8652
rect 4372 8598 4396 8650
rect 4396 8598 4428 8650
rect 4476 8598 4520 8650
rect 4520 8598 4532 8650
rect 4372 8596 4428 8598
rect 4476 8596 4532 8598
rect 4580 8596 4636 8652
rect 4684 8650 4740 8652
rect 4788 8650 4844 8652
rect 4684 8598 4696 8650
rect 4696 8598 4740 8650
rect 4788 8598 4820 8650
rect 4820 8598 4844 8650
rect 4684 8596 4740 8598
rect 4788 8596 4844 8598
rect 4892 8596 4948 8652
rect 4268 7028 4324 7084
rect 4372 7082 4428 7084
rect 4476 7082 4532 7084
rect 4372 7030 4396 7082
rect 4396 7030 4428 7082
rect 4476 7030 4520 7082
rect 4520 7030 4532 7082
rect 4372 7028 4428 7030
rect 4476 7028 4532 7030
rect 4580 7028 4636 7084
rect 4684 7082 4740 7084
rect 4788 7082 4844 7084
rect 4684 7030 4696 7082
rect 4696 7030 4740 7082
rect 4788 7030 4820 7082
rect 4820 7030 4844 7082
rect 4684 7028 4740 7030
rect 4788 7028 4844 7030
rect 4892 7028 4948 7084
rect 1708 6300 1764 6356
rect 2268 6076 2324 6132
rect 2268 5794 2324 5796
rect 2268 5742 2270 5794
rect 2270 5742 2322 5794
rect 2322 5742 2324 5794
rect 2268 5740 2324 5742
rect 4268 5460 4324 5516
rect 4372 5514 4428 5516
rect 4476 5514 4532 5516
rect 4372 5462 4396 5514
rect 4396 5462 4428 5514
rect 4476 5462 4520 5514
rect 4520 5462 4532 5514
rect 4372 5460 4428 5462
rect 4476 5460 4532 5462
rect 4580 5460 4636 5516
rect 4684 5514 4740 5516
rect 4788 5514 4844 5516
rect 4684 5462 4696 5514
rect 4696 5462 4740 5514
rect 4788 5462 4820 5514
rect 4820 5462 4844 5514
rect 4684 5460 4740 5462
rect 4788 5460 4844 5462
rect 4892 5460 4948 5516
rect 1820 5234 1876 5236
rect 1820 5182 1822 5234
rect 1822 5182 1874 5234
rect 1874 5182 1876 5234
rect 1820 5180 1876 5182
rect 4268 3892 4324 3948
rect 4372 3946 4428 3948
rect 4476 3946 4532 3948
rect 4372 3894 4396 3946
rect 4396 3894 4428 3946
rect 4476 3894 4520 3946
rect 4520 3894 4532 3946
rect 4372 3892 4428 3894
rect 4476 3892 4532 3894
rect 4580 3892 4636 3948
rect 4684 3946 4740 3948
rect 4788 3946 4844 3948
rect 4684 3894 4696 3946
rect 4696 3894 4740 3946
rect 4788 3894 4820 3946
rect 4820 3894 4844 3946
rect 4684 3892 4740 3894
rect 4788 3892 4844 3894
rect 4892 3892 4948 3948
rect 7308 19906 7364 19908
rect 7308 19854 7310 19906
rect 7310 19854 7362 19906
rect 7362 19854 7364 19906
rect 7308 19852 7364 19854
rect 8768 18788 8824 18844
rect 8872 18842 8928 18844
rect 8976 18842 9032 18844
rect 8872 18790 8896 18842
rect 8896 18790 8928 18842
rect 8976 18790 9020 18842
rect 9020 18790 9032 18842
rect 8872 18788 8928 18790
rect 8976 18788 9032 18790
rect 9080 18788 9136 18844
rect 9184 18842 9240 18844
rect 9288 18842 9344 18844
rect 9184 18790 9196 18842
rect 9196 18790 9240 18842
rect 9288 18790 9320 18842
rect 9320 18790 9344 18842
rect 9184 18788 9240 18790
rect 9288 18788 9344 18790
rect 9392 18788 9448 18844
rect 8768 17220 8824 17276
rect 8872 17274 8928 17276
rect 8976 17274 9032 17276
rect 8872 17222 8896 17274
rect 8896 17222 8928 17274
rect 8976 17222 9020 17274
rect 9020 17222 9032 17274
rect 8872 17220 8928 17222
rect 8976 17220 9032 17222
rect 9080 17220 9136 17276
rect 9184 17274 9240 17276
rect 9288 17274 9344 17276
rect 9184 17222 9196 17274
rect 9196 17222 9240 17274
rect 9288 17222 9320 17274
rect 9320 17222 9344 17274
rect 9184 17220 9240 17222
rect 9288 17220 9344 17222
rect 9392 17220 9448 17276
rect 8768 15652 8824 15708
rect 8872 15706 8928 15708
rect 8976 15706 9032 15708
rect 8872 15654 8896 15706
rect 8896 15654 8928 15706
rect 8976 15654 9020 15706
rect 9020 15654 9032 15706
rect 8872 15652 8928 15654
rect 8976 15652 9032 15654
rect 9080 15652 9136 15708
rect 9184 15706 9240 15708
rect 9288 15706 9344 15708
rect 9184 15654 9196 15706
rect 9196 15654 9240 15706
rect 9288 15654 9320 15706
rect 9320 15654 9344 15706
rect 9184 15652 9240 15654
rect 9288 15652 9344 15654
rect 9392 15652 9448 15708
rect 8768 14084 8824 14140
rect 8872 14138 8928 14140
rect 8976 14138 9032 14140
rect 8872 14086 8896 14138
rect 8896 14086 8928 14138
rect 8976 14086 9020 14138
rect 9020 14086 9032 14138
rect 8872 14084 8928 14086
rect 8976 14084 9032 14086
rect 9080 14084 9136 14140
rect 9184 14138 9240 14140
rect 9288 14138 9344 14140
rect 9184 14086 9196 14138
rect 9196 14086 9240 14138
rect 9288 14086 9320 14138
rect 9320 14086 9344 14138
rect 9184 14084 9240 14086
rect 9288 14084 9344 14086
rect 9392 14084 9448 14140
rect 12236 42530 12292 42532
rect 12236 42478 12238 42530
rect 12238 42478 12290 42530
rect 12290 42478 12292 42530
rect 12236 42476 12292 42478
rect 12908 42530 12964 42532
rect 12908 42478 12910 42530
rect 12910 42478 12962 42530
rect 12962 42478 12964 42530
rect 12908 42476 12964 42478
rect 13268 43092 13324 43148
rect 13372 43146 13428 43148
rect 13476 43146 13532 43148
rect 13372 43094 13396 43146
rect 13396 43094 13428 43146
rect 13476 43094 13520 43146
rect 13520 43094 13532 43146
rect 13372 43092 13428 43094
rect 13476 43092 13532 43094
rect 13580 43092 13636 43148
rect 13684 43146 13740 43148
rect 13788 43146 13844 43148
rect 13684 43094 13696 43146
rect 13696 43094 13740 43146
rect 13788 43094 13820 43146
rect 13820 43094 13844 43146
rect 13684 43092 13740 43094
rect 13788 43092 13844 43094
rect 13892 43092 13948 43148
rect 13580 42924 13636 42980
rect 13244 42812 13300 42868
rect 14028 42812 14084 42868
rect 13804 42754 13860 42756
rect 13804 42702 13806 42754
rect 13806 42702 13858 42754
rect 13858 42702 13860 42754
rect 13804 42700 13860 42702
rect 13804 42476 13860 42532
rect 15148 42700 15204 42756
rect 14700 42642 14756 42644
rect 14700 42590 14702 42642
rect 14702 42590 14754 42642
rect 14754 42590 14756 42642
rect 14700 42588 14756 42590
rect 17768 48580 17824 48636
rect 17872 48634 17928 48636
rect 17976 48634 18032 48636
rect 17872 48582 17896 48634
rect 17896 48582 17928 48634
rect 17976 48582 18020 48634
rect 18020 48582 18032 48634
rect 17872 48580 17928 48582
rect 17976 48580 18032 48582
rect 18080 48580 18136 48636
rect 18184 48634 18240 48636
rect 18288 48634 18344 48636
rect 18184 48582 18196 48634
rect 18196 48582 18240 48634
rect 18288 48582 18320 48634
rect 18320 48582 18344 48634
rect 18184 48580 18240 48582
rect 18288 48580 18344 48582
rect 18392 48580 18448 48636
rect 19852 48354 19908 48356
rect 19852 48302 19854 48354
rect 19854 48302 19906 48354
rect 19906 48302 19908 48354
rect 19852 48300 19908 48302
rect 20300 48300 20356 48356
rect 15820 48242 15876 48244
rect 15820 48190 15822 48242
rect 15822 48190 15874 48242
rect 15874 48190 15876 48242
rect 15820 48188 15876 48190
rect 20860 50482 20916 50484
rect 20860 50430 20862 50482
rect 20862 50430 20914 50482
rect 20914 50430 20916 50482
rect 20860 50428 20916 50430
rect 25564 49810 25620 49812
rect 25564 49758 25566 49810
rect 25566 49758 25618 49810
rect 25618 49758 25620 49810
rect 25564 49756 25620 49758
rect 26908 52050 26964 52052
rect 26908 51998 26910 52050
rect 26910 51998 26962 52050
rect 26962 51998 26964 52050
rect 26908 51996 26964 51998
rect 27020 51938 27076 51940
rect 27020 51886 27022 51938
rect 27022 51886 27074 51938
rect 27074 51886 27076 51938
rect 27020 51884 27076 51886
rect 27692 52892 27748 52948
rect 29260 53340 29316 53396
rect 30828 53618 30884 53620
rect 30828 53566 30830 53618
rect 30830 53566 30882 53618
rect 30882 53566 30884 53618
rect 30828 53564 30884 53566
rect 40268 55636 40324 55692
rect 40372 55690 40428 55692
rect 40476 55690 40532 55692
rect 40372 55638 40396 55690
rect 40396 55638 40428 55690
rect 40476 55638 40520 55690
rect 40520 55638 40532 55690
rect 40372 55636 40428 55638
rect 40476 55636 40532 55638
rect 40580 55636 40636 55692
rect 40684 55690 40740 55692
rect 40788 55690 40844 55692
rect 40684 55638 40696 55690
rect 40696 55638 40740 55690
rect 40788 55638 40820 55690
rect 40820 55638 40844 55690
rect 40684 55636 40740 55638
rect 40788 55636 40844 55638
rect 40892 55636 40948 55692
rect 33180 55298 33236 55300
rect 33180 55246 33182 55298
rect 33182 55246 33234 55298
rect 33234 55246 33236 55298
rect 33180 55244 33236 55246
rect 33628 55298 33684 55300
rect 33628 55246 33630 55298
rect 33630 55246 33682 55298
rect 33682 55246 33684 55298
rect 33628 55244 33684 55246
rect 32060 53564 32116 53620
rect 29596 53116 29652 53172
rect 29372 53004 29428 53060
rect 28028 52834 28084 52836
rect 28028 52782 28030 52834
rect 28030 52782 28082 52834
rect 28082 52782 28084 52834
rect 28028 52780 28084 52782
rect 28812 52946 28868 52948
rect 28812 52894 28814 52946
rect 28814 52894 28866 52946
rect 28866 52894 28868 52946
rect 28812 52892 28868 52894
rect 28588 52780 28644 52836
rect 28588 52444 28644 52500
rect 28476 52386 28532 52388
rect 28476 52334 28478 52386
rect 28478 52334 28530 52386
rect 28530 52334 28532 52386
rect 28476 52332 28532 52334
rect 28364 52274 28420 52276
rect 28364 52222 28366 52274
rect 28366 52222 28418 52274
rect 28418 52222 28420 52274
rect 28364 52220 28420 52222
rect 29260 52274 29316 52276
rect 29260 52222 29262 52274
rect 29262 52222 29314 52274
rect 29314 52222 29316 52274
rect 29260 52220 29316 52222
rect 28140 52162 28196 52164
rect 28140 52110 28142 52162
rect 28142 52110 28194 52162
rect 28194 52110 28196 52162
rect 28140 52108 28196 52110
rect 28812 52108 28868 52164
rect 27804 52050 27860 52052
rect 27804 51998 27806 52050
rect 27806 51998 27858 52050
rect 27858 51998 27860 52050
rect 27804 51996 27860 51998
rect 26768 51716 26824 51772
rect 26872 51770 26928 51772
rect 26976 51770 27032 51772
rect 26872 51718 26896 51770
rect 26896 51718 26928 51770
rect 26976 51718 27020 51770
rect 27020 51718 27032 51770
rect 26872 51716 26928 51718
rect 26976 51716 27032 51718
rect 27080 51716 27136 51772
rect 27184 51770 27240 51772
rect 27288 51770 27344 51772
rect 27184 51718 27196 51770
rect 27196 51718 27240 51770
rect 27288 51718 27320 51770
rect 27320 51718 27344 51770
rect 27184 51716 27240 51718
rect 27288 51716 27344 51718
rect 27392 51716 27448 51772
rect 29932 53506 29988 53508
rect 29932 53454 29934 53506
rect 29934 53454 29986 53506
rect 29986 53454 29988 53506
rect 29932 53452 29988 53454
rect 29820 53058 29876 53060
rect 29820 53006 29822 53058
rect 29822 53006 29874 53058
rect 29874 53006 29876 53058
rect 29820 53004 29876 53006
rect 26768 50148 26824 50204
rect 26872 50202 26928 50204
rect 26976 50202 27032 50204
rect 26872 50150 26896 50202
rect 26896 50150 26928 50202
rect 26976 50150 27020 50202
rect 27020 50150 27032 50202
rect 26872 50148 26928 50150
rect 26976 50148 27032 50150
rect 27080 50148 27136 50204
rect 27184 50202 27240 50204
rect 27288 50202 27344 50204
rect 27184 50150 27196 50202
rect 27196 50150 27240 50202
rect 27288 50150 27320 50202
rect 27320 50150 27344 50202
rect 27184 50148 27240 50150
rect 27288 50148 27344 50150
rect 27392 50148 27448 50204
rect 26348 49756 26404 49812
rect 29484 50316 29540 50372
rect 30716 53506 30772 53508
rect 30716 53454 30718 53506
rect 30718 53454 30770 53506
rect 30770 53454 30772 53506
rect 30716 53452 30772 53454
rect 31276 53506 31332 53508
rect 31276 53454 31278 53506
rect 31278 53454 31330 53506
rect 31330 53454 31332 53506
rect 31276 53452 31332 53454
rect 30156 53340 30212 53396
rect 31164 53004 31220 53060
rect 30156 52668 30212 52724
rect 30156 52162 30212 52164
rect 30156 52110 30158 52162
rect 30158 52110 30210 52162
rect 30210 52110 30212 52162
rect 30156 52108 30212 52110
rect 30828 52108 30884 52164
rect 31276 52946 31332 52948
rect 31276 52894 31278 52946
rect 31278 52894 31330 52946
rect 31330 52894 31332 52946
rect 31276 52892 31332 52894
rect 31948 52892 32004 52948
rect 31268 52500 31324 52556
rect 31372 52554 31428 52556
rect 31476 52554 31532 52556
rect 31372 52502 31396 52554
rect 31396 52502 31428 52554
rect 31476 52502 31520 52554
rect 31520 52502 31532 52554
rect 31372 52500 31428 52502
rect 31476 52500 31532 52502
rect 31580 52500 31636 52556
rect 31684 52554 31740 52556
rect 31788 52554 31844 52556
rect 31684 52502 31696 52554
rect 31696 52502 31740 52554
rect 31788 52502 31820 52554
rect 31820 52502 31844 52554
rect 31684 52500 31740 52502
rect 31788 52500 31844 52502
rect 31892 52500 31948 52556
rect 31052 52332 31108 52388
rect 32172 52668 32228 52724
rect 33964 53788 34020 53844
rect 33740 53058 33796 53060
rect 33740 53006 33742 53058
rect 33742 53006 33794 53058
rect 33794 53006 33796 53058
rect 33740 53004 33796 53006
rect 32172 52332 32228 52388
rect 31276 52220 31332 52276
rect 31268 50932 31324 50988
rect 31372 50986 31428 50988
rect 31476 50986 31532 50988
rect 31372 50934 31396 50986
rect 31396 50934 31428 50986
rect 31476 50934 31520 50986
rect 31520 50934 31532 50986
rect 31372 50932 31428 50934
rect 31476 50932 31532 50934
rect 31580 50932 31636 50988
rect 31684 50986 31740 50988
rect 31788 50986 31844 50988
rect 31684 50934 31696 50986
rect 31696 50934 31740 50986
rect 31788 50934 31820 50986
rect 31820 50934 31844 50986
rect 31684 50932 31740 50934
rect 31788 50932 31844 50934
rect 31892 50932 31948 50988
rect 32956 52162 33012 52164
rect 32956 52110 32958 52162
rect 32958 52110 33010 52162
rect 33010 52110 33012 52162
rect 32956 52108 33012 52110
rect 35768 54852 35824 54908
rect 35872 54906 35928 54908
rect 35976 54906 36032 54908
rect 35872 54854 35896 54906
rect 35896 54854 35928 54906
rect 35976 54854 36020 54906
rect 36020 54854 36032 54906
rect 35872 54852 35928 54854
rect 35976 54852 36032 54854
rect 36080 54852 36136 54908
rect 36184 54906 36240 54908
rect 36288 54906 36344 54908
rect 36184 54854 36196 54906
rect 36196 54854 36240 54906
rect 36288 54854 36320 54906
rect 36320 54854 36344 54906
rect 36184 54852 36240 54854
rect 36288 54852 36344 54854
rect 36392 54852 36448 54908
rect 34412 53506 34468 53508
rect 34412 53454 34414 53506
rect 34414 53454 34466 53506
rect 34466 53454 34468 53506
rect 34412 53452 34468 53454
rect 34300 52946 34356 52948
rect 34300 52894 34302 52946
rect 34302 52894 34354 52946
rect 34354 52894 34356 52946
rect 34300 52892 34356 52894
rect 34300 52668 34356 52724
rect 34636 53506 34692 53508
rect 34636 53454 34638 53506
rect 34638 53454 34690 53506
rect 34690 53454 34692 53506
rect 34636 53452 34692 53454
rect 34412 52444 34468 52500
rect 35084 53788 35140 53844
rect 35644 53788 35700 53844
rect 35420 53564 35476 53620
rect 35196 53452 35252 53508
rect 37100 55298 37156 55300
rect 37100 55246 37102 55298
rect 37102 55246 37154 55298
rect 37154 55246 37156 55298
rect 37100 55244 37156 55246
rect 39788 55298 39844 55300
rect 39788 55246 39790 55298
rect 39790 55246 39842 55298
rect 39842 55246 39844 55298
rect 39788 55244 39844 55246
rect 38892 54460 38948 54516
rect 36540 53676 36596 53732
rect 36764 53788 36820 53844
rect 35868 53618 35924 53620
rect 35868 53566 35870 53618
rect 35870 53566 35922 53618
rect 35922 53566 35924 53618
rect 35868 53564 35924 53566
rect 34972 52444 35028 52500
rect 36204 53506 36260 53508
rect 36204 53454 36206 53506
rect 36206 53454 36258 53506
rect 36258 53454 36260 53506
rect 36204 53452 36260 53454
rect 36540 53452 36596 53508
rect 35768 53284 35824 53340
rect 35872 53338 35928 53340
rect 35976 53338 36032 53340
rect 35872 53286 35896 53338
rect 35896 53286 35928 53338
rect 35976 53286 36020 53338
rect 36020 53286 36032 53338
rect 35872 53284 35928 53286
rect 35976 53284 36032 53286
rect 36080 53284 36136 53340
rect 36184 53338 36240 53340
rect 36288 53338 36344 53340
rect 36184 53286 36196 53338
rect 36196 53286 36240 53338
rect 36288 53286 36320 53338
rect 36320 53286 36344 53338
rect 36184 53284 36240 53286
rect 36288 53284 36344 53286
rect 36392 53284 36448 53340
rect 35532 53170 35588 53172
rect 35532 53118 35534 53170
rect 35534 53118 35586 53170
rect 35586 53118 35588 53170
rect 35532 53116 35588 53118
rect 35868 53170 35924 53172
rect 35868 53118 35870 53170
rect 35870 53118 35922 53170
rect 35922 53118 35924 53170
rect 35868 53116 35924 53118
rect 35420 52892 35476 52948
rect 35644 52780 35700 52836
rect 36988 53340 37044 53396
rect 36988 53170 37044 53172
rect 36988 53118 36990 53170
rect 36990 53118 37042 53170
rect 37042 53118 37044 53170
rect 36988 53116 37044 53118
rect 38220 53730 38276 53732
rect 38220 53678 38222 53730
rect 38222 53678 38274 53730
rect 38274 53678 38276 53730
rect 38220 53676 38276 53678
rect 37212 52892 37268 52948
rect 36540 52834 36596 52836
rect 36540 52782 36542 52834
rect 36542 52782 36594 52834
rect 36594 52782 36596 52834
rect 36540 52780 36596 52782
rect 35644 52556 35700 52612
rect 35756 52668 35812 52724
rect 35308 52332 35364 52388
rect 40236 54514 40292 54516
rect 40236 54462 40238 54514
rect 40238 54462 40290 54514
rect 40290 54462 40292 54514
rect 40236 54460 40292 54462
rect 39900 54402 39956 54404
rect 39900 54350 39902 54402
rect 39902 54350 39954 54402
rect 39954 54350 39956 54402
rect 39900 54348 39956 54350
rect 39228 53676 39284 53732
rect 38332 53116 38388 53172
rect 41916 54572 41972 54628
rect 40268 54068 40324 54124
rect 40372 54122 40428 54124
rect 40476 54122 40532 54124
rect 40372 54070 40396 54122
rect 40396 54070 40428 54122
rect 40476 54070 40520 54122
rect 40520 54070 40532 54122
rect 40372 54068 40428 54070
rect 40476 54068 40532 54070
rect 40580 54068 40636 54124
rect 40684 54122 40740 54124
rect 40788 54122 40844 54124
rect 40684 54070 40696 54122
rect 40696 54070 40740 54122
rect 40788 54070 40820 54122
rect 40820 54070 40844 54122
rect 40684 54068 40740 54070
rect 40788 54068 40844 54070
rect 40892 54068 40948 54124
rect 39452 53340 39508 53396
rect 40124 53788 40180 53844
rect 39564 53228 39620 53284
rect 37324 52556 37380 52612
rect 38444 52834 38500 52836
rect 38444 52782 38446 52834
rect 38446 52782 38498 52834
rect 38498 52782 38500 52834
rect 38444 52780 38500 52782
rect 35308 52108 35364 52164
rect 36204 52162 36260 52164
rect 36204 52110 36206 52162
rect 36206 52110 36258 52162
rect 36258 52110 36260 52162
rect 36204 52108 36260 52110
rect 34188 51996 34244 52052
rect 29932 50316 29988 50372
rect 22268 49364 22324 49420
rect 22372 49418 22428 49420
rect 22476 49418 22532 49420
rect 22372 49366 22396 49418
rect 22396 49366 22428 49418
rect 22476 49366 22520 49418
rect 22520 49366 22532 49418
rect 22372 49364 22428 49366
rect 22476 49364 22532 49366
rect 22580 49364 22636 49420
rect 22684 49418 22740 49420
rect 22788 49418 22844 49420
rect 22684 49366 22696 49418
rect 22696 49366 22740 49418
rect 22788 49366 22820 49418
rect 22820 49366 22844 49418
rect 22684 49364 22740 49366
rect 22788 49364 22844 49366
rect 22892 49364 22948 49420
rect 16492 47964 16548 48020
rect 16492 47180 16548 47236
rect 17276 47292 17332 47348
rect 17612 47180 17668 47236
rect 18172 47234 18228 47236
rect 18172 47182 18174 47234
rect 18174 47182 18226 47234
rect 18226 47182 18228 47234
rect 18172 47180 18228 47182
rect 20748 47964 20804 48020
rect 20748 47404 20804 47460
rect 26768 48580 26824 48636
rect 26872 48634 26928 48636
rect 26976 48634 27032 48636
rect 26872 48582 26896 48634
rect 26896 48582 26928 48634
rect 26976 48582 27020 48634
rect 27020 48582 27032 48634
rect 26872 48580 26928 48582
rect 26976 48580 27032 48582
rect 27080 48580 27136 48636
rect 27184 48634 27240 48636
rect 27288 48634 27344 48636
rect 27184 48582 27196 48634
rect 27196 48582 27240 48634
rect 27288 48582 27320 48634
rect 27320 48582 27344 48634
rect 27184 48580 27240 48582
rect 27288 48580 27344 48582
rect 27392 48580 27448 48636
rect 21084 48130 21140 48132
rect 21084 48078 21086 48130
rect 21086 48078 21138 48130
rect 21138 48078 21140 48130
rect 21084 48076 21140 48078
rect 22092 48130 22148 48132
rect 22092 48078 22094 48130
rect 22094 48078 22146 48130
rect 22146 48078 22148 48130
rect 22092 48076 22148 48078
rect 21420 48018 21476 48020
rect 21420 47966 21422 48018
rect 21422 47966 21474 48018
rect 21474 47966 21476 48018
rect 21420 47964 21476 47966
rect 21756 47458 21812 47460
rect 21756 47406 21758 47458
rect 21758 47406 21810 47458
rect 21810 47406 21812 47458
rect 21756 47404 21812 47406
rect 20524 47180 20580 47236
rect 22268 47796 22324 47852
rect 22372 47850 22428 47852
rect 22476 47850 22532 47852
rect 22372 47798 22396 47850
rect 22396 47798 22428 47850
rect 22476 47798 22520 47850
rect 22520 47798 22532 47850
rect 22372 47796 22428 47798
rect 22476 47796 22532 47798
rect 22580 47796 22636 47852
rect 22684 47850 22740 47852
rect 22788 47850 22844 47852
rect 22684 47798 22696 47850
rect 22696 47798 22740 47850
rect 22788 47798 22820 47850
rect 22820 47798 22844 47850
rect 22684 47796 22740 47798
rect 22788 47796 22844 47798
rect 22892 47796 22948 47852
rect 22092 47180 22148 47236
rect 17768 47012 17824 47068
rect 17872 47066 17928 47068
rect 17976 47066 18032 47068
rect 17872 47014 17896 47066
rect 17896 47014 17928 47066
rect 17976 47014 18020 47066
rect 18020 47014 18032 47066
rect 17872 47012 17928 47014
rect 17976 47012 18032 47014
rect 18080 47012 18136 47068
rect 18184 47066 18240 47068
rect 18288 47066 18344 47068
rect 18184 47014 18196 47066
rect 18196 47014 18240 47066
rect 18288 47014 18320 47066
rect 18320 47014 18344 47066
rect 18184 47012 18240 47014
rect 18288 47012 18344 47014
rect 18392 47012 18448 47068
rect 20972 47068 21028 47124
rect 21532 47068 21588 47124
rect 17612 46508 17668 46564
rect 17768 45444 17824 45500
rect 17872 45498 17928 45500
rect 17976 45498 18032 45500
rect 17872 45446 17896 45498
rect 17896 45446 17928 45498
rect 17976 45446 18020 45498
rect 18020 45446 18032 45498
rect 17872 45444 17928 45446
rect 17976 45444 18032 45446
rect 18080 45444 18136 45500
rect 18184 45498 18240 45500
rect 18288 45498 18344 45500
rect 18184 45446 18196 45498
rect 18196 45446 18240 45498
rect 18288 45446 18320 45498
rect 18320 45446 18344 45498
rect 18184 45444 18240 45446
rect 18288 45444 18344 45446
rect 18392 45444 18448 45500
rect 17388 45164 17444 45220
rect 16492 45106 16548 45108
rect 16492 45054 16494 45106
rect 16494 45054 16546 45106
rect 16546 45054 16548 45106
rect 16492 45052 16548 45054
rect 16156 44882 16212 44884
rect 16156 44830 16158 44882
rect 16158 44830 16210 44882
rect 16210 44830 16212 44882
rect 16156 44828 16212 44830
rect 19628 45218 19684 45220
rect 19628 45166 19630 45218
rect 19630 45166 19682 45218
rect 19682 45166 19684 45218
rect 19628 45164 19684 45166
rect 17388 44156 17444 44212
rect 17612 44828 17668 44884
rect 20076 44380 20132 44436
rect 21420 44492 21476 44548
rect 17948 44098 18004 44100
rect 17948 44046 17950 44098
rect 17950 44046 18002 44098
rect 18002 44046 18004 44098
rect 17948 44044 18004 44046
rect 17768 43876 17824 43932
rect 17872 43930 17928 43932
rect 17976 43930 18032 43932
rect 17872 43878 17896 43930
rect 17896 43878 17928 43930
rect 17976 43878 18020 43930
rect 18020 43878 18032 43930
rect 17872 43876 17928 43878
rect 17976 43876 18032 43878
rect 18080 43876 18136 43932
rect 18184 43930 18240 43932
rect 18288 43930 18344 43932
rect 18184 43878 18196 43930
rect 18196 43878 18240 43930
rect 18288 43878 18320 43930
rect 18320 43878 18344 43930
rect 18184 43876 18240 43878
rect 18288 43876 18344 43878
rect 18392 43876 18448 43932
rect 20748 43596 20804 43652
rect 20748 42812 20804 42868
rect 18956 42754 19012 42756
rect 18956 42702 18958 42754
rect 18958 42702 19010 42754
rect 19010 42702 19012 42754
rect 18956 42700 19012 42702
rect 19516 42754 19572 42756
rect 19516 42702 19518 42754
rect 19518 42702 19570 42754
rect 19570 42702 19572 42754
rect 19516 42700 19572 42702
rect 20188 42754 20244 42756
rect 20188 42702 20190 42754
rect 20190 42702 20242 42754
rect 20242 42702 20244 42754
rect 20188 42700 20244 42702
rect 15596 42588 15652 42644
rect 19404 42642 19460 42644
rect 19404 42590 19406 42642
rect 19406 42590 19458 42642
rect 19458 42590 19460 42642
rect 19404 42588 19460 42590
rect 14364 42476 14420 42532
rect 15260 42530 15316 42532
rect 15260 42478 15262 42530
rect 15262 42478 15314 42530
rect 15314 42478 15316 42530
rect 15260 42476 15316 42478
rect 16940 42476 16996 42532
rect 16380 41916 16436 41972
rect 17768 42308 17824 42364
rect 17872 42362 17928 42364
rect 17976 42362 18032 42364
rect 17872 42310 17896 42362
rect 17896 42310 17928 42362
rect 17976 42310 18020 42362
rect 18020 42310 18032 42362
rect 17872 42308 17928 42310
rect 17976 42308 18032 42310
rect 18080 42308 18136 42364
rect 18184 42362 18240 42364
rect 18288 42362 18344 42364
rect 18184 42310 18196 42362
rect 18196 42310 18240 42362
rect 18288 42310 18320 42362
rect 18320 42310 18344 42362
rect 18184 42308 18240 42310
rect 18288 42308 18344 42310
rect 18392 42308 18448 42364
rect 17500 41970 17556 41972
rect 17500 41918 17502 41970
rect 17502 41918 17554 41970
rect 17554 41918 17556 41970
rect 17500 41916 17556 41918
rect 19740 41970 19796 41972
rect 19740 41918 19742 41970
rect 19742 41918 19794 41970
rect 19794 41918 19796 41970
rect 19740 41916 19796 41918
rect 13268 41524 13324 41580
rect 13372 41578 13428 41580
rect 13476 41578 13532 41580
rect 13372 41526 13396 41578
rect 13396 41526 13428 41578
rect 13476 41526 13520 41578
rect 13520 41526 13532 41578
rect 13372 41524 13428 41526
rect 13476 41524 13532 41526
rect 13580 41524 13636 41580
rect 13684 41578 13740 41580
rect 13788 41578 13844 41580
rect 13684 41526 13696 41578
rect 13696 41526 13740 41578
rect 13788 41526 13820 41578
rect 13820 41526 13844 41578
rect 13684 41524 13740 41526
rect 13788 41524 13844 41526
rect 13892 41524 13948 41580
rect 13132 41356 13188 41412
rect 12348 40908 12404 40964
rect 16940 40348 16996 40404
rect 13580 40124 13636 40180
rect 16828 40124 16884 40180
rect 12460 39900 12516 39956
rect 13268 39956 13324 40012
rect 13372 40010 13428 40012
rect 13476 40010 13532 40012
rect 13372 39958 13396 40010
rect 13396 39958 13428 40010
rect 13476 39958 13520 40010
rect 13520 39958 13532 40010
rect 13372 39956 13428 39958
rect 13476 39956 13532 39958
rect 13580 39956 13636 40012
rect 13684 40010 13740 40012
rect 13788 40010 13844 40012
rect 13684 39958 13696 40010
rect 13696 39958 13740 40010
rect 13788 39958 13820 40010
rect 13820 39958 13844 40010
rect 13684 39956 13740 39958
rect 13788 39956 13844 39958
rect 13892 39956 13948 40012
rect 15484 39564 15540 39620
rect 12796 39506 12852 39508
rect 12796 39454 12798 39506
rect 12798 39454 12850 39506
rect 12850 39454 12852 39506
rect 12796 39452 12852 39454
rect 13468 39506 13524 39508
rect 13468 39454 13470 39506
rect 13470 39454 13522 39506
rect 13522 39454 13524 39506
rect 13468 39452 13524 39454
rect 11788 39340 11844 39396
rect 10556 37378 10612 37380
rect 10556 37326 10558 37378
rect 10558 37326 10610 37378
rect 10610 37326 10612 37378
rect 10556 37324 10612 37326
rect 11340 36876 11396 36932
rect 11564 36258 11620 36260
rect 11564 36206 11566 36258
rect 11566 36206 11618 36258
rect 11618 36206 11620 36258
rect 11564 36204 11620 36206
rect 13356 39340 13412 39396
rect 14140 39394 14196 39396
rect 14140 39342 14142 39394
rect 14142 39342 14194 39394
rect 14194 39342 14196 39394
rect 14140 39340 14196 39342
rect 13268 38388 13324 38444
rect 13372 38442 13428 38444
rect 13476 38442 13532 38444
rect 13372 38390 13396 38442
rect 13396 38390 13428 38442
rect 13476 38390 13520 38442
rect 13520 38390 13532 38442
rect 13372 38388 13428 38390
rect 13476 38388 13532 38390
rect 13580 38388 13636 38444
rect 13684 38442 13740 38444
rect 13788 38442 13844 38444
rect 13684 38390 13696 38442
rect 13696 38390 13740 38442
rect 13788 38390 13820 38442
rect 13820 38390 13844 38442
rect 13684 38388 13740 38390
rect 13788 38388 13844 38390
rect 13892 38388 13948 38444
rect 11900 36988 11956 37044
rect 13268 36820 13324 36876
rect 13372 36874 13428 36876
rect 13476 36874 13532 36876
rect 13372 36822 13396 36874
rect 13396 36822 13428 36874
rect 13476 36822 13520 36874
rect 13520 36822 13532 36874
rect 13372 36820 13428 36822
rect 13476 36820 13532 36822
rect 13580 36820 13636 36876
rect 13684 36874 13740 36876
rect 13788 36874 13844 36876
rect 13684 36822 13696 36874
rect 13696 36822 13740 36874
rect 13788 36822 13820 36874
rect 13820 36822 13844 36874
rect 13684 36820 13740 36822
rect 13788 36820 13844 36822
rect 13892 36820 13948 36876
rect 12348 36482 12404 36484
rect 12348 36430 12350 36482
rect 12350 36430 12402 36482
rect 12402 36430 12404 36482
rect 12348 36428 12404 36430
rect 16268 39058 16324 39060
rect 16268 39006 16270 39058
rect 16270 39006 16322 39058
rect 16322 39006 16324 39058
rect 16268 39004 16324 39006
rect 16828 38722 16884 38724
rect 16828 38670 16830 38722
rect 16830 38670 16882 38722
rect 16882 38670 16884 38722
rect 16828 38668 16884 38670
rect 17612 41692 17668 41748
rect 24108 47068 24164 47124
rect 24892 47234 24948 47236
rect 24892 47182 24894 47234
rect 24894 47182 24946 47234
rect 24946 47182 24948 47234
rect 24892 47180 24948 47182
rect 26768 47012 26824 47068
rect 26872 47066 26928 47068
rect 26976 47066 27032 47068
rect 26872 47014 26896 47066
rect 26896 47014 26928 47066
rect 26976 47014 27020 47066
rect 27020 47014 27032 47066
rect 26872 47012 26928 47014
rect 26976 47012 27032 47014
rect 27080 47012 27136 47068
rect 27184 47066 27240 47068
rect 27288 47066 27344 47068
rect 27184 47014 27196 47066
rect 27196 47014 27240 47066
rect 27288 47014 27320 47066
rect 27320 47014 27344 47066
rect 27184 47012 27240 47014
rect 27288 47012 27344 47014
rect 27392 47012 27448 47068
rect 24892 46844 24948 46900
rect 22268 46228 22324 46284
rect 22372 46282 22428 46284
rect 22476 46282 22532 46284
rect 22372 46230 22396 46282
rect 22396 46230 22428 46282
rect 22476 46230 22520 46282
rect 22520 46230 22532 46282
rect 22372 46228 22428 46230
rect 22476 46228 22532 46230
rect 22580 46228 22636 46284
rect 22684 46282 22740 46284
rect 22788 46282 22844 46284
rect 22684 46230 22696 46282
rect 22696 46230 22740 46282
rect 22788 46230 22820 46282
rect 22820 46230 22844 46282
rect 22684 46228 22740 46230
rect 22788 46228 22844 46230
rect 22892 46228 22948 46284
rect 26124 46674 26180 46676
rect 26124 46622 26126 46674
rect 26126 46622 26178 46674
rect 26178 46622 26180 46674
rect 26124 46620 26180 46622
rect 26908 46620 26964 46676
rect 27244 46396 27300 46452
rect 29036 49810 29092 49812
rect 29036 49758 29038 49810
rect 29038 49758 29090 49810
rect 29090 49758 29092 49810
rect 29036 49756 29092 49758
rect 29932 49644 29988 49700
rect 31948 49698 32004 49700
rect 31948 49646 31950 49698
rect 31950 49646 32002 49698
rect 32002 49646 32004 49698
rect 31948 49644 32004 49646
rect 31268 49364 31324 49420
rect 31372 49418 31428 49420
rect 31476 49418 31532 49420
rect 31372 49366 31396 49418
rect 31396 49366 31428 49418
rect 31476 49366 31520 49418
rect 31520 49366 31532 49418
rect 31372 49364 31428 49366
rect 31476 49364 31532 49366
rect 31580 49364 31636 49420
rect 31684 49418 31740 49420
rect 31788 49418 31844 49420
rect 31684 49366 31696 49418
rect 31696 49366 31740 49418
rect 31788 49366 31820 49418
rect 31820 49366 31844 49418
rect 31684 49364 31740 49366
rect 31788 49364 31844 49366
rect 31892 49364 31948 49420
rect 29260 49138 29316 49140
rect 29260 49086 29262 49138
rect 29262 49086 29314 49138
rect 29314 49086 29316 49138
rect 29260 49084 29316 49086
rect 31268 47796 31324 47852
rect 31372 47850 31428 47852
rect 31476 47850 31532 47852
rect 31372 47798 31396 47850
rect 31396 47798 31428 47850
rect 31476 47798 31520 47850
rect 31520 47798 31532 47850
rect 31372 47796 31428 47798
rect 31476 47796 31532 47798
rect 31580 47796 31636 47852
rect 31684 47850 31740 47852
rect 31788 47850 31844 47852
rect 31684 47798 31696 47850
rect 31696 47798 31740 47850
rect 31788 47798 31820 47850
rect 31820 47798 31844 47850
rect 31684 47796 31740 47798
rect 31788 47796 31844 47798
rect 31892 47796 31948 47852
rect 30380 47516 30436 47572
rect 26768 45444 26824 45500
rect 26872 45498 26928 45500
rect 26976 45498 27032 45500
rect 26872 45446 26896 45498
rect 26896 45446 26928 45498
rect 26976 45446 27020 45498
rect 27020 45446 27032 45498
rect 26872 45444 26928 45446
rect 26976 45444 27032 45446
rect 27080 45444 27136 45500
rect 27184 45498 27240 45500
rect 27288 45498 27344 45500
rect 27184 45446 27196 45498
rect 27196 45446 27240 45498
rect 27288 45446 27320 45498
rect 27320 45446 27344 45498
rect 27184 45444 27240 45446
rect 27288 45444 27344 45446
rect 27392 45444 27448 45500
rect 31612 47516 31668 47572
rect 29148 46562 29204 46564
rect 29148 46510 29150 46562
rect 29150 46510 29202 46562
rect 29202 46510 29204 46562
rect 29148 46508 29204 46510
rect 29820 46562 29876 46564
rect 29820 46510 29822 46562
rect 29822 46510 29874 46562
rect 29874 46510 29876 46562
rect 29820 46508 29876 46510
rect 29484 46450 29540 46452
rect 29484 46398 29486 46450
rect 29486 46398 29538 46450
rect 29538 46398 29540 46450
rect 29484 46396 29540 46398
rect 28588 45724 28644 45780
rect 23436 45218 23492 45220
rect 23436 45166 23438 45218
rect 23438 45166 23490 45218
rect 23490 45166 23492 45218
rect 23436 45164 23492 45166
rect 22268 44660 22324 44716
rect 22372 44714 22428 44716
rect 22476 44714 22532 44716
rect 22372 44662 22396 44714
rect 22396 44662 22428 44714
rect 22476 44662 22520 44714
rect 22520 44662 22532 44714
rect 22372 44660 22428 44662
rect 22476 44660 22532 44662
rect 22580 44660 22636 44716
rect 22684 44714 22740 44716
rect 22788 44714 22844 44716
rect 22684 44662 22696 44714
rect 22696 44662 22740 44714
rect 22788 44662 22820 44714
rect 22820 44662 22844 44714
rect 22684 44660 22740 44662
rect 22788 44660 22844 44662
rect 22892 44660 22948 44716
rect 22540 44434 22596 44436
rect 22540 44382 22542 44434
rect 22542 44382 22594 44434
rect 22594 44382 22596 44434
rect 22540 44380 22596 44382
rect 22204 44044 22260 44100
rect 23100 44098 23156 44100
rect 23100 44046 23102 44098
rect 23102 44046 23154 44098
rect 23154 44046 23156 44098
rect 23100 44044 23156 44046
rect 24220 44044 24276 44100
rect 26768 43876 26824 43932
rect 26872 43930 26928 43932
rect 26976 43930 27032 43932
rect 26872 43878 26896 43930
rect 26896 43878 26928 43930
rect 26976 43878 27020 43930
rect 27020 43878 27032 43930
rect 26872 43876 26928 43878
rect 26976 43876 27032 43878
rect 27080 43876 27136 43932
rect 27184 43930 27240 43932
rect 27288 43930 27344 43932
rect 27184 43878 27196 43930
rect 27196 43878 27240 43930
rect 27288 43878 27320 43930
rect 27320 43878 27344 43930
rect 27184 43876 27240 43878
rect 27288 43876 27344 43878
rect 27392 43876 27448 43932
rect 21756 43596 21812 43652
rect 22268 43092 22324 43148
rect 22372 43146 22428 43148
rect 22476 43146 22532 43148
rect 22372 43094 22396 43146
rect 22396 43094 22428 43146
rect 22476 43094 22520 43146
rect 22520 43094 22532 43146
rect 22372 43092 22428 43094
rect 22476 43092 22532 43094
rect 22580 43092 22636 43148
rect 22684 43146 22740 43148
rect 22788 43146 22844 43148
rect 22684 43094 22696 43146
rect 22696 43094 22740 43146
rect 22788 43094 22820 43146
rect 22820 43094 22844 43146
rect 22684 43092 22740 43094
rect 22788 43092 22844 43094
rect 22892 43092 22948 43148
rect 21868 42700 21924 42756
rect 27244 43260 27300 43316
rect 28252 42812 28308 42868
rect 26236 42588 26292 42644
rect 26908 42642 26964 42644
rect 26908 42590 26910 42642
rect 26910 42590 26962 42642
rect 26962 42590 26964 42642
rect 26908 42588 26964 42590
rect 26768 42308 26824 42364
rect 26872 42362 26928 42364
rect 26976 42362 27032 42364
rect 26872 42310 26896 42362
rect 26896 42310 26928 42362
rect 26976 42310 27020 42362
rect 27020 42310 27032 42362
rect 26872 42308 26928 42310
rect 26976 42308 27032 42310
rect 27080 42308 27136 42364
rect 27184 42362 27240 42364
rect 27288 42362 27344 42364
rect 27184 42310 27196 42362
rect 27196 42310 27240 42362
rect 27288 42310 27320 42362
rect 27320 42310 27344 42362
rect 27184 42308 27240 42310
rect 27288 42308 27344 42310
rect 27392 42308 27448 42364
rect 21868 42028 21924 42084
rect 21532 41916 21588 41972
rect 21980 41916 22036 41972
rect 18508 41020 18564 41076
rect 17768 40740 17824 40796
rect 17872 40794 17928 40796
rect 17976 40794 18032 40796
rect 17872 40742 17896 40794
rect 17896 40742 17928 40794
rect 17976 40742 18020 40794
rect 18020 40742 18032 40794
rect 17872 40740 17928 40742
rect 17976 40740 18032 40742
rect 18080 40740 18136 40796
rect 18184 40794 18240 40796
rect 18288 40794 18344 40796
rect 18184 40742 18196 40794
rect 18196 40742 18240 40794
rect 18288 40742 18320 40794
rect 18320 40742 18344 40794
rect 18184 40740 18240 40742
rect 18288 40740 18344 40742
rect 18392 40740 18448 40796
rect 19068 41074 19124 41076
rect 19068 41022 19070 41074
rect 19070 41022 19122 41074
rect 19122 41022 19124 41074
rect 19068 41020 19124 41022
rect 21084 40572 21140 40628
rect 17500 40402 17556 40404
rect 17500 40350 17502 40402
rect 17502 40350 17554 40402
rect 17554 40350 17556 40402
rect 17500 40348 17556 40350
rect 17768 39172 17824 39228
rect 17872 39226 17928 39228
rect 17976 39226 18032 39228
rect 17872 39174 17896 39226
rect 17896 39174 17928 39226
rect 17976 39174 18020 39226
rect 18020 39174 18032 39226
rect 17872 39172 17928 39174
rect 17976 39172 18032 39174
rect 18080 39172 18136 39228
rect 18184 39226 18240 39228
rect 18288 39226 18344 39228
rect 18184 39174 18196 39226
rect 18196 39174 18240 39226
rect 18288 39174 18320 39226
rect 18320 39174 18344 39226
rect 18184 39172 18240 39174
rect 18288 39172 18344 39174
rect 18392 39172 18448 39228
rect 17500 39058 17556 39060
rect 17500 39006 17502 39058
rect 17502 39006 17554 39058
rect 17554 39006 17556 39058
rect 17500 39004 17556 39006
rect 24444 42082 24500 42084
rect 24444 42030 24446 42082
rect 24446 42030 24498 42082
rect 24498 42030 24500 42082
rect 24444 42028 24500 42030
rect 23548 41916 23604 41972
rect 22268 41524 22324 41580
rect 22372 41578 22428 41580
rect 22476 41578 22532 41580
rect 22372 41526 22396 41578
rect 22396 41526 22428 41578
rect 22476 41526 22520 41578
rect 22520 41526 22532 41578
rect 22372 41524 22428 41526
rect 22476 41524 22532 41526
rect 22580 41524 22636 41580
rect 22684 41578 22740 41580
rect 22788 41578 22844 41580
rect 22684 41526 22696 41578
rect 22696 41526 22740 41578
rect 22788 41526 22820 41578
rect 22820 41526 22844 41578
rect 22684 41524 22740 41526
rect 22788 41524 22844 41526
rect 22892 41524 22948 41580
rect 21980 40626 22036 40628
rect 21980 40574 21982 40626
rect 21982 40574 22034 40626
rect 22034 40574 22036 40626
rect 21980 40572 22036 40574
rect 22652 41020 22708 41076
rect 22988 40626 23044 40628
rect 22988 40574 22990 40626
rect 22990 40574 23042 40626
rect 23042 40574 23044 40626
rect 22988 40572 23044 40574
rect 26768 40740 26824 40796
rect 26872 40794 26928 40796
rect 26976 40794 27032 40796
rect 26872 40742 26896 40794
rect 26896 40742 26928 40794
rect 26976 40742 27020 40794
rect 27020 40742 27032 40794
rect 26872 40740 26928 40742
rect 26976 40740 27032 40742
rect 27080 40740 27136 40796
rect 27184 40794 27240 40796
rect 27288 40794 27344 40796
rect 27184 40742 27196 40794
rect 27196 40742 27240 40794
rect 27288 40742 27320 40794
rect 27320 40742 27344 40794
rect 27184 40740 27240 40742
rect 27288 40740 27344 40742
rect 27392 40740 27448 40796
rect 29260 45778 29316 45780
rect 29260 45726 29262 45778
rect 29262 45726 29314 45778
rect 29314 45726 29316 45778
rect 29260 45724 29316 45726
rect 30604 45778 30660 45780
rect 30604 45726 30606 45778
rect 30606 45726 30658 45778
rect 30658 45726 30660 45778
rect 30604 45724 30660 45726
rect 31268 46228 31324 46284
rect 31372 46282 31428 46284
rect 31476 46282 31532 46284
rect 31372 46230 31396 46282
rect 31396 46230 31428 46282
rect 31476 46230 31520 46282
rect 31520 46230 31532 46282
rect 31372 46228 31428 46230
rect 31476 46228 31532 46230
rect 31580 46228 31636 46284
rect 31684 46282 31740 46284
rect 31788 46282 31844 46284
rect 31684 46230 31696 46282
rect 31696 46230 31740 46282
rect 31788 46230 31820 46282
rect 31820 46230 31844 46282
rect 31684 46228 31740 46230
rect 31788 46228 31844 46230
rect 31892 46228 31948 46284
rect 31500 46060 31556 46116
rect 32844 49196 32900 49252
rect 32284 49084 32340 49140
rect 37996 51996 38052 52052
rect 35768 51716 35824 51772
rect 35872 51770 35928 51772
rect 35976 51770 36032 51772
rect 35872 51718 35896 51770
rect 35896 51718 35928 51770
rect 35976 51718 36020 51770
rect 36020 51718 36032 51770
rect 35872 51716 35928 51718
rect 35976 51716 36032 51718
rect 36080 51716 36136 51772
rect 36184 51770 36240 51772
rect 36288 51770 36344 51772
rect 36184 51718 36196 51770
rect 36196 51718 36240 51770
rect 36288 51718 36320 51770
rect 36320 51718 36344 51770
rect 36184 51716 36240 51718
rect 36288 51716 36344 51718
rect 36392 51716 36448 51772
rect 38892 51996 38948 52052
rect 39228 52556 39284 52612
rect 38668 51548 38724 51604
rect 36540 51324 36596 51380
rect 38444 51378 38500 51380
rect 38444 51326 38446 51378
rect 38446 51326 38498 51378
rect 38498 51326 38500 51378
rect 38444 51324 38500 51326
rect 39116 51324 39172 51380
rect 39564 51996 39620 52052
rect 39564 51436 39620 51492
rect 42588 54460 42644 54516
rect 41468 53788 41524 53844
rect 40908 53228 40964 53284
rect 41132 52946 41188 52948
rect 41132 52894 41134 52946
rect 41134 52894 41186 52946
rect 41186 52894 41188 52946
rect 41132 52892 41188 52894
rect 40124 52556 40180 52612
rect 40268 52500 40324 52556
rect 40372 52554 40428 52556
rect 40476 52554 40532 52556
rect 40372 52502 40396 52554
rect 40396 52502 40428 52554
rect 40476 52502 40520 52554
rect 40520 52502 40532 52554
rect 40372 52500 40428 52502
rect 40476 52500 40532 52502
rect 40580 52500 40636 52556
rect 40684 52554 40740 52556
rect 40788 52554 40844 52556
rect 40684 52502 40696 52554
rect 40696 52502 40740 52554
rect 40788 52502 40820 52554
rect 40820 52502 40844 52554
rect 40684 52500 40740 52502
rect 40788 52500 40844 52502
rect 40892 52500 40948 52556
rect 41468 52444 41524 52500
rect 41692 52668 41748 52724
rect 41916 53004 41972 53060
rect 41580 52332 41636 52388
rect 39676 51548 39732 51604
rect 40124 51548 40180 51604
rect 39900 50594 39956 50596
rect 39900 50542 39902 50594
rect 39902 50542 39954 50594
rect 39954 50542 39956 50594
rect 39900 50540 39956 50542
rect 33740 50428 33796 50484
rect 32508 47180 32564 47236
rect 33628 47234 33684 47236
rect 33628 47182 33630 47234
rect 33630 47182 33682 47234
rect 33682 47182 33684 47234
rect 33628 47180 33684 47182
rect 33292 46674 33348 46676
rect 33292 46622 33294 46674
rect 33294 46622 33346 46674
rect 33346 46622 33348 46674
rect 33292 46620 33348 46622
rect 32172 46060 32228 46116
rect 30604 44380 30660 44436
rect 29260 43538 29316 43540
rect 29260 43486 29262 43538
rect 29262 43486 29314 43538
rect 29314 43486 29316 43538
rect 29260 43484 29316 43486
rect 29932 43538 29988 43540
rect 29932 43486 29934 43538
rect 29934 43486 29986 43538
rect 29986 43486 29988 43538
rect 29932 43484 29988 43486
rect 31268 44660 31324 44716
rect 31372 44714 31428 44716
rect 31476 44714 31532 44716
rect 31372 44662 31396 44714
rect 31396 44662 31428 44714
rect 31476 44662 31520 44714
rect 31520 44662 31532 44714
rect 31372 44660 31428 44662
rect 31476 44660 31532 44662
rect 31580 44660 31636 44716
rect 31684 44714 31740 44716
rect 31788 44714 31844 44716
rect 31684 44662 31696 44714
rect 31696 44662 31740 44714
rect 31788 44662 31820 44714
rect 31820 44662 31844 44714
rect 31684 44660 31740 44662
rect 31788 44660 31844 44662
rect 31892 44660 31948 44716
rect 31052 44434 31108 44436
rect 31052 44382 31054 44434
rect 31054 44382 31106 44434
rect 31106 44382 31108 44434
rect 31052 44380 31108 44382
rect 31948 43708 32004 43764
rect 29596 43314 29652 43316
rect 29596 43262 29598 43314
rect 29598 43262 29650 43314
rect 29650 43262 29652 43314
rect 29596 43260 29652 43262
rect 28588 42812 28644 42868
rect 29372 42866 29428 42868
rect 29372 42814 29374 42866
rect 29374 42814 29426 42866
rect 29426 42814 29428 42866
rect 29372 42812 29428 42814
rect 22268 39956 22324 40012
rect 22372 40010 22428 40012
rect 22476 40010 22532 40012
rect 22372 39958 22396 40010
rect 22396 39958 22428 40010
rect 22476 39958 22520 40010
rect 22520 39958 22532 40010
rect 22372 39956 22428 39958
rect 22476 39956 22532 39958
rect 22580 39956 22636 40012
rect 22684 40010 22740 40012
rect 22788 40010 22844 40012
rect 22684 39958 22696 40010
rect 22696 39958 22740 40010
rect 22788 39958 22820 40010
rect 22820 39958 22844 40010
rect 22684 39956 22740 39958
rect 22788 39956 22844 39958
rect 22892 39956 22948 40012
rect 28252 40236 28308 40292
rect 26796 40124 26852 40180
rect 26768 39172 26824 39228
rect 26872 39226 26928 39228
rect 26976 39226 27032 39228
rect 26872 39174 26896 39226
rect 26896 39174 26928 39226
rect 26976 39174 27020 39226
rect 27020 39174 27032 39226
rect 26872 39172 26928 39174
rect 26976 39172 27032 39174
rect 27080 39172 27136 39228
rect 27184 39226 27240 39228
rect 27288 39226 27344 39228
rect 27184 39174 27196 39226
rect 27196 39174 27240 39226
rect 27288 39174 27320 39226
rect 27320 39174 27344 39226
rect 27184 39172 27240 39174
rect 27288 39172 27344 39174
rect 27392 39172 27448 39228
rect 16156 36316 16212 36372
rect 15372 35698 15428 35700
rect 15372 35646 15374 35698
rect 15374 35646 15426 35698
rect 15426 35646 15428 35698
rect 15372 35644 15428 35646
rect 17276 38220 17332 38276
rect 20188 37772 20244 37828
rect 17768 37604 17824 37660
rect 17872 37658 17928 37660
rect 17976 37658 18032 37660
rect 17872 37606 17896 37658
rect 17896 37606 17928 37658
rect 17976 37606 18020 37658
rect 18020 37606 18032 37658
rect 17872 37604 17928 37606
rect 17976 37604 18032 37606
rect 18080 37604 18136 37660
rect 18184 37658 18240 37660
rect 18288 37658 18344 37660
rect 18184 37606 18196 37658
rect 18196 37606 18240 37658
rect 18288 37606 18320 37658
rect 18320 37606 18344 37658
rect 18184 37604 18240 37606
rect 18288 37604 18344 37606
rect 18392 37604 18448 37660
rect 18396 37490 18452 37492
rect 18396 37438 18398 37490
rect 18398 37438 18450 37490
rect 18450 37438 18452 37490
rect 18396 37436 18452 37438
rect 19740 37436 19796 37492
rect 19628 36876 19684 36932
rect 17612 36652 17668 36708
rect 17500 36316 17556 36372
rect 18620 36652 18676 36708
rect 18508 36370 18564 36372
rect 18508 36318 18510 36370
rect 18510 36318 18562 36370
rect 18562 36318 18564 36370
rect 18508 36316 18564 36318
rect 17768 36036 17824 36092
rect 17872 36090 17928 36092
rect 17976 36090 18032 36092
rect 17872 36038 17896 36090
rect 17896 36038 17928 36090
rect 17976 36038 18020 36090
rect 18020 36038 18032 36090
rect 17872 36036 17928 36038
rect 17976 36036 18032 36038
rect 18080 36036 18136 36092
rect 18184 36090 18240 36092
rect 18288 36090 18344 36092
rect 18184 36038 18196 36090
rect 18196 36038 18240 36090
rect 18288 36038 18320 36090
rect 18320 36038 18344 36090
rect 18184 36036 18240 36038
rect 18288 36036 18344 36038
rect 18392 36036 18448 36092
rect 18956 36706 19012 36708
rect 18956 36654 18958 36706
rect 18958 36654 19010 36706
rect 19010 36654 19012 36706
rect 18956 36652 19012 36654
rect 20748 37996 20804 38052
rect 20524 37660 20580 37716
rect 20524 36876 20580 36932
rect 20748 36988 20804 37044
rect 30380 40796 30436 40852
rect 30156 40460 30212 40516
rect 28924 40402 28980 40404
rect 28924 40350 28926 40402
rect 28926 40350 28978 40402
rect 28978 40350 28980 40402
rect 28924 40348 28980 40350
rect 29596 40402 29652 40404
rect 29596 40350 29598 40402
rect 29598 40350 29650 40402
rect 29650 40350 29652 40402
rect 29596 40348 29652 40350
rect 31948 43372 32004 43428
rect 32060 43596 32116 43652
rect 31724 43260 31780 43316
rect 31268 43092 31324 43148
rect 31372 43146 31428 43148
rect 31476 43146 31532 43148
rect 31372 43094 31396 43146
rect 31396 43094 31428 43146
rect 31476 43094 31520 43146
rect 31520 43094 31532 43146
rect 31372 43092 31428 43094
rect 31476 43092 31532 43094
rect 31580 43092 31636 43148
rect 31684 43146 31740 43148
rect 31788 43146 31844 43148
rect 31684 43094 31696 43146
rect 31696 43094 31740 43146
rect 31788 43094 31820 43146
rect 31820 43094 31844 43146
rect 31684 43092 31740 43094
rect 31788 43092 31844 43094
rect 31892 43092 31948 43148
rect 31612 42924 31668 42980
rect 30604 40460 30660 40516
rect 30828 42812 30884 42868
rect 29036 40236 29092 40292
rect 29260 40178 29316 40180
rect 29260 40126 29262 40178
rect 29262 40126 29314 40178
rect 29314 40126 29316 40178
rect 29260 40124 29316 40126
rect 22268 38388 22324 38444
rect 22372 38442 22428 38444
rect 22476 38442 22532 38444
rect 22372 38390 22396 38442
rect 22396 38390 22428 38442
rect 22476 38390 22520 38442
rect 22520 38390 22532 38442
rect 22372 38388 22428 38390
rect 22476 38388 22532 38390
rect 22580 38388 22636 38444
rect 22684 38442 22740 38444
rect 22788 38442 22844 38444
rect 22684 38390 22696 38442
rect 22696 38390 22740 38442
rect 22788 38390 22820 38442
rect 22820 38390 22844 38442
rect 22684 38388 22740 38390
rect 22788 38388 22844 38390
rect 22892 38388 22948 38444
rect 21868 38050 21924 38052
rect 21868 37998 21870 38050
rect 21870 37998 21922 38050
rect 21922 37998 21924 38050
rect 21868 37996 21924 37998
rect 21644 37660 21700 37716
rect 21308 37266 21364 37268
rect 21308 37214 21310 37266
rect 21310 37214 21362 37266
rect 21362 37214 21364 37266
rect 21308 37212 21364 37214
rect 21084 36988 21140 37044
rect 25004 37826 25060 37828
rect 25004 37774 25006 37826
rect 25006 37774 25058 37826
rect 25058 37774 25060 37826
rect 25004 37772 25060 37774
rect 25004 37212 25060 37268
rect 26768 37604 26824 37660
rect 26872 37658 26928 37660
rect 26976 37658 27032 37660
rect 26872 37606 26896 37658
rect 26896 37606 26928 37658
rect 26976 37606 27020 37658
rect 27020 37606 27032 37658
rect 26872 37604 26928 37606
rect 26976 37604 27032 37606
rect 27080 37604 27136 37660
rect 27184 37658 27240 37660
rect 27288 37658 27344 37660
rect 27184 37606 27196 37658
rect 27196 37606 27240 37658
rect 27288 37606 27320 37658
rect 27320 37606 27344 37658
rect 27184 37604 27240 37606
rect 27288 37604 27344 37606
rect 27392 37604 27448 37660
rect 24220 36988 24276 37044
rect 22268 36820 22324 36876
rect 22372 36874 22428 36876
rect 22476 36874 22532 36876
rect 22372 36822 22396 36874
rect 22396 36822 22428 36874
rect 22476 36822 22520 36874
rect 22520 36822 22532 36874
rect 22372 36820 22428 36822
rect 22476 36820 22532 36822
rect 22580 36820 22636 36876
rect 22684 36874 22740 36876
rect 22788 36874 22844 36876
rect 22684 36822 22696 36874
rect 22696 36822 22740 36874
rect 22788 36822 22820 36874
rect 22820 36822 22844 36874
rect 22684 36820 22740 36822
rect 22788 36820 22844 36822
rect 22892 36820 22948 36876
rect 20748 36652 20804 36708
rect 16716 35644 16772 35700
rect 13268 35252 13324 35308
rect 13372 35306 13428 35308
rect 13476 35306 13532 35308
rect 13372 35254 13396 35306
rect 13396 35254 13428 35306
rect 13476 35254 13520 35306
rect 13520 35254 13532 35306
rect 13372 35252 13428 35254
rect 13476 35252 13532 35254
rect 13580 35252 13636 35308
rect 13684 35306 13740 35308
rect 13788 35306 13844 35308
rect 13684 35254 13696 35306
rect 13696 35254 13740 35306
rect 13788 35254 13820 35306
rect 13820 35254 13844 35306
rect 13684 35252 13740 35254
rect 13788 35252 13844 35254
rect 13892 35252 13948 35308
rect 12012 34188 12068 34244
rect 14028 34242 14084 34244
rect 14028 34190 14030 34242
rect 14030 34190 14082 34242
rect 14082 34190 14084 34242
rect 14028 34188 14084 34190
rect 12012 33628 12068 33684
rect 13244 34076 13300 34132
rect 13268 33684 13324 33740
rect 13372 33738 13428 33740
rect 13476 33738 13532 33740
rect 13372 33686 13396 33738
rect 13396 33686 13428 33738
rect 13476 33686 13520 33738
rect 13520 33686 13532 33738
rect 13372 33684 13428 33686
rect 13476 33684 13532 33686
rect 13580 33684 13636 33740
rect 13684 33738 13740 33740
rect 13788 33738 13844 33740
rect 13684 33686 13696 33738
rect 13696 33686 13740 33738
rect 13788 33686 13820 33738
rect 13820 33686 13844 33738
rect 13684 33684 13740 33686
rect 13788 33684 13844 33686
rect 13892 33684 13948 33740
rect 17768 34468 17824 34524
rect 17872 34522 17928 34524
rect 17976 34522 18032 34524
rect 17872 34470 17896 34522
rect 17896 34470 17928 34522
rect 17976 34470 18020 34522
rect 18020 34470 18032 34522
rect 17872 34468 17928 34470
rect 17976 34468 18032 34470
rect 18080 34468 18136 34524
rect 18184 34522 18240 34524
rect 18288 34522 18344 34524
rect 18184 34470 18196 34522
rect 18196 34470 18240 34522
rect 18288 34470 18320 34522
rect 18320 34470 18344 34522
rect 18184 34468 18240 34470
rect 18288 34468 18344 34470
rect 18392 34468 18448 34524
rect 19516 33964 19572 34020
rect 14588 33458 14644 33460
rect 14588 33406 14590 33458
rect 14590 33406 14642 33458
rect 14642 33406 14644 33458
rect 14588 33404 14644 33406
rect 19068 33458 19124 33460
rect 19068 33406 19070 33458
rect 19070 33406 19122 33458
rect 19122 33406 19124 33458
rect 19068 33404 19124 33406
rect 15372 33292 15428 33348
rect 12348 32674 12404 32676
rect 12348 32622 12350 32674
rect 12350 32622 12402 32674
rect 12402 32622 12404 32674
rect 12348 32620 12404 32622
rect 14588 32284 14644 32340
rect 13268 32116 13324 32172
rect 13372 32170 13428 32172
rect 13476 32170 13532 32172
rect 13372 32118 13396 32170
rect 13396 32118 13428 32170
rect 13476 32118 13520 32170
rect 13520 32118 13532 32170
rect 13372 32116 13428 32118
rect 13476 32116 13532 32118
rect 13580 32116 13636 32172
rect 13684 32170 13740 32172
rect 13788 32170 13844 32172
rect 13684 32118 13696 32170
rect 13696 32118 13740 32170
rect 13788 32118 13820 32170
rect 13820 32118 13844 32170
rect 13684 32116 13740 32118
rect 13788 32116 13844 32118
rect 13892 32116 13948 32172
rect 15148 32674 15204 32676
rect 15148 32622 15150 32674
rect 15150 32622 15202 32674
rect 15202 32622 15204 32674
rect 15148 32620 15204 32622
rect 13268 30548 13324 30604
rect 13372 30602 13428 30604
rect 13476 30602 13532 30604
rect 13372 30550 13396 30602
rect 13396 30550 13428 30602
rect 13476 30550 13520 30602
rect 13520 30550 13532 30602
rect 13372 30548 13428 30550
rect 13476 30548 13532 30550
rect 13580 30548 13636 30604
rect 13684 30602 13740 30604
rect 13788 30602 13844 30604
rect 13684 30550 13696 30602
rect 13696 30550 13740 30602
rect 13788 30550 13820 30602
rect 13820 30550 13844 30602
rect 13684 30548 13740 30550
rect 13788 30548 13844 30550
rect 13892 30548 13948 30604
rect 14700 30098 14756 30100
rect 14700 30046 14702 30098
rect 14702 30046 14754 30098
rect 14754 30046 14756 30098
rect 14700 30044 14756 30046
rect 12012 29986 12068 29988
rect 12012 29934 12014 29986
rect 12014 29934 12066 29986
rect 12066 29934 12068 29986
rect 12012 29932 12068 29934
rect 13020 29314 13076 29316
rect 13020 29262 13022 29314
rect 13022 29262 13074 29314
rect 13074 29262 13076 29314
rect 13020 29260 13076 29262
rect 13268 28980 13324 29036
rect 13372 29034 13428 29036
rect 13476 29034 13532 29036
rect 13372 28982 13396 29034
rect 13396 28982 13428 29034
rect 13476 28982 13520 29034
rect 13520 28982 13532 29034
rect 13372 28980 13428 28982
rect 13476 28980 13532 28982
rect 13580 28980 13636 29036
rect 13684 29034 13740 29036
rect 13788 29034 13844 29036
rect 13684 28982 13696 29034
rect 13696 28982 13740 29034
rect 13788 28982 13820 29034
rect 13820 28982 13844 29034
rect 13684 28980 13740 28982
rect 13788 28980 13844 28982
rect 13892 28980 13948 29036
rect 13020 28028 13076 28084
rect 12236 27858 12292 27860
rect 12236 27806 12238 27858
rect 12238 27806 12290 27858
rect 12290 27806 12292 27858
rect 12236 27804 12292 27806
rect 13804 28028 13860 28084
rect 10556 24892 10612 24948
rect 10780 24108 10836 24164
rect 11116 25394 11172 25396
rect 11116 25342 11118 25394
rect 11118 25342 11170 25394
rect 11170 25342 11172 25394
rect 11116 25340 11172 25342
rect 13268 27412 13324 27468
rect 13372 27466 13428 27468
rect 13476 27466 13532 27468
rect 13372 27414 13396 27466
rect 13396 27414 13428 27466
rect 13476 27414 13520 27466
rect 13520 27414 13532 27466
rect 13372 27412 13428 27414
rect 13476 27412 13532 27414
rect 13580 27412 13636 27468
rect 13684 27466 13740 27468
rect 13788 27466 13844 27468
rect 13684 27414 13696 27466
rect 13696 27414 13740 27466
rect 13788 27414 13820 27466
rect 13820 27414 13844 27466
rect 13684 27412 13740 27414
rect 13788 27412 13844 27414
rect 13892 27412 13948 27468
rect 16156 32620 16212 32676
rect 15484 32284 15540 32340
rect 20300 35810 20356 35812
rect 20300 35758 20302 35810
rect 20302 35758 20354 35810
rect 20354 35758 20356 35810
rect 20300 35756 20356 35758
rect 22268 35252 22324 35308
rect 22372 35306 22428 35308
rect 22476 35306 22532 35308
rect 22372 35254 22396 35306
rect 22396 35254 22428 35306
rect 22476 35254 22520 35306
rect 22520 35254 22532 35306
rect 22372 35252 22428 35254
rect 22476 35252 22532 35254
rect 22580 35252 22636 35308
rect 22684 35306 22740 35308
rect 22788 35306 22844 35308
rect 22684 35254 22696 35306
rect 22696 35254 22740 35306
rect 22788 35254 22820 35306
rect 22820 35254 22844 35306
rect 22684 35252 22740 35254
rect 22788 35252 22844 35254
rect 22892 35252 22948 35308
rect 20972 34748 21028 34804
rect 28364 38050 28420 38052
rect 28364 37998 28366 38050
rect 28366 37998 28418 38050
rect 28418 37998 28420 38050
rect 28364 37996 28420 37998
rect 28476 37938 28532 37940
rect 28476 37886 28478 37938
rect 28478 37886 28530 37938
rect 28530 37886 28532 37938
rect 28476 37884 28532 37886
rect 29932 38108 29988 38164
rect 31164 42866 31220 42868
rect 31164 42814 31166 42866
rect 31166 42814 31218 42866
rect 31218 42814 31220 42866
rect 31164 42812 31220 42814
rect 31268 41524 31324 41580
rect 31372 41578 31428 41580
rect 31476 41578 31532 41580
rect 31372 41526 31396 41578
rect 31396 41526 31428 41578
rect 31476 41526 31520 41578
rect 31520 41526 31532 41578
rect 31372 41524 31428 41526
rect 31476 41524 31532 41526
rect 31580 41524 31636 41580
rect 31684 41578 31740 41580
rect 31788 41578 31844 41580
rect 31684 41526 31696 41578
rect 31696 41526 31740 41578
rect 31788 41526 31820 41578
rect 31820 41526 31844 41578
rect 31684 41524 31740 41526
rect 31788 41524 31844 41526
rect 31892 41524 31948 41580
rect 30940 40514 30996 40516
rect 30940 40462 30942 40514
rect 30942 40462 30994 40514
rect 30994 40462 30996 40514
rect 30940 40460 30996 40462
rect 31612 40796 31668 40852
rect 35768 50148 35824 50204
rect 35872 50202 35928 50204
rect 35976 50202 36032 50204
rect 35872 50150 35896 50202
rect 35896 50150 35928 50202
rect 35976 50150 36020 50202
rect 36020 50150 36032 50202
rect 35872 50148 35928 50150
rect 35976 50148 36032 50150
rect 36080 50148 36136 50204
rect 36184 50202 36240 50204
rect 36288 50202 36344 50204
rect 36184 50150 36196 50202
rect 36196 50150 36240 50202
rect 36288 50150 36320 50202
rect 36320 50150 36344 50202
rect 36184 50148 36240 50150
rect 36288 50148 36344 50150
rect 36392 50148 36448 50204
rect 37660 49922 37716 49924
rect 37660 49870 37662 49922
rect 37662 49870 37714 49922
rect 37714 49870 37716 49922
rect 37660 49868 37716 49870
rect 38444 49810 38500 49812
rect 38444 49758 38446 49810
rect 38446 49758 38498 49810
rect 38498 49758 38500 49810
rect 38444 49756 38500 49758
rect 39004 49698 39060 49700
rect 39004 49646 39006 49698
rect 39006 49646 39058 49698
rect 39058 49646 39060 49698
rect 39004 49644 39060 49646
rect 35532 49532 35588 49588
rect 35084 49196 35140 49252
rect 34748 47516 34804 47572
rect 34636 47292 34692 47348
rect 33964 46620 34020 46676
rect 34524 46620 34580 46676
rect 33740 45778 33796 45780
rect 33740 45726 33742 45778
rect 33742 45726 33794 45778
rect 33794 45726 33796 45778
rect 33740 45724 33796 45726
rect 33068 43650 33124 43652
rect 33068 43598 33070 43650
rect 33070 43598 33122 43650
rect 33122 43598 33124 43650
rect 33068 43596 33124 43598
rect 33740 43820 33796 43876
rect 32508 43426 32564 43428
rect 32508 43374 32510 43426
rect 32510 43374 32562 43426
rect 32562 43374 32564 43426
rect 32508 43372 32564 43374
rect 34188 42924 34244 42980
rect 32172 40796 32228 40852
rect 33292 40796 33348 40852
rect 33404 40908 33460 40964
rect 31268 39956 31324 40012
rect 31372 40010 31428 40012
rect 31476 40010 31532 40012
rect 31372 39958 31396 40010
rect 31396 39958 31428 40010
rect 31476 39958 31520 40010
rect 31520 39958 31532 40010
rect 31372 39956 31428 39958
rect 31476 39956 31532 39958
rect 31580 39956 31636 40012
rect 31684 40010 31740 40012
rect 31788 40010 31844 40012
rect 31684 39958 31696 40010
rect 31696 39958 31740 40010
rect 31788 39958 31820 40010
rect 31820 39958 31844 40010
rect 31684 39956 31740 39958
rect 31788 39956 31844 39958
rect 31892 39956 31948 40012
rect 31836 39788 31892 39844
rect 34972 46508 35028 46564
rect 35756 49138 35812 49140
rect 35756 49086 35758 49138
rect 35758 49086 35810 49138
rect 35810 49086 35812 49138
rect 35756 49084 35812 49086
rect 38668 49084 38724 49140
rect 35768 48580 35824 48636
rect 35872 48634 35928 48636
rect 35976 48634 36032 48636
rect 35872 48582 35896 48634
rect 35896 48582 35928 48634
rect 35976 48582 36020 48634
rect 36020 48582 36032 48634
rect 35872 48580 35928 48582
rect 35976 48580 36032 48582
rect 36080 48580 36136 48636
rect 36184 48634 36240 48636
rect 36288 48634 36344 48636
rect 36184 48582 36196 48634
rect 36196 48582 36240 48634
rect 36288 48582 36320 48634
rect 36320 48582 36344 48634
rect 36184 48580 36240 48582
rect 36288 48580 36344 48582
rect 36392 48580 36448 48636
rect 35644 47516 35700 47572
rect 35084 45724 35140 45780
rect 35084 44380 35140 44436
rect 34860 44156 34916 44212
rect 35308 47292 35364 47348
rect 40908 51490 40964 51492
rect 40908 51438 40910 51490
rect 40910 51438 40962 51490
rect 40962 51438 40964 51490
rect 40908 51436 40964 51438
rect 40268 50932 40324 50988
rect 40372 50986 40428 50988
rect 40476 50986 40532 50988
rect 40372 50934 40396 50986
rect 40396 50934 40428 50986
rect 40476 50934 40520 50986
rect 40520 50934 40532 50986
rect 40372 50932 40428 50934
rect 40476 50932 40532 50934
rect 40580 50932 40636 50988
rect 40684 50986 40740 50988
rect 40788 50986 40844 50988
rect 40684 50934 40696 50986
rect 40696 50934 40740 50986
rect 40788 50934 40820 50986
rect 40820 50934 40844 50986
rect 40684 50932 40740 50934
rect 40788 50932 40844 50934
rect 40892 50932 40948 50988
rect 39900 49084 39956 49140
rect 39900 48466 39956 48468
rect 39900 48414 39902 48466
rect 39902 48414 39954 48466
rect 39954 48414 39956 48466
rect 39900 48412 39956 48414
rect 40012 47964 40068 48020
rect 37660 47346 37716 47348
rect 37660 47294 37662 47346
rect 37662 47294 37714 47346
rect 37714 47294 37716 47346
rect 37660 47292 37716 47294
rect 39116 47292 39172 47348
rect 35768 47012 35824 47068
rect 35872 47066 35928 47068
rect 35976 47066 36032 47068
rect 35872 47014 35896 47066
rect 35896 47014 35928 47066
rect 35976 47014 36020 47066
rect 36020 47014 36032 47066
rect 35872 47012 35928 47014
rect 35976 47012 36032 47014
rect 36080 47012 36136 47068
rect 36184 47066 36240 47068
rect 36288 47066 36344 47068
rect 36184 47014 36196 47066
rect 36196 47014 36240 47066
rect 36288 47014 36320 47066
rect 36320 47014 36344 47066
rect 36184 47012 36240 47014
rect 36288 47012 36344 47014
rect 36392 47012 36448 47068
rect 38556 46956 38612 47012
rect 35644 46674 35700 46676
rect 35644 46622 35646 46674
rect 35646 46622 35698 46674
rect 35698 46622 35700 46674
rect 35644 46620 35700 46622
rect 36764 46060 36820 46116
rect 35768 45444 35824 45500
rect 35872 45498 35928 45500
rect 35976 45498 36032 45500
rect 35872 45446 35896 45498
rect 35896 45446 35928 45498
rect 35976 45446 36020 45498
rect 36020 45446 36032 45498
rect 35872 45444 35928 45446
rect 35976 45444 36032 45446
rect 36080 45444 36136 45500
rect 36184 45498 36240 45500
rect 36288 45498 36344 45500
rect 36184 45446 36196 45498
rect 36196 45446 36240 45498
rect 36288 45446 36320 45498
rect 36320 45446 36344 45498
rect 36184 45444 36240 45446
rect 36288 45444 36344 45446
rect 36392 45444 36448 45500
rect 35980 44434 36036 44436
rect 35980 44382 35982 44434
rect 35982 44382 36034 44434
rect 36034 44382 36036 44434
rect 35980 44380 36036 44382
rect 38220 46732 38276 46788
rect 39004 46060 39060 46116
rect 38556 45778 38612 45780
rect 38556 45726 38558 45778
rect 38558 45726 38610 45778
rect 38610 45726 38612 45778
rect 38556 45724 38612 45726
rect 35532 44156 35588 44212
rect 34188 40962 34244 40964
rect 34188 40910 34190 40962
rect 34190 40910 34242 40962
rect 34242 40910 34244 40962
rect 34188 40908 34244 40910
rect 33740 40572 33796 40628
rect 33068 39788 33124 39844
rect 35196 43538 35252 43540
rect 35196 43486 35198 43538
rect 35198 43486 35250 43538
rect 35250 43486 35252 43538
rect 35196 43484 35252 43486
rect 35084 42978 35140 42980
rect 35084 42926 35086 42978
rect 35086 42926 35138 42978
rect 35138 42926 35140 42978
rect 35084 42924 35140 42926
rect 35768 43876 35824 43932
rect 35872 43930 35928 43932
rect 35976 43930 36032 43932
rect 35872 43878 35896 43930
rect 35896 43878 35928 43930
rect 35976 43878 36020 43930
rect 36020 43878 36032 43930
rect 35872 43876 35928 43878
rect 35976 43876 36032 43878
rect 36080 43876 36136 43932
rect 36184 43930 36240 43932
rect 36288 43930 36344 43932
rect 36184 43878 36196 43930
rect 36196 43878 36240 43930
rect 36288 43878 36320 43930
rect 36320 43878 36344 43930
rect 36184 43876 36240 43878
rect 36288 43876 36344 43878
rect 36392 43876 36448 43932
rect 38444 45612 38500 45668
rect 40012 46396 40068 46452
rect 39340 45724 39396 45780
rect 38556 45388 38612 45444
rect 35308 41186 35364 41188
rect 35308 41134 35310 41186
rect 35310 41134 35362 41186
rect 35362 41134 35364 41186
rect 35308 41132 35364 41134
rect 34972 40908 35028 40964
rect 34860 40460 34916 40516
rect 35196 40796 35252 40852
rect 35196 39004 35252 39060
rect 31268 38388 31324 38444
rect 31372 38442 31428 38444
rect 31476 38442 31532 38444
rect 31372 38390 31396 38442
rect 31396 38390 31428 38442
rect 31476 38390 31520 38442
rect 31520 38390 31532 38442
rect 31372 38388 31428 38390
rect 31476 38388 31532 38390
rect 31580 38388 31636 38444
rect 31684 38442 31740 38444
rect 31788 38442 31844 38444
rect 31684 38390 31696 38442
rect 31696 38390 31740 38442
rect 31788 38390 31820 38442
rect 31820 38390 31844 38442
rect 31684 38388 31740 38390
rect 31788 38388 31844 38390
rect 31892 38388 31948 38444
rect 33404 38220 33460 38276
rect 30156 37996 30212 38052
rect 32956 37938 33012 37940
rect 32956 37886 32958 37938
rect 32958 37886 33010 37938
rect 33010 37886 33012 37938
rect 32956 37884 33012 37886
rect 29148 37324 29204 37380
rect 29820 37324 29876 37380
rect 27692 37212 27748 37268
rect 29708 37266 29764 37268
rect 29708 37214 29710 37266
rect 29710 37214 29762 37266
rect 29762 37214 29764 37266
rect 29708 37212 29764 37214
rect 29148 36988 29204 37044
rect 26768 36036 26824 36092
rect 26872 36090 26928 36092
rect 26976 36090 27032 36092
rect 26872 36038 26896 36090
rect 26896 36038 26928 36090
rect 26976 36038 27020 36090
rect 27020 36038 27032 36090
rect 26872 36036 26928 36038
rect 26976 36036 27032 36038
rect 27080 36036 27136 36092
rect 27184 36090 27240 36092
rect 27288 36090 27344 36092
rect 27184 36038 27196 36090
rect 27196 36038 27240 36090
rect 27288 36038 27320 36090
rect 27320 36038 27344 36090
rect 27184 36036 27240 36038
rect 27288 36036 27344 36038
rect 27392 36036 27448 36092
rect 24892 34802 24948 34804
rect 24892 34750 24894 34802
rect 24894 34750 24946 34802
rect 24946 34750 24948 34802
rect 24892 34748 24948 34750
rect 19628 33404 19684 33460
rect 17768 32900 17824 32956
rect 17872 32954 17928 32956
rect 17976 32954 18032 32956
rect 17872 32902 17896 32954
rect 17896 32902 17928 32954
rect 17976 32902 18020 32954
rect 18020 32902 18032 32954
rect 17872 32900 17928 32902
rect 17976 32900 18032 32902
rect 18080 32900 18136 32956
rect 18184 32954 18240 32956
rect 18288 32954 18344 32956
rect 18184 32902 18196 32954
rect 18196 32902 18240 32954
rect 18288 32902 18320 32954
rect 18320 32902 18344 32954
rect 18184 32900 18240 32902
rect 18288 32900 18344 32902
rect 18392 32900 18448 32956
rect 20300 32674 20356 32676
rect 20300 32622 20302 32674
rect 20302 32622 20354 32674
rect 20354 32622 20356 32674
rect 20300 32620 20356 32622
rect 22268 33684 22324 33740
rect 22372 33738 22428 33740
rect 22476 33738 22532 33740
rect 22372 33686 22396 33738
rect 22396 33686 22428 33738
rect 22476 33686 22520 33738
rect 22520 33686 22532 33738
rect 22372 33684 22428 33686
rect 22476 33684 22532 33686
rect 22580 33684 22636 33740
rect 22684 33738 22740 33740
rect 22788 33738 22844 33740
rect 22684 33686 22696 33738
rect 22696 33686 22740 33738
rect 22788 33686 22820 33738
rect 22820 33686 22844 33738
rect 22684 33684 22740 33686
rect 22788 33684 22844 33686
rect 22892 33684 22948 33740
rect 23436 32674 23492 32676
rect 23436 32622 23438 32674
rect 23438 32622 23490 32674
rect 23490 32622 23492 32674
rect 23436 32620 23492 32622
rect 26768 34468 26824 34524
rect 26872 34522 26928 34524
rect 26976 34522 27032 34524
rect 26872 34470 26896 34522
rect 26896 34470 26928 34522
rect 26976 34470 27020 34522
rect 27020 34470 27032 34522
rect 26872 34468 26928 34470
rect 26976 34468 27032 34470
rect 27080 34468 27136 34524
rect 27184 34522 27240 34524
rect 27288 34522 27344 34524
rect 27184 34470 27196 34522
rect 27196 34470 27240 34522
rect 27288 34470 27320 34522
rect 27320 34470 27344 34522
rect 27184 34468 27240 34470
rect 27288 34468 27344 34470
rect 27392 34468 27448 34524
rect 26768 32900 26824 32956
rect 26872 32954 26928 32956
rect 26976 32954 27032 32956
rect 26872 32902 26896 32954
rect 26896 32902 26928 32954
rect 26976 32902 27020 32954
rect 27020 32902 27032 32954
rect 26872 32900 26928 32902
rect 26976 32900 27032 32902
rect 27080 32900 27136 32956
rect 27184 32954 27240 32956
rect 27288 32954 27344 32956
rect 27184 32902 27196 32954
rect 27196 32902 27240 32954
rect 27288 32902 27320 32954
rect 27320 32902 27344 32954
rect 27184 32900 27240 32902
rect 27288 32900 27344 32902
rect 27392 32900 27448 32956
rect 20412 32284 20468 32340
rect 24220 32338 24276 32340
rect 24220 32286 24222 32338
rect 24222 32286 24274 32338
rect 24274 32286 24276 32338
rect 24220 32284 24276 32286
rect 22268 32116 22324 32172
rect 22372 32170 22428 32172
rect 22476 32170 22532 32172
rect 22372 32118 22396 32170
rect 22396 32118 22428 32170
rect 22476 32118 22520 32170
rect 22520 32118 22532 32170
rect 22372 32116 22428 32118
rect 22476 32116 22532 32118
rect 22580 32116 22636 32172
rect 22684 32170 22740 32172
rect 22788 32170 22844 32172
rect 22684 32118 22696 32170
rect 22696 32118 22740 32170
rect 22788 32118 22820 32170
rect 22820 32118 22844 32170
rect 22684 32116 22740 32118
rect 22788 32116 22844 32118
rect 22892 32116 22948 32172
rect 16716 31612 16772 31668
rect 18060 31666 18116 31668
rect 18060 31614 18062 31666
rect 18062 31614 18114 31666
rect 18114 31614 18116 31666
rect 18060 31612 18116 31614
rect 17500 31554 17556 31556
rect 17500 31502 17502 31554
rect 17502 31502 17554 31554
rect 17554 31502 17556 31554
rect 17500 31500 17556 31502
rect 15932 30322 15988 30324
rect 15932 30270 15934 30322
rect 15934 30270 15986 30322
rect 15986 30270 15988 30322
rect 15932 30268 15988 30270
rect 16828 30268 16884 30324
rect 16268 30098 16324 30100
rect 16268 30046 16270 30098
rect 16270 30046 16322 30098
rect 16322 30046 16324 30098
rect 16268 30044 16324 30046
rect 16156 29260 16212 29316
rect 16940 28812 16996 28868
rect 15148 27804 15204 27860
rect 17388 28028 17444 28084
rect 15148 27132 15204 27188
rect 18396 31554 18452 31556
rect 18396 31502 18398 31554
rect 18398 31502 18450 31554
rect 18450 31502 18452 31554
rect 18396 31500 18452 31502
rect 19964 31500 20020 31556
rect 17768 31332 17824 31388
rect 17872 31386 17928 31388
rect 17976 31386 18032 31388
rect 17872 31334 17896 31386
rect 17896 31334 17928 31386
rect 17976 31334 18020 31386
rect 18020 31334 18032 31386
rect 17872 31332 17928 31334
rect 17976 31332 18032 31334
rect 18080 31332 18136 31388
rect 18184 31386 18240 31388
rect 18288 31386 18344 31388
rect 18184 31334 18196 31386
rect 18196 31334 18240 31386
rect 18288 31334 18320 31386
rect 18320 31334 18344 31386
rect 18184 31332 18240 31334
rect 18288 31332 18344 31334
rect 18392 31332 18448 31388
rect 20412 30994 20468 30996
rect 20412 30942 20414 30994
rect 20414 30942 20466 30994
rect 20466 30942 20468 30994
rect 20412 30940 20468 30942
rect 21644 30994 21700 30996
rect 21644 30942 21646 30994
rect 21646 30942 21698 30994
rect 21698 30942 21700 30994
rect 21644 30940 21700 30942
rect 22268 30548 22324 30604
rect 22372 30602 22428 30604
rect 22476 30602 22532 30604
rect 22372 30550 22396 30602
rect 22396 30550 22428 30602
rect 22476 30550 22520 30602
rect 22520 30550 22532 30602
rect 22372 30548 22428 30550
rect 22476 30548 22532 30550
rect 22580 30548 22636 30604
rect 22684 30602 22740 30604
rect 22788 30602 22844 30604
rect 22684 30550 22696 30602
rect 22696 30550 22740 30602
rect 22788 30550 22820 30602
rect 22820 30550 22844 30602
rect 22684 30548 22740 30550
rect 22788 30548 22844 30550
rect 22892 30548 22948 30604
rect 19964 30268 20020 30324
rect 21532 30044 21588 30100
rect 17768 29764 17824 29820
rect 17872 29818 17928 29820
rect 17976 29818 18032 29820
rect 17872 29766 17896 29818
rect 17896 29766 17928 29818
rect 17976 29766 18020 29818
rect 18020 29766 18032 29818
rect 17872 29764 17928 29766
rect 17976 29764 18032 29766
rect 18080 29764 18136 29820
rect 18184 29818 18240 29820
rect 18288 29818 18344 29820
rect 18184 29766 18196 29818
rect 18196 29766 18240 29818
rect 18288 29766 18320 29818
rect 18320 29766 18344 29818
rect 18184 29764 18240 29766
rect 18288 29764 18344 29766
rect 18392 29764 18448 29820
rect 22428 30044 22484 30100
rect 23996 30044 24052 30100
rect 17724 29426 17780 29428
rect 17724 29374 17726 29426
rect 17726 29374 17778 29426
rect 17778 29374 17780 29426
rect 17724 29372 17780 29374
rect 18956 29426 19012 29428
rect 18956 29374 18958 29426
rect 18958 29374 19010 29426
rect 19010 29374 19012 29426
rect 18956 29372 19012 29374
rect 21980 28700 22036 28756
rect 17768 28196 17824 28252
rect 17872 28250 17928 28252
rect 17976 28250 18032 28252
rect 17872 28198 17896 28250
rect 17896 28198 17928 28250
rect 17976 28198 18020 28250
rect 18020 28198 18032 28250
rect 17872 28196 17928 28198
rect 17976 28196 18032 28198
rect 18080 28196 18136 28252
rect 18184 28250 18240 28252
rect 18288 28250 18344 28252
rect 18184 28198 18196 28250
rect 18196 28198 18240 28250
rect 18288 28198 18320 28250
rect 18320 28198 18344 28250
rect 18184 28196 18240 28198
rect 18288 28196 18344 28198
rect 18392 28196 18448 28252
rect 16604 26962 16660 26964
rect 16604 26910 16606 26962
rect 16606 26910 16658 26962
rect 16658 26910 16660 26962
rect 16604 26908 16660 26910
rect 20748 27186 20804 27188
rect 20748 27134 20750 27186
rect 20750 27134 20802 27186
rect 20802 27134 20804 27186
rect 20748 27132 20804 27134
rect 21980 27132 22036 27188
rect 21756 27074 21812 27076
rect 21756 27022 21758 27074
rect 21758 27022 21810 27074
rect 21810 27022 21812 27074
rect 21756 27020 21812 27022
rect 17612 26908 17668 26964
rect 12012 26796 12068 26852
rect 22268 28980 22324 29036
rect 22372 29034 22428 29036
rect 22476 29034 22532 29036
rect 22372 28982 22396 29034
rect 22396 28982 22428 29034
rect 22476 28982 22520 29034
rect 22520 28982 22532 29034
rect 22372 28980 22428 28982
rect 22476 28980 22532 28982
rect 22580 28980 22636 29036
rect 22684 29034 22740 29036
rect 22788 29034 22844 29036
rect 22684 28982 22696 29034
rect 22696 28982 22740 29034
rect 22788 28982 22820 29034
rect 22820 28982 22844 29034
rect 22684 28980 22740 28982
rect 22788 28980 22844 28982
rect 22892 28980 22948 29036
rect 24220 28754 24276 28756
rect 24220 28702 24222 28754
rect 24222 28702 24274 28754
rect 24274 28702 24276 28754
rect 24220 28700 24276 28702
rect 24444 28588 24500 28644
rect 25452 30156 25508 30212
rect 25452 28700 25508 28756
rect 24668 27804 24724 27860
rect 22268 27412 22324 27468
rect 22372 27466 22428 27468
rect 22476 27466 22532 27468
rect 22372 27414 22396 27466
rect 22396 27414 22428 27466
rect 22476 27414 22520 27466
rect 22520 27414 22532 27466
rect 22372 27412 22428 27414
rect 22476 27412 22532 27414
rect 22580 27412 22636 27468
rect 22684 27466 22740 27468
rect 22788 27466 22844 27468
rect 22684 27414 22696 27466
rect 22696 27414 22740 27466
rect 22788 27414 22820 27466
rect 22820 27414 22844 27466
rect 22684 27412 22740 27414
rect 22788 27412 22844 27414
rect 22892 27412 22948 27468
rect 23100 27020 23156 27076
rect 17768 26628 17824 26684
rect 17872 26682 17928 26684
rect 17976 26682 18032 26684
rect 17872 26630 17896 26682
rect 17896 26630 17928 26682
rect 17976 26630 18020 26682
rect 18020 26630 18032 26682
rect 17872 26628 17928 26630
rect 17976 26628 18032 26630
rect 18080 26628 18136 26684
rect 18184 26682 18240 26684
rect 18288 26682 18344 26684
rect 18184 26630 18196 26682
rect 18196 26630 18240 26682
rect 18288 26630 18320 26682
rect 18320 26630 18344 26682
rect 18184 26628 18240 26630
rect 18288 26628 18344 26630
rect 18392 26628 18448 26684
rect 17612 26460 17668 26516
rect 19180 26514 19236 26516
rect 19180 26462 19182 26514
rect 19182 26462 19234 26514
rect 19234 26462 19236 26514
rect 19180 26460 19236 26462
rect 19628 26460 19684 26516
rect 13268 25844 13324 25900
rect 13372 25898 13428 25900
rect 13476 25898 13532 25900
rect 13372 25846 13396 25898
rect 13396 25846 13428 25898
rect 13476 25846 13520 25898
rect 13520 25846 13532 25898
rect 13372 25844 13428 25846
rect 13476 25844 13532 25846
rect 13580 25844 13636 25900
rect 13684 25898 13740 25900
rect 13788 25898 13844 25900
rect 13684 25846 13696 25898
rect 13696 25846 13740 25898
rect 13788 25846 13820 25898
rect 13820 25846 13844 25898
rect 13684 25844 13740 25846
rect 13788 25844 13844 25846
rect 13892 25844 13948 25900
rect 16156 25676 16212 25732
rect 11340 25228 11396 25284
rect 11564 25340 11620 25396
rect 10220 23266 10276 23268
rect 10220 23214 10222 23266
rect 10222 23214 10274 23266
rect 10274 23214 10276 23266
rect 10220 23212 10276 23214
rect 9884 22204 9940 22260
rect 10780 22258 10836 22260
rect 10780 22206 10782 22258
rect 10782 22206 10834 22258
rect 10834 22206 10836 22258
rect 10780 22204 10836 22206
rect 12348 25394 12404 25396
rect 12348 25342 12350 25394
rect 12350 25342 12402 25394
rect 12402 25342 12404 25394
rect 12348 25340 12404 25342
rect 12684 25282 12740 25284
rect 12684 25230 12686 25282
rect 12686 25230 12738 25282
rect 12738 25230 12740 25282
rect 12684 25228 12740 25230
rect 15148 25228 15204 25284
rect 11900 24946 11956 24948
rect 11900 24894 11902 24946
rect 11902 24894 11954 24946
rect 11954 24894 11956 24946
rect 11900 24892 11956 24894
rect 13244 24892 13300 24948
rect 13268 24276 13324 24332
rect 13372 24330 13428 24332
rect 13476 24330 13532 24332
rect 13372 24278 13396 24330
rect 13396 24278 13428 24330
rect 13476 24278 13520 24330
rect 13520 24278 13532 24330
rect 13372 24276 13428 24278
rect 13476 24276 13532 24278
rect 13580 24276 13636 24332
rect 13684 24330 13740 24332
rect 13788 24330 13844 24332
rect 13684 24278 13696 24330
rect 13696 24278 13740 24330
rect 13788 24278 13820 24330
rect 13820 24278 13844 24330
rect 13684 24276 13740 24278
rect 13788 24276 13844 24278
rect 13892 24276 13948 24332
rect 15148 23996 15204 24052
rect 12460 23714 12516 23716
rect 12460 23662 12462 23714
rect 12462 23662 12514 23714
rect 12514 23662 12516 23714
rect 12460 23660 12516 23662
rect 11676 22146 11732 22148
rect 11676 22094 11678 22146
rect 11678 22094 11730 22146
rect 11730 22094 11732 22146
rect 11676 22092 11732 22094
rect 15596 23660 15652 23716
rect 17768 25060 17824 25116
rect 17872 25114 17928 25116
rect 17976 25114 18032 25116
rect 17872 25062 17896 25114
rect 17896 25062 17928 25114
rect 17976 25062 18020 25114
rect 18020 25062 18032 25114
rect 17872 25060 17928 25062
rect 17976 25060 18032 25062
rect 18080 25060 18136 25116
rect 18184 25114 18240 25116
rect 18288 25114 18344 25116
rect 18184 25062 18196 25114
rect 18196 25062 18240 25114
rect 18288 25062 18320 25114
rect 18320 25062 18344 25114
rect 18184 25060 18240 25062
rect 18288 25060 18344 25062
rect 18392 25060 18448 25116
rect 16380 23996 16436 24052
rect 17768 23492 17824 23548
rect 17872 23546 17928 23548
rect 17976 23546 18032 23548
rect 17872 23494 17896 23546
rect 17896 23494 17928 23546
rect 17976 23494 18020 23546
rect 18020 23494 18032 23546
rect 17872 23492 17928 23494
rect 17976 23492 18032 23494
rect 18080 23492 18136 23548
rect 18184 23546 18240 23548
rect 18288 23546 18344 23548
rect 18184 23494 18196 23546
rect 18196 23494 18240 23546
rect 18288 23494 18320 23546
rect 18320 23494 18344 23546
rect 18184 23492 18240 23494
rect 18288 23492 18344 23494
rect 18392 23492 18448 23548
rect 13268 22708 13324 22764
rect 13372 22762 13428 22764
rect 13476 22762 13532 22764
rect 13372 22710 13396 22762
rect 13396 22710 13428 22762
rect 13476 22710 13520 22762
rect 13520 22710 13532 22762
rect 13372 22708 13428 22710
rect 13476 22708 13532 22710
rect 13580 22708 13636 22764
rect 13684 22762 13740 22764
rect 13788 22762 13844 22764
rect 13684 22710 13696 22762
rect 13696 22710 13740 22762
rect 13788 22710 13820 22762
rect 13820 22710 13844 22762
rect 13684 22708 13740 22710
rect 13788 22708 13844 22710
rect 13892 22708 13948 22764
rect 14588 22146 14644 22148
rect 14588 22094 14590 22146
rect 14590 22094 14642 22146
rect 14642 22094 14644 22146
rect 14588 22092 14644 22094
rect 12460 21756 12516 21812
rect 13020 21810 13076 21812
rect 13020 21758 13022 21810
rect 13022 21758 13074 21810
rect 13074 21758 13076 21810
rect 13020 21756 13076 21758
rect 14812 21756 14868 21812
rect 13804 21698 13860 21700
rect 13804 21646 13806 21698
rect 13806 21646 13858 21698
rect 13858 21646 13860 21698
rect 13804 21644 13860 21646
rect 10668 21586 10724 21588
rect 10668 21534 10670 21586
rect 10670 21534 10722 21586
rect 10722 21534 10724 21586
rect 10668 21532 10724 21534
rect 14364 21586 14420 21588
rect 14364 21534 14366 21586
rect 14366 21534 14418 21586
rect 14418 21534 14420 21586
rect 14364 21532 14420 21534
rect 13268 21140 13324 21196
rect 13372 21194 13428 21196
rect 13476 21194 13532 21196
rect 13372 21142 13396 21194
rect 13396 21142 13428 21194
rect 13476 21142 13520 21194
rect 13520 21142 13532 21194
rect 13372 21140 13428 21142
rect 13476 21140 13532 21142
rect 13580 21140 13636 21196
rect 13684 21194 13740 21196
rect 13788 21194 13844 21196
rect 13684 21142 13696 21194
rect 13696 21142 13740 21194
rect 13788 21142 13820 21194
rect 13820 21142 13844 21194
rect 13684 21140 13740 21142
rect 13788 21140 13844 21142
rect 13892 21140 13948 21196
rect 14588 20748 14644 20804
rect 17768 21924 17824 21980
rect 17872 21978 17928 21980
rect 17976 21978 18032 21980
rect 17872 21926 17896 21978
rect 17896 21926 17928 21978
rect 17976 21926 18020 21978
rect 18020 21926 18032 21978
rect 17872 21924 17928 21926
rect 17976 21924 18032 21926
rect 18080 21924 18136 21980
rect 18184 21978 18240 21980
rect 18288 21978 18344 21980
rect 18184 21926 18196 21978
rect 18196 21926 18240 21978
rect 18288 21926 18320 21978
rect 18320 21926 18344 21978
rect 18184 21924 18240 21926
rect 18288 21924 18344 21926
rect 18392 21924 18448 21980
rect 15596 21756 15652 21812
rect 15148 21698 15204 21700
rect 15148 21646 15150 21698
rect 15150 21646 15202 21698
rect 15202 21646 15204 21698
rect 15148 21644 15204 21646
rect 16156 21586 16212 21588
rect 16156 21534 16158 21586
rect 16158 21534 16210 21586
rect 16210 21534 16212 21586
rect 16156 21532 16212 21534
rect 15820 20860 15876 20916
rect 16828 20860 16884 20916
rect 19292 23714 19348 23716
rect 19292 23662 19294 23714
rect 19294 23662 19346 23714
rect 19346 23662 19348 23714
rect 19292 23660 19348 23662
rect 19628 23212 19684 23268
rect 22316 26514 22372 26516
rect 22316 26462 22318 26514
rect 22318 26462 22370 26514
rect 22370 26462 22372 26514
rect 22316 26460 22372 26462
rect 23100 26514 23156 26516
rect 23100 26462 23102 26514
rect 23102 26462 23154 26514
rect 23154 26462 23156 26514
rect 23100 26460 23156 26462
rect 22268 25844 22324 25900
rect 22372 25898 22428 25900
rect 22476 25898 22532 25900
rect 22372 25846 22396 25898
rect 22396 25846 22428 25898
rect 22476 25846 22520 25898
rect 22520 25846 22532 25898
rect 22372 25844 22428 25846
rect 22476 25844 22532 25846
rect 22580 25844 22636 25900
rect 22684 25898 22740 25900
rect 22788 25898 22844 25900
rect 22684 25846 22696 25898
rect 22696 25846 22740 25898
rect 22788 25846 22820 25898
rect 22820 25846 22844 25898
rect 22684 25844 22740 25846
rect 22788 25844 22844 25846
rect 22892 25844 22948 25900
rect 25676 27858 25732 27860
rect 25676 27806 25678 27858
rect 25678 27806 25730 27858
rect 25730 27806 25732 27858
rect 25676 27804 25732 27806
rect 25676 25618 25732 25620
rect 25676 25566 25678 25618
rect 25678 25566 25730 25618
rect 25730 25566 25732 25618
rect 25676 25564 25732 25566
rect 25340 25452 25396 25508
rect 22268 24276 22324 24332
rect 22372 24330 22428 24332
rect 22476 24330 22532 24332
rect 22372 24278 22396 24330
rect 22396 24278 22428 24330
rect 22476 24278 22520 24330
rect 22520 24278 22532 24330
rect 22372 24276 22428 24278
rect 22476 24276 22532 24278
rect 22580 24276 22636 24332
rect 22684 24330 22740 24332
rect 22788 24330 22844 24332
rect 22684 24278 22696 24330
rect 22696 24278 22740 24330
rect 22788 24278 22820 24330
rect 22820 24278 22844 24330
rect 22684 24276 22740 24278
rect 22788 24276 22844 24278
rect 22892 24276 22948 24332
rect 20300 23266 20356 23268
rect 20300 23214 20302 23266
rect 20302 23214 20354 23266
rect 20354 23214 20356 23266
rect 20300 23212 20356 23214
rect 21420 23660 21476 23716
rect 21644 23660 21700 23716
rect 21756 23212 21812 23268
rect 20076 21756 20132 21812
rect 15260 20802 15316 20804
rect 15260 20750 15262 20802
rect 15262 20750 15314 20802
rect 15314 20750 15316 20802
rect 15260 20748 15316 20750
rect 10444 20076 10500 20132
rect 18396 20914 18452 20916
rect 18396 20862 18398 20914
rect 18398 20862 18450 20914
rect 18450 20862 18452 20914
rect 18396 20860 18452 20862
rect 17836 20636 17892 20692
rect 18732 20636 18788 20692
rect 17768 20356 17824 20412
rect 17872 20410 17928 20412
rect 17976 20410 18032 20412
rect 17872 20358 17896 20410
rect 17896 20358 17928 20410
rect 17976 20358 18020 20410
rect 18020 20358 18032 20410
rect 17872 20356 17928 20358
rect 17976 20356 18032 20358
rect 18080 20356 18136 20412
rect 18184 20410 18240 20412
rect 18288 20410 18344 20412
rect 18184 20358 18196 20410
rect 18196 20358 18240 20410
rect 18288 20358 18320 20410
rect 18320 20358 18344 20410
rect 18184 20356 18240 20358
rect 18288 20356 18344 20358
rect 18392 20356 18448 20412
rect 22540 23714 22596 23716
rect 22540 23662 22542 23714
rect 22542 23662 22594 23714
rect 22594 23662 22596 23714
rect 22540 23660 22596 23662
rect 22204 23100 22260 23156
rect 23436 23266 23492 23268
rect 23436 23214 23438 23266
rect 23438 23214 23490 23266
rect 23490 23214 23492 23266
rect 23436 23212 23492 23214
rect 23100 23100 23156 23156
rect 24220 23154 24276 23156
rect 24220 23102 24222 23154
rect 24222 23102 24274 23154
rect 24274 23102 24276 23154
rect 24220 23100 24276 23102
rect 22268 22708 22324 22764
rect 22372 22762 22428 22764
rect 22476 22762 22532 22764
rect 22372 22710 22396 22762
rect 22396 22710 22428 22762
rect 22476 22710 22520 22762
rect 22520 22710 22532 22762
rect 22372 22708 22428 22710
rect 22476 22708 22532 22710
rect 22580 22708 22636 22764
rect 22684 22762 22740 22764
rect 22788 22762 22844 22764
rect 22684 22710 22696 22762
rect 22696 22710 22740 22762
rect 22788 22710 22820 22762
rect 22820 22710 22844 22762
rect 22684 22708 22740 22710
rect 22788 22708 22844 22710
rect 22892 22708 22948 22764
rect 23100 21756 23156 21812
rect 22268 21140 22324 21196
rect 22372 21194 22428 21196
rect 22476 21194 22532 21196
rect 22372 21142 22396 21194
rect 22396 21142 22428 21194
rect 22476 21142 22520 21194
rect 22520 21142 22532 21194
rect 22372 21140 22428 21142
rect 22476 21140 22532 21142
rect 22580 21140 22636 21196
rect 22684 21194 22740 21196
rect 22788 21194 22844 21196
rect 22684 21142 22696 21194
rect 22696 21142 22740 21194
rect 22788 21142 22820 21194
rect 22820 21142 22844 21194
rect 22684 21140 22740 21142
rect 22788 21140 22844 21142
rect 22892 21140 22948 21196
rect 22988 20802 23044 20804
rect 22988 20750 22990 20802
rect 22990 20750 23042 20802
rect 23042 20750 23044 20802
rect 22988 20748 23044 20750
rect 24220 20802 24276 20804
rect 24220 20750 24222 20802
rect 24222 20750 24274 20802
rect 24274 20750 24276 20802
rect 24220 20748 24276 20750
rect 22428 20636 22484 20692
rect 23436 20690 23492 20692
rect 23436 20638 23438 20690
rect 23438 20638 23490 20690
rect 23490 20638 23492 20690
rect 23436 20636 23492 20638
rect 23996 20690 24052 20692
rect 23996 20638 23998 20690
rect 23998 20638 24050 20690
rect 24050 20638 24052 20690
rect 23996 20636 24052 20638
rect 24556 20578 24612 20580
rect 24556 20526 24558 20578
rect 24558 20526 24610 20578
rect 24610 20526 24612 20578
rect 24556 20524 24612 20526
rect 25340 20524 25396 20580
rect 17500 19852 17556 19908
rect 13268 19572 13324 19628
rect 13372 19626 13428 19628
rect 13476 19626 13532 19628
rect 13372 19574 13396 19626
rect 13396 19574 13428 19626
rect 13476 19574 13520 19626
rect 13520 19574 13532 19626
rect 13372 19572 13428 19574
rect 13476 19572 13532 19574
rect 13580 19572 13636 19628
rect 13684 19626 13740 19628
rect 13788 19626 13844 19628
rect 13684 19574 13696 19626
rect 13696 19574 13740 19626
rect 13788 19574 13820 19626
rect 13820 19574 13844 19626
rect 13684 19572 13740 19574
rect 13788 19572 13844 19574
rect 13892 19572 13948 19628
rect 18508 19404 18564 19460
rect 22268 19572 22324 19628
rect 22372 19626 22428 19628
rect 22476 19626 22532 19628
rect 22372 19574 22396 19626
rect 22396 19574 22428 19626
rect 22476 19574 22520 19626
rect 22520 19574 22532 19626
rect 22372 19572 22428 19574
rect 22476 19572 22532 19574
rect 22580 19572 22636 19628
rect 22684 19626 22740 19628
rect 22788 19626 22844 19628
rect 22684 19574 22696 19626
rect 22696 19574 22740 19626
rect 22788 19574 22820 19626
rect 22820 19574 22844 19626
rect 22684 19572 22740 19574
rect 22788 19572 22844 19574
rect 22892 19572 22948 19628
rect 19292 19404 19348 19460
rect 17768 18788 17824 18844
rect 17872 18842 17928 18844
rect 17976 18842 18032 18844
rect 17872 18790 17896 18842
rect 17896 18790 17928 18842
rect 17976 18790 18020 18842
rect 18020 18790 18032 18842
rect 17872 18788 17928 18790
rect 17976 18788 18032 18790
rect 18080 18788 18136 18844
rect 18184 18842 18240 18844
rect 18288 18842 18344 18844
rect 18184 18790 18196 18842
rect 18196 18790 18240 18842
rect 18288 18790 18320 18842
rect 18320 18790 18344 18842
rect 18184 18788 18240 18790
rect 18288 18788 18344 18790
rect 18392 18788 18448 18844
rect 13268 18004 13324 18060
rect 13372 18058 13428 18060
rect 13476 18058 13532 18060
rect 13372 18006 13396 18058
rect 13396 18006 13428 18058
rect 13476 18006 13520 18058
rect 13520 18006 13532 18058
rect 13372 18004 13428 18006
rect 13476 18004 13532 18006
rect 13580 18004 13636 18060
rect 13684 18058 13740 18060
rect 13788 18058 13844 18060
rect 13684 18006 13696 18058
rect 13696 18006 13740 18058
rect 13788 18006 13820 18058
rect 13820 18006 13844 18058
rect 13684 18004 13740 18006
rect 13788 18004 13844 18006
rect 13892 18004 13948 18060
rect 22268 18004 22324 18060
rect 22372 18058 22428 18060
rect 22476 18058 22532 18060
rect 22372 18006 22396 18058
rect 22396 18006 22428 18058
rect 22476 18006 22520 18058
rect 22520 18006 22532 18058
rect 22372 18004 22428 18006
rect 22476 18004 22532 18006
rect 22580 18004 22636 18060
rect 22684 18058 22740 18060
rect 22788 18058 22844 18060
rect 22684 18006 22696 18058
rect 22696 18006 22740 18058
rect 22788 18006 22820 18058
rect 22820 18006 22844 18058
rect 22684 18004 22740 18006
rect 22788 18004 22844 18006
rect 22892 18004 22948 18060
rect 17768 17220 17824 17276
rect 17872 17274 17928 17276
rect 17976 17274 18032 17276
rect 17872 17222 17896 17274
rect 17896 17222 17928 17274
rect 17976 17222 18020 17274
rect 18020 17222 18032 17274
rect 17872 17220 17928 17222
rect 17976 17220 18032 17222
rect 18080 17220 18136 17276
rect 18184 17274 18240 17276
rect 18288 17274 18344 17276
rect 18184 17222 18196 17274
rect 18196 17222 18240 17274
rect 18288 17222 18320 17274
rect 18320 17222 18344 17274
rect 18184 17220 18240 17222
rect 18288 17220 18344 17222
rect 18392 17220 18448 17276
rect 13268 16436 13324 16492
rect 13372 16490 13428 16492
rect 13476 16490 13532 16492
rect 13372 16438 13396 16490
rect 13396 16438 13428 16490
rect 13476 16438 13520 16490
rect 13520 16438 13532 16490
rect 13372 16436 13428 16438
rect 13476 16436 13532 16438
rect 13580 16436 13636 16492
rect 13684 16490 13740 16492
rect 13788 16490 13844 16492
rect 13684 16438 13696 16490
rect 13696 16438 13740 16490
rect 13788 16438 13820 16490
rect 13820 16438 13844 16490
rect 13684 16436 13740 16438
rect 13788 16436 13844 16438
rect 13892 16436 13948 16492
rect 22268 16436 22324 16492
rect 22372 16490 22428 16492
rect 22476 16490 22532 16492
rect 22372 16438 22396 16490
rect 22396 16438 22428 16490
rect 22476 16438 22520 16490
rect 22520 16438 22532 16490
rect 22372 16436 22428 16438
rect 22476 16436 22532 16438
rect 22580 16436 22636 16492
rect 22684 16490 22740 16492
rect 22788 16490 22844 16492
rect 22684 16438 22696 16490
rect 22696 16438 22740 16490
rect 22788 16438 22820 16490
rect 22820 16438 22844 16490
rect 22684 16436 22740 16438
rect 22788 16436 22844 16438
rect 22892 16436 22948 16492
rect 17768 15652 17824 15708
rect 17872 15706 17928 15708
rect 17976 15706 18032 15708
rect 17872 15654 17896 15706
rect 17896 15654 17928 15706
rect 17976 15654 18020 15706
rect 18020 15654 18032 15706
rect 17872 15652 17928 15654
rect 17976 15652 18032 15654
rect 18080 15652 18136 15708
rect 18184 15706 18240 15708
rect 18288 15706 18344 15708
rect 18184 15654 18196 15706
rect 18196 15654 18240 15706
rect 18288 15654 18320 15706
rect 18320 15654 18344 15706
rect 18184 15652 18240 15654
rect 18288 15652 18344 15654
rect 18392 15652 18448 15708
rect 13268 14868 13324 14924
rect 13372 14922 13428 14924
rect 13476 14922 13532 14924
rect 13372 14870 13396 14922
rect 13396 14870 13428 14922
rect 13476 14870 13520 14922
rect 13520 14870 13532 14922
rect 13372 14868 13428 14870
rect 13476 14868 13532 14870
rect 13580 14868 13636 14924
rect 13684 14922 13740 14924
rect 13788 14922 13844 14924
rect 13684 14870 13696 14922
rect 13696 14870 13740 14922
rect 13788 14870 13820 14922
rect 13820 14870 13844 14922
rect 13684 14868 13740 14870
rect 13788 14868 13844 14870
rect 13892 14868 13948 14924
rect 22268 14868 22324 14924
rect 22372 14922 22428 14924
rect 22476 14922 22532 14924
rect 22372 14870 22396 14922
rect 22396 14870 22428 14922
rect 22476 14870 22520 14922
rect 22520 14870 22532 14922
rect 22372 14868 22428 14870
rect 22476 14868 22532 14870
rect 22580 14868 22636 14924
rect 22684 14922 22740 14924
rect 22788 14922 22844 14924
rect 22684 14870 22696 14922
rect 22696 14870 22740 14922
rect 22788 14870 22820 14922
rect 22820 14870 22844 14922
rect 22684 14868 22740 14870
rect 22788 14868 22844 14870
rect 22892 14868 22948 14924
rect 20748 14476 20804 14532
rect 21420 14530 21476 14532
rect 21420 14478 21422 14530
rect 21422 14478 21474 14530
rect 21474 14478 21476 14530
rect 21420 14476 21476 14478
rect 17768 14084 17824 14140
rect 17872 14138 17928 14140
rect 17976 14138 18032 14140
rect 17872 14086 17896 14138
rect 17896 14086 17928 14138
rect 17976 14086 18020 14138
rect 18020 14086 18032 14138
rect 17872 14084 17928 14086
rect 17976 14084 18032 14086
rect 18080 14084 18136 14140
rect 18184 14138 18240 14140
rect 18288 14138 18344 14140
rect 18184 14086 18196 14138
rect 18196 14086 18240 14138
rect 18288 14086 18320 14138
rect 18320 14086 18344 14138
rect 18184 14084 18240 14086
rect 18288 14084 18344 14086
rect 18392 14084 18448 14140
rect 9660 13916 9716 13972
rect 13268 13300 13324 13356
rect 13372 13354 13428 13356
rect 13476 13354 13532 13356
rect 13372 13302 13396 13354
rect 13396 13302 13428 13354
rect 13476 13302 13520 13354
rect 13520 13302 13532 13354
rect 13372 13300 13428 13302
rect 13476 13300 13532 13302
rect 13580 13300 13636 13356
rect 13684 13354 13740 13356
rect 13788 13354 13844 13356
rect 13684 13302 13696 13354
rect 13696 13302 13740 13354
rect 13788 13302 13820 13354
rect 13820 13302 13844 13354
rect 13684 13300 13740 13302
rect 13788 13300 13844 13302
rect 13892 13300 13948 13356
rect 8768 12516 8824 12572
rect 8872 12570 8928 12572
rect 8976 12570 9032 12572
rect 8872 12518 8896 12570
rect 8896 12518 8928 12570
rect 8976 12518 9020 12570
rect 9020 12518 9032 12570
rect 8872 12516 8928 12518
rect 8976 12516 9032 12518
rect 9080 12516 9136 12572
rect 9184 12570 9240 12572
rect 9288 12570 9344 12572
rect 9184 12518 9196 12570
rect 9196 12518 9240 12570
rect 9288 12518 9320 12570
rect 9320 12518 9344 12570
rect 9184 12516 9240 12518
rect 9288 12516 9344 12518
rect 9392 12516 9448 12572
rect 17768 12516 17824 12572
rect 17872 12570 17928 12572
rect 17976 12570 18032 12572
rect 17872 12518 17896 12570
rect 17896 12518 17928 12570
rect 17976 12518 18020 12570
rect 18020 12518 18032 12570
rect 17872 12516 17928 12518
rect 17976 12516 18032 12518
rect 18080 12516 18136 12572
rect 18184 12570 18240 12572
rect 18288 12570 18344 12572
rect 18184 12518 18196 12570
rect 18196 12518 18240 12570
rect 18288 12518 18320 12570
rect 18320 12518 18344 12570
rect 18184 12516 18240 12518
rect 18288 12516 18344 12518
rect 18392 12516 18448 12572
rect 13268 11732 13324 11788
rect 13372 11786 13428 11788
rect 13476 11786 13532 11788
rect 13372 11734 13396 11786
rect 13396 11734 13428 11786
rect 13476 11734 13520 11786
rect 13520 11734 13532 11786
rect 13372 11732 13428 11734
rect 13476 11732 13532 11734
rect 13580 11732 13636 11788
rect 13684 11786 13740 11788
rect 13788 11786 13844 11788
rect 13684 11734 13696 11786
rect 13696 11734 13740 11786
rect 13788 11734 13820 11786
rect 13820 11734 13844 11786
rect 13684 11732 13740 11734
rect 13788 11732 13844 11734
rect 13892 11732 13948 11788
rect 8768 10948 8824 11004
rect 8872 11002 8928 11004
rect 8976 11002 9032 11004
rect 8872 10950 8896 11002
rect 8896 10950 8928 11002
rect 8976 10950 9020 11002
rect 9020 10950 9032 11002
rect 8872 10948 8928 10950
rect 8976 10948 9032 10950
rect 9080 10948 9136 11004
rect 9184 11002 9240 11004
rect 9288 11002 9344 11004
rect 9184 10950 9196 11002
rect 9196 10950 9240 11002
rect 9288 10950 9320 11002
rect 9320 10950 9344 11002
rect 9184 10948 9240 10950
rect 9288 10948 9344 10950
rect 9392 10948 9448 11004
rect 17768 10948 17824 11004
rect 17872 11002 17928 11004
rect 17976 11002 18032 11004
rect 17872 10950 17896 11002
rect 17896 10950 17928 11002
rect 17976 10950 18020 11002
rect 18020 10950 18032 11002
rect 17872 10948 17928 10950
rect 17976 10948 18032 10950
rect 18080 10948 18136 11004
rect 18184 11002 18240 11004
rect 18288 11002 18344 11004
rect 18184 10950 18196 11002
rect 18196 10950 18240 11002
rect 18288 10950 18320 11002
rect 18320 10950 18344 11002
rect 18184 10948 18240 10950
rect 18288 10948 18344 10950
rect 18392 10948 18448 11004
rect 13268 10164 13324 10220
rect 13372 10218 13428 10220
rect 13476 10218 13532 10220
rect 13372 10166 13396 10218
rect 13396 10166 13428 10218
rect 13476 10166 13520 10218
rect 13520 10166 13532 10218
rect 13372 10164 13428 10166
rect 13476 10164 13532 10166
rect 13580 10164 13636 10220
rect 13684 10218 13740 10220
rect 13788 10218 13844 10220
rect 13684 10166 13696 10218
rect 13696 10166 13740 10218
rect 13788 10166 13820 10218
rect 13820 10166 13844 10218
rect 13684 10164 13740 10166
rect 13788 10164 13844 10166
rect 13892 10164 13948 10220
rect 8768 9380 8824 9436
rect 8872 9434 8928 9436
rect 8976 9434 9032 9436
rect 8872 9382 8896 9434
rect 8896 9382 8928 9434
rect 8976 9382 9020 9434
rect 9020 9382 9032 9434
rect 8872 9380 8928 9382
rect 8976 9380 9032 9382
rect 9080 9380 9136 9436
rect 9184 9434 9240 9436
rect 9288 9434 9344 9436
rect 9184 9382 9196 9434
rect 9196 9382 9240 9434
rect 9288 9382 9320 9434
rect 9320 9382 9344 9434
rect 9184 9380 9240 9382
rect 9288 9380 9344 9382
rect 9392 9380 9448 9436
rect 17768 9380 17824 9436
rect 17872 9434 17928 9436
rect 17976 9434 18032 9436
rect 17872 9382 17896 9434
rect 17896 9382 17928 9434
rect 17976 9382 18020 9434
rect 18020 9382 18032 9434
rect 17872 9380 17928 9382
rect 17976 9380 18032 9382
rect 18080 9380 18136 9436
rect 18184 9434 18240 9436
rect 18288 9434 18344 9436
rect 18184 9382 18196 9434
rect 18196 9382 18240 9434
rect 18288 9382 18320 9434
rect 18320 9382 18344 9434
rect 18184 9380 18240 9382
rect 18288 9380 18344 9382
rect 18392 9380 18448 9436
rect 13268 8596 13324 8652
rect 13372 8650 13428 8652
rect 13476 8650 13532 8652
rect 13372 8598 13396 8650
rect 13396 8598 13428 8650
rect 13476 8598 13520 8650
rect 13520 8598 13532 8650
rect 13372 8596 13428 8598
rect 13476 8596 13532 8598
rect 13580 8596 13636 8652
rect 13684 8650 13740 8652
rect 13788 8650 13844 8652
rect 13684 8598 13696 8650
rect 13696 8598 13740 8650
rect 13788 8598 13820 8650
rect 13820 8598 13844 8650
rect 13684 8596 13740 8598
rect 13788 8596 13844 8598
rect 13892 8596 13948 8652
rect 8768 7812 8824 7868
rect 8872 7866 8928 7868
rect 8976 7866 9032 7868
rect 8872 7814 8896 7866
rect 8896 7814 8928 7866
rect 8976 7814 9020 7866
rect 9020 7814 9032 7866
rect 8872 7812 8928 7814
rect 8976 7812 9032 7814
rect 9080 7812 9136 7868
rect 9184 7866 9240 7868
rect 9288 7866 9344 7868
rect 9184 7814 9196 7866
rect 9196 7814 9240 7866
rect 9288 7814 9320 7866
rect 9320 7814 9344 7866
rect 9184 7812 9240 7814
rect 9288 7812 9344 7814
rect 9392 7812 9448 7868
rect 17768 7812 17824 7868
rect 17872 7866 17928 7868
rect 17976 7866 18032 7868
rect 17872 7814 17896 7866
rect 17896 7814 17928 7866
rect 17976 7814 18020 7866
rect 18020 7814 18032 7866
rect 17872 7812 17928 7814
rect 17976 7812 18032 7814
rect 18080 7812 18136 7868
rect 18184 7866 18240 7868
rect 18288 7866 18344 7868
rect 18184 7814 18196 7866
rect 18196 7814 18240 7866
rect 18288 7814 18320 7866
rect 18320 7814 18344 7866
rect 18184 7812 18240 7814
rect 18288 7812 18344 7814
rect 18392 7812 18448 7868
rect 13268 7028 13324 7084
rect 13372 7082 13428 7084
rect 13476 7082 13532 7084
rect 13372 7030 13396 7082
rect 13396 7030 13428 7082
rect 13476 7030 13520 7082
rect 13520 7030 13532 7082
rect 13372 7028 13428 7030
rect 13476 7028 13532 7030
rect 13580 7028 13636 7084
rect 13684 7082 13740 7084
rect 13788 7082 13844 7084
rect 13684 7030 13696 7082
rect 13696 7030 13740 7082
rect 13788 7030 13820 7082
rect 13820 7030 13844 7082
rect 13684 7028 13740 7030
rect 13788 7028 13844 7030
rect 13892 7028 13948 7084
rect 8768 6244 8824 6300
rect 8872 6298 8928 6300
rect 8976 6298 9032 6300
rect 8872 6246 8896 6298
rect 8896 6246 8928 6298
rect 8976 6246 9020 6298
rect 9020 6246 9032 6298
rect 8872 6244 8928 6246
rect 8976 6244 9032 6246
rect 9080 6244 9136 6300
rect 9184 6298 9240 6300
rect 9288 6298 9344 6300
rect 9184 6246 9196 6298
rect 9196 6246 9240 6298
rect 9288 6246 9320 6298
rect 9320 6246 9344 6298
rect 9184 6244 9240 6246
rect 9288 6244 9344 6246
rect 9392 6244 9448 6300
rect 17768 6244 17824 6300
rect 17872 6298 17928 6300
rect 17976 6298 18032 6300
rect 17872 6246 17896 6298
rect 17896 6246 17928 6298
rect 17976 6246 18020 6298
rect 18020 6246 18032 6298
rect 17872 6244 17928 6246
rect 17976 6244 18032 6246
rect 18080 6244 18136 6300
rect 18184 6298 18240 6300
rect 18288 6298 18344 6300
rect 18184 6246 18196 6298
rect 18196 6246 18240 6298
rect 18288 6246 18320 6298
rect 18320 6246 18344 6298
rect 18184 6244 18240 6246
rect 18288 6244 18344 6246
rect 18392 6244 18448 6300
rect 13268 5460 13324 5516
rect 13372 5514 13428 5516
rect 13476 5514 13532 5516
rect 13372 5462 13396 5514
rect 13396 5462 13428 5514
rect 13476 5462 13520 5514
rect 13520 5462 13532 5514
rect 13372 5460 13428 5462
rect 13476 5460 13532 5462
rect 13580 5460 13636 5516
rect 13684 5514 13740 5516
rect 13788 5514 13844 5516
rect 13684 5462 13696 5514
rect 13696 5462 13740 5514
rect 13788 5462 13820 5514
rect 13820 5462 13844 5514
rect 13684 5460 13740 5462
rect 13788 5460 13844 5462
rect 13892 5460 13948 5516
rect 8768 4676 8824 4732
rect 8872 4730 8928 4732
rect 8976 4730 9032 4732
rect 8872 4678 8896 4730
rect 8896 4678 8928 4730
rect 8976 4678 9020 4730
rect 9020 4678 9032 4730
rect 8872 4676 8928 4678
rect 8976 4676 9032 4678
rect 9080 4676 9136 4732
rect 9184 4730 9240 4732
rect 9288 4730 9344 4732
rect 9184 4678 9196 4730
rect 9196 4678 9240 4730
rect 9288 4678 9320 4730
rect 9320 4678 9344 4730
rect 9184 4676 9240 4678
rect 9288 4676 9344 4678
rect 9392 4676 9448 4732
rect 17768 4676 17824 4732
rect 17872 4730 17928 4732
rect 17976 4730 18032 4732
rect 17872 4678 17896 4730
rect 17896 4678 17928 4730
rect 17976 4678 18020 4730
rect 18020 4678 18032 4730
rect 17872 4676 17928 4678
rect 17976 4676 18032 4678
rect 18080 4676 18136 4732
rect 18184 4730 18240 4732
rect 18288 4730 18344 4732
rect 18184 4678 18196 4730
rect 18196 4678 18240 4730
rect 18288 4678 18320 4730
rect 18320 4678 18344 4730
rect 18184 4676 18240 4678
rect 18288 4676 18344 4678
rect 18392 4676 18448 4732
rect 22268 13300 22324 13356
rect 22372 13354 22428 13356
rect 22476 13354 22532 13356
rect 22372 13302 22396 13354
rect 22396 13302 22428 13354
rect 22476 13302 22520 13354
rect 22520 13302 22532 13354
rect 22372 13300 22428 13302
rect 22476 13300 22532 13302
rect 22580 13300 22636 13356
rect 22684 13354 22740 13356
rect 22788 13354 22844 13356
rect 22684 13302 22696 13354
rect 22696 13302 22740 13354
rect 22788 13302 22820 13354
rect 22820 13302 22844 13354
rect 22684 13300 22740 13302
rect 22788 13300 22844 13302
rect 22892 13300 22948 13356
rect 22268 11732 22324 11788
rect 22372 11786 22428 11788
rect 22476 11786 22532 11788
rect 22372 11734 22396 11786
rect 22396 11734 22428 11786
rect 22476 11734 22520 11786
rect 22520 11734 22532 11786
rect 22372 11732 22428 11734
rect 22476 11732 22532 11734
rect 22580 11732 22636 11788
rect 22684 11786 22740 11788
rect 22788 11786 22844 11788
rect 22684 11734 22696 11786
rect 22696 11734 22740 11786
rect 22788 11734 22820 11786
rect 22820 11734 22844 11786
rect 22684 11732 22740 11734
rect 22788 11732 22844 11734
rect 22892 11732 22948 11788
rect 27132 31778 27188 31780
rect 27132 31726 27134 31778
rect 27134 31726 27186 31778
rect 27186 31726 27188 31778
rect 27132 31724 27188 31726
rect 26460 31500 26516 31556
rect 27468 31554 27524 31556
rect 27468 31502 27470 31554
rect 27470 31502 27522 31554
rect 27522 31502 27524 31554
rect 27468 31500 27524 31502
rect 26768 31332 26824 31388
rect 26872 31386 26928 31388
rect 26976 31386 27032 31388
rect 26872 31334 26896 31386
rect 26896 31334 26928 31386
rect 26976 31334 27020 31386
rect 27020 31334 27032 31386
rect 26872 31332 26928 31334
rect 26976 31332 27032 31334
rect 27080 31332 27136 31388
rect 27184 31386 27240 31388
rect 27288 31386 27344 31388
rect 27184 31334 27196 31386
rect 27196 31334 27240 31386
rect 27288 31334 27320 31386
rect 27320 31334 27344 31386
rect 27184 31332 27240 31334
rect 27288 31332 27344 31334
rect 27392 31332 27448 31388
rect 26236 30210 26292 30212
rect 26236 30158 26238 30210
rect 26238 30158 26290 30210
rect 26290 30158 26292 30210
rect 26236 30156 26292 30158
rect 27244 30210 27300 30212
rect 27244 30158 27246 30210
rect 27246 30158 27298 30210
rect 27298 30158 27300 30210
rect 27244 30156 27300 30158
rect 26768 29764 26824 29820
rect 26872 29818 26928 29820
rect 26976 29818 27032 29820
rect 26872 29766 26896 29818
rect 26896 29766 26928 29818
rect 26976 29766 27020 29818
rect 27020 29766 27032 29818
rect 26872 29764 26928 29766
rect 26976 29764 27032 29766
rect 27080 29764 27136 29820
rect 27184 29818 27240 29820
rect 27288 29818 27344 29820
rect 27184 29766 27196 29818
rect 27196 29766 27240 29818
rect 27288 29766 27320 29818
rect 27320 29766 27344 29818
rect 27184 29764 27240 29766
rect 27288 29764 27344 29766
rect 27392 29764 27448 29820
rect 26572 29596 26628 29652
rect 25900 28754 25956 28756
rect 25900 28702 25902 28754
rect 25902 28702 25954 28754
rect 25954 28702 25956 28754
rect 25900 28700 25956 28702
rect 26236 28642 26292 28644
rect 26236 28590 26238 28642
rect 26238 28590 26290 28642
rect 26290 28590 26292 28642
rect 26236 28588 26292 28590
rect 26796 28642 26852 28644
rect 26796 28590 26798 28642
rect 26798 28590 26850 28642
rect 26850 28590 26852 28642
rect 26796 28588 26852 28590
rect 26768 28196 26824 28252
rect 26872 28250 26928 28252
rect 26976 28250 27032 28252
rect 26872 28198 26896 28250
rect 26896 28198 26928 28250
rect 26976 28198 27020 28250
rect 27020 28198 27032 28250
rect 26872 28196 26928 28198
rect 26976 28196 27032 28198
rect 27080 28196 27136 28252
rect 27184 28250 27240 28252
rect 27288 28250 27344 28252
rect 27184 28198 27196 28250
rect 27196 28198 27240 28250
rect 27288 28198 27320 28250
rect 27320 28198 27344 28250
rect 27184 28196 27240 28198
rect 27288 28196 27344 28198
rect 27392 28196 27448 28252
rect 26768 26628 26824 26684
rect 26872 26682 26928 26684
rect 26976 26682 27032 26684
rect 26872 26630 26896 26682
rect 26896 26630 26928 26682
rect 26976 26630 27020 26682
rect 27020 26630 27032 26682
rect 26872 26628 26928 26630
rect 26976 26628 27032 26630
rect 27080 26628 27136 26684
rect 27184 26682 27240 26684
rect 27288 26682 27344 26684
rect 27184 26630 27196 26682
rect 27196 26630 27240 26682
rect 27288 26630 27320 26682
rect 27320 26630 27344 26682
rect 27184 26628 27240 26630
rect 27288 26628 27344 26630
rect 27392 26628 27448 26684
rect 26460 26290 26516 26292
rect 26460 26238 26462 26290
rect 26462 26238 26514 26290
rect 26514 26238 26516 26290
rect 26460 26236 26516 26238
rect 26124 25564 26180 25620
rect 26236 25506 26292 25508
rect 26236 25454 26238 25506
rect 26238 25454 26290 25506
rect 26290 25454 26292 25506
rect 26236 25452 26292 25454
rect 26460 25228 26516 25284
rect 27244 26236 27300 26292
rect 29036 32396 29092 32452
rect 29932 36988 29988 37044
rect 30044 36204 30100 36260
rect 31724 36988 31780 37044
rect 31268 36820 31324 36876
rect 31372 36874 31428 36876
rect 31476 36874 31532 36876
rect 31372 36822 31396 36874
rect 31396 36822 31428 36874
rect 31476 36822 31520 36874
rect 31520 36822 31532 36874
rect 31372 36820 31428 36822
rect 31476 36820 31532 36822
rect 31580 36820 31636 36876
rect 31684 36874 31740 36876
rect 31788 36874 31844 36876
rect 31684 36822 31696 36874
rect 31696 36822 31740 36874
rect 31788 36822 31820 36874
rect 31820 36822 31844 36874
rect 31684 36820 31740 36822
rect 31788 36820 31844 36822
rect 31892 36820 31948 36876
rect 31612 36652 31668 36708
rect 34860 37938 34916 37940
rect 34860 37886 34862 37938
rect 34862 37886 34914 37938
rect 34914 37886 34916 37938
rect 34860 37884 34916 37886
rect 34860 37436 34916 37492
rect 35420 40402 35476 40404
rect 35420 40350 35422 40402
rect 35422 40350 35474 40402
rect 35474 40350 35476 40402
rect 35420 40348 35476 40350
rect 35868 42924 35924 42980
rect 35768 42308 35824 42364
rect 35872 42362 35928 42364
rect 35976 42362 36032 42364
rect 35872 42310 35896 42362
rect 35896 42310 35928 42362
rect 35976 42310 36020 42362
rect 36020 42310 36032 42362
rect 35872 42308 35928 42310
rect 35976 42308 36032 42310
rect 36080 42308 36136 42364
rect 36184 42362 36240 42364
rect 36288 42362 36344 42364
rect 36184 42310 36196 42362
rect 36196 42310 36240 42362
rect 36288 42310 36320 42362
rect 36320 42310 36344 42362
rect 36184 42308 36240 42310
rect 36288 42308 36344 42310
rect 36392 42308 36448 42364
rect 35868 41186 35924 41188
rect 35868 41134 35870 41186
rect 35870 41134 35922 41186
rect 35922 41134 35924 41186
rect 35868 41132 35924 41134
rect 37100 41020 37156 41076
rect 35768 40740 35824 40796
rect 35872 40794 35928 40796
rect 35976 40794 36032 40796
rect 35872 40742 35896 40794
rect 35896 40742 35928 40794
rect 35976 40742 36020 40794
rect 36020 40742 36032 40794
rect 35872 40740 35928 40742
rect 35976 40740 36032 40742
rect 36080 40740 36136 40796
rect 36184 40794 36240 40796
rect 36288 40794 36344 40796
rect 36184 40742 36196 40794
rect 36196 40742 36240 40794
rect 36288 40742 36320 40794
rect 36320 40742 36344 40794
rect 36184 40740 36240 40742
rect 36288 40740 36344 40742
rect 36392 40740 36448 40796
rect 36092 40460 36148 40516
rect 36540 39618 36596 39620
rect 36540 39566 36542 39618
rect 36542 39566 36594 39618
rect 36594 39566 36596 39618
rect 36540 39564 36596 39566
rect 36204 39506 36260 39508
rect 36204 39454 36206 39506
rect 36206 39454 36258 39506
rect 36258 39454 36260 39506
rect 36204 39452 36260 39454
rect 35868 39394 35924 39396
rect 35868 39342 35870 39394
rect 35870 39342 35922 39394
rect 35922 39342 35924 39394
rect 35868 39340 35924 39342
rect 36316 39394 36372 39396
rect 36316 39342 36318 39394
rect 36318 39342 36370 39394
rect 36370 39342 36372 39394
rect 36316 39340 36372 39342
rect 35768 39172 35824 39228
rect 35872 39226 35928 39228
rect 35976 39226 36032 39228
rect 35872 39174 35896 39226
rect 35896 39174 35928 39226
rect 35976 39174 36020 39226
rect 36020 39174 36032 39226
rect 35872 39172 35928 39174
rect 35976 39172 36032 39174
rect 36080 39172 36136 39228
rect 36184 39226 36240 39228
rect 36288 39226 36344 39228
rect 36184 39174 36196 39226
rect 36196 39174 36240 39226
rect 36288 39174 36320 39226
rect 36320 39174 36344 39226
rect 36184 39172 36240 39174
rect 36288 39172 36344 39174
rect 36392 39172 36448 39228
rect 35644 38668 35700 38724
rect 35084 37266 35140 37268
rect 35084 37214 35086 37266
rect 35086 37214 35138 37266
rect 35138 37214 35140 37266
rect 35084 37212 35140 37214
rect 35768 37604 35824 37660
rect 35872 37658 35928 37660
rect 35976 37658 36032 37660
rect 35872 37606 35896 37658
rect 35896 37606 35928 37658
rect 35976 37606 36020 37658
rect 36020 37606 36032 37658
rect 35872 37604 35928 37606
rect 35976 37604 36032 37606
rect 36080 37604 36136 37660
rect 36184 37658 36240 37660
rect 36288 37658 36344 37660
rect 36184 37606 36196 37658
rect 36196 37606 36240 37658
rect 36288 37606 36320 37658
rect 36320 37606 36344 37658
rect 36184 37604 36240 37606
rect 36288 37604 36344 37606
rect 36392 37604 36448 37660
rect 38444 43372 38500 43428
rect 39900 45666 39956 45668
rect 39900 45614 39902 45666
rect 39902 45614 39954 45666
rect 39954 45614 39956 45666
rect 39900 45612 39956 45614
rect 38780 42028 38836 42084
rect 35644 37100 35700 37156
rect 34300 36988 34356 37044
rect 35084 36988 35140 37044
rect 36876 37100 36932 37156
rect 36988 39506 37044 39508
rect 36988 39454 36990 39506
rect 36990 39454 37042 39506
rect 37042 39454 37044 39506
rect 36988 39452 37044 39454
rect 37324 39618 37380 39620
rect 37324 39566 37326 39618
rect 37326 39566 37378 39618
rect 37378 39566 37380 39618
rect 37324 39564 37380 39566
rect 35756 36988 35812 37044
rect 36876 36652 36932 36708
rect 36764 36316 36820 36372
rect 31164 36258 31220 36260
rect 31164 36206 31166 36258
rect 31166 36206 31218 36258
rect 31218 36206 31220 36258
rect 31164 36204 31220 36206
rect 34300 36258 34356 36260
rect 34300 36206 34302 36258
rect 34302 36206 34354 36258
rect 34354 36206 34356 36258
rect 34300 36204 34356 36206
rect 35768 36036 35824 36092
rect 35872 36090 35928 36092
rect 35976 36090 36032 36092
rect 35872 36038 35896 36090
rect 35896 36038 35928 36090
rect 35976 36038 36020 36090
rect 36020 36038 36032 36090
rect 35872 36036 35928 36038
rect 35976 36036 36032 36038
rect 36080 36036 36136 36092
rect 36184 36090 36240 36092
rect 36288 36090 36344 36092
rect 36184 36038 36196 36090
rect 36196 36038 36240 36090
rect 36288 36038 36320 36090
rect 36320 36038 36344 36090
rect 36184 36036 36240 36038
rect 36288 36036 36344 36038
rect 36392 36036 36448 36092
rect 29708 33852 29764 33908
rect 36764 35922 36820 35924
rect 36764 35870 36766 35922
rect 36766 35870 36818 35922
rect 36818 35870 36820 35922
rect 36764 35868 36820 35870
rect 35868 35644 35924 35700
rect 31268 35252 31324 35308
rect 31372 35306 31428 35308
rect 31476 35306 31532 35308
rect 31372 35254 31396 35306
rect 31396 35254 31428 35306
rect 31476 35254 31520 35306
rect 31520 35254 31532 35306
rect 31372 35252 31428 35254
rect 31476 35252 31532 35254
rect 31580 35252 31636 35308
rect 31684 35306 31740 35308
rect 31788 35306 31844 35308
rect 31684 35254 31696 35306
rect 31696 35254 31740 35306
rect 31788 35254 31820 35306
rect 31820 35254 31844 35306
rect 31684 35252 31740 35254
rect 31788 35252 31844 35254
rect 31892 35252 31948 35308
rect 36652 35698 36708 35700
rect 36652 35646 36654 35698
rect 36654 35646 36706 35698
rect 36706 35646 36708 35698
rect 36652 35644 36708 35646
rect 35308 35026 35364 35028
rect 35308 34974 35310 35026
rect 35310 34974 35362 35026
rect 35362 34974 35364 35026
rect 35308 34972 35364 34974
rect 30940 34636 30996 34692
rect 30044 32508 30100 32564
rect 30156 33964 30212 34020
rect 31388 34018 31444 34020
rect 31388 33966 31390 34018
rect 31390 33966 31442 34018
rect 31442 33966 31444 34018
rect 31388 33964 31444 33966
rect 32172 34018 32228 34020
rect 32172 33966 32174 34018
rect 32174 33966 32226 34018
rect 32226 33966 32228 34018
rect 32172 33964 32228 33966
rect 33404 33964 33460 34020
rect 31268 33684 31324 33740
rect 31372 33738 31428 33740
rect 31476 33738 31532 33740
rect 31372 33686 31396 33738
rect 31396 33686 31428 33738
rect 31476 33686 31520 33738
rect 31520 33686 31532 33738
rect 31372 33684 31428 33686
rect 31476 33684 31532 33686
rect 31580 33684 31636 33740
rect 31684 33738 31740 33740
rect 31788 33738 31844 33740
rect 31684 33686 31696 33738
rect 31696 33686 31740 33738
rect 31788 33686 31820 33738
rect 31820 33686 31844 33738
rect 31684 33684 31740 33686
rect 31788 33684 31844 33686
rect 31892 33684 31948 33740
rect 30156 32450 30212 32452
rect 30156 32398 30158 32450
rect 30158 32398 30210 32450
rect 30210 32398 30212 32450
rect 30156 32396 30212 32398
rect 28140 31724 28196 31780
rect 27916 30716 27972 30772
rect 28812 28588 28868 28644
rect 28252 28476 28308 28532
rect 28812 27634 28868 27636
rect 28812 27582 28814 27634
rect 28814 27582 28866 27634
rect 28866 27582 28868 27634
rect 28812 27580 28868 27582
rect 26908 25506 26964 25508
rect 26908 25454 26910 25506
rect 26910 25454 26962 25506
rect 26962 25454 26964 25506
rect 26908 25452 26964 25454
rect 27692 25282 27748 25284
rect 27692 25230 27694 25282
rect 27694 25230 27746 25282
rect 27746 25230 27748 25282
rect 27692 25228 27748 25230
rect 26768 25060 26824 25116
rect 26872 25114 26928 25116
rect 26976 25114 27032 25116
rect 26872 25062 26896 25114
rect 26896 25062 26928 25114
rect 26976 25062 27020 25114
rect 27020 25062 27032 25114
rect 26872 25060 26928 25062
rect 26976 25060 27032 25062
rect 27080 25060 27136 25116
rect 27184 25114 27240 25116
rect 27288 25114 27344 25116
rect 27184 25062 27196 25114
rect 27196 25062 27240 25114
rect 27288 25062 27320 25114
rect 27320 25062 27344 25114
rect 27184 25060 27240 25062
rect 27288 25060 27344 25062
rect 27392 25060 27448 25116
rect 26348 23378 26404 23380
rect 26348 23326 26350 23378
rect 26350 23326 26402 23378
rect 26402 23326 26404 23378
rect 26348 23324 26404 23326
rect 26768 23492 26824 23548
rect 26872 23546 26928 23548
rect 26976 23546 27032 23548
rect 26872 23494 26896 23546
rect 26896 23494 26928 23546
rect 26976 23494 27020 23546
rect 27020 23494 27032 23546
rect 26872 23492 26928 23494
rect 26976 23492 27032 23494
rect 27080 23492 27136 23548
rect 27184 23546 27240 23548
rect 27288 23546 27344 23548
rect 27184 23494 27196 23546
rect 27196 23494 27240 23546
rect 27288 23494 27320 23546
rect 27320 23494 27344 23546
rect 27184 23492 27240 23494
rect 27288 23492 27344 23494
rect 27392 23492 27448 23548
rect 27132 23324 27188 23380
rect 26768 21924 26824 21980
rect 26872 21978 26928 21980
rect 26976 21978 27032 21980
rect 26872 21926 26896 21978
rect 26896 21926 26928 21978
rect 26976 21926 27020 21978
rect 27020 21926 27032 21978
rect 26872 21924 26928 21926
rect 26976 21924 27032 21926
rect 27080 21924 27136 21980
rect 27184 21978 27240 21980
rect 27288 21978 27344 21980
rect 27184 21926 27196 21978
rect 27196 21926 27240 21978
rect 27288 21926 27320 21978
rect 27320 21926 27344 21978
rect 27184 21924 27240 21926
rect 27288 21924 27344 21926
rect 27392 21924 27448 21980
rect 27020 21474 27076 21476
rect 27020 21422 27022 21474
rect 27022 21422 27074 21474
rect 27074 21422 27076 21474
rect 27020 21420 27076 21422
rect 26572 20972 26628 21028
rect 27356 20972 27412 21028
rect 26768 20356 26824 20412
rect 26872 20410 26928 20412
rect 26976 20410 27032 20412
rect 26872 20358 26896 20410
rect 26896 20358 26928 20410
rect 26976 20358 27020 20410
rect 27020 20358 27032 20410
rect 26872 20356 26928 20358
rect 26976 20356 27032 20358
rect 27080 20356 27136 20412
rect 27184 20410 27240 20412
rect 27288 20410 27344 20412
rect 27184 20358 27196 20410
rect 27196 20358 27240 20410
rect 27288 20358 27320 20410
rect 27320 20358 27344 20410
rect 27184 20356 27240 20358
rect 27288 20356 27344 20358
rect 27392 20356 27448 20412
rect 27804 20076 27860 20132
rect 26768 18788 26824 18844
rect 26872 18842 26928 18844
rect 26976 18842 27032 18844
rect 26872 18790 26896 18842
rect 26896 18790 26928 18842
rect 26976 18790 27020 18842
rect 27020 18790 27032 18842
rect 26872 18788 26928 18790
rect 26976 18788 27032 18790
rect 27080 18788 27136 18844
rect 27184 18842 27240 18844
rect 27288 18842 27344 18844
rect 27184 18790 27196 18842
rect 27196 18790 27240 18842
rect 27288 18790 27320 18842
rect 27320 18790 27344 18842
rect 27184 18788 27240 18790
rect 27288 18788 27344 18790
rect 27392 18788 27448 18844
rect 26768 17220 26824 17276
rect 26872 17274 26928 17276
rect 26976 17274 27032 17276
rect 26872 17222 26896 17274
rect 26896 17222 26928 17274
rect 26976 17222 27020 17274
rect 27020 17222 27032 17274
rect 26872 17220 26928 17222
rect 26976 17220 27032 17222
rect 27080 17220 27136 17276
rect 27184 17274 27240 17276
rect 27288 17274 27344 17276
rect 27184 17222 27196 17274
rect 27196 17222 27240 17274
rect 27288 17222 27320 17274
rect 27320 17222 27344 17274
rect 27184 17220 27240 17222
rect 27288 17220 27344 17222
rect 27392 17220 27448 17276
rect 26768 15652 26824 15708
rect 26872 15706 26928 15708
rect 26976 15706 27032 15708
rect 26872 15654 26896 15706
rect 26896 15654 26928 15706
rect 26976 15654 27020 15706
rect 27020 15654 27032 15706
rect 26872 15652 26928 15654
rect 26976 15652 27032 15654
rect 27080 15652 27136 15708
rect 27184 15706 27240 15708
rect 27288 15706 27344 15708
rect 27184 15654 27196 15706
rect 27196 15654 27240 15706
rect 27288 15654 27320 15706
rect 27320 15654 27344 15706
rect 27184 15652 27240 15654
rect 27288 15652 27344 15654
rect 27392 15652 27448 15708
rect 27692 14306 27748 14308
rect 27692 14254 27694 14306
rect 27694 14254 27746 14306
rect 27746 14254 27748 14306
rect 27692 14252 27748 14254
rect 26768 14084 26824 14140
rect 26872 14138 26928 14140
rect 26976 14138 27032 14140
rect 26872 14086 26896 14138
rect 26896 14086 26928 14138
rect 26976 14086 27020 14138
rect 27020 14086 27032 14138
rect 26872 14084 26928 14086
rect 26976 14084 27032 14086
rect 27080 14084 27136 14140
rect 27184 14138 27240 14140
rect 27288 14138 27344 14140
rect 27184 14086 27196 14138
rect 27196 14086 27240 14138
rect 27288 14086 27320 14138
rect 27320 14086 27344 14138
rect 27184 14084 27240 14086
rect 27288 14084 27344 14086
rect 27392 14084 27448 14140
rect 26768 12516 26824 12572
rect 26872 12570 26928 12572
rect 26976 12570 27032 12572
rect 26872 12518 26896 12570
rect 26896 12518 26928 12570
rect 26976 12518 27020 12570
rect 27020 12518 27032 12570
rect 26872 12516 26928 12518
rect 26976 12516 27032 12518
rect 27080 12516 27136 12572
rect 27184 12570 27240 12572
rect 27288 12570 27344 12572
rect 27184 12518 27196 12570
rect 27196 12518 27240 12570
rect 27288 12518 27320 12570
rect 27320 12518 27344 12570
rect 27184 12516 27240 12518
rect 27288 12516 27344 12518
rect 27392 12516 27448 12572
rect 25788 11116 25844 11172
rect 26768 10948 26824 11004
rect 26872 11002 26928 11004
rect 26976 11002 27032 11004
rect 26872 10950 26896 11002
rect 26896 10950 26928 11002
rect 26976 10950 27020 11002
rect 27020 10950 27032 11002
rect 26872 10948 26928 10950
rect 26976 10948 27032 10950
rect 27080 10948 27136 11004
rect 27184 11002 27240 11004
rect 27288 11002 27344 11004
rect 27184 10950 27196 11002
rect 27196 10950 27240 11002
rect 27288 10950 27320 11002
rect 27320 10950 27344 11002
rect 27184 10948 27240 10950
rect 27288 10948 27344 10950
rect 27392 10948 27448 11004
rect 22268 10164 22324 10220
rect 22372 10218 22428 10220
rect 22476 10218 22532 10220
rect 22372 10166 22396 10218
rect 22396 10166 22428 10218
rect 22476 10166 22520 10218
rect 22520 10166 22532 10218
rect 22372 10164 22428 10166
rect 22476 10164 22532 10166
rect 22580 10164 22636 10220
rect 22684 10218 22740 10220
rect 22788 10218 22844 10220
rect 22684 10166 22696 10218
rect 22696 10166 22740 10218
rect 22788 10166 22820 10218
rect 22820 10166 22844 10218
rect 22684 10164 22740 10166
rect 22788 10164 22844 10166
rect 22892 10164 22948 10220
rect 28252 25452 28308 25508
rect 28588 24892 28644 24948
rect 28588 22258 28644 22260
rect 28588 22206 28590 22258
rect 28590 22206 28642 22258
rect 28642 22206 28644 22258
rect 28588 22204 28644 22206
rect 28364 21756 28420 21812
rect 29932 30770 29988 30772
rect 29932 30718 29934 30770
rect 29934 30718 29986 30770
rect 29986 30718 29988 30770
rect 29932 30716 29988 30718
rect 29596 28700 29652 28756
rect 29260 28476 29316 28532
rect 29148 28364 29204 28420
rect 30044 28588 30100 28644
rect 29932 27244 29988 27300
rect 29484 27186 29540 27188
rect 29484 27134 29486 27186
rect 29486 27134 29538 27186
rect 29538 27134 29540 27186
rect 29484 27132 29540 27134
rect 29708 26908 29764 26964
rect 32508 33122 32564 33124
rect 32508 33070 32510 33122
rect 32510 33070 32562 33122
rect 32562 33070 32564 33122
rect 32508 33068 32564 33070
rect 32508 32396 32564 32452
rect 31268 32116 31324 32172
rect 31372 32170 31428 32172
rect 31476 32170 31532 32172
rect 31372 32118 31396 32170
rect 31396 32118 31428 32170
rect 31476 32118 31520 32170
rect 31520 32118 31532 32170
rect 31372 32116 31428 32118
rect 31476 32116 31532 32118
rect 31580 32116 31636 32172
rect 31684 32170 31740 32172
rect 31788 32170 31844 32172
rect 31684 32118 31696 32170
rect 31696 32118 31740 32170
rect 31788 32118 31820 32170
rect 31820 32118 31844 32170
rect 31684 32116 31740 32118
rect 31788 32116 31844 32118
rect 31892 32116 31948 32172
rect 30604 31836 30660 31892
rect 32172 30940 32228 30996
rect 31724 30882 31780 30884
rect 31724 30830 31726 30882
rect 31726 30830 31778 30882
rect 31778 30830 31780 30882
rect 31724 30828 31780 30830
rect 31268 30548 31324 30604
rect 31372 30602 31428 30604
rect 31476 30602 31532 30604
rect 31372 30550 31396 30602
rect 31396 30550 31428 30602
rect 31476 30550 31520 30602
rect 31520 30550 31532 30602
rect 31372 30548 31428 30550
rect 31476 30548 31532 30550
rect 31580 30548 31636 30604
rect 31684 30602 31740 30604
rect 31788 30602 31844 30604
rect 31684 30550 31696 30602
rect 31696 30550 31740 30602
rect 31788 30550 31820 30602
rect 31820 30550 31844 30602
rect 31684 30548 31740 30550
rect 31788 30548 31844 30550
rect 31892 30548 31948 30604
rect 30268 30210 30324 30212
rect 30268 30158 30270 30210
rect 30270 30158 30322 30210
rect 30322 30158 30324 30210
rect 30268 30156 30324 30158
rect 30268 28700 30324 28756
rect 30940 30156 30996 30212
rect 33180 30828 33236 30884
rect 32732 30210 32788 30212
rect 32732 30158 32734 30210
rect 32734 30158 32786 30210
rect 32786 30158 32788 30210
rect 32732 30156 32788 30158
rect 33068 30156 33124 30212
rect 31268 28980 31324 29036
rect 31372 29034 31428 29036
rect 31476 29034 31532 29036
rect 31372 28982 31396 29034
rect 31396 28982 31428 29034
rect 31476 28982 31520 29034
rect 31520 28982 31532 29034
rect 31372 28980 31428 28982
rect 31476 28980 31532 28982
rect 31580 28980 31636 29036
rect 31684 29034 31740 29036
rect 31788 29034 31844 29036
rect 31684 28982 31696 29034
rect 31696 28982 31740 29034
rect 31788 28982 31820 29034
rect 31820 28982 31844 29034
rect 31684 28980 31740 28982
rect 31788 28980 31844 28982
rect 31892 28980 31948 29036
rect 32060 28476 32116 28532
rect 30940 28418 30996 28420
rect 30940 28366 30942 28418
rect 30942 28366 30994 28418
rect 30994 28366 30996 28418
rect 30940 28364 30996 28366
rect 32060 28140 32116 28196
rect 33180 29596 33236 29652
rect 33068 28140 33124 28196
rect 31268 27412 31324 27468
rect 31372 27466 31428 27468
rect 31476 27466 31532 27468
rect 31372 27414 31396 27466
rect 31396 27414 31428 27466
rect 31476 27414 31520 27466
rect 31520 27414 31532 27466
rect 31372 27412 31428 27414
rect 31476 27412 31532 27414
rect 31580 27412 31636 27468
rect 31684 27466 31740 27468
rect 31788 27466 31844 27468
rect 31684 27414 31696 27466
rect 31696 27414 31740 27466
rect 31788 27414 31820 27466
rect 31820 27414 31844 27466
rect 31684 27412 31740 27414
rect 31788 27412 31844 27414
rect 31892 27412 31948 27468
rect 30380 27132 30436 27188
rect 30492 27244 30548 27300
rect 30156 26908 30212 26964
rect 32060 27244 32116 27300
rect 32620 27244 32676 27300
rect 31164 27074 31220 27076
rect 31164 27022 31166 27074
rect 31166 27022 31218 27074
rect 31218 27022 31220 27074
rect 31164 27020 31220 27022
rect 32060 27020 32116 27076
rect 35532 34300 35588 34356
rect 35308 33852 35364 33908
rect 35756 34802 35812 34804
rect 35756 34750 35758 34802
rect 35758 34750 35810 34802
rect 35810 34750 35812 34802
rect 35756 34748 35812 34750
rect 37100 37826 37156 37828
rect 37100 37774 37102 37826
rect 37102 37774 37154 37826
rect 37154 37774 37156 37826
rect 37100 37772 37156 37774
rect 37324 37436 37380 37492
rect 38556 40572 38612 40628
rect 37996 37378 38052 37380
rect 37996 37326 37998 37378
rect 37998 37326 38050 37378
rect 38050 37326 38052 37378
rect 37996 37324 38052 37326
rect 38332 38220 38388 38276
rect 38444 37996 38500 38052
rect 39004 40626 39060 40628
rect 39004 40574 39006 40626
rect 39006 40574 39058 40626
rect 39058 40574 39060 40626
rect 39004 40572 39060 40574
rect 39564 41970 39620 41972
rect 39564 41918 39566 41970
rect 39566 41918 39618 41970
rect 39618 41918 39620 41970
rect 39564 41916 39620 41918
rect 39900 40908 39956 40964
rect 37100 36428 37156 36484
rect 37324 36482 37380 36484
rect 37324 36430 37326 36482
rect 37326 36430 37378 36482
rect 37378 36430 37380 36482
rect 37324 36428 37380 36430
rect 39228 37324 39284 37380
rect 39116 37154 39172 37156
rect 39116 37102 39118 37154
rect 39118 37102 39170 37154
rect 39170 37102 39172 37154
rect 39116 37100 39172 37102
rect 37660 36370 37716 36372
rect 37660 36318 37662 36370
rect 37662 36318 37714 36370
rect 37714 36318 37716 36370
rect 37660 36316 37716 36318
rect 37324 35922 37380 35924
rect 37324 35870 37326 35922
rect 37326 35870 37378 35922
rect 37378 35870 37380 35922
rect 37324 35868 37380 35870
rect 36988 35644 37044 35700
rect 37212 34860 37268 34916
rect 36204 34636 36260 34692
rect 35768 34468 35824 34524
rect 35872 34522 35928 34524
rect 35976 34522 36032 34524
rect 35872 34470 35896 34522
rect 35896 34470 35928 34522
rect 35976 34470 36020 34522
rect 36020 34470 36032 34522
rect 35872 34468 35928 34470
rect 35976 34468 36032 34470
rect 36080 34468 36136 34524
rect 36184 34522 36240 34524
rect 36288 34522 36344 34524
rect 36184 34470 36196 34522
rect 36196 34470 36240 34522
rect 36288 34470 36320 34522
rect 36320 34470 36344 34522
rect 36184 34468 36240 34470
rect 36288 34468 36344 34470
rect 36392 34468 36448 34524
rect 36988 34524 37044 34580
rect 38668 34914 38724 34916
rect 38668 34862 38670 34914
rect 38670 34862 38722 34914
rect 38722 34862 38724 34914
rect 38668 34860 38724 34862
rect 38892 35084 38948 35140
rect 39788 37266 39844 37268
rect 39788 37214 39790 37266
rect 39790 37214 39842 37266
rect 39842 37214 39844 37266
rect 39788 37212 39844 37214
rect 39564 37100 39620 37156
rect 39340 35698 39396 35700
rect 39340 35646 39342 35698
rect 39342 35646 39394 35698
rect 39394 35646 39396 35698
rect 39340 35644 39396 35646
rect 39116 34748 39172 34804
rect 39900 35084 39956 35140
rect 36428 34076 36484 34132
rect 38444 33516 38500 33572
rect 35868 33068 35924 33124
rect 35768 32900 35824 32956
rect 35872 32954 35928 32956
rect 35976 32954 36032 32956
rect 35872 32902 35896 32954
rect 35896 32902 35928 32954
rect 35976 32902 36020 32954
rect 36020 32902 36032 32954
rect 35872 32900 35928 32902
rect 35976 32900 36032 32902
rect 36080 32900 36136 32956
rect 36184 32954 36240 32956
rect 36288 32954 36344 32956
rect 36184 32902 36196 32954
rect 36196 32902 36240 32954
rect 36288 32902 36320 32954
rect 36320 32902 36344 32954
rect 36184 32900 36240 32902
rect 36288 32900 36344 32902
rect 36392 32900 36448 32956
rect 35980 32674 36036 32676
rect 35980 32622 35982 32674
rect 35982 32622 36034 32674
rect 36034 32622 36036 32674
rect 35980 32620 36036 32622
rect 35868 31666 35924 31668
rect 35868 31614 35870 31666
rect 35870 31614 35922 31666
rect 35922 31614 35924 31666
rect 35868 31612 35924 31614
rect 36316 31666 36372 31668
rect 36316 31614 36318 31666
rect 36318 31614 36370 31666
rect 36370 31614 36372 31666
rect 36316 31612 36372 31614
rect 36540 31666 36596 31668
rect 36540 31614 36542 31666
rect 36542 31614 36594 31666
rect 36594 31614 36596 31666
rect 36540 31612 36596 31614
rect 35768 31332 35824 31388
rect 35872 31386 35928 31388
rect 35976 31386 36032 31388
rect 35872 31334 35896 31386
rect 35896 31334 35928 31386
rect 35976 31334 36020 31386
rect 36020 31334 36032 31386
rect 35872 31332 35928 31334
rect 35976 31332 36032 31334
rect 36080 31332 36136 31388
rect 36184 31386 36240 31388
rect 36288 31386 36344 31388
rect 36184 31334 36196 31386
rect 36196 31334 36240 31386
rect 36288 31334 36320 31386
rect 36320 31334 36344 31386
rect 36184 31332 36240 31334
rect 36288 31332 36344 31334
rect 36392 31332 36448 31388
rect 33516 30994 33572 30996
rect 33516 30942 33518 30994
rect 33518 30942 33570 30994
rect 33570 30942 33572 30994
rect 33516 30940 33572 30942
rect 35868 30156 35924 30212
rect 35768 29764 35824 29820
rect 35872 29818 35928 29820
rect 35976 29818 36032 29820
rect 35872 29766 35896 29818
rect 35896 29766 35928 29818
rect 35976 29766 36020 29818
rect 36020 29766 36032 29818
rect 35872 29764 35928 29766
rect 35976 29764 36032 29766
rect 36080 29764 36136 29820
rect 36184 29818 36240 29820
rect 36288 29818 36344 29820
rect 36184 29766 36196 29818
rect 36196 29766 36240 29818
rect 36288 29766 36320 29818
rect 36320 29766 36344 29818
rect 36184 29764 36240 29766
rect 36288 29764 36344 29766
rect 36392 29764 36448 29820
rect 39564 34412 39620 34468
rect 40796 50594 40852 50596
rect 40796 50542 40798 50594
rect 40798 50542 40850 50594
rect 40850 50542 40852 50594
rect 40796 50540 40852 50542
rect 40460 50482 40516 50484
rect 40460 50430 40462 50482
rect 40462 50430 40514 50482
rect 40514 50430 40516 50482
rect 40460 50428 40516 50430
rect 41580 51436 41636 51492
rect 41692 52444 41748 52500
rect 44768 56420 44824 56476
rect 44872 56474 44928 56476
rect 44976 56474 45032 56476
rect 44872 56422 44896 56474
rect 44896 56422 44928 56474
rect 44976 56422 45020 56474
rect 45020 56422 45032 56474
rect 44872 56420 44928 56422
rect 44976 56420 45032 56422
rect 45080 56420 45136 56476
rect 45184 56474 45240 56476
rect 45288 56474 45344 56476
rect 45184 56422 45196 56474
rect 45196 56422 45240 56474
rect 45288 56422 45320 56474
rect 45320 56422 45344 56474
rect 45184 56420 45240 56422
rect 45288 56420 45344 56422
rect 45392 56420 45448 56476
rect 53768 56420 53824 56476
rect 53872 56474 53928 56476
rect 53976 56474 54032 56476
rect 53872 56422 53896 56474
rect 53896 56422 53928 56474
rect 53976 56422 54020 56474
rect 54020 56422 54032 56474
rect 53872 56420 53928 56422
rect 53976 56420 54032 56422
rect 54080 56420 54136 56476
rect 54184 56474 54240 56476
rect 54288 56474 54344 56476
rect 54184 56422 54196 56474
rect 54196 56422 54240 56474
rect 54288 56422 54320 56474
rect 54320 56422 54344 56474
rect 54184 56420 54240 56422
rect 54288 56420 54344 56422
rect 54392 56420 54448 56476
rect 62768 56420 62824 56476
rect 62872 56474 62928 56476
rect 62976 56474 63032 56476
rect 62872 56422 62896 56474
rect 62896 56422 62928 56474
rect 62976 56422 63020 56474
rect 63020 56422 63032 56474
rect 62872 56420 62928 56422
rect 62976 56420 63032 56422
rect 63080 56420 63136 56476
rect 63184 56474 63240 56476
rect 63288 56474 63344 56476
rect 63184 56422 63196 56474
rect 63196 56422 63240 56474
rect 63288 56422 63320 56474
rect 63320 56422 63344 56474
rect 63184 56420 63240 56422
rect 63288 56420 63344 56422
rect 63392 56420 63448 56476
rect 71768 56420 71824 56476
rect 71872 56474 71928 56476
rect 71976 56474 72032 56476
rect 71872 56422 71896 56474
rect 71896 56422 71928 56474
rect 71976 56422 72020 56474
rect 72020 56422 72032 56474
rect 71872 56420 71928 56422
rect 71976 56420 72032 56422
rect 72080 56420 72136 56476
rect 72184 56474 72240 56476
rect 72288 56474 72344 56476
rect 72184 56422 72196 56474
rect 72196 56422 72240 56474
rect 72288 56422 72320 56474
rect 72320 56422 72344 56474
rect 72184 56420 72240 56422
rect 72288 56420 72344 56422
rect 72392 56420 72448 56476
rect 80768 56420 80824 56476
rect 80872 56474 80928 56476
rect 80976 56474 81032 56476
rect 80872 56422 80896 56474
rect 80896 56422 80928 56474
rect 80976 56422 81020 56474
rect 81020 56422 81032 56474
rect 80872 56420 80928 56422
rect 80976 56420 81032 56422
rect 81080 56420 81136 56476
rect 81184 56474 81240 56476
rect 81288 56474 81344 56476
rect 81184 56422 81196 56474
rect 81196 56422 81240 56474
rect 81288 56422 81320 56474
rect 81320 56422 81344 56474
rect 81184 56420 81240 56422
rect 81288 56420 81344 56422
rect 81392 56420 81448 56476
rect 68348 56252 68404 56308
rect 69020 56252 69076 56308
rect 49268 55636 49324 55692
rect 49372 55690 49428 55692
rect 49476 55690 49532 55692
rect 49372 55638 49396 55690
rect 49396 55638 49428 55690
rect 49476 55638 49520 55690
rect 49520 55638 49532 55690
rect 49372 55636 49428 55638
rect 49476 55636 49532 55638
rect 49580 55636 49636 55692
rect 49684 55690 49740 55692
rect 49788 55690 49844 55692
rect 49684 55638 49696 55690
rect 49696 55638 49740 55690
rect 49788 55638 49820 55690
rect 49820 55638 49844 55690
rect 49684 55636 49740 55638
rect 49788 55636 49844 55638
rect 49892 55636 49948 55692
rect 67116 56028 67172 56084
rect 58268 55636 58324 55692
rect 58372 55690 58428 55692
rect 58476 55690 58532 55692
rect 58372 55638 58396 55690
rect 58396 55638 58428 55690
rect 58476 55638 58520 55690
rect 58520 55638 58532 55690
rect 58372 55636 58428 55638
rect 58476 55636 58532 55638
rect 58580 55636 58636 55692
rect 58684 55690 58740 55692
rect 58788 55690 58844 55692
rect 58684 55638 58696 55690
rect 58696 55638 58740 55690
rect 58788 55638 58820 55690
rect 58820 55638 58844 55690
rect 58684 55636 58740 55638
rect 58788 55636 58844 55638
rect 58892 55636 58948 55692
rect 43596 55244 43652 55300
rect 43260 54348 43316 54404
rect 43260 54124 43316 54180
rect 42700 52892 42756 52948
rect 42028 52668 42084 52724
rect 41692 51324 41748 51380
rect 42028 52108 42084 52164
rect 43260 52108 43316 52164
rect 42252 51378 42308 51380
rect 42252 51326 42254 51378
rect 42254 51326 42306 51378
rect 42306 51326 42308 51378
rect 42252 51324 42308 51326
rect 41132 49868 41188 49924
rect 43708 55298 43764 55300
rect 43708 55246 43710 55298
rect 43710 55246 43762 55298
rect 43762 55246 43764 55298
rect 43708 55244 43764 55246
rect 44268 55298 44324 55300
rect 44268 55246 44270 55298
rect 44270 55246 44322 55298
rect 44322 55246 44324 55298
rect 44268 55244 44324 55246
rect 45164 55298 45220 55300
rect 45164 55246 45166 55298
rect 45166 55246 45218 55298
rect 45218 55246 45220 55298
rect 45164 55244 45220 55246
rect 45948 55186 46004 55188
rect 45948 55134 45950 55186
rect 45950 55134 46002 55186
rect 46002 55134 46004 55186
rect 45948 55132 46004 55134
rect 44768 54852 44824 54908
rect 44872 54906 44928 54908
rect 44976 54906 45032 54908
rect 44872 54854 44896 54906
rect 44896 54854 44928 54906
rect 44976 54854 45020 54906
rect 45020 54854 45032 54906
rect 44872 54852 44928 54854
rect 44976 54852 45032 54854
rect 45080 54852 45136 54908
rect 45184 54906 45240 54908
rect 45288 54906 45344 54908
rect 45184 54854 45196 54906
rect 45196 54854 45240 54906
rect 45288 54854 45320 54906
rect 45320 54854 45344 54906
rect 45184 54852 45240 54854
rect 45288 54852 45344 54854
rect 45392 54852 45448 54908
rect 47740 54684 47796 54740
rect 44156 54572 44212 54628
rect 44604 54626 44660 54628
rect 44604 54574 44606 54626
rect 44606 54574 44658 54626
rect 44658 54574 44660 54626
rect 44604 54572 44660 54574
rect 48860 55132 48916 55188
rect 47964 54626 48020 54628
rect 47964 54574 47966 54626
rect 47966 54574 48018 54626
rect 48018 54574 48020 54626
rect 47964 54572 48020 54574
rect 44156 54402 44212 54404
rect 44156 54350 44158 54402
rect 44158 54350 44210 54402
rect 44210 54350 44212 54402
rect 44156 54348 44212 54350
rect 44940 54290 44996 54292
rect 44940 54238 44942 54290
rect 44942 54238 44994 54290
rect 44994 54238 44996 54290
rect 44940 54236 44996 54238
rect 44828 54124 44884 54180
rect 44940 53730 44996 53732
rect 44940 53678 44942 53730
rect 44942 53678 44994 53730
rect 44994 53678 44996 53730
rect 44940 53676 44996 53678
rect 43708 52108 43764 52164
rect 43820 53004 43876 53060
rect 46732 53900 46788 53956
rect 45948 53676 46004 53732
rect 44768 53284 44824 53340
rect 44872 53338 44928 53340
rect 44976 53338 45032 53340
rect 44872 53286 44896 53338
rect 44896 53286 44928 53338
rect 44976 53286 45020 53338
rect 45020 53286 45032 53338
rect 44872 53284 44928 53286
rect 44976 53284 45032 53286
rect 45080 53284 45136 53340
rect 45184 53338 45240 53340
rect 45288 53338 45344 53340
rect 45184 53286 45196 53338
rect 45196 53286 45240 53338
rect 45288 53286 45320 53338
rect 45320 53286 45344 53338
rect 45184 53284 45240 53286
rect 45288 53284 45344 53286
rect 45392 53284 45448 53340
rect 45500 53058 45556 53060
rect 45500 53006 45502 53058
rect 45502 53006 45554 53058
rect 45554 53006 45556 53058
rect 45500 53004 45556 53006
rect 43932 52444 43988 52500
rect 44716 52556 44772 52612
rect 46060 53004 46116 53060
rect 45612 52556 45668 52612
rect 46172 52444 46228 52500
rect 45948 52162 46004 52164
rect 45948 52110 45950 52162
rect 45950 52110 46002 52162
rect 46002 52110 46004 52162
rect 45948 52108 46004 52110
rect 46620 52108 46676 52164
rect 46396 51996 46452 52052
rect 46172 51884 46228 51940
rect 44768 51716 44824 51772
rect 44872 51770 44928 51772
rect 44976 51770 45032 51772
rect 44872 51718 44896 51770
rect 44896 51718 44928 51770
rect 44976 51718 45020 51770
rect 45020 51718 45032 51770
rect 44872 51716 44928 51718
rect 44976 51716 45032 51718
rect 45080 51716 45136 51772
rect 45184 51770 45240 51772
rect 45288 51770 45344 51772
rect 45184 51718 45196 51770
rect 45196 51718 45240 51770
rect 45288 51718 45320 51770
rect 45320 51718 45344 51770
rect 45184 51716 45240 51718
rect 45288 51716 45344 51718
rect 45392 51716 45448 51772
rect 44604 51548 44660 51604
rect 43596 50764 43652 50820
rect 46396 51378 46452 51380
rect 46396 51326 46398 51378
rect 46398 51326 46450 51378
rect 46450 51326 46452 51378
rect 46396 51324 46452 51326
rect 45500 50594 45556 50596
rect 45500 50542 45502 50594
rect 45502 50542 45554 50594
rect 45554 50542 45556 50594
rect 45500 50540 45556 50542
rect 46172 50594 46228 50596
rect 46172 50542 46174 50594
rect 46174 50542 46226 50594
rect 46226 50542 46228 50594
rect 46172 50540 46228 50542
rect 43596 50428 43652 50484
rect 46060 50482 46116 50484
rect 46060 50430 46062 50482
rect 46062 50430 46114 50482
rect 46114 50430 46116 50482
rect 46060 50428 46116 50430
rect 44768 50148 44824 50204
rect 44872 50202 44928 50204
rect 44976 50202 45032 50204
rect 44872 50150 44896 50202
rect 44896 50150 44928 50202
rect 44976 50150 45020 50202
rect 45020 50150 45032 50202
rect 44872 50148 44928 50150
rect 44976 50148 45032 50150
rect 45080 50148 45136 50204
rect 45184 50202 45240 50204
rect 45288 50202 45344 50204
rect 45184 50150 45196 50202
rect 45196 50150 45240 50202
rect 45288 50150 45320 50202
rect 45320 50150 45344 50202
rect 45184 50148 45240 50150
rect 45288 50148 45344 50150
rect 45392 50148 45448 50204
rect 42252 49644 42308 49700
rect 40268 49364 40324 49420
rect 40372 49418 40428 49420
rect 40476 49418 40532 49420
rect 40372 49366 40396 49418
rect 40396 49366 40428 49418
rect 40476 49366 40520 49418
rect 40520 49366 40532 49418
rect 40372 49364 40428 49366
rect 40476 49364 40532 49366
rect 40580 49364 40636 49420
rect 40684 49418 40740 49420
rect 40788 49418 40844 49420
rect 40684 49366 40696 49418
rect 40696 49366 40740 49418
rect 40788 49366 40820 49418
rect 40820 49366 40844 49418
rect 40684 49364 40740 49366
rect 40788 49364 40844 49366
rect 40892 49364 40948 49420
rect 41020 48466 41076 48468
rect 41020 48414 41022 48466
rect 41022 48414 41074 48466
rect 41074 48414 41076 48466
rect 41020 48412 41076 48414
rect 40460 48018 40516 48020
rect 40460 47966 40462 48018
rect 40462 47966 40514 48018
rect 40514 47966 40516 48018
rect 40460 47964 40516 47966
rect 40268 47796 40324 47852
rect 40372 47850 40428 47852
rect 40476 47850 40532 47852
rect 40372 47798 40396 47850
rect 40396 47798 40428 47850
rect 40476 47798 40520 47850
rect 40520 47798 40532 47850
rect 40372 47796 40428 47798
rect 40476 47796 40532 47798
rect 40580 47796 40636 47852
rect 40684 47850 40740 47852
rect 40788 47850 40844 47852
rect 40684 47798 40696 47850
rect 40696 47798 40740 47850
rect 40788 47798 40820 47850
rect 40820 47798 40844 47850
rect 40684 47796 40740 47798
rect 40788 47796 40844 47798
rect 40892 47796 40948 47852
rect 41020 47068 41076 47124
rect 40236 46508 40292 46564
rect 41020 46562 41076 46564
rect 41020 46510 41022 46562
rect 41022 46510 41074 46562
rect 41074 46510 41076 46562
rect 41020 46508 41076 46510
rect 40268 46228 40324 46284
rect 40372 46282 40428 46284
rect 40476 46282 40532 46284
rect 40372 46230 40396 46282
rect 40396 46230 40428 46282
rect 40476 46230 40520 46282
rect 40520 46230 40532 46282
rect 40372 46228 40428 46230
rect 40476 46228 40532 46230
rect 40580 46228 40636 46284
rect 40684 46282 40740 46284
rect 40788 46282 40844 46284
rect 40684 46230 40696 46282
rect 40696 46230 40740 46282
rect 40788 46230 40820 46282
rect 40820 46230 40844 46282
rect 40684 46228 40740 46230
rect 40788 46228 40844 46230
rect 40892 46228 40948 46284
rect 40684 45890 40740 45892
rect 40684 45838 40686 45890
rect 40686 45838 40738 45890
rect 40738 45838 40740 45890
rect 40684 45836 40740 45838
rect 40236 45778 40292 45780
rect 40236 45726 40238 45778
rect 40238 45726 40290 45778
rect 40290 45726 40292 45778
rect 40236 45724 40292 45726
rect 41020 45724 41076 45780
rect 40268 44660 40324 44716
rect 40372 44714 40428 44716
rect 40476 44714 40532 44716
rect 40372 44662 40396 44714
rect 40396 44662 40428 44714
rect 40476 44662 40520 44714
rect 40520 44662 40532 44714
rect 40372 44660 40428 44662
rect 40476 44660 40532 44662
rect 40580 44660 40636 44716
rect 40684 44714 40740 44716
rect 40788 44714 40844 44716
rect 40684 44662 40696 44714
rect 40696 44662 40740 44714
rect 40788 44662 40820 44714
rect 40820 44662 40844 44714
rect 40684 44660 40740 44662
rect 40788 44660 40844 44662
rect 40892 44660 40948 44716
rect 40908 44156 40964 44212
rect 40268 43092 40324 43148
rect 40372 43146 40428 43148
rect 40476 43146 40532 43148
rect 40372 43094 40396 43146
rect 40396 43094 40428 43146
rect 40476 43094 40520 43146
rect 40520 43094 40532 43146
rect 40372 43092 40428 43094
rect 40476 43092 40532 43094
rect 40580 43092 40636 43148
rect 40684 43146 40740 43148
rect 40788 43146 40844 43148
rect 40684 43094 40696 43146
rect 40696 43094 40740 43146
rect 40788 43094 40820 43146
rect 40820 43094 40844 43146
rect 40684 43092 40740 43094
rect 40788 43092 40844 43094
rect 40892 43092 40948 43148
rect 41020 41916 41076 41972
rect 40268 41524 40324 41580
rect 40372 41578 40428 41580
rect 40476 41578 40532 41580
rect 40372 41526 40396 41578
rect 40396 41526 40428 41578
rect 40476 41526 40520 41578
rect 40520 41526 40532 41578
rect 40372 41524 40428 41526
rect 40476 41524 40532 41526
rect 40580 41524 40636 41580
rect 40684 41578 40740 41580
rect 40788 41578 40844 41580
rect 40684 41526 40696 41578
rect 40696 41526 40740 41578
rect 40788 41526 40820 41578
rect 40820 41526 40844 41578
rect 40684 41524 40740 41526
rect 40788 41524 40844 41526
rect 40892 41524 40948 41580
rect 40348 40290 40404 40292
rect 40348 40238 40350 40290
rect 40350 40238 40402 40290
rect 40402 40238 40404 40290
rect 40348 40236 40404 40238
rect 40268 39956 40324 40012
rect 40372 40010 40428 40012
rect 40476 40010 40532 40012
rect 40372 39958 40396 40010
rect 40396 39958 40428 40010
rect 40476 39958 40520 40010
rect 40520 39958 40532 40010
rect 40372 39956 40428 39958
rect 40476 39956 40532 39958
rect 40580 39956 40636 40012
rect 40684 40010 40740 40012
rect 40788 40010 40844 40012
rect 40684 39958 40696 40010
rect 40696 39958 40740 40010
rect 40788 39958 40820 40010
rect 40820 39958 40844 40010
rect 40684 39956 40740 39958
rect 40788 39956 40844 39958
rect 40892 39956 40948 40012
rect 40268 38388 40324 38444
rect 40372 38442 40428 38444
rect 40476 38442 40532 38444
rect 40372 38390 40396 38442
rect 40396 38390 40428 38442
rect 40476 38390 40520 38442
rect 40520 38390 40532 38442
rect 40372 38388 40428 38390
rect 40476 38388 40532 38390
rect 40580 38388 40636 38444
rect 40684 38442 40740 38444
rect 40788 38442 40844 38444
rect 40684 38390 40696 38442
rect 40696 38390 40740 38442
rect 40788 38390 40820 38442
rect 40820 38390 40844 38442
rect 40684 38388 40740 38390
rect 40788 38388 40844 38390
rect 40892 38388 40948 38444
rect 40460 37548 40516 37604
rect 41020 37266 41076 37268
rect 41020 37214 41022 37266
rect 41022 37214 41074 37266
rect 41074 37214 41076 37266
rect 41020 37212 41076 37214
rect 40268 36820 40324 36876
rect 40372 36874 40428 36876
rect 40476 36874 40532 36876
rect 40372 36822 40396 36874
rect 40396 36822 40428 36874
rect 40476 36822 40520 36874
rect 40520 36822 40532 36874
rect 40372 36820 40428 36822
rect 40476 36820 40532 36822
rect 40580 36820 40636 36876
rect 40684 36874 40740 36876
rect 40788 36874 40844 36876
rect 40684 36822 40696 36874
rect 40696 36822 40740 36874
rect 40788 36822 40820 36874
rect 40820 36822 40844 36874
rect 40684 36820 40740 36822
rect 40788 36820 40844 36822
rect 40892 36820 40948 36876
rect 40268 35252 40324 35308
rect 40372 35306 40428 35308
rect 40476 35306 40532 35308
rect 40372 35254 40396 35306
rect 40396 35254 40428 35306
rect 40476 35254 40520 35306
rect 40520 35254 40532 35306
rect 40372 35252 40428 35254
rect 40476 35252 40532 35254
rect 40580 35252 40636 35308
rect 40684 35306 40740 35308
rect 40788 35306 40844 35308
rect 40684 35254 40696 35306
rect 40696 35254 40740 35306
rect 40788 35254 40820 35306
rect 40820 35254 40844 35306
rect 40684 35252 40740 35254
rect 40788 35252 40844 35254
rect 40892 35252 40948 35308
rect 40796 34972 40852 35028
rect 40124 34412 40180 34468
rect 41804 47068 41860 47124
rect 41580 46508 41636 46564
rect 41356 45106 41412 45108
rect 41356 45054 41358 45106
rect 41358 45054 41410 45106
rect 41410 45054 41412 45106
rect 41356 45052 41412 45054
rect 41468 41244 41524 41300
rect 41916 45836 41972 45892
rect 41916 45276 41972 45332
rect 42140 44940 42196 44996
rect 41804 44156 41860 44212
rect 42140 41244 42196 41300
rect 41580 40514 41636 40516
rect 41580 40462 41582 40514
rect 41582 40462 41634 40514
rect 41634 40462 41636 40514
rect 41580 40460 41636 40462
rect 42028 41074 42084 41076
rect 42028 41022 42030 41074
rect 42030 41022 42082 41074
rect 42082 41022 42084 41074
rect 42028 41020 42084 41022
rect 41244 40236 41300 40292
rect 41244 38556 41300 38612
rect 41244 37548 41300 37604
rect 41356 38220 41412 38276
rect 41468 37826 41524 37828
rect 41468 37774 41470 37826
rect 41470 37774 41522 37826
rect 41522 37774 41524 37826
rect 41468 37772 41524 37774
rect 42812 49532 42868 49588
rect 44768 48580 44824 48636
rect 44872 48634 44928 48636
rect 44976 48634 45032 48636
rect 44872 48582 44896 48634
rect 44896 48582 44928 48634
rect 44976 48582 45020 48634
rect 45020 48582 45032 48634
rect 44872 48580 44928 48582
rect 44976 48580 45032 48582
rect 45080 48580 45136 48636
rect 45184 48634 45240 48636
rect 45288 48634 45344 48636
rect 45184 48582 45196 48634
rect 45196 48582 45240 48634
rect 45288 48582 45320 48634
rect 45320 48582 45344 48634
rect 45184 48580 45240 48582
rect 45288 48580 45344 48582
rect 45392 48580 45448 48636
rect 43260 47458 43316 47460
rect 43260 47406 43262 47458
rect 43262 47406 43314 47458
rect 43314 47406 43316 47458
rect 43260 47404 43316 47406
rect 42812 46956 42868 47012
rect 43708 47404 43764 47460
rect 43596 45164 43652 45220
rect 42700 44994 42756 44996
rect 42700 44942 42702 44994
rect 42702 44942 42754 44994
rect 42754 44942 42756 44994
rect 42700 44940 42756 44942
rect 42364 44156 42420 44212
rect 42364 41916 42420 41972
rect 42364 41298 42420 41300
rect 42364 41246 42366 41298
rect 42366 41246 42418 41298
rect 42418 41246 42420 41298
rect 42364 41244 42420 41246
rect 42700 40514 42756 40516
rect 42700 40462 42702 40514
rect 42702 40462 42754 40514
rect 42754 40462 42756 40514
rect 42700 40460 42756 40462
rect 42588 39340 42644 39396
rect 42028 38274 42084 38276
rect 42028 38222 42030 38274
rect 42030 38222 42082 38274
rect 42082 38222 42084 38274
rect 42028 38220 42084 38222
rect 41916 37772 41972 37828
rect 41916 37548 41972 37604
rect 41692 37324 41748 37380
rect 42028 37266 42084 37268
rect 42028 37214 42030 37266
rect 42030 37214 42082 37266
rect 42082 37214 42084 37266
rect 42028 37212 42084 37214
rect 41692 36988 41748 37044
rect 41244 34860 41300 34916
rect 39228 33516 39284 33572
rect 38556 32284 38612 32340
rect 40268 33684 40324 33740
rect 40372 33738 40428 33740
rect 40476 33738 40532 33740
rect 40372 33686 40396 33738
rect 40396 33686 40428 33738
rect 40476 33686 40520 33738
rect 40520 33686 40532 33738
rect 40372 33684 40428 33686
rect 40476 33684 40532 33686
rect 40580 33684 40636 33740
rect 40684 33738 40740 33740
rect 40788 33738 40844 33740
rect 40684 33686 40696 33738
rect 40696 33686 40740 33738
rect 40788 33686 40820 33738
rect 40820 33686 40844 33738
rect 40684 33684 40740 33686
rect 40788 33684 40844 33686
rect 40892 33684 40948 33740
rect 39900 32732 39956 32788
rect 36876 31164 36932 31220
rect 37100 30716 37156 30772
rect 36988 30156 37044 30212
rect 36652 29596 36708 29652
rect 34860 27970 34916 27972
rect 34860 27918 34862 27970
rect 34862 27918 34914 27970
rect 34914 27918 34916 27970
rect 34860 27916 34916 27918
rect 35196 27916 35252 27972
rect 35768 28196 35824 28252
rect 35872 28250 35928 28252
rect 35976 28250 36032 28252
rect 35872 28198 35896 28250
rect 35896 28198 35928 28250
rect 35976 28198 36020 28250
rect 36020 28198 36032 28250
rect 35872 28196 35928 28198
rect 35976 28196 36032 28198
rect 36080 28196 36136 28252
rect 36184 28250 36240 28252
rect 36288 28250 36344 28252
rect 36184 28198 36196 28250
rect 36196 28198 36240 28250
rect 36288 28198 36320 28250
rect 36320 28198 36344 28250
rect 36184 28196 36240 28198
rect 36288 28196 36344 28198
rect 36392 28196 36448 28252
rect 35196 26908 35252 26964
rect 31268 25844 31324 25900
rect 31372 25898 31428 25900
rect 31476 25898 31532 25900
rect 31372 25846 31396 25898
rect 31396 25846 31428 25898
rect 31476 25846 31520 25898
rect 31520 25846 31532 25898
rect 31372 25844 31428 25846
rect 31476 25844 31532 25846
rect 31580 25844 31636 25900
rect 31684 25898 31740 25900
rect 31788 25898 31844 25900
rect 31684 25846 31696 25898
rect 31696 25846 31740 25898
rect 31788 25846 31820 25898
rect 31820 25846 31844 25898
rect 31684 25844 31740 25846
rect 31788 25844 31844 25846
rect 31892 25844 31948 25900
rect 33068 25394 33124 25396
rect 33068 25342 33070 25394
rect 33070 25342 33122 25394
rect 33122 25342 33124 25394
rect 33068 25340 33124 25342
rect 30492 25004 30548 25060
rect 30156 24946 30212 24948
rect 30156 24894 30158 24946
rect 30158 24894 30210 24946
rect 30210 24894 30212 24946
rect 30156 24892 30212 24894
rect 29372 24780 29428 24836
rect 32060 25004 32116 25060
rect 30492 24834 30548 24836
rect 30492 24782 30494 24834
rect 30494 24782 30546 24834
rect 30546 24782 30548 24834
rect 30492 24780 30548 24782
rect 31268 24276 31324 24332
rect 31372 24330 31428 24332
rect 31476 24330 31532 24332
rect 31372 24278 31396 24330
rect 31396 24278 31428 24330
rect 31476 24278 31520 24330
rect 31520 24278 31532 24330
rect 31372 24276 31428 24278
rect 31476 24276 31532 24278
rect 31580 24276 31636 24332
rect 31684 24330 31740 24332
rect 31788 24330 31844 24332
rect 31684 24278 31696 24330
rect 31696 24278 31740 24330
rect 31788 24278 31820 24330
rect 31820 24278 31844 24330
rect 31684 24276 31740 24278
rect 31788 24276 31844 24278
rect 31892 24276 31948 24332
rect 32620 23826 32676 23828
rect 32620 23774 32622 23826
rect 32622 23774 32674 23826
rect 32674 23774 32676 23826
rect 32620 23772 32676 23774
rect 33068 23826 33124 23828
rect 33068 23774 33070 23826
rect 33070 23774 33122 23826
rect 33122 23774 33124 23826
rect 33068 23772 33124 23774
rect 30268 22930 30324 22932
rect 30268 22878 30270 22930
rect 30270 22878 30322 22930
rect 30322 22878 30324 22930
rect 30268 22876 30324 22878
rect 29708 22204 29764 22260
rect 29036 21756 29092 21812
rect 29372 21420 29428 21476
rect 29148 20972 29204 21028
rect 32284 23324 32340 23380
rect 32620 23324 32676 23380
rect 31268 22708 31324 22764
rect 31372 22762 31428 22764
rect 31476 22762 31532 22764
rect 31372 22710 31396 22762
rect 31396 22710 31428 22762
rect 31476 22710 31520 22762
rect 31520 22710 31532 22762
rect 31372 22708 31428 22710
rect 31476 22708 31532 22710
rect 31580 22708 31636 22764
rect 31684 22762 31740 22764
rect 31788 22762 31844 22764
rect 31684 22710 31696 22762
rect 31696 22710 31740 22762
rect 31788 22710 31820 22762
rect 31820 22710 31844 22762
rect 31684 22708 31740 22710
rect 31788 22708 31844 22710
rect 31892 22708 31948 22764
rect 30604 21756 30660 21812
rect 30156 21026 30212 21028
rect 30156 20974 30158 21026
rect 30158 20974 30210 21026
rect 30210 20974 30212 21026
rect 30156 20972 30212 20974
rect 28588 20802 28644 20804
rect 28588 20750 28590 20802
rect 28590 20750 28642 20802
rect 28642 20750 28644 20802
rect 28588 20748 28644 20750
rect 28588 20188 28644 20244
rect 28476 20130 28532 20132
rect 28476 20078 28478 20130
rect 28478 20078 28530 20130
rect 28530 20078 28532 20130
rect 28476 20076 28532 20078
rect 29372 20130 29428 20132
rect 29372 20078 29374 20130
rect 29374 20078 29426 20130
rect 29426 20078 29428 20130
rect 29372 20076 29428 20078
rect 31948 21810 32004 21812
rect 31948 21758 31950 21810
rect 31950 21758 32002 21810
rect 32002 21758 32004 21810
rect 31948 21756 32004 21758
rect 32508 21362 32564 21364
rect 32508 21310 32510 21362
rect 32510 21310 32562 21362
rect 32562 21310 32564 21362
rect 32508 21308 32564 21310
rect 31268 21140 31324 21196
rect 31372 21194 31428 21196
rect 31476 21194 31532 21196
rect 31372 21142 31396 21194
rect 31396 21142 31428 21194
rect 31476 21142 31520 21194
rect 31520 21142 31532 21194
rect 31372 21140 31428 21142
rect 31476 21140 31532 21142
rect 31580 21140 31636 21196
rect 31684 21194 31740 21196
rect 31788 21194 31844 21196
rect 31684 21142 31696 21194
rect 31696 21142 31740 21194
rect 31788 21142 31820 21194
rect 31820 21142 31844 21194
rect 31684 21140 31740 21142
rect 31788 21140 31844 21142
rect 31892 21140 31948 21196
rect 33068 21644 33124 21700
rect 32620 20748 32676 20804
rect 30604 20076 30660 20132
rect 31268 19572 31324 19628
rect 31372 19626 31428 19628
rect 31476 19626 31532 19628
rect 31372 19574 31396 19626
rect 31396 19574 31428 19626
rect 31476 19574 31520 19626
rect 31520 19574 31532 19626
rect 31372 19572 31428 19574
rect 31476 19572 31532 19574
rect 31580 19572 31636 19628
rect 31684 19626 31740 19628
rect 31788 19626 31844 19628
rect 31684 19574 31696 19626
rect 31696 19574 31740 19626
rect 31788 19574 31820 19626
rect 31820 19574 31844 19626
rect 31684 19572 31740 19574
rect 31788 19572 31844 19574
rect 31892 19572 31948 19628
rect 31268 18004 31324 18060
rect 31372 18058 31428 18060
rect 31476 18058 31532 18060
rect 31372 18006 31396 18058
rect 31396 18006 31428 18058
rect 31476 18006 31520 18058
rect 31520 18006 31532 18058
rect 31372 18004 31428 18006
rect 31476 18004 31532 18006
rect 31580 18004 31636 18060
rect 31684 18058 31740 18060
rect 31788 18058 31844 18060
rect 31684 18006 31696 18058
rect 31696 18006 31740 18058
rect 31788 18006 31820 18058
rect 31820 18006 31844 18058
rect 31684 18004 31740 18006
rect 31788 18004 31844 18006
rect 31892 18004 31948 18060
rect 31268 16436 31324 16492
rect 31372 16490 31428 16492
rect 31476 16490 31532 16492
rect 31372 16438 31396 16490
rect 31396 16438 31428 16490
rect 31476 16438 31520 16490
rect 31520 16438 31532 16490
rect 31372 16436 31428 16438
rect 31476 16436 31532 16438
rect 31580 16436 31636 16492
rect 31684 16490 31740 16492
rect 31788 16490 31844 16492
rect 31684 16438 31696 16490
rect 31696 16438 31740 16490
rect 31788 16438 31820 16490
rect 31820 16438 31844 16490
rect 31684 16436 31740 16438
rect 31788 16436 31844 16438
rect 31892 16436 31948 16492
rect 31268 14868 31324 14924
rect 31372 14922 31428 14924
rect 31476 14922 31532 14924
rect 31372 14870 31396 14922
rect 31396 14870 31428 14922
rect 31476 14870 31520 14922
rect 31520 14870 31532 14922
rect 31372 14868 31428 14870
rect 31476 14868 31532 14870
rect 31580 14868 31636 14924
rect 31684 14922 31740 14924
rect 31788 14922 31844 14924
rect 31684 14870 31696 14922
rect 31696 14870 31740 14922
rect 31788 14870 31820 14922
rect 31820 14870 31844 14922
rect 31684 14868 31740 14870
rect 31788 14868 31844 14870
rect 31892 14868 31948 14924
rect 31268 13300 31324 13356
rect 31372 13354 31428 13356
rect 31476 13354 31532 13356
rect 31372 13302 31396 13354
rect 31396 13302 31428 13354
rect 31476 13302 31520 13354
rect 31520 13302 31532 13354
rect 31372 13300 31428 13302
rect 31476 13300 31532 13302
rect 31580 13300 31636 13356
rect 31684 13354 31740 13356
rect 31788 13354 31844 13356
rect 31684 13302 31696 13354
rect 31696 13302 31740 13354
rect 31788 13302 31820 13354
rect 31820 13302 31844 13354
rect 31684 13300 31740 13302
rect 31788 13300 31844 13302
rect 31892 13300 31948 13356
rect 34188 25340 34244 25396
rect 34076 25282 34132 25284
rect 34076 25230 34078 25282
rect 34078 25230 34130 25282
rect 34130 25230 34132 25282
rect 34076 25228 34132 25230
rect 33852 24668 33908 24724
rect 34860 25340 34916 25396
rect 34972 25228 35028 25284
rect 33628 23324 33684 23380
rect 33628 22370 33684 22372
rect 33628 22318 33630 22370
rect 33630 22318 33682 22370
rect 33682 22318 33684 22370
rect 33628 22316 33684 22318
rect 33404 22092 33460 22148
rect 34188 22146 34244 22148
rect 34188 22094 34190 22146
rect 34190 22094 34242 22146
rect 34242 22094 34244 22146
rect 34188 22092 34244 22094
rect 33628 21308 33684 21364
rect 33740 20802 33796 20804
rect 33740 20750 33742 20802
rect 33742 20750 33794 20802
rect 33794 20750 33796 20802
rect 33740 20748 33796 20750
rect 34412 20636 34468 20692
rect 34748 24668 34804 24724
rect 34636 22316 34692 22372
rect 33292 12236 33348 12292
rect 30940 12012 30996 12068
rect 28028 9548 28084 9604
rect 28476 9660 28532 9716
rect 26768 9380 26824 9436
rect 26872 9434 26928 9436
rect 26976 9434 27032 9436
rect 26872 9382 26896 9434
rect 26896 9382 26928 9434
rect 26976 9382 27020 9434
rect 27020 9382 27032 9434
rect 26872 9380 26928 9382
rect 26976 9380 27032 9382
rect 27080 9380 27136 9436
rect 27184 9434 27240 9436
rect 27288 9434 27344 9436
rect 27184 9382 27196 9434
rect 27196 9382 27240 9434
rect 27288 9382 27320 9434
rect 27320 9382 27344 9434
rect 27184 9380 27240 9382
rect 27288 9380 27344 9382
rect 27392 9380 27448 9436
rect 22268 8596 22324 8652
rect 22372 8650 22428 8652
rect 22476 8650 22532 8652
rect 22372 8598 22396 8650
rect 22396 8598 22428 8650
rect 22476 8598 22520 8650
rect 22520 8598 22532 8650
rect 22372 8596 22428 8598
rect 22476 8596 22532 8598
rect 22580 8596 22636 8652
rect 22684 8650 22740 8652
rect 22788 8650 22844 8652
rect 22684 8598 22696 8650
rect 22696 8598 22740 8650
rect 22788 8598 22820 8650
rect 22820 8598 22844 8650
rect 22684 8596 22740 8598
rect 22788 8596 22844 8598
rect 22892 8596 22948 8652
rect 26768 7812 26824 7868
rect 26872 7866 26928 7868
rect 26976 7866 27032 7868
rect 26872 7814 26896 7866
rect 26896 7814 26928 7866
rect 26976 7814 27020 7866
rect 27020 7814 27032 7866
rect 26872 7812 26928 7814
rect 26976 7812 27032 7814
rect 27080 7812 27136 7868
rect 27184 7866 27240 7868
rect 27288 7866 27344 7868
rect 27184 7814 27196 7866
rect 27196 7814 27240 7866
rect 27288 7814 27320 7866
rect 27320 7814 27344 7866
rect 27184 7812 27240 7814
rect 27288 7812 27344 7814
rect 27392 7812 27448 7868
rect 22268 7028 22324 7084
rect 22372 7082 22428 7084
rect 22476 7082 22532 7084
rect 22372 7030 22396 7082
rect 22396 7030 22428 7082
rect 22476 7030 22520 7082
rect 22520 7030 22532 7082
rect 22372 7028 22428 7030
rect 22476 7028 22532 7030
rect 22580 7028 22636 7084
rect 22684 7082 22740 7084
rect 22788 7082 22844 7084
rect 22684 7030 22696 7082
rect 22696 7030 22740 7082
rect 22788 7030 22820 7082
rect 22820 7030 22844 7082
rect 22684 7028 22740 7030
rect 22788 7028 22844 7030
rect 22892 7028 22948 7084
rect 25116 6690 25172 6692
rect 25116 6638 25118 6690
rect 25118 6638 25170 6690
rect 25170 6638 25172 6690
rect 25116 6636 25172 6638
rect 25900 6690 25956 6692
rect 25900 6638 25902 6690
rect 25902 6638 25954 6690
rect 25954 6638 25956 6690
rect 25900 6636 25956 6638
rect 22268 5460 22324 5516
rect 22372 5514 22428 5516
rect 22476 5514 22532 5516
rect 22372 5462 22396 5514
rect 22396 5462 22428 5514
rect 22476 5462 22520 5514
rect 22520 5462 22532 5514
rect 22372 5460 22428 5462
rect 22476 5460 22532 5462
rect 22580 5460 22636 5516
rect 22684 5514 22740 5516
rect 22788 5514 22844 5516
rect 22684 5462 22696 5514
rect 22696 5462 22740 5514
rect 22788 5462 22820 5514
rect 22820 5462 22844 5514
rect 22684 5460 22740 5462
rect 22788 5460 22844 5462
rect 22892 5460 22948 5516
rect 20748 4060 20804 4116
rect 13268 3892 13324 3948
rect 13372 3946 13428 3948
rect 13476 3946 13532 3948
rect 13372 3894 13396 3946
rect 13396 3894 13428 3946
rect 13476 3894 13520 3946
rect 13520 3894 13532 3946
rect 13372 3892 13428 3894
rect 13476 3892 13532 3894
rect 13580 3892 13636 3948
rect 13684 3946 13740 3948
rect 13788 3946 13844 3948
rect 13684 3894 13696 3946
rect 13696 3894 13740 3946
rect 13788 3894 13820 3946
rect 13820 3894 13844 3946
rect 13684 3892 13740 3894
rect 13788 3892 13844 3894
rect 13892 3892 13948 3948
rect 22268 3892 22324 3948
rect 22372 3946 22428 3948
rect 22476 3946 22532 3948
rect 22372 3894 22396 3946
rect 22396 3894 22428 3946
rect 22476 3894 22520 3946
rect 22520 3894 22532 3946
rect 22372 3892 22428 3894
rect 22476 3892 22532 3894
rect 22580 3892 22636 3948
rect 22684 3946 22740 3948
rect 22788 3946 22844 3948
rect 22684 3894 22696 3946
rect 22696 3894 22740 3946
rect 22788 3894 22820 3946
rect 22820 3894 22844 3946
rect 22684 3892 22740 3894
rect 22788 3892 22844 3894
rect 22892 3892 22948 3948
rect 28364 6690 28420 6692
rect 28364 6638 28366 6690
rect 28366 6638 28418 6690
rect 28418 6638 28420 6690
rect 28364 6636 28420 6638
rect 26796 6412 26852 6468
rect 26768 6244 26824 6300
rect 26872 6298 26928 6300
rect 26976 6298 27032 6300
rect 26872 6246 26896 6298
rect 26896 6246 26928 6298
rect 26976 6246 27020 6298
rect 27020 6246 27032 6298
rect 26872 6244 26928 6246
rect 26976 6244 27032 6246
rect 27080 6244 27136 6300
rect 27184 6298 27240 6300
rect 27288 6298 27344 6300
rect 27184 6246 27196 6298
rect 27196 6246 27240 6298
rect 27288 6246 27320 6298
rect 27320 6246 27344 6298
rect 27184 6244 27240 6246
rect 27288 6244 27344 6246
rect 27392 6244 27448 6300
rect 26572 5234 26628 5236
rect 26572 5182 26574 5234
rect 26574 5182 26626 5234
rect 26626 5182 26628 5234
rect 26572 5180 26628 5182
rect 27916 5068 27972 5124
rect 30044 8988 30100 9044
rect 29372 6466 29428 6468
rect 29372 6414 29374 6466
rect 29374 6414 29426 6466
rect 29426 6414 29428 6466
rect 29372 6412 29428 6414
rect 30716 6636 30772 6692
rect 30156 4956 30212 5012
rect 26768 4676 26824 4732
rect 26872 4730 26928 4732
rect 26976 4730 27032 4732
rect 26872 4678 26896 4730
rect 26896 4678 26928 4730
rect 26976 4678 27020 4730
rect 27020 4678 27032 4730
rect 26872 4676 26928 4678
rect 26976 4676 27032 4678
rect 27080 4676 27136 4732
rect 27184 4730 27240 4732
rect 27288 4730 27344 4732
rect 27184 4678 27196 4730
rect 27196 4678 27240 4730
rect 27288 4678 27320 4730
rect 27320 4678 27344 4730
rect 27184 4676 27240 4678
rect 27288 4676 27344 4678
rect 27392 4676 27448 4732
rect 30156 4450 30212 4452
rect 30156 4398 30158 4450
rect 30158 4398 30210 4450
rect 30210 4398 30212 4450
rect 30156 4396 30212 4398
rect 31268 11732 31324 11788
rect 31372 11786 31428 11788
rect 31476 11786 31532 11788
rect 31372 11734 31396 11786
rect 31396 11734 31428 11786
rect 31476 11734 31520 11786
rect 31520 11734 31532 11786
rect 31372 11732 31428 11734
rect 31476 11732 31532 11734
rect 31580 11732 31636 11788
rect 31684 11786 31740 11788
rect 31788 11786 31844 11788
rect 31684 11734 31696 11786
rect 31696 11734 31740 11786
rect 31788 11734 31820 11786
rect 31820 11734 31844 11786
rect 31684 11732 31740 11734
rect 31788 11732 31844 11734
rect 31892 11732 31948 11788
rect 31164 11394 31220 11396
rect 31164 11342 31166 11394
rect 31166 11342 31218 11394
rect 31218 11342 31220 11394
rect 31164 11340 31220 11342
rect 31268 10164 31324 10220
rect 31372 10218 31428 10220
rect 31476 10218 31532 10220
rect 31372 10166 31396 10218
rect 31396 10166 31428 10218
rect 31476 10166 31520 10218
rect 31520 10166 31532 10218
rect 31372 10164 31428 10166
rect 31476 10164 31532 10166
rect 31580 10164 31636 10220
rect 31684 10218 31740 10220
rect 31788 10218 31844 10220
rect 31684 10166 31696 10218
rect 31696 10166 31740 10218
rect 31788 10166 31820 10218
rect 31820 10166 31844 10218
rect 31684 10164 31740 10166
rect 31788 10164 31844 10166
rect 31892 10164 31948 10220
rect 31948 9714 32004 9716
rect 31948 9662 31950 9714
rect 31950 9662 32002 9714
rect 32002 9662 32004 9714
rect 31948 9660 32004 9662
rect 31836 9042 31892 9044
rect 31836 8990 31838 9042
rect 31838 8990 31890 9042
rect 31890 8990 31892 9042
rect 31836 8988 31892 8990
rect 31268 8596 31324 8652
rect 31372 8650 31428 8652
rect 31476 8650 31532 8652
rect 31372 8598 31396 8650
rect 31396 8598 31428 8650
rect 31476 8598 31520 8650
rect 31520 8598 31532 8650
rect 31372 8596 31428 8598
rect 31476 8596 31532 8598
rect 31580 8596 31636 8652
rect 31684 8650 31740 8652
rect 31788 8650 31844 8652
rect 31684 8598 31696 8650
rect 31696 8598 31740 8650
rect 31788 8598 31820 8650
rect 31820 8598 31844 8650
rect 31684 8596 31740 8598
rect 31788 8596 31844 8598
rect 31892 8596 31948 8652
rect 32508 7474 32564 7476
rect 32508 7422 32510 7474
rect 32510 7422 32562 7474
rect 32562 7422 32564 7474
rect 32508 7420 32564 7422
rect 31268 7028 31324 7084
rect 31372 7082 31428 7084
rect 31476 7082 31532 7084
rect 31372 7030 31396 7082
rect 31396 7030 31428 7082
rect 31476 7030 31520 7082
rect 31520 7030 31532 7082
rect 31372 7028 31428 7030
rect 31476 7028 31532 7030
rect 31580 7028 31636 7084
rect 31684 7082 31740 7084
rect 31788 7082 31844 7084
rect 31684 7030 31696 7082
rect 31696 7030 31740 7082
rect 31788 7030 31820 7082
rect 31820 7030 31844 7082
rect 31684 7028 31740 7030
rect 31788 7028 31844 7030
rect 31892 7028 31948 7084
rect 33516 6748 33572 6804
rect 33740 6188 33796 6244
rect 33404 5852 33460 5908
rect 31268 5460 31324 5516
rect 31372 5514 31428 5516
rect 31476 5514 31532 5516
rect 31372 5462 31396 5514
rect 31396 5462 31428 5514
rect 31476 5462 31520 5514
rect 31520 5462 31532 5514
rect 31372 5460 31428 5462
rect 31476 5460 31532 5462
rect 31580 5460 31636 5516
rect 31684 5514 31740 5516
rect 31788 5514 31844 5516
rect 31684 5462 31696 5514
rect 31696 5462 31740 5514
rect 31788 5462 31820 5514
rect 31820 5462 31844 5514
rect 31684 5460 31740 5462
rect 31788 5460 31844 5462
rect 31892 5460 31948 5516
rect 33292 5292 33348 5348
rect 25900 3724 25956 3780
rect 28812 3724 28868 3780
rect 32508 4284 32564 4340
rect 31268 3892 31324 3948
rect 31372 3946 31428 3948
rect 31476 3946 31532 3948
rect 31372 3894 31396 3946
rect 31396 3894 31428 3946
rect 31476 3894 31520 3946
rect 31520 3894 31532 3946
rect 31372 3892 31428 3894
rect 31476 3892 31532 3894
rect 31580 3892 31636 3948
rect 31684 3946 31740 3948
rect 31788 3946 31844 3948
rect 31684 3894 31696 3946
rect 31696 3894 31740 3946
rect 31788 3894 31820 3946
rect 31820 3894 31844 3946
rect 31684 3892 31740 3894
rect 31788 3892 31844 3894
rect 31892 3892 31948 3948
rect 17836 3666 17892 3668
rect 17836 3614 17838 3666
rect 17838 3614 17890 3666
rect 17890 3614 17892 3666
rect 17836 3612 17892 3614
rect 31724 3554 31780 3556
rect 31724 3502 31726 3554
rect 31726 3502 31778 3554
rect 31778 3502 31780 3554
rect 31724 3500 31780 3502
rect 33068 4172 33124 4228
rect 34300 8146 34356 8148
rect 34300 8094 34302 8146
rect 34302 8094 34354 8146
rect 34354 8094 34356 8146
rect 34300 8092 34356 8094
rect 34636 7586 34692 7588
rect 34636 7534 34638 7586
rect 34638 7534 34690 7586
rect 34690 7534 34692 7586
rect 34636 7532 34692 7534
rect 33852 6076 33908 6132
rect 33964 6748 34020 6804
rect 33852 5906 33908 5908
rect 33852 5854 33854 5906
rect 33854 5854 33906 5906
rect 33906 5854 33908 5906
rect 33852 5852 33908 5854
rect 34748 6860 34804 6916
rect 34412 6578 34468 6580
rect 34412 6526 34414 6578
rect 34414 6526 34466 6578
rect 34466 6526 34468 6578
rect 34412 6524 34468 6526
rect 34300 6188 34356 6244
rect 38892 31500 38948 31556
rect 39788 32620 39844 32676
rect 41244 33852 41300 33908
rect 41468 34412 41524 34468
rect 41020 32786 41076 32788
rect 41020 32734 41022 32786
rect 41022 32734 41074 32786
rect 41074 32734 41076 32786
rect 41020 32732 41076 32734
rect 41468 32620 41524 32676
rect 40236 32562 40292 32564
rect 40236 32510 40238 32562
rect 40238 32510 40290 32562
rect 40290 32510 40292 32562
rect 40236 32508 40292 32510
rect 39900 32284 39956 32340
rect 39788 31500 39844 31556
rect 37324 28700 37380 28756
rect 37996 27970 38052 27972
rect 37996 27918 37998 27970
rect 37998 27918 38050 27970
rect 38050 27918 38052 27970
rect 37996 27916 38052 27918
rect 37548 27186 37604 27188
rect 37548 27134 37550 27186
rect 37550 27134 37602 27186
rect 37602 27134 37604 27186
rect 37548 27132 37604 27134
rect 38108 27186 38164 27188
rect 38108 27134 38110 27186
rect 38110 27134 38162 27186
rect 38162 27134 38164 27186
rect 38108 27132 38164 27134
rect 36988 26850 37044 26852
rect 36988 26798 36990 26850
rect 36990 26798 37042 26850
rect 37042 26798 37044 26850
rect 36988 26796 37044 26798
rect 35768 26628 35824 26684
rect 35872 26682 35928 26684
rect 35976 26682 36032 26684
rect 35872 26630 35896 26682
rect 35896 26630 35928 26682
rect 35976 26630 36020 26682
rect 36020 26630 36032 26682
rect 35872 26628 35928 26630
rect 35976 26628 36032 26630
rect 36080 26628 36136 26684
rect 36184 26682 36240 26684
rect 36288 26682 36344 26684
rect 36184 26630 36196 26682
rect 36196 26630 36240 26682
rect 36288 26630 36320 26682
rect 36320 26630 36344 26682
rect 36184 26628 36240 26630
rect 36288 26628 36344 26630
rect 36392 26628 36448 26684
rect 35768 25060 35824 25116
rect 35872 25114 35928 25116
rect 35976 25114 36032 25116
rect 35872 25062 35896 25114
rect 35896 25062 35928 25114
rect 35976 25062 36020 25114
rect 36020 25062 36032 25114
rect 35872 25060 35928 25062
rect 35976 25060 36032 25062
rect 36080 25060 36136 25116
rect 36184 25114 36240 25116
rect 36288 25114 36344 25116
rect 36184 25062 36196 25114
rect 36196 25062 36240 25114
rect 36288 25062 36320 25114
rect 36320 25062 36344 25114
rect 36184 25060 36240 25062
rect 36288 25060 36344 25062
rect 36392 25060 36448 25116
rect 38780 30156 38836 30212
rect 38780 27132 38836 27188
rect 35196 24780 35252 24836
rect 35868 24834 35924 24836
rect 35868 24782 35870 24834
rect 35870 24782 35922 24834
rect 35922 24782 35924 24834
rect 35868 24780 35924 24782
rect 36652 24722 36708 24724
rect 36652 24670 36654 24722
rect 36654 24670 36706 24722
rect 36706 24670 36708 24722
rect 36652 24668 36708 24670
rect 35768 23492 35824 23548
rect 35872 23546 35928 23548
rect 35976 23546 36032 23548
rect 35872 23494 35896 23546
rect 35896 23494 35928 23546
rect 35976 23494 36020 23546
rect 36020 23494 36032 23546
rect 35872 23492 35928 23494
rect 35976 23492 36032 23494
rect 36080 23492 36136 23548
rect 36184 23546 36240 23548
rect 36288 23546 36344 23548
rect 36184 23494 36196 23546
rect 36196 23494 36240 23546
rect 36288 23494 36320 23546
rect 36320 23494 36344 23546
rect 36184 23492 36240 23494
rect 36288 23492 36344 23494
rect 36392 23492 36448 23548
rect 38108 24108 38164 24164
rect 37996 23324 38052 23380
rect 38108 22482 38164 22484
rect 38108 22430 38110 22482
rect 38110 22430 38162 22482
rect 38162 22430 38164 22482
rect 38108 22428 38164 22430
rect 35768 21924 35824 21980
rect 35872 21978 35928 21980
rect 35976 21978 36032 21980
rect 35872 21926 35896 21978
rect 35896 21926 35928 21978
rect 35976 21926 36020 21978
rect 36020 21926 36032 21978
rect 35872 21924 35928 21926
rect 35976 21924 36032 21926
rect 36080 21924 36136 21980
rect 36184 21978 36240 21980
rect 36288 21978 36344 21980
rect 36184 21926 36196 21978
rect 36196 21926 36240 21978
rect 36288 21926 36320 21978
rect 36320 21926 36344 21978
rect 36184 21924 36240 21926
rect 36288 21924 36344 21926
rect 36392 21924 36448 21980
rect 36204 21698 36260 21700
rect 36204 21646 36206 21698
rect 36206 21646 36258 21698
rect 36258 21646 36260 21698
rect 36204 21644 36260 21646
rect 36988 20636 37044 20692
rect 35768 20356 35824 20412
rect 35872 20410 35928 20412
rect 35976 20410 36032 20412
rect 35872 20358 35896 20410
rect 35896 20358 35928 20410
rect 35976 20358 36020 20410
rect 36020 20358 36032 20410
rect 35872 20356 35928 20358
rect 35976 20356 36032 20358
rect 36080 20356 36136 20412
rect 36184 20410 36240 20412
rect 36288 20410 36344 20412
rect 36184 20358 36196 20410
rect 36196 20358 36240 20410
rect 36288 20358 36320 20410
rect 36320 20358 36344 20410
rect 36184 20356 36240 20358
rect 36288 20356 36344 20358
rect 36392 20356 36448 20412
rect 35768 18788 35824 18844
rect 35872 18842 35928 18844
rect 35976 18842 36032 18844
rect 35872 18790 35896 18842
rect 35896 18790 35928 18842
rect 35976 18790 36020 18842
rect 36020 18790 36032 18842
rect 35872 18788 35928 18790
rect 35976 18788 36032 18790
rect 36080 18788 36136 18844
rect 36184 18842 36240 18844
rect 36288 18842 36344 18844
rect 36184 18790 36196 18842
rect 36196 18790 36240 18842
rect 36288 18790 36320 18842
rect 36320 18790 36344 18842
rect 36184 18788 36240 18790
rect 36288 18788 36344 18790
rect 36392 18788 36448 18844
rect 35768 17220 35824 17276
rect 35872 17274 35928 17276
rect 35976 17274 36032 17276
rect 35872 17222 35896 17274
rect 35896 17222 35928 17274
rect 35976 17222 36020 17274
rect 36020 17222 36032 17274
rect 35872 17220 35928 17222
rect 35976 17220 36032 17222
rect 36080 17220 36136 17276
rect 36184 17274 36240 17276
rect 36288 17274 36344 17276
rect 36184 17222 36196 17274
rect 36196 17222 36240 17274
rect 36288 17222 36320 17274
rect 36320 17222 36344 17274
rect 36184 17220 36240 17222
rect 36288 17220 36344 17222
rect 36392 17220 36448 17276
rect 35768 15652 35824 15708
rect 35872 15706 35928 15708
rect 35976 15706 36032 15708
rect 35872 15654 35896 15706
rect 35896 15654 35928 15706
rect 35976 15654 36020 15706
rect 36020 15654 36032 15706
rect 35872 15652 35928 15654
rect 35976 15652 36032 15654
rect 36080 15652 36136 15708
rect 36184 15706 36240 15708
rect 36288 15706 36344 15708
rect 36184 15654 36196 15706
rect 36196 15654 36240 15706
rect 36288 15654 36320 15706
rect 36320 15654 36344 15706
rect 36184 15652 36240 15654
rect 36288 15652 36344 15654
rect 36392 15652 36448 15708
rect 39228 24498 39284 24500
rect 39228 24446 39230 24498
rect 39230 24446 39282 24498
rect 39282 24446 39284 24498
rect 39228 24444 39284 24446
rect 40268 32116 40324 32172
rect 40372 32170 40428 32172
rect 40476 32170 40532 32172
rect 40372 32118 40396 32170
rect 40396 32118 40428 32170
rect 40476 32118 40520 32170
rect 40520 32118 40532 32170
rect 40372 32116 40428 32118
rect 40476 32116 40532 32118
rect 40580 32116 40636 32172
rect 40684 32170 40740 32172
rect 40788 32170 40844 32172
rect 40684 32118 40696 32170
rect 40696 32118 40740 32170
rect 40788 32118 40820 32170
rect 40820 32118 40844 32170
rect 40684 32116 40740 32118
rect 40788 32116 40844 32118
rect 40892 32116 40948 32172
rect 41468 31778 41524 31780
rect 41468 31726 41470 31778
rect 41470 31726 41522 31778
rect 41522 31726 41524 31778
rect 41468 31724 41524 31726
rect 41580 32732 41636 32788
rect 43260 44156 43316 44212
rect 43260 43650 43316 43652
rect 43260 43598 43262 43650
rect 43262 43598 43314 43650
rect 43314 43598 43316 43650
rect 43260 43596 43316 43598
rect 43596 38892 43652 38948
rect 42364 38108 42420 38164
rect 42700 37154 42756 37156
rect 42700 37102 42702 37154
rect 42702 37102 42754 37154
rect 42754 37102 42756 37154
rect 42700 37100 42756 37102
rect 43372 37772 43428 37828
rect 43372 37378 43428 37380
rect 43372 37326 43374 37378
rect 43374 37326 43426 37378
rect 43426 37326 43428 37378
rect 43372 37324 43428 37326
rect 43036 37100 43092 37156
rect 42924 36204 42980 36260
rect 41804 32284 41860 32340
rect 42364 32732 42420 32788
rect 41692 31948 41748 32004
rect 40684 31500 40740 31556
rect 40268 30548 40324 30604
rect 40372 30602 40428 30604
rect 40476 30602 40532 30604
rect 40372 30550 40396 30602
rect 40396 30550 40428 30602
rect 40476 30550 40520 30602
rect 40520 30550 40532 30602
rect 40372 30548 40428 30550
rect 40476 30548 40532 30550
rect 40580 30548 40636 30604
rect 40684 30602 40740 30604
rect 40788 30602 40844 30604
rect 40684 30550 40696 30602
rect 40696 30550 40740 30602
rect 40788 30550 40820 30602
rect 40820 30550 40844 30602
rect 40684 30548 40740 30550
rect 40788 30548 40844 30550
rect 40892 30548 40948 30604
rect 40012 29708 40068 29764
rect 41692 29148 41748 29204
rect 40268 28980 40324 29036
rect 40372 29034 40428 29036
rect 40476 29034 40532 29036
rect 40372 28982 40396 29034
rect 40396 28982 40428 29034
rect 40476 28982 40520 29034
rect 40520 28982 40532 29034
rect 40372 28980 40428 28982
rect 40476 28980 40532 28982
rect 40580 28980 40636 29036
rect 40684 29034 40740 29036
rect 40788 29034 40844 29036
rect 40684 28982 40696 29034
rect 40696 28982 40740 29034
rect 40788 28982 40820 29034
rect 40820 28982 40844 29034
rect 40684 28980 40740 28982
rect 40788 28980 40844 28982
rect 40892 28980 40948 29036
rect 40268 27412 40324 27468
rect 40372 27466 40428 27468
rect 40476 27466 40532 27468
rect 40372 27414 40396 27466
rect 40396 27414 40428 27466
rect 40476 27414 40520 27466
rect 40520 27414 40532 27466
rect 40372 27412 40428 27414
rect 40476 27412 40532 27414
rect 40580 27412 40636 27468
rect 40684 27466 40740 27468
rect 40788 27466 40844 27468
rect 40684 27414 40696 27466
rect 40696 27414 40740 27466
rect 40788 27414 40820 27466
rect 40820 27414 40844 27466
rect 40684 27412 40740 27414
rect 40788 27412 40844 27414
rect 40892 27412 40948 27468
rect 38780 23548 38836 23604
rect 38668 22876 38724 22932
rect 38556 22428 38612 22484
rect 39004 21532 39060 21588
rect 40268 25844 40324 25900
rect 40372 25898 40428 25900
rect 40476 25898 40532 25900
rect 40372 25846 40396 25898
rect 40396 25846 40428 25898
rect 40476 25846 40520 25898
rect 40520 25846 40532 25898
rect 40372 25844 40428 25846
rect 40476 25844 40532 25846
rect 40580 25844 40636 25900
rect 40684 25898 40740 25900
rect 40788 25898 40844 25900
rect 40684 25846 40696 25898
rect 40696 25846 40740 25898
rect 40788 25846 40820 25898
rect 40820 25846 40844 25898
rect 40684 25844 40740 25846
rect 40788 25844 40844 25846
rect 40892 25844 40948 25900
rect 41580 24780 41636 24836
rect 40124 24444 40180 24500
rect 40268 24276 40324 24332
rect 40372 24330 40428 24332
rect 40476 24330 40532 24332
rect 40372 24278 40396 24330
rect 40396 24278 40428 24330
rect 40476 24278 40520 24330
rect 40520 24278 40532 24330
rect 40372 24276 40428 24278
rect 40476 24276 40532 24278
rect 40580 24276 40636 24332
rect 40684 24330 40740 24332
rect 40788 24330 40844 24332
rect 40684 24278 40696 24330
rect 40696 24278 40740 24330
rect 40788 24278 40820 24330
rect 40820 24278 40844 24330
rect 40684 24276 40740 24278
rect 40788 24276 40844 24278
rect 40892 24276 40948 24332
rect 40236 23660 40292 23716
rect 40012 23548 40068 23604
rect 41580 23548 41636 23604
rect 40268 22708 40324 22764
rect 40372 22762 40428 22764
rect 40476 22762 40532 22764
rect 40372 22710 40396 22762
rect 40396 22710 40428 22762
rect 40476 22710 40520 22762
rect 40520 22710 40532 22762
rect 40372 22708 40428 22710
rect 40476 22708 40532 22710
rect 40580 22708 40636 22764
rect 40684 22762 40740 22764
rect 40788 22762 40844 22764
rect 40684 22710 40696 22762
rect 40696 22710 40740 22762
rect 40788 22710 40820 22762
rect 40820 22710 40844 22762
rect 40684 22708 40740 22710
rect 40788 22708 40844 22710
rect 40892 22708 40948 22764
rect 39900 21756 39956 21812
rect 39004 20972 39060 21028
rect 39228 20802 39284 20804
rect 39228 20750 39230 20802
rect 39230 20750 39282 20802
rect 39282 20750 39284 20802
rect 39228 20748 39284 20750
rect 40268 21140 40324 21196
rect 40372 21194 40428 21196
rect 40476 21194 40532 21196
rect 40372 21142 40396 21194
rect 40396 21142 40428 21194
rect 40476 21142 40520 21194
rect 40520 21142 40532 21194
rect 40372 21140 40428 21142
rect 40476 21140 40532 21142
rect 40580 21140 40636 21196
rect 40684 21194 40740 21196
rect 40788 21194 40844 21196
rect 40684 21142 40696 21194
rect 40696 21142 40740 21194
rect 40788 21142 40820 21194
rect 40820 21142 40844 21194
rect 40684 21140 40740 21142
rect 40788 21140 40844 21142
rect 40892 21140 40948 21196
rect 40124 20748 40180 20804
rect 40236 20188 40292 20244
rect 40460 20018 40516 20020
rect 40460 19966 40462 20018
rect 40462 19966 40514 20018
rect 40514 19966 40516 20018
rect 40460 19964 40516 19966
rect 40268 19572 40324 19628
rect 40372 19626 40428 19628
rect 40476 19626 40532 19628
rect 40372 19574 40396 19626
rect 40396 19574 40428 19626
rect 40476 19574 40520 19626
rect 40520 19574 40532 19626
rect 40372 19572 40428 19574
rect 40476 19572 40532 19574
rect 40580 19572 40636 19628
rect 40684 19626 40740 19628
rect 40788 19626 40844 19628
rect 40684 19574 40696 19626
rect 40696 19574 40740 19626
rect 40788 19574 40820 19626
rect 40820 19574 40844 19626
rect 40684 19572 40740 19574
rect 40788 19572 40844 19574
rect 40892 19572 40948 19628
rect 40012 19234 40068 19236
rect 40012 19182 40014 19234
rect 40014 19182 40066 19234
rect 40066 19182 40068 19234
rect 40012 19180 40068 19182
rect 42924 32732 42980 32788
rect 42364 32002 42420 32004
rect 42364 31950 42366 32002
rect 42366 31950 42418 32002
rect 42418 31950 42420 32002
rect 42364 31948 42420 31950
rect 42700 31724 42756 31780
rect 43372 31724 43428 31780
rect 42140 30210 42196 30212
rect 42140 30158 42142 30210
rect 42142 30158 42194 30210
rect 42194 30158 42196 30210
rect 42140 30156 42196 30158
rect 42476 30044 42532 30100
rect 43596 30098 43652 30100
rect 43596 30046 43598 30098
rect 43598 30046 43650 30098
rect 43650 30046 43652 30098
rect 43596 30044 43652 30046
rect 46060 47346 46116 47348
rect 46060 47294 46062 47346
rect 46062 47294 46114 47346
rect 46114 47294 46116 47346
rect 46060 47292 46116 47294
rect 44768 47012 44824 47068
rect 44872 47066 44928 47068
rect 44976 47066 45032 47068
rect 44872 47014 44896 47066
rect 44896 47014 44928 47066
rect 44976 47014 45020 47066
rect 45020 47014 45032 47066
rect 44872 47012 44928 47014
rect 44976 47012 45032 47014
rect 45080 47012 45136 47068
rect 45184 47066 45240 47068
rect 45288 47066 45344 47068
rect 45184 47014 45196 47066
rect 45196 47014 45240 47066
rect 45288 47014 45320 47066
rect 45320 47014 45344 47066
rect 45184 47012 45240 47014
rect 45288 47012 45344 47014
rect 45392 47012 45448 47068
rect 44768 45444 44824 45500
rect 44872 45498 44928 45500
rect 44976 45498 45032 45500
rect 44872 45446 44896 45498
rect 44896 45446 44928 45498
rect 44976 45446 45020 45498
rect 45020 45446 45032 45498
rect 44872 45444 44928 45446
rect 44976 45444 45032 45446
rect 45080 45444 45136 45500
rect 45184 45498 45240 45500
rect 45288 45498 45344 45500
rect 45184 45446 45196 45498
rect 45196 45446 45240 45498
rect 45288 45446 45320 45498
rect 45320 45446 45344 45498
rect 45184 45444 45240 45446
rect 45288 45444 45344 45446
rect 45392 45444 45448 45500
rect 44492 45330 44548 45332
rect 44492 45278 44494 45330
rect 44494 45278 44546 45330
rect 44546 45278 44548 45330
rect 44492 45276 44548 45278
rect 45276 45276 45332 45332
rect 43820 45218 43876 45220
rect 43820 45166 43822 45218
rect 43822 45166 43874 45218
rect 43874 45166 43876 45218
rect 43820 45164 43876 45166
rect 44768 43876 44824 43932
rect 44872 43930 44928 43932
rect 44976 43930 45032 43932
rect 44872 43878 44896 43930
rect 44896 43878 44928 43930
rect 44976 43878 45020 43930
rect 45020 43878 45032 43930
rect 44872 43876 44928 43878
rect 44976 43876 45032 43878
rect 45080 43876 45136 43932
rect 45184 43930 45240 43932
rect 45288 43930 45344 43932
rect 45184 43878 45196 43930
rect 45196 43878 45240 43930
rect 45288 43878 45320 43930
rect 45320 43878 45344 43930
rect 45184 43876 45240 43878
rect 45288 43876 45344 43878
rect 45392 43876 45448 43932
rect 46060 44268 46116 44324
rect 45836 43596 45892 43652
rect 46396 43650 46452 43652
rect 46396 43598 46398 43650
rect 46398 43598 46450 43650
rect 46450 43598 46452 43650
rect 46396 43596 46452 43598
rect 44768 42308 44824 42364
rect 44872 42362 44928 42364
rect 44976 42362 45032 42364
rect 44872 42310 44896 42362
rect 44896 42310 44928 42362
rect 44976 42310 45020 42362
rect 45020 42310 45032 42362
rect 44872 42308 44928 42310
rect 44976 42308 45032 42310
rect 45080 42308 45136 42364
rect 45184 42362 45240 42364
rect 45288 42362 45344 42364
rect 45184 42310 45196 42362
rect 45196 42310 45240 42362
rect 45288 42310 45320 42362
rect 45320 42310 45344 42362
rect 45184 42308 45240 42310
rect 45288 42308 45344 42310
rect 45392 42308 45448 42364
rect 44492 41970 44548 41972
rect 44492 41918 44494 41970
rect 44494 41918 44546 41970
rect 44546 41918 44548 41970
rect 44492 41916 44548 41918
rect 44268 41132 44324 41188
rect 45276 41186 45332 41188
rect 45276 41134 45278 41186
rect 45278 41134 45330 41186
rect 45330 41134 45332 41186
rect 45276 41132 45332 41134
rect 44768 40740 44824 40796
rect 44872 40794 44928 40796
rect 44976 40794 45032 40796
rect 44872 40742 44896 40794
rect 44896 40742 44928 40794
rect 44976 40742 45020 40794
rect 45020 40742 45032 40794
rect 44872 40740 44928 40742
rect 44976 40740 45032 40742
rect 45080 40740 45136 40796
rect 45184 40794 45240 40796
rect 45288 40794 45344 40796
rect 45184 40742 45196 40794
rect 45196 40742 45240 40794
rect 45288 40742 45320 40794
rect 45320 40742 45344 40794
rect 45184 40740 45240 40742
rect 45288 40740 45344 40742
rect 45392 40740 45448 40796
rect 45948 40514 46004 40516
rect 45948 40462 45950 40514
rect 45950 40462 46002 40514
rect 46002 40462 46004 40514
rect 45948 40460 46004 40462
rect 44768 39172 44824 39228
rect 44872 39226 44928 39228
rect 44976 39226 45032 39228
rect 44872 39174 44896 39226
rect 44896 39174 44928 39226
rect 44976 39174 45020 39226
rect 45020 39174 45032 39226
rect 44872 39172 44928 39174
rect 44976 39172 45032 39174
rect 45080 39172 45136 39228
rect 45184 39226 45240 39228
rect 45288 39226 45344 39228
rect 45184 39174 45196 39226
rect 45196 39174 45240 39226
rect 45288 39174 45320 39226
rect 45320 39174 45344 39226
rect 45184 39172 45240 39174
rect 45288 39172 45344 39174
rect 45392 39172 45448 39228
rect 43820 38946 43876 38948
rect 43820 38894 43822 38946
rect 43822 38894 43874 38946
rect 43874 38894 43876 38946
rect 43820 38892 43876 38894
rect 44492 38556 44548 38612
rect 45276 38556 45332 38612
rect 44768 37604 44824 37660
rect 44872 37658 44928 37660
rect 44976 37658 45032 37660
rect 44872 37606 44896 37658
rect 44896 37606 44928 37658
rect 44976 37606 45020 37658
rect 45020 37606 45032 37658
rect 44872 37604 44928 37606
rect 44976 37604 45032 37606
rect 45080 37604 45136 37660
rect 45184 37658 45240 37660
rect 45288 37658 45344 37660
rect 45184 37606 45196 37658
rect 45196 37606 45240 37658
rect 45288 37606 45320 37658
rect 45320 37606 45344 37658
rect 45184 37604 45240 37606
rect 45288 37604 45344 37606
rect 45392 37604 45448 37660
rect 45612 37212 45668 37268
rect 44156 37100 44212 37156
rect 44044 36204 44100 36260
rect 44768 36036 44824 36092
rect 44872 36090 44928 36092
rect 44976 36090 45032 36092
rect 44872 36038 44896 36090
rect 44896 36038 44928 36090
rect 44976 36038 45020 36090
rect 45020 36038 45032 36090
rect 44872 36036 44928 36038
rect 44976 36036 45032 36038
rect 45080 36036 45136 36092
rect 45184 36090 45240 36092
rect 45288 36090 45344 36092
rect 45184 36038 45196 36090
rect 45196 36038 45240 36090
rect 45288 36038 45320 36090
rect 45320 36038 45344 36090
rect 45184 36036 45240 36038
rect 45288 36036 45344 36038
rect 45392 36036 45448 36092
rect 45052 35586 45108 35588
rect 45052 35534 45054 35586
rect 45054 35534 45106 35586
rect 45106 35534 45108 35586
rect 45052 35532 45108 35534
rect 44604 34748 44660 34804
rect 44940 34802 44996 34804
rect 44940 34750 44942 34802
rect 44942 34750 44994 34802
rect 44994 34750 44996 34802
rect 44940 34748 44996 34750
rect 45388 34636 45444 34692
rect 44768 34468 44824 34524
rect 44872 34522 44928 34524
rect 44976 34522 45032 34524
rect 44872 34470 44896 34522
rect 44896 34470 44928 34522
rect 44976 34470 45020 34522
rect 45020 34470 45032 34522
rect 44872 34468 44928 34470
rect 44976 34468 45032 34470
rect 45080 34468 45136 34524
rect 45184 34522 45240 34524
rect 45288 34522 45344 34524
rect 45184 34470 45196 34522
rect 45196 34470 45240 34522
rect 45288 34470 45320 34522
rect 45320 34470 45344 34522
rect 45184 34468 45240 34470
rect 45288 34468 45344 34470
rect 45392 34468 45448 34524
rect 44156 33516 44212 33572
rect 43820 32562 43876 32564
rect 43820 32510 43822 32562
rect 43822 32510 43874 32562
rect 43874 32510 43876 32562
rect 43820 32508 43876 32510
rect 43820 31500 43876 31556
rect 44044 31836 44100 31892
rect 43708 29932 43764 29988
rect 43260 29260 43316 29316
rect 42140 29202 42196 29204
rect 42140 29150 42142 29202
rect 42142 29150 42194 29202
rect 42194 29150 42196 29202
rect 42140 29148 42196 29150
rect 44044 30156 44100 30212
rect 44156 30268 44212 30324
rect 44156 29708 44212 29764
rect 44156 29538 44212 29540
rect 44156 29486 44158 29538
rect 44158 29486 44210 29538
rect 44210 29486 44212 29538
rect 44156 29484 44212 29486
rect 44604 33516 44660 33572
rect 44492 32396 44548 32452
rect 44716 33404 44772 33460
rect 44940 33852 44996 33908
rect 51772 55020 51828 55076
rect 49756 54626 49812 54628
rect 49756 54574 49758 54626
rect 49758 54574 49810 54626
rect 49810 54574 49812 54626
rect 49756 54572 49812 54574
rect 48748 54514 48804 54516
rect 48748 54462 48750 54514
rect 48750 54462 48802 54514
rect 48802 54462 48804 54514
rect 48748 54460 48804 54462
rect 48076 54402 48132 54404
rect 48076 54350 48078 54402
rect 48078 54350 48130 54402
rect 48130 54350 48132 54402
rect 48076 54348 48132 54350
rect 47292 53116 47348 53172
rect 47740 53452 47796 53508
rect 47740 52556 47796 52612
rect 47180 52274 47236 52276
rect 47180 52222 47182 52274
rect 47182 52222 47234 52274
rect 47234 52222 47236 52274
rect 47180 52220 47236 52222
rect 48188 52892 48244 52948
rect 52780 55074 52836 55076
rect 52780 55022 52782 55074
rect 52782 55022 52834 55074
rect 52834 55022 52836 55074
rect 52780 55020 52836 55022
rect 52668 54460 52724 54516
rect 53116 55074 53172 55076
rect 53116 55022 53118 55074
rect 53118 55022 53170 55074
rect 53170 55022 53172 55074
rect 53116 55020 53172 55022
rect 53768 54852 53824 54908
rect 53872 54906 53928 54908
rect 53976 54906 54032 54908
rect 53872 54854 53896 54906
rect 53896 54854 53928 54906
rect 53976 54854 54020 54906
rect 54020 54854 54032 54906
rect 53872 54852 53928 54854
rect 53976 54852 54032 54854
rect 54080 54852 54136 54908
rect 54184 54906 54240 54908
rect 54288 54906 54344 54908
rect 54184 54854 54196 54906
rect 54196 54854 54240 54906
rect 54288 54854 54320 54906
rect 54320 54854 54344 54906
rect 54184 54852 54240 54854
rect 54288 54852 54344 54854
rect 54392 54852 54448 54908
rect 52892 54348 52948 54404
rect 49268 54068 49324 54124
rect 49372 54122 49428 54124
rect 49476 54122 49532 54124
rect 49372 54070 49396 54122
rect 49396 54070 49428 54122
rect 49476 54070 49520 54122
rect 49520 54070 49532 54122
rect 49372 54068 49428 54070
rect 49476 54068 49532 54070
rect 49580 54068 49636 54124
rect 49684 54122 49740 54124
rect 49788 54122 49844 54124
rect 49684 54070 49696 54122
rect 49696 54070 49740 54122
rect 49788 54070 49820 54122
rect 49820 54070 49844 54122
rect 49684 54068 49740 54070
rect 49788 54068 49844 54070
rect 49892 54068 49948 54124
rect 50092 53676 50148 53732
rect 46956 51996 47012 52052
rect 46732 51884 46788 51940
rect 49420 52946 49476 52948
rect 49420 52894 49422 52946
rect 49422 52894 49474 52946
rect 49474 52894 49476 52946
rect 49420 52892 49476 52894
rect 49084 52780 49140 52836
rect 49980 52722 50036 52724
rect 49980 52670 49982 52722
rect 49982 52670 50034 52722
rect 50034 52670 50036 52722
rect 49980 52668 50036 52670
rect 49084 52556 49140 52612
rect 48748 52444 48804 52500
rect 48300 52274 48356 52276
rect 48300 52222 48302 52274
rect 48302 52222 48354 52274
rect 48354 52222 48356 52274
rect 48300 52220 48356 52222
rect 49268 52500 49324 52556
rect 49372 52554 49428 52556
rect 49476 52554 49532 52556
rect 49372 52502 49396 52554
rect 49396 52502 49428 52554
rect 49476 52502 49520 52554
rect 49520 52502 49532 52554
rect 49372 52500 49428 52502
rect 49476 52500 49532 52502
rect 49580 52500 49636 52556
rect 49684 52554 49740 52556
rect 49788 52554 49844 52556
rect 49684 52502 49696 52554
rect 49696 52502 49740 52554
rect 49788 52502 49820 52554
rect 49820 52502 49844 52554
rect 49684 52500 49740 52502
rect 49788 52500 49844 52502
rect 49892 52500 49948 52556
rect 50204 53116 50260 53172
rect 50428 53564 50484 53620
rect 50204 52444 50260 52500
rect 49756 52386 49812 52388
rect 49756 52334 49758 52386
rect 49758 52334 49810 52386
rect 49810 52334 49812 52386
rect 49756 52332 49812 52334
rect 49644 52162 49700 52164
rect 49644 52110 49646 52162
rect 49646 52110 49698 52162
rect 49698 52110 49700 52162
rect 49644 52108 49700 52110
rect 47852 51884 47908 51940
rect 46732 51378 46788 51380
rect 46732 51326 46734 51378
rect 46734 51326 46786 51378
rect 46786 51326 46788 51378
rect 46732 51324 46788 51326
rect 47404 51378 47460 51380
rect 47404 51326 47406 51378
rect 47406 51326 47458 51378
rect 47458 51326 47460 51378
rect 47404 51324 47460 51326
rect 49268 50932 49324 50988
rect 49372 50986 49428 50988
rect 49476 50986 49532 50988
rect 49372 50934 49396 50986
rect 49396 50934 49428 50986
rect 49476 50934 49520 50986
rect 49520 50934 49532 50986
rect 49372 50932 49428 50934
rect 49476 50932 49532 50934
rect 49580 50932 49636 50988
rect 49684 50986 49740 50988
rect 49788 50986 49844 50988
rect 49684 50934 49696 50986
rect 49696 50934 49740 50986
rect 49788 50934 49820 50986
rect 49820 50934 49844 50986
rect 49684 50932 49740 50934
rect 49788 50932 49844 50934
rect 49892 50932 49948 50988
rect 49084 50482 49140 50484
rect 49084 50430 49086 50482
rect 49086 50430 49138 50482
rect 49138 50430 49140 50482
rect 49084 50428 49140 50430
rect 50428 52332 50484 52388
rect 50316 49868 50372 49924
rect 50428 50540 50484 50596
rect 52892 54124 52948 54180
rect 51212 53676 51268 53732
rect 50764 53452 50820 53508
rect 51100 53452 51156 53508
rect 50876 53116 50932 53172
rect 50764 52444 50820 52500
rect 51660 53564 51716 53620
rect 55580 54514 55636 54516
rect 55580 54462 55582 54514
rect 55582 54462 55634 54514
rect 55634 54462 55636 54514
rect 55580 54460 55636 54462
rect 54236 54124 54292 54180
rect 53900 53676 53956 53732
rect 53768 53284 53824 53340
rect 53872 53338 53928 53340
rect 53976 53338 54032 53340
rect 53872 53286 53896 53338
rect 53896 53286 53928 53338
rect 53976 53286 54020 53338
rect 54020 53286 54032 53338
rect 53872 53284 53928 53286
rect 53976 53284 54032 53286
rect 54080 53284 54136 53340
rect 54184 53338 54240 53340
rect 54288 53338 54344 53340
rect 54184 53286 54196 53338
rect 54196 53286 54240 53338
rect 54288 53286 54320 53338
rect 54320 53286 54344 53338
rect 54184 53284 54240 53286
rect 54288 53284 54344 53286
rect 54392 53284 54448 53340
rect 55580 52946 55636 52948
rect 55580 52894 55582 52946
rect 55582 52894 55634 52946
rect 55634 52894 55636 52946
rect 55580 52892 55636 52894
rect 54460 52780 54516 52836
rect 52444 52332 52500 52388
rect 53340 52332 53396 52388
rect 52108 52220 52164 52276
rect 53788 52274 53844 52276
rect 53788 52222 53790 52274
rect 53790 52222 53842 52274
rect 53842 52222 53844 52274
rect 53788 52220 53844 52222
rect 54348 52220 54404 52276
rect 55132 52834 55188 52836
rect 55132 52782 55134 52834
rect 55134 52782 55186 52834
rect 55186 52782 55188 52834
rect 55132 52780 55188 52782
rect 55132 52332 55188 52388
rect 55020 52220 55076 52276
rect 55692 52108 55748 52164
rect 57596 55074 57652 55076
rect 57596 55022 57598 55074
rect 57598 55022 57650 55074
rect 57650 55022 57652 55074
rect 57596 55020 57652 55022
rect 56812 54460 56868 54516
rect 56028 53452 56084 53508
rect 56140 54236 56196 54292
rect 56028 52668 56084 52724
rect 56812 54236 56868 54292
rect 56364 53506 56420 53508
rect 56364 53454 56366 53506
rect 56366 53454 56418 53506
rect 56418 53454 56420 53506
rect 56364 53452 56420 53454
rect 56476 53228 56532 53284
rect 57708 54572 57764 54628
rect 57820 54796 57876 54852
rect 57820 54402 57876 54404
rect 57820 54350 57822 54402
rect 57822 54350 57874 54402
rect 57874 54350 57876 54402
rect 57820 54348 57876 54350
rect 57484 54236 57540 54292
rect 57372 53788 57428 53844
rect 58380 54572 58436 54628
rect 60508 55020 60564 55076
rect 59164 54684 59220 54740
rect 58380 54236 58436 54292
rect 58268 54068 58324 54124
rect 58372 54122 58428 54124
rect 58476 54122 58532 54124
rect 58372 54070 58396 54122
rect 58396 54070 58428 54122
rect 58476 54070 58520 54122
rect 58520 54070 58532 54122
rect 58372 54068 58428 54070
rect 58476 54068 58532 54070
rect 58580 54068 58636 54124
rect 58684 54122 58740 54124
rect 58788 54122 58844 54124
rect 58684 54070 58696 54122
rect 58696 54070 58740 54122
rect 58788 54070 58820 54122
rect 58820 54070 58844 54122
rect 58684 54068 58740 54070
rect 58788 54068 58844 54070
rect 58892 54068 58948 54124
rect 58044 53788 58100 53844
rect 57820 53564 57876 53620
rect 57148 53004 57204 53060
rect 56588 52892 56644 52948
rect 56924 52668 56980 52724
rect 56812 52332 56868 52388
rect 55804 51996 55860 52052
rect 53768 51716 53824 51772
rect 53872 51770 53928 51772
rect 53976 51770 54032 51772
rect 53872 51718 53896 51770
rect 53896 51718 53928 51770
rect 53976 51718 54020 51770
rect 54020 51718 54032 51770
rect 53872 51716 53928 51718
rect 53976 51716 54032 51718
rect 54080 51716 54136 51772
rect 54184 51770 54240 51772
rect 54288 51770 54344 51772
rect 54184 51718 54196 51770
rect 54196 51718 54240 51770
rect 54288 51718 54320 51770
rect 54320 51718 54344 51770
rect 54184 51716 54240 51718
rect 54288 51716 54344 51718
rect 54392 51716 54448 51772
rect 56476 51996 56532 52052
rect 56812 52162 56868 52164
rect 56812 52110 56814 52162
rect 56814 52110 56866 52162
rect 56866 52110 56868 52162
rect 56812 52108 56868 52110
rect 57372 52668 57428 52724
rect 57484 53340 57540 53396
rect 57260 52332 57316 52388
rect 57708 53116 57764 53172
rect 54796 51212 54852 51268
rect 53768 50148 53824 50204
rect 53872 50202 53928 50204
rect 53976 50202 54032 50204
rect 53872 50150 53896 50202
rect 53896 50150 53928 50202
rect 53976 50150 54020 50202
rect 54020 50150 54032 50202
rect 53872 50148 53928 50150
rect 53976 50148 54032 50150
rect 54080 50148 54136 50204
rect 54184 50202 54240 50204
rect 54288 50202 54344 50204
rect 54184 50150 54196 50202
rect 54196 50150 54240 50202
rect 54288 50150 54320 50202
rect 54320 50150 54344 50202
rect 54184 50148 54240 50150
rect 54288 50148 54344 50150
rect 54392 50148 54448 50204
rect 51548 49922 51604 49924
rect 51548 49870 51550 49922
rect 51550 49870 51602 49922
rect 51602 49870 51604 49922
rect 51548 49868 51604 49870
rect 59500 54572 59556 54628
rect 59276 54236 59332 54292
rect 58044 53228 58100 53284
rect 58940 52946 58996 52948
rect 58940 52894 58942 52946
rect 58942 52894 58994 52946
rect 58994 52894 58996 52946
rect 58940 52892 58996 52894
rect 57932 52444 57988 52500
rect 58268 52500 58324 52556
rect 58372 52554 58428 52556
rect 58476 52554 58532 52556
rect 58372 52502 58396 52554
rect 58396 52502 58428 52554
rect 58476 52502 58520 52554
rect 58520 52502 58532 52554
rect 58372 52500 58428 52502
rect 58476 52500 58532 52502
rect 58580 52500 58636 52556
rect 58684 52554 58740 52556
rect 58788 52554 58844 52556
rect 58684 52502 58696 52554
rect 58696 52502 58740 52554
rect 58788 52502 58820 52554
rect 58820 52502 58844 52554
rect 58684 52500 58740 52502
rect 58788 52500 58844 52502
rect 58892 52500 58948 52556
rect 58492 52386 58548 52388
rect 58492 52334 58494 52386
rect 58494 52334 58546 52386
rect 58546 52334 58548 52386
rect 58492 52332 58548 52334
rect 58156 52220 58212 52276
rect 49268 49364 49324 49420
rect 49372 49418 49428 49420
rect 49476 49418 49532 49420
rect 49372 49366 49396 49418
rect 49396 49366 49428 49418
rect 49476 49366 49520 49418
rect 49520 49366 49532 49418
rect 49372 49364 49428 49366
rect 49476 49364 49532 49366
rect 49580 49364 49636 49420
rect 49684 49418 49740 49420
rect 49788 49418 49844 49420
rect 49684 49366 49696 49418
rect 49696 49366 49740 49418
rect 49788 49366 49820 49418
rect 49820 49366 49844 49418
rect 49684 49364 49740 49366
rect 49788 49364 49844 49366
rect 49892 49364 49948 49420
rect 53768 48580 53824 48636
rect 53872 48634 53928 48636
rect 53976 48634 54032 48636
rect 53872 48582 53896 48634
rect 53896 48582 53928 48634
rect 53976 48582 54020 48634
rect 54020 48582 54032 48634
rect 53872 48580 53928 48582
rect 53976 48580 54032 48582
rect 54080 48580 54136 48636
rect 54184 48634 54240 48636
rect 54288 48634 54344 48636
rect 54184 48582 54196 48634
rect 54196 48582 54240 48634
rect 54288 48582 54320 48634
rect 54320 48582 54344 48634
rect 54184 48580 54240 48582
rect 54288 48580 54344 48582
rect 54392 48580 54448 48636
rect 52332 48466 52388 48468
rect 52332 48414 52334 48466
rect 52334 48414 52386 48466
rect 52386 48414 52388 48466
rect 52332 48412 52388 48414
rect 52668 48412 52724 48468
rect 47740 47964 47796 48020
rect 47404 47458 47460 47460
rect 47404 47406 47406 47458
rect 47406 47406 47458 47458
rect 47458 47406 47460 47458
rect 47404 47404 47460 47406
rect 49268 47796 49324 47852
rect 49372 47850 49428 47852
rect 49476 47850 49532 47852
rect 49372 47798 49396 47850
rect 49396 47798 49428 47850
rect 49476 47798 49520 47850
rect 49520 47798 49532 47850
rect 49372 47796 49428 47798
rect 49476 47796 49532 47798
rect 49580 47796 49636 47852
rect 49684 47850 49740 47852
rect 49788 47850 49844 47852
rect 49684 47798 49696 47850
rect 49696 47798 49740 47850
rect 49788 47798 49820 47850
rect 49820 47798 49844 47850
rect 49684 47796 49740 47798
rect 49788 47796 49844 47798
rect 49892 47796 49948 47852
rect 48188 47516 48244 47572
rect 46956 47346 47012 47348
rect 46956 47294 46958 47346
rect 46958 47294 47010 47346
rect 47010 47294 47012 47346
rect 46956 47292 47012 47294
rect 47404 45836 47460 45892
rect 48748 47570 48804 47572
rect 48748 47518 48750 47570
rect 48750 47518 48802 47570
rect 48802 47518 48804 47570
rect 48748 47516 48804 47518
rect 50092 47516 50148 47572
rect 48860 47404 48916 47460
rect 47516 45612 47572 45668
rect 47516 45052 47572 45108
rect 46060 37772 46116 37828
rect 46396 37378 46452 37380
rect 46396 37326 46398 37378
rect 46398 37326 46450 37378
rect 46450 37326 46452 37378
rect 46396 37324 46452 37326
rect 47180 44268 47236 44324
rect 48076 44322 48132 44324
rect 48076 44270 48078 44322
rect 48078 44270 48130 44322
rect 48130 44270 48132 44322
rect 48076 44268 48132 44270
rect 47740 44210 47796 44212
rect 47740 44158 47742 44210
rect 47742 44158 47794 44210
rect 47794 44158 47796 44210
rect 47740 44156 47796 44158
rect 47628 43596 47684 43652
rect 48636 44210 48692 44212
rect 48636 44158 48638 44210
rect 48638 44158 48690 44210
rect 48690 44158 48692 44210
rect 48636 44156 48692 44158
rect 49196 47458 49252 47460
rect 49196 47406 49198 47458
rect 49198 47406 49250 47458
rect 49250 47406 49252 47458
rect 49196 47404 49252 47406
rect 49268 46228 49324 46284
rect 49372 46282 49428 46284
rect 49476 46282 49532 46284
rect 49372 46230 49396 46282
rect 49396 46230 49428 46282
rect 49476 46230 49520 46282
rect 49520 46230 49532 46282
rect 49372 46228 49428 46230
rect 49476 46228 49532 46230
rect 49580 46228 49636 46284
rect 49684 46282 49740 46284
rect 49788 46282 49844 46284
rect 49684 46230 49696 46282
rect 49696 46230 49740 46282
rect 49788 46230 49820 46282
rect 49820 46230 49844 46282
rect 49684 46228 49740 46230
rect 49788 46228 49844 46230
rect 49892 46228 49948 46284
rect 49196 45890 49252 45892
rect 49196 45838 49198 45890
rect 49198 45838 49250 45890
rect 49250 45838 49252 45890
rect 49196 45836 49252 45838
rect 49268 44660 49324 44716
rect 49372 44714 49428 44716
rect 49476 44714 49532 44716
rect 49372 44662 49396 44714
rect 49396 44662 49428 44714
rect 49476 44662 49520 44714
rect 49520 44662 49532 44714
rect 49372 44660 49428 44662
rect 49476 44660 49532 44662
rect 49580 44660 49636 44716
rect 49684 44714 49740 44716
rect 49788 44714 49844 44716
rect 49684 44662 49696 44714
rect 49696 44662 49740 44714
rect 49788 44662 49820 44714
rect 49820 44662 49844 44714
rect 49684 44660 49740 44662
rect 49788 44660 49844 44662
rect 49892 44660 49948 44716
rect 51436 46898 51492 46900
rect 51436 46846 51438 46898
rect 51438 46846 51490 46898
rect 51490 46846 51492 46898
rect 51436 46844 51492 46846
rect 52444 46844 52500 46900
rect 52220 46450 52276 46452
rect 52220 46398 52222 46450
rect 52222 46398 52274 46450
rect 52274 46398 52276 46450
rect 52220 46396 52276 46398
rect 52444 45388 52500 45444
rect 50316 45276 50372 45332
rect 48972 44156 49028 44212
rect 48412 40460 48468 40516
rect 47740 38946 47796 38948
rect 47740 38894 47742 38946
rect 47742 38894 47794 38946
rect 47794 38894 47796 38946
rect 47740 38892 47796 38894
rect 47180 37772 47236 37828
rect 45948 36092 46004 36148
rect 46396 36092 46452 36148
rect 46508 35532 46564 35588
rect 46620 35474 46676 35476
rect 46620 35422 46622 35474
rect 46622 35422 46674 35474
rect 46674 35422 46676 35474
rect 46620 35420 46676 35422
rect 46284 35308 46340 35364
rect 46620 35196 46676 35252
rect 46060 34914 46116 34916
rect 46060 34862 46062 34914
rect 46062 34862 46114 34914
rect 46114 34862 46116 34914
rect 46060 34860 46116 34862
rect 46284 34188 46340 34244
rect 44940 33068 44996 33124
rect 45164 33346 45220 33348
rect 45164 33294 45166 33346
rect 45166 33294 45218 33346
rect 45218 33294 45220 33346
rect 45164 33292 45220 33294
rect 44768 32900 44824 32956
rect 44872 32954 44928 32956
rect 44976 32954 45032 32956
rect 44872 32902 44896 32954
rect 44896 32902 44928 32954
rect 44976 32902 45020 32954
rect 45020 32902 45032 32954
rect 44872 32900 44928 32902
rect 44976 32900 45032 32902
rect 45080 32900 45136 32956
rect 45184 32954 45240 32956
rect 45288 32954 45344 32956
rect 45184 32902 45196 32954
rect 45196 32902 45240 32954
rect 45288 32902 45320 32954
rect 45320 32902 45344 32954
rect 45184 32900 45240 32902
rect 45288 32900 45344 32902
rect 45392 32900 45448 32956
rect 45612 31948 45668 32004
rect 44828 31778 44884 31780
rect 44828 31726 44830 31778
rect 44830 31726 44882 31778
rect 44882 31726 44884 31778
rect 44828 31724 44884 31726
rect 45388 31500 45444 31556
rect 44768 31332 44824 31388
rect 44872 31386 44928 31388
rect 44976 31386 45032 31388
rect 44872 31334 44896 31386
rect 44896 31334 44928 31386
rect 44976 31334 45020 31386
rect 45020 31334 45032 31386
rect 44872 31332 44928 31334
rect 44976 31332 45032 31334
rect 45080 31332 45136 31388
rect 45184 31386 45240 31388
rect 45288 31386 45344 31388
rect 45184 31334 45196 31386
rect 45196 31334 45240 31386
rect 45288 31334 45320 31386
rect 45320 31334 45344 31386
rect 45184 31332 45240 31334
rect 45288 31332 45344 31334
rect 45392 31332 45448 31388
rect 45052 30940 45108 30996
rect 44492 30268 44548 30324
rect 44604 30044 44660 30100
rect 45052 30210 45108 30212
rect 45052 30158 45054 30210
rect 45054 30158 45106 30210
rect 45106 30158 45108 30210
rect 45052 30156 45108 30158
rect 44940 30044 44996 30100
rect 45948 33458 46004 33460
rect 45948 33406 45950 33458
rect 45950 33406 46002 33458
rect 46002 33406 46004 33458
rect 45948 33404 46004 33406
rect 45836 31948 45892 32004
rect 46172 33292 46228 33348
rect 46620 34972 46676 35028
rect 48076 38220 48132 38276
rect 48188 38050 48244 38052
rect 48188 37998 48190 38050
rect 48190 37998 48242 38050
rect 48242 37998 48244 38050
rect 48188 37996 48244 37998
rect 48412 37996 48468 38052
rect 48748 37772 48804 37828
rect 47740 35810 47796 35812
rect 47740 35758 47742 35810
rect 47742 35758 47794 35810
rect 47794 35758 47796 35810
rect 47740 35756 47796 35758
rect 47068 35532 47124 35588
rect 47180 35420 47236 35476
rect 47068 34748 47124 34804
rect 46844 34636 46900 34692
rect 46620 34188 46676 34244
rect 46396 33122 46452 33124
rect 46396 33070 46398 33122
rect 46398 33070 46450 33122
rect 46450 33070 46452 33122
rect 46396 33068 46452 33070
rect 46172 31948 46228 32004
rect 46396 31836 46452 31892
rect 45724 30940 45780 30996
rect 46284 30828 46340 30884
rect 45724 30156 45780 30212
rect 44768 29764 44824 29820
rect 44872 29818 44928 29820
rect 44976 29818 45032 29820
rect 44872 29766 44896 29818
rect 44896 29766 44928 29818
rect 44976 29766 45020 29818
rect 45020 29766 45032 29818
rect 44872 29764 44928 29766
rect 44976 29764 45032 29766
rect 45080 29764 45136 29820
rect 45184 29818 45240 29820
rect 45288 29818 45344 29820
rect 45184 29766 45196 29818
rect 45196 29766 45240 29818
rect 45288 29766 45320 29818
rect 45320 29766 45344 29818
rect 45184 29764 45240 29766
rect 45288 29764 45344 29766
rect 45392 29764 45448 29820
rect 44716 29426 44772 29428
rect 44716 29374 44718 29426
rect 44718 29374 44770 29426
rect 44770 29374 44772 29426
rect 44716 29372 44772 29374
rect 44044 29260 44100 29316
rect 45500 29426 45556 29428
rect 45500 29374 45502 29426
rect 45502 29374 45554 29426
rect 45554 29374 45556 29426
rect 45500 29372 45556 29374
rect 43148 25506 43204 25508
rect 43148 25454 43150 25506
rect 43150 25454 43202 25506
rect 43202 25454 43204 25506
rect 43148 25452 43204 25454
rect 42700 25282 42756 25284
rect 42700 25230 42702 25282
rect 42702 25230 42754 25282
rect 42754 25230 42756 25282
rect 42700 25228 42756 25230
rect 43260 25340 43316 25396
rect 43820 25394 43876 25396
rect 43820 25342 43822 25394
rect 43822 25342 43874 25394
rect 43874 25342 43876 25394
rect 43820 25340 43876 25342
rect 43932 25116 43988 25172
rect 43932 24780 43988 24836
rect 42364 23714 42420 23716
rect 42364 23662 42366 23714
rect 42366 23662 42418 23714
rect 42418 23662 42420 23714
rect 42364 23660 42420 23662
rect 43372 21810 43428 21812
rect 43372 21758 43374 21810
rect 43374 21758 43426 21810
rect 43426 21758 43428 21810
rect 43372 21756 43428 21758
rect 42924 21532 42980 21588
rect 42140 20972 42196 21028
rect 43820 21810 43876 21812
rect 43820 21758 43822 21810
rect 43822 21758 43874 21810
rect 43874 21758 43876 21810
rect 43820 21756 43876 21758
rect 43596 21420 43652 21476
rect 43820 21362 43876 21364
rect 43820 21310 43822 21362
rect 43822 21310 43874 21362
rect 43874 21310 43876 21362
rect 43820 21308 43876 21310
rect 43932 20690 43988 20692
rect 43932 20638 43934 20690
rect 43934 20638 43986 20690
rect 43986 20638 43988 20690
rect 43932 20636 43988 20638
rect 44380 28642 44436 28644
rect 44380 28590 44382 28642
rect 44382 28590 44434 28642
rect 44434 28590 44436 28642
rect 44380 28588 44436 28590
rect 44768 28196 44824 28252
rect 44872 28250 44928 28252
rect 44976 28250 45032 28252
rect 44872 28198 44896 28250
rect 44896 28198 44928 28250
rect 44976 28198 45020 28250
rect 45020 28198 45032 28250
rect 44872 28196 44928 28198
rect 44976 28196 45032 28198
rect 45080 28196 45136 28252
rect 45184 28250 45240 28252
rect 45288 28250 45344 28252
rect 45184 28198 45196 28250
rect 45196 28198 45240 28250
rect 45288 28198 45320 28250
rect 45320 28198 45344 28250
rect 45184 28196 45240 28198
rect 45288 28196 45344 28198
rect 45392 28196 45448 28252
rect 46172 30044 46228 30100
rect 46508 30156 46564 30212
rect 46396 29484 46452 29540
rect 46060 29426 46116 29428
rect 46060 29374 46062 29426
rect 46062 29374 46114 29426
rect 46114 29374 46116 29426
rect 46060 29372 46116 29374
rect 45836 29260 45892 29316
rect 45836 28642 45892 28644
rect 45836 28590 45838 28642
rect 45838 28590 45890 28642
rect 45890 28590 45892 28642
rect 45836 28588 45892 28590
rect 46396 27692 46452 27748
rect 44768 26628 44824 26684
rect 44872 26682 44928 26684
rect 44976 26682 45032 26684
rect 44872 26630 44896 26682
rect 44896 26630 44928 26682
rect 44976 26630 45020 26682
rect 45020 26630 45032 26682
rect 44872 26628 44928 26630
rect 44976 26628 45032 26630
rect 45080 26628 45136 26684
rect 45184 26682 45240 26684
rect 45288 26682 45344 26684
rect 45184 26630 45196 26682
rect 45196 26630 45240 26682
rect 45288 26630 45320 26682
rect 45320 26630 45344 26682
rect 45184 26628 45240 26630
rect 45288 26628 45344 26630
rect 45392 26628 45448 26684
rect 45276 25340 45332 25396
rect 44268 25116 44324 25172
rect 44768 25060 44824 25116
rect 44872 25114 44928 25116
rect 44976 25114 45032 25116
rect 44872 25062 44896 25114
rect 44896 25062 44928 25114
rect 44976 25062 45020 25114
rect 45020 25062 45032 25114
rect 44872 25060 44928 25062
rect 44976 25060 45032 25062
rect 45080 25060 45136 25116
rect 45184 25114 45240 25116
rect 45288 25114 45344 25116
rect 45184 25062 45196 25114
rect 45196 25062 45240 25114
rect 45288 25062 45320 25114
rect 45320 25062 45344 25114
rect 45184 25060 45240 25062
rect 45288 25060 45344 25062
rect 45392 25060 45448 25116
rect 44156 20578 44212 20580
rect 44156 20526 44158 20578
rect 44158 20526 44210 20578
rect 44210 20526 44212 20578
rect 44156 20524 44212 20526
rect 44268 19234 44324 19236
rect 44268 19182 44270 19234
rect 44270 19182 44322 19234
rect 44322 19182 44324 19234
rect 44268 19180 44324 19182
rect 40268 18004 40324 18060
rect 40372 18058 40428 18060
rect 40476 18058 40532 18060
rect 40372 18006 40396 18058
rect 40396 18006 40428 18058
rect 40476 18006 40520 18058
rect 40520 18006 40532 18058
rect 40372 18004 40428 18006
rect 40476 18004 40532 18006
rect 40580 18004 40636 18060
rect 40684 18058 40740 18060
rect 40788 18058 40844 18060
rect 40684 18006 40696 18058
rect 40696 18006 40740 18058
rect 40788 18006 40820 18058
rect 40820 18006 40844 18058
rect 40684 18004 40740 18006
rect 40788 18004 40844 18006
rect 40892 18004 40948 18060
rect 40268 16436 40324 16492
rect 40372 16490 40428 16492
rect 40476 16490 40532 16492
rect 40372 16438 40396 16490
rect 40396 16438 40428 16490
rect 40476 16438 40520 16490
rect 40520 16438 40532 16490
rect 40372 16436 40428 16438
rect 40476 16436 40532 16438
rect 40580 16436 40636 16492
rect 40684 16490 40740 16492
rect 40788 16490 40844 16492
rect 40684 16438 40696 16490
rect 40696 16438 40740 16490
rect 40788 16438 40820 16490
rect 40820 16438 40844 16490
rect 40684 16436 40740 16438
rect 40788 16436 40844 16438
rect 40892 16436 40948 16492
rect 41244 15148 41300 15204
rect 35768 14084 35824 14140
rect 35872 14138 35928 14140
rect 35976 14138 36032 14140
rect 35872 14086 35896 14138
rect 35896 14086 35928 14138
rect 35976 14086 36020 14138
rect 36020 14086 36032 14138
rect 35872 14084 35928 14086
rect 35976 14084 36032 14086
rect 36080 14084 36136 14140
rect 36184 14138 36240 14140
rect 36288 14138 36344 14140
rect 36184 14086 36196 14138
rect 36196 14086 36240 14138
rect 36288 14086 36320 14138
rect 36320 14086 36344 14138
rect 36184 14084 36240 14086
rect 36288 14084 36344 14086
rect 36392 14084 36448 14140
rect 35768 12516 35824 12572
rect 35872 12570 35928 12572
rect 35976 12570 36032 12572
rect 35872 12518 35896 12570
rect 35896 12518 35928 12570
rect 35976 12518 36020 12570
rect 36020 12518 36032 12570
rect 35872 12516 35928 12518
rect 35976 12516 36032 12518
rect 36080 12516 36136 12572
rect 36184 12570 36240 12572
rect 36288 12570 36344 12572
rect 36184 12518 36196 12570
rect 36196 12518 36240 12570
rect 36288 12518 36320 12570
rect 36320 12518 36344 12570
rect 36184 12516 36240 12518
rect 36288 12516 36344 12518
rect 36392 12516 36448 12572
rect 35768 10948 35824 11004
rect 35872 11002 35928 11004
rect 35976 11002 36032 11004
rect 35872 10950 35896 11002
rect 35896 10950 35928 11002
rect 35976 10950 36020 11002
rect 36020 10950 36032 11002
rect 35872 10948 35928 10950
rect 35976 10948 36032 10950
rect 36080 10948 36136 11004
rect 36184 11002 36240 11004
rect 36288 11002 36344 11004
rect 36184 10950 36196 11002
rect 36196 10950 36240 11002
rect 36288 10950 36320 11002
rect 36320 10950 36344 11002
rect 36184 10948 36240 10950
rect 36288 10948 36344 10950
rect 36392 10948 36448 11004
rect 35308 8988 35364 9044
rect 34972 6300 35028 6356
rect 35084 7420 35140 7476
rect 34076 5180 34132 5236
rect 33852 4956 33908 5012
rect 33852 4338 33908 4340
rect 33852 4286 33854 4338
rect 33854 4286 33906 4338
rect 33906 4286 33908 4338
rect 33852 4284 33908 4286
rect 33292 3724 33348 3780
rect 32508 3500 32564 3556
rect 8768 3108 8824 3164
rect 8872 3162 8928 3164
rect 8976 3162 9032 3164
rect 8872 3110 8896 3162
rect 8896 3110 8928 3162
rect 8976 3110 9020 3162
rect 9020 3110 9032 3162
rect 8872 3108 8928 3110
rect 8976 3108 9032 3110
rect 9080 3108 9136 3164
rect 9184 3162 9240 3164
rect 9288 3162 9344 3164
rect 9184 3110 9196 3162
rect 9196 3110 9240 3162
rect 9288 3110 9320 3162
rect 9320 3110 9344 3162
rect 9184 3108 9240 3110
rect 9288 3108 9344 3110
rect 9392 3108 9448 3164
rect 17768 3108 17824 3164
rect 17872 3162 17928 3164
rect 17976 3162 18032 3164
rect 17872 3110 17896 3162
rect 17896 3110 17928 3162
rect 17976 3110 18020 3162
rect 18020 3110 18032 3162
rect 17872 3108 17928 3110
rect 17976 3108 18032 3110
rect 18080 3108 18136 3164
rect 18184 3162 18240 3164
rect 18288 3162 18344 3164
rect 18184 3110 18196 3162
rect 18196 3110 18240 3162
rect 18288 3110 18320 3162
rect 18320 3110 18344 3162
rect 18184 3108 18240 3110
rect 18288 3108 18344 3110
rect 18392 3108 18448 3164
rect 26768 3108 26824 3164
rect 26872 3162 26928 3164
rect 26976 3162 27032 3164
rect 26872 3110 26896 3162
rect 26896 3110 26928 3162
rect 26976 3110 27020 3162
rect 27020 3110 27032 3162
rect 26872 3108 26928 3110
rect 26976 3108 27032 3110
rect 27080 3108 27136 3164
rect 27184 3162 27240 3164
rect 27288 3162 27344 3164
rect 27184 3110 27196 3162
rect 27196 3110 27240 3162
rect 27288 3110 27320 3162
rect 27320 3110 27344 3162
rect 27184 3108 27240 3110
rect 27288 3108 27344 3110
rect 27392 3108 27448 3164
rect 34188 4284 34244 4340
rect 34972 5404 35028 5460
rect 34412 5234 34468 5236
rect 34412 5182 34414 5234
rect 34414 5182 34466 5234
rect 34466 5182 34468 5234
rect 34412 5180 34468 5182
rect 35532 9660 35588 9716
rect 35768 9380 35824 9436
rect 35872 9434 35928 9436
rect 35976 9434 36032 9436
rect 35872 9382 35896 9434
rect 35896 9382 35928 9434
rect 35976 9382 36020 9434
rect 36020 9382 36032 9434
rect 35872 9380 35928 9382
rect 35976 9380 36032 9382
rect 36080 9380 36136 9436
rect 36184 9434 36240 9436
rect 36288 9434 36344 9436
rect 36184 9382 36196 9434
rect 36196 9382 36240 9434
rect 36288 9382 36320 9434
rect 36320 9382 36344 9434
rect 36184 9380 36240 9382
rect 36288 9380 36344 9382
rect 36392 9380 36448 9436
rect 36428 9212 36484 9268
rect 35768 7812 35824 7868
rect 35872 7866 35928 7868
rect 35976 7866 36032 7868
rect 35872 7814 35896 7866
rect 35896 7814 35928 7866
rect 35976 7814 36020 7866
rect 36020 7814 36032 7866
rect 35872 7812 35928 7814
rect 35976 7812 36032 7814
rect 36080 7812 36136 7868
rect 36184 7866 36240 7868
rect 36288 7866 36344 7868
rect 36184 7814 36196 7866
rect 36196 7814 36240 7866
rect 36288 7814 36320 7866
rect 36320 7814 36344 7866
rect 36184 7812 36240 7814
rect 36288 7812 36344 7814
rect 36392 7812 36448 7868
rect 37660 11228 37716 11284
rect 37212 9212 37268 9268
rect 37436 9772 37492 9828
rect 37212 7532 37268 7588
rect 37436 8092 37492 8148
rect 37324 6914 37380 6916
rect 37324 6862 37326 6914
rect 37326 6862 37378 6914
rect 37378 6862 37380 6914
rect 37324 6860 37380 6862
rect 35768 6244 35824 6300
rect 35872 6298 35928 6300
rect 35976 6298 36032 6300
rect 35872 6246 35896 6298
rect 35896 6246 35928 6298
rect 35976 6246 36020 6298
rect 36020 6246 36032 6298
rect 35872 6244 35928 6246
rect 35976 6244 36032 6246
rect 36080 6244 36136 6300
rect 36184 6298 36240 6300
rect 36288 6298 36344 6300
rect 36184 6246 36196 6298
rect 36196 6246 36240 6298
rect 36288 6246 36320 6298
rect 36320 6246 36344 6298
rect 36184 6244 36240 6246
rect 36288 6244 36344 6246
rect 36392 6244 36448 6300
rect 35644 6018 35700 6020
rect 35644 5966 35646 6018
rect 35646 5966 35698 6018
rect 35698 5966 35700 6018
rect 35644 5964 35700 5966
rect 36540 5404 36596 5460
rect 35420 5292 35476 5348
rect 36428 5292 36484 5348
rect 34748 5068 34804 5124
rect 34636 4338 34692 4340
rect 34636 4286 34638 4338
rect 34638 4286 34690 4338
rect 34690 4286 34692 4338
rect 34636 4284 34692 4286
rect 35768 4676 35824 4732
rect 35872 4730 35928 4732
rect 35976 4730 36032 4732
rect 35872 4678 35896 4730
rect 35896 4678 35928 4730
rect 35976 4678 36020 4730
rect 36020 4678 36032 4730
rect 35872 4676 35928 4678
rect 35976 4676 36032 4678
rect 36080 4676 36136 4732
rect 36184 4730 36240 4732
rect 36288 4730 36344 4732
rect 36184 4678 36196 4730
rect 36196 4678 36240 4730
rect 36288 4678 36320 4730
rect 36320 4678 36344 4730
rect 36184 4676 36240 4678
rect 36288 4676 36344 4678
rect 36392 4676 36448 4732
rect 35196 4284 35252 4340
rect 37996 5404 38052 5460
rect 40268 14868 40324 14924
rect 40372 14922 40428 14924
rect 40476 14922 40532 14924
rect 40372 14870 40396 14922
rect 40396 14870 40428 14922
rect 40476 14870 40520 14922
rect 40520 14870 40532 14922
rect 40372 14868 40428 14870
rect 40476 14868 40532 14870
rect 40580 14868 40636 14924
rect 40684 14922 40740 14924
rect 40788 14922 40844 14924
rect 40684 14870 40696 14922
rect 40696 14870 40740 14922
rect 40788 14870 40820 14922
rect 40820 14870 40844 14922
rect 40684 14868 40740 14870
rect 40788 14868 40844 14870
rect 40892 14868 40948 14924
rect 40268 13300 40324 13356
rect 40372 13354 40428 13356
rect 40476 13354 40532 13356
rect 40372 13302 40396 13354
rect 40396 13302 40428 13354
rect 40476 13302 40520 13354
rect 40520 13302 40532 13354
rect 40372 13300 40428 13302
rect 40476 13300 40532 13302
rect 40580 13300 40636 13356
rect 40684 13354 40740 13356
rect 40788 13354 40844 13356
rect 40684 13302 40696 13354
rect 40696 13302 40740 13354
rect 40788 13302 40820 13354
rect 40820 13302 40844 13354
rect 40684 13300 40740 13302
rect 40788 13300 40844 13302
rect 40892 13300 40948 13356
rect 39004 11394 39060 11396
rect 39004 11342 39006 11394
rect 39006 11342 39058 11394
rect 39058 11342 39060 11394
rect 39004 11340 39060 11342
rect 39004 9826 39060 9828
rect 39004 9774 39006 9826
rect 39006 9774 39058 9826
rect 39058 9774 39060 9826
rect 39004 9772 39060 9774
rect 40268 11732 40324 11788
rect 40372 11786 40428 11788
rect 40476 11786 40532 11788
rect 40372 11734 40396 11786
rect 40396 11734 40428 11786
rect 40476 11734 40520 11786
rect 40520 11734 40532 11786
rect 40372 11732 40428 11734
rect 40476 11732 40532 11734
rect 40580 11732 40636 11788
rect 40684 11786 40740 11788
rect 40788 11786 40844 11788
rect 40684 11734 40696 11786
rect 40696 11734 40740 11786
rect 40788 11734 40820 11786
rect 40820 11734 40844 11786
rect 40684 11732 40740 11734
rect 40788 11732 40844 11734
rect 40892 11732 40948 11788
rect 41020 11282 41076 11284
rect 41020 11230 41022 11282
rect 41022 11230 41074 11282
rect 41074 11230 41076 11282
rect 41020 11228 41076 11230
rect 40268 10164 40324 10220
rect 40372 10218 40428 10220
rect 40476 10218 40532 10220
rect 40372 10166 40396 10218
rect 40396 10166 40428 10218
rect 40476 10166 40520 10218
rect 40520 10166 40532 10218
rect 40372 10164 40428 10166
rect 40476 10164 40532 10166
rect 40580 10164 40636 10220
rect 40684 10218 40740 10220
rect 40788 10218 40844 10220
rect 40684 10166 40696 10218
rect 40696 10166 40740 10218
rect 40788 10166 40820 10218
rect 40820 10166 40844 10218
rect 40684 10164 40740 10166
rect 40788 10164 40844 10166
rect 40892 10164 40948 10220
rect 40012 9660 40068 9716
rect 41020 9714 41076 9716
rect 41020 9662 41022 9714
rect 41022 9662 41074 9714
rect 41074 9662 41076 9714
rect 41020 9660 41076 9662
rect 40268 8596 40324 8652
rect 40372 8650 40428 8652
rect 40476 8650 40532 8652
rect 40372 8598 40396 8650
rect 40396 8598 40428 8650
rect 40476 8598 40520 8650
rect 40520 8598 40532 8650
rect 40372 8596 40428 8598
rect 40476 8596 40532 8598
rect 40580 8596 40636 8652
rect 40684 8650 40740 8652
rect 40788 8650 40844 8652
rect 40684 8598 40696 8650
rect 40696 8598 40740 8650
rect 40788 8598 40820 8650
rect 40820 8598 40844 8650
rect 40684 8596 40740 8598
rect 40788 8596 40844 8598
rect 40892 8596 40948 8652
rect 38332 7362 38388 7364
rect 38332 7310 38334 7362
rect 38334 7310 38386 7362
rect 38386 7310 38388 7362
rect 38332 7308 38388 7310
rect 41020 7196 41076 7252
rect 40268 7028 40324 7084
rect 40372 7082 40428 7084
rect 40476 7082 40532 7084
rect 40372 7030 40396 7082
rect 40396 7030 40428 7082
rect 40476 7030 40520 7082
rect 40520 7030 40532 7082
rect 40372 7028 40428 7030
rect 40476 7028 40532 7030
rect 40580 7028 40636 7084
rect 40684 7082 40740 7084
rect 40788 7082 40844 7084
rect 40684 7030 40696 7082
rect 40696 7030 40740 7082
rect 40788 7030 40820 7082
rect 40820 7030 40844 7082
rect 40684 7028 40740 7030
rect 40788 7028 40844 7030
rect 40892 7028 40948 7084
rect 40124 6748 40180 6804
rect 40908 6636 40964 6692
rect 38780 5404 38836 5460
rect 38332 4450 38388 4452
rect 38332 4398 38334 4450
rect 38334 4398 38386 4450
rect 38386 4398 38388 4450
rect 38332 4396 38388 4398
rect 38220 3836 38276 3892
rect 34748 3554 34804 3556
rect 34748 3502 34750 3554
rect 34750 3502 34802 3554
rect 34802 3502 34804 3554
rect 34748 3500 34804 3502
rect 36092 3554 36148 3556
rect 36092 3502 36094 3554
rect 36094 3502 36146 3554
rect 36146 3502 36148 3554
rect 36092 3500 36148 3502
rect 37436 3554 37492 3556
rect 37436 3502 37438 3554
rect 37438 3502 37490 3554
rect 37490 3502 37492 3554
rect 37436 3500 37492 3502
rect 37884 3554 37940 3556
rect 37884 3502 37886 3554
rect 37886 3502 37938 3554
rect 37938 3502 37940 3554
rect 37884 3500 37940 3502
rect 38332 3554 38388 3556
rect 38332 3502 38334 3554
rect 38334 3502 38386 3554
rect 38386 3502 38388 3554
rect 38332 3500 38388 3502
rect 38668 3612 38724 3668
rect 38780 4060 38836 4116
rect 39228 4956 39284 5012
rect 39116 3724 39172 3780
rect 40268 5460 40324 5516
rect 40372 5514 40428 5516
rect 40476 5514 40532 5516
rect 40372 5462 40396 5514
rect 40396 5462 40428 5514
rect 40476 5462 40520 5514
rect 40520 5462 40532 5514
rect 40372 5460 40428 5462
rect 40476 5460 40532 5462
rect 40580 5460 40636 5516
rect 40684 5514 40740 5516
rect 40788 5514 40844 5516
rect 40684 5462 40696 5514
rect 40696 5462 40740 5514
rect 40788 5462 40820 5514
rect 40820 5462 40844 5514
rect 40684 5460 40740 5462
rect 40788 5460 40844 5462
rect 40892 5460 40948 5516
rect 41132 4620 41188 4676
rect 41244 6524 41300 6580
rect 40124 4508 40180 4564
rect 40236 4338 40292 4340
rect 40236 4286 40238 4338
rect 40238 4286 40290 4338
rect 40290 4286 40292 4338
rect 40236 4284 40292 4286
rect 41132 4172 41188 4228
rect 40268 3892 40324 3948
rect 40372 3946 40428 3948
rect 40476 3946 40532 3948
rect 40372 3894 40396 3946
rect 40396 3894 40428 3946
rect 40476 3894 40520 3946
rect 40520 3894 40532 3946
rect 40372 3892 40428 3894
rect 40476 3892 40532 3894
rect 40580 3892 40636 3948
rect 40684 3946 40740 3948
rect 40788 3946 40844 3948
rect 40684 3894 40696 3946
rect 40696 3894 40740 3946
rect 40788 3894 40820 3946
rect 40820 3894 40844 3946
rect 40684 3892 40740 3894
rect 40788 3892 40844 3894
rect 40892 3892 40948 3948
rect 41020 3778 41076 3780
rect 41020 3726 41022 3778
rect 41022 3726 41074 3778
rect 41074 3726 41076 3778
rect 41020 3724 41076 3726
rect 40908 3666 40964 3668
rect 40908 3614 40910 3666
rect 40910 3614 40962 3666
rect 40962 3614 40964 3666
rect 40908 3612 40964 3614
rect 40348 3554 40404 3556
rect 40348 3502 40350 3554
rect 40350 3502 40402 3554
rect 40402 3502 40404 3554
rect 40348 3500 40404 3502
rect 38556 3388 38612 3444
rect 39004 3388 39060 3444
rect 35768 3108 35824 3164
rect 35872 3162 35928 3164
rect 35976 3162 36032 3164
rect 35872 3110 35896 3162
rect 35896 3110 35928 3162
rect 35976 3110 36020 3162
rect 36020 3110 36032 3162
rect 35872 3108 35928 3110
rect 35976 3108 36032 3110
rect 36080 3108 36136 3164
rect 36184 3162 36240 3164
rect 36288 3162 36344 3164
rect 36184 3110 36196 3162
rect 36196 3110 36240 3162
rect 36288 3110 36320 3162
rect 36320 3110 36344 3162
rect 36184 3108 36240 3110
rect 36288 3108 36344 3110
rect 36392 3108 36448 3164
rect 39788 3442 39844 3444
rect 39788 3390 39790 3442
rect 39790 3390 39842 3442
rect 39842 3390 39844 3442
rect 39788 3388 39844 3390
rect 41468 6412 41524 6468
rect 41692 6130 41748 6132
rect 41692 6078 41694 6130
rect 41694 6078 41746 6130
rect 41746 6078 41748 6130
rect 41692 6076 41748 6078
rect 41580 4844 41636 4900
rect 41692 5180 41748 5236
rect 41468 4732 41524 4788
rect 41468 3724 41524 3780
rect 41580 4620 41636 4676
rect 43036 15148 43092 15204
rect 44768 23492 44824 23548
rect 44872 23546 44928 23548
rect 44976 23546 45032 23548
rect 44872 23494 44896 23546
rect 44896 23494 44928 23546
rect 44976 23494 45020 23546
rect 45020 23494 45032 23546
rect 44872 23492 44928 23494
rect 44976 23492 45032 23494
rect 45080 23492 45136 23548
rect 45184 23546 45240 23548
rect 45288 23546 45344 23548
rect 45184 23494 45196 23546
rect 45196 23494 45240 23546
rect 45288 23494 45320 23546
rect 45320 23494 45344 23546
rect 45184 23492 45240 23494
rect 45288 23492 45344 23494
rect 45392 23492 45448 23548
rect 45164 23154 45220 23156
rect 45164 23102 45166 23154
rect 45166 23102 45218 23154
rect 45218 23102 45220 23154
rect 45164 23100 45220 23102
rect 46060 23100 46116 23156
rect 44768 21924 44824 21980
rect 44872 21978 44928 21980
rect 44976 21978 45032 21980
rect 44872 21926 44896 21978
rect 44896 21926 44928 21978
rect 44976 21926 45020 21978
rect 45020 21926 45032 21978
rect 44872 21924 44928 21926
rect 44976 21924 45032 21926
rect 45080 21924 45136 21980
rect 45184 21978 45240 21980
rect 45288 21978 45344 21980
rect 45184 21926 45196 21978
rect 45196 21926 45240 21978
rect 45288 21926 45320 21978
rect 45320 21926 45344 21978
rect 45184 21924 45240 21926
rect 45288 21924 45344 21926
rect 45392 21924 45448 21980
rect 46284 22540 46340 22596
rect 45612 21420 45668 21476
rect 44768 20356 44824 20412
rect 44872 20410 44928 20412
rect 44976 20410 45032 20412
rect 44872 20358 44896 20410
rect 44896 20358 44928 20410
rect 44976 20358 45020 20410
rect 45020 20358 45032 20410
rect 44872 20356 44928 20358
rect 44976 20356 45032 20358
rect 45080 20356 45136 20412
rect 45184 20410 45240 20412
rect 45288 20410 45344 20412
rect 45184 20358 45196 20410
rect 45196 20358 45240 20410
rect 45288 20358 45320 20410
rect 45320 20358 45344 20410
rect 45184 20356 45240 20358
rect 45288 20356 45344 20358
rect 45392 20356 45448 20412
rect 44768 18788 44824 18844
rect 44872 18842 44928 18844
rect 44976 18842 45032 18844
rect 44872 18790 44896 18842
rect 44896 18790 44928 18842
rect 44976 18790 45020 18842
rect 45020 18790 45032 18842
rect 44872 18788 44928 18790
rect 44976 18788 45032 18790
rect 45080 18788 45136 18844
rect 45184 18842 45240 18844
rect 45288 18842 45344 18844
rect 45184 18790 45196 18842
rect 45196 18790 45240 18842
rect 45288 18790 45320 18842
rect 45320 18790 45344 18842
rect 45184 18788 45240 18790
rect 45288 18788 45344 18790
rect 45392 18788 45448 18844
rect 44768 17220 44824 17276
rect 44872 17274 44928 17276
rect 44976 17274 45032 17276
rect 44872 17222 44896 17274
rect 44896 17222 44928 17274
rect 44976 17222 45020 17274
rect 45020 17222 45032 17274
rect 44872 17220 44928 17222
rect 44976 17220 45032 17222
rect 45080 17220 45136 17276
rect 45184 17274 45240 17276
rect 45288 17274 45344 17276
rect 45184 17222 45196 17274
rect 45196 17222 45240 17274
rect 45288 17222 45320 17274
rect 45320 17222 45344 17274
rect 45184 17220 45240 17222
rect 45288 17220 45344 17222
rect 45392 17220 45448 17276
rect 44768 15652 44824 15708
rect 44872 15706 44928 15708
rect 44976 15706 45032 15708
rect 44872 15654 44896 15706
rect 44896 15654 44928 15706
rect 44976 15654 45020 15706
rect 45020 15654 45032 15706
rect 44872 15652 44928 15654
rect 44976 15652 45032 15654
rect 45080 15652 45136 15708
rect 45184 15706 45240 15708
rect 45288 15706 45344 15708
rect 45184 15654 45196 15706
rect 45196 15654 45240 15706
rect 45288 15654 45320 15706
rect 45320 15654 45344 15706
rect 45184 15652 45240 15654
rect 45288 15652 45344 15654
rect 45392 15652 45448 15708
rect 42476 9324 42532 9380
rect 42140 7474 42196 7476
rect 42140 7422 42142 7474
rect 42142 7422 42194 7474
rect 42194 7422 42196 7474
rect 42140 7420 42196 7422
rect 41916 6748 41972 6804
rect 42028 6076 42084 6132
rect 41804 4172 41860 4228
rect 41916 5068 41972 5124
rect 42700 8930 42756 8932
rect 42700 8878 42702 8930
rect 42702 8878 42754 8930
rect 42754 8878 42756 8930
rect 42700 8876 42756 8878
rect 43036 11228 43092 11284
rect 42364 7250 42420 7252
rect 42364 7198 42366 7250
rect 42366 7198 42418 7250
rect 42418 7198 42420 7250
rect 42364 7196 42420 7198
rect 42588 6130 42644 6132
rect 42588 6078 42590 6130
rect 42590 6078 42642 6130
rect 42642 6078 42644 6130
rect 42588 6076 42644 6078
rect 42252 5234 42308 5236
rect 42252 5182 42254 5234
rect 42254 5182 42306 5234
rect 42306 5182 42308 5234
rect 42252 5180 42308 5182
rect 42476 4956 42532 5012
rect 42140 4732 42196 4788
rect 42364 4508 42420 4564
rect 42028 4060 42084 4116
rect 42252 3724 42308 3780
rect 41580 3554 41636 3556
rect 41580 3502 41582 3554
rect 41582 3502 41634 3554
rect 41634 3502 41636 3554
rect 41580 3500 41636 3502
rect 42588 3724 42644 3780
rect 42588 3442 42644 3444
rect 42588 3390 42590 3442
rect 42590 3390 42642 3442
rect 42642 3390 42644 3442
rect 42588 3388 42644 3390
rect 42924 5180 42980 5236
rect 42812 5122 42868 5124
rect 42812 5070 42814 5122
rect 42814 5070 42866 5122
rect 42866 5070 42868 5122
rect 42812 5068 42868 5070
rect 43708 9324 43764 9380
rect 43148 4396 43204 4452
rect 43484 4844 43540 4900
rect 43036 3500 43092 3556
rect 44268 14364 44324 14420
rect 44156 8876 44212 8932
rect 44044 8146 44100 8148
rect 44044 8094 44046 8146
rect 44046 8094 44098 8146
rect 44098 8094 44100 8146
rect 44044 8092 44100 8094
rect 44380 12066 44436 12068
rect 44380 12014 44382 12066
rect 44382 12014 44434 12066
rect 44434 12014 44436 12066
rect 44380 12012 44436 12014
rect 43820 4284 43876 4340
rect 44156 7308 44212 7364
rect 47404 34130 47460 34132
rect 47404 34078 47406 34130
rect 47406 34078 47458 34130
rect 47458 34078 47460 34130
rect 47404 34076 47460 34078
rect 47852 33404 47908 33460
rect 49868 44044 49924 44100
rect 49268 43092 49324 43148
rect 49372 43146 49428 43148
rect 49476 43146 49532 43148
rect 49372 43094 49396 43146
rect 49396 43094 49428 43146
rect 49476 43094 49520 43146
rect 49520 43094 49532 43146
rect 49372 43092 49428 43094
rect 49476 43092 49532 43094
rect 49580 43092 49636 43148
rect 49684 43146 49740 43148
rect 49788 43146 49844 43148
rect 49684 43094 49696 43146
rect 49696 43094 49740 43146
rect 49788 43094 49820 43146
rect 49820 43094 49844 43146
rect 49684 43092 49740 43094
rect 49788 43092 49844 43094
rect 49892 43092 49948 43148
rect 49644 42082 49700 42084
rect 49644 42030 49646 42082
rect 49646 42030 49698 42082
rect 49698 42030 49700 42082
rect 49644 42028 49700 42030
rect 49268 41524 49324 41580
rect 49372 41578 49428 41580
rect 49476 41578 49532 41580
rect 49372 41526 49396 41578
rect 49396 41526 49428 41578
rect 49476 41526 49520 41578
rect 49520 41526 49532 41578
rect 49372 41524 49428 41526
rect 49476 41524 49532 41526
rect 49580 41524 49636 41580
rect 49684 41578 49740 41580
rect 49788 41578 49844 41580
rect 49684 41526 49696 41578
rect 49696 41526 49740 41578
rect 49788 41526 49820 41578
rect 49820 41526 49844 41578
rect 49684 41524 49740 41526
rect 49788 41524 49844 41526
rect 49892 41524 49948 41580
rect 49532 41020 49588 41076
rect 51100 41804 51156 41860
rect 50988 41074 51044 41076
rect 50988 41022 50990 41074
rect 50990 41022 51042 41074
rect 51042 41022 51044 41074
rect 50988 41020 51044 41022
rect 49420 40402 49476 40404
rect 49420 40350 49422 40402
rect 49422 40350 49474 40402
rect 49474 40350 49476 40402
rect 49420 40348 49476 40350
rect 50092 40402 50148 40404
rect 50092 40350 50094 40402
rect 50094 40350 50146 40402
rect 50146 40350 50148 40402
rect 50092 40348 50148 40350
rect 49268 39956 49324 40012
rect 49372 40010 49428 40012
rect 49476 40010 49532 40012
rect 49372 39958 49396 40010
rect 49396 39958 49428 40010
rect 49476 39958 49520 40010
rect 49520 39958 49532 40010
rect 49372 39956 49428 39958
rect 49476 39956 49532 39958
rect 49580 39956 49636 40012
rect 49684 40010 49740 40012
rect 49788 40010 49844 40012
rect 49684 39958 49696 40010
rect 49696 39958 49740 40010
rect 49788 39958 49820 40010
rect 49820 39958 49844 40010
rect 49684 39956 49740 39958
rect 49788 39956 49844 39958
rect 49892 39956 49948 40012
rect 49084 38892 49140 38948
rect 48972 37154 49028 37156
rect 48972 37102 48974 37154
rect 48974 37102 49026 37154
rect 49026 37102 49028 37154
rect 48972 37100 49028 37102
rect 49268 38388 49324 38444
rect 49372 38442 49428 38444
rect 49476 38442 49532 38444
rect 49372 38390 49396 38442
rect 49396 38390 49428 38442
rect 49476 38390 49520 38442
rect 49520 38390 49532 38442
rect 49372 38388 49428 38390
rect 49476 38388 49532 38390
rect 49580 38388 49636 38444
rect 49684 38442 49740 38444
rect 49788 38442 49844 38444
rect 49684 38390 49696 38442
rect 49696 38390 49740 38442
rect 49788 38390 49820 38442
rect 49820 38390 49844 38442
rect 49684 38388 49740 38390
rect 49788 38388 49844 38390
rect 49892 38388 49948 38444
rect 49756 38050 49812 38052
rect 49756 37998 49758 38050
rect 49758 37998 49810 38050
rect 49810 37998 49812 38050
rect 49756 37996 49812 37998
rect 50652 40348 50708 40404
rect 50204 38220 50260 38276
rect 50540 39004 50596 39060
rect 48412 34802 48468 34804
rect 48412 34750 48414 34802
rect 48414 34750 48466 34802
rect 48466 34750 48468 34802
rect 48412 34748 48468 34750
rect 48524 34076 48580 34132
rect 49268 36820 49324 36876
rect 49372 36874 49428 36876
rect 49476 36874 49532 36876
rect 49372 36822 49396 36874
rect 49396 36822 49428 36874
rect 49476 36822 49520 36874
rect 49520 36822 49532 36874
rect 49372 36820 49428 36822
rect 49476 36820 49532 36822
rect 49580 36820 49636 36876
rect 49684 36874 49740 36876
rect 49788 36874 49844 36876
rect 49684 36822 49696 36874
rect 49696 36822 49740 36874
rect 49788 36822 49820 36874
rect 49820 36822 49844 36874
rect 49684 36820 49740 36822
rect 49788 36820 49844 36822
rect 49892 36820 49948 36876
rect 50204 36876 50260 36932
rect 50316 37100 50372 37156
rect 49084 35756 49140 35812
rect 49756 36540 49812 36596
rect 50428 37100 50484 37156
rect 50876 36594 50932 36596
rect 50876 36542 50878 36594
rect 50878 36542 50930 36594
rect 50930 36542 50932 36594
rect 50876 36540 50932 36542
rect 51996 44210 52052 44212
rect 51996 44158 51998 44210
rect 51998 44158 52050 44210
rect 52050 44158 52052 44210
rect 51996 44156 52052 44158
rect 53228 48466 53284 48468
rect 53228 48414 53230 48466
rect 53230 48414 53282 48466
rect 53282 48414 53284 48466
rect 53228 48412 53284 48414
rect 54460 48412 54516 48468
rect 54460 47292 54516 47348
rect 53768 47012 53824 47068
rect 53872 47066 53928 47068
rect 53976 47066 54032 47068
rect 53872 47014 53896 47066
rect 53896 47014 53928 47066
rect 53976 47014 54020 47066
rect 54020 47014 54032 47066
rect 53872 47012 53928 47014
rect 53976 47012 54032 47014
rect 54080 47012 54136 47068
rect 54184 47066 54240 47068
rect 54288 47066 54344 47068
rect 54184 47014 54196 47066
rect 54196 47014 54240 47066
rect 54288 47014 54320 47066
rect 54320 47014 54344 47066
rect 54184 47012 54240 47014
rect 54288 47012 54344 47014
rect 54392 47012 54448 47068
rect 53564 46844 53620 46900
rect 52892 46396 52948 46452
rect 54124 46620 54180 46676
rect 54572 46620 54628 46676
rect 54236 46562 54292 46564
rect 54236 46510 54238 46562
rect 54238 46510 54290 46562
rect 54290 46510 54292 46562
rect 54236 46508 54292 46510
rect 54124 45836 54180 45892
rect 54460 45666 54516 45668
rect 54460 45614 54462 45666
rect 54462 45614 54514 45666
rect 54514 45614 54516 45666
rect 54460 45612 54516 45614
rect 53768 45444 53824 45500
rect 53872 45498 53928 45500
rect 53976 45498 54032 45500
rect 53872 45446 53896 45498
rect 53896 45446 53928 45498
rect 53976 45446 54020 45498
rect 54020 45446 54032 45498
rect 53872 45444 53928 45446
rect 53976 45444 54032 45446
rect 54080 45444 54136 45500
rect 54184 45498 54240 45500
rect 54288 45498 54344 45500
rect 54184 45446 54196 45498
rect 54196 45446 54240 45498
rect 54288 45446 54320 45498
rect 54320 45446 54344 45498
rect 54184 45444 54240 45446
rect 54288 45444 54344 45446
rect 54392 45444 54448 45500
rect 53452 45388 53508 45444
rect 54908 46172 54964 46228
rect 55020 45890 55076 45892
rect 55020 45838 55022 45890
rect 55022 45838 55074 45890
rect 55074 45838 55076 45890
rect 55020 45836 55076 45838
rect 53564 44828 53620 44884
rect 52892 44098 52948 44100
rect 52892 44046 52894 44098
rect 52894 44046 52946 44098
rect 52946 44046 52948 44098
rect 52892 44044 52948 44046
rect 52780 43650 52836 43652
rect 52780 43598 52782 43650
rect 52782 43598 52834 43650
rect 52834 43598 52836 43650
rect 52780 43596 52836 43598
rect 52220 39340 52276 39396
rect 52556 39340 52612 39396
rect 51548 38162 51604 38164
rect 51548 38110 51550 38162
rect 51550 38110 51602 38162
rect 51602 38110 51604 38162
rect 51548 38108 51604 38110
rect 53228 43596 53284 43652
rect 55020 45612 55076 45668
rect 54908 44828 54964 44884
rect 54124 44268 54180 44324
rect 54572 44210 54628 44212
rect 54572 44158 54574 44210
rect 54574 44158 54626 44210
rect 54626 44158 54628 44210
rect 54572 44156 54628 44158
rect 53768 43876 53824 43932
rect 53872 43930 53928 43932
rect 53976 43930 54032 43932
rect 53872 43878 53896 43930
rect 53896 43878 53928 43930
rect 53976 43878 54020 43930
rect 54020 43878 54032 43930
rect 53872 43876 53928 43878
rect 53976 43876 54032 43878
rect 54080 43876 54136 43932
rect 54184 43930 54240 43932
rect 54288 43930 54344 43932
rect 54184 43878 54196 43930
rect 54196 43878 54240 43930
rect 54288 43878 54320 43930
rect 54320 43878 54344 43930
rect 54184 43876 54240 43878
rect 54288 43876 54344 43878
rect 54392 43876 54448 43932
rect 53900 43650 53956 43652
rect 53900 43598 53902 43650
rect 53902 43598 53954 43650
rect 53954 43598 53956 43650
rect 53900 43596 53956 43598
rect 53768 42308 53824 42364
rect 53872 42362 53928 42364
rect 53976 42362 54032 42364
rect 53872 42310 53896 42362
rect 53896 42310 53928 42362
rect 53976 42310 54020 42362
rect 54020 42310 54032 42362
rect 53872 42308 53928 42310
rect 53976 42308 54032 42310
rect 54080 42308 54136 42364
rect 54184 42362 54240 42364
rect 54288 42362 54344 42364
rect 54184 42310 54196 42362
rect 54196 42310 54240 42362
rect 54288 42310 54320 42362
rect 54320 42310 54344 42362
rect 54184 42308 54240 42310
rect 54288 42308 54344 42310
rect 54392 42308 54448 42364
rect 54796 44268 54852 44324
rect 53788 41858 53844 41860
rect 53788 41806 53790 41858
rect 53790 41806 53842 41858
rect 53842 41806 53844 41858
rect 53788 41804 53844 41806
rect 53340 41356 53396 41412
rect 53564 41020 53620 41076
rect 53228 40460 53284 40516
rect 53116 40402 53172 40404
rect 53116 40350 53118 40402
rect 53118 40350 53170 40402
rect 53170 40350 53172 40402
rect 53116 40348 53172 40350
rect 53768 40740 53824 40796
rect 53872 40794 53928 40796
rect 53976 40794 54032 40796
rect 53872 40742 53896 40794
rect 53896 40742 53928 40794
rect 53976 40742 54020 40794
rect 54020 40742 54032 40794
rect 53872 40740 53928 40742
rect 53976 40740 54032 40742
rect 54080 40740 54136 40796
rect 54184 40794 54240 40796
rect 54288 40794 54344 40796
rect 54184 40742 54196 40794
rect 54196 40742 54240 40794
rect 54288 40742 54320 40794
rect 54320 40742 54344 40794
rect 54184 40740 54240 40742
rect 54288 40740 54344 40742
rect 54392 40740 54448 40796
rect 54684 41020 54740 41076
rect 52892 39058 52948 39060
rect 52892 39006 52894 39058
rect 52894 39006 52946 39058
rect 52946 39006 52948 39058
rect 52892 39004 52948 39006
rect 51212 37154 51268 37156
rect 51212 37102 51214 37154
rect 51214 37102 51266 37154
rect 51266 37102 51268 37154
rect 51212 37100 51268 37102
rect 51100 36988 51156 37044
rect 49268 35252 49324 35308
rect 49372 35306 49428 35308
rect 49476 35306 49532 35308
rect 49372 35254 49396 35306
rect 49396 35254 49428 35306
rect 49476 35254 49520 35306
rect 49520 35254 49532 35306
rect 49372 35252 49428 35254
rect 49476 35252 49532 35254
rect 49580 35252 49636 35308
rect 49684 35306 49740 35308
rect 49788 35306 49844 35308
rect 49684 35254 49696 35306
rect 49696 35254 49740 35306
rect 49788 35254 49820 35306
rect 49820 35254 49844 35306
rect 49684 35252 49740 35254
rect 49788 35252 49844 35254
rect 49892 35252 49948 35308
rect 48972 34636 49028 34692
rect 49084 34748 49140 34804
rect 48860 33404 48916 33460
rect 48748 33180 48804 33236
rect 49308 34636 49364 34692
rect 49868 34636 49924 34692
rect 50316 35084 50372 35140
rect 51436 36876 51492 36932
rect 52108 36876 52164 36932
rect 51996 36764 52052 36820
rect 51548 36092 51604 36148
rect 52556 37996 52612 38052
rect 50316 34748 50372 34804
rect 50988 34972 51044 35028
rect 50428 34636 50484 34692
rect 51100 34636 51156 34692
rect 52108 35026 52164 35028
rect 52108 34974 52110 35026
rect 52110 34974 52162 35026
rect 52162 34974 52164 35026
rect 52108 34972 52164 34974
rect 51660 34636 51716 34692
rect 49756 34130 49812 34132
rect 49756 34078 49758 34130
rect 49758 34078 49810 34130
rect 49810 34078 49812 34130
rect 49756 34076 49812 34078
rect 50092 34130 50148 34132
rect 50092 34078 50094 34130
rect 50094 34078 50146 34130
rect 50146 34078 50148 34130
rect 50092 34076 50148 34078
rect 49268 33684 49324 33740
rect 49372 33738 49428 33740
rect 49476 33738 49532 33740
rect 49372 33686 49396 33738
rect 49396 33686 49428 33738
rect 49476 33686 49520 33738
rect 49520 33686 49532 33738
rect 49372 33684 49428 33686
rect 49476 33684 49532 33686
rect 49580 33684 49636 33740
rect 49684 33738 49740 33740
rect 49788 33738 49844 33740
rect 49684 33686 49696 33738
rect 49696 33686 49740 33738
rect 49788 33686 49820 33738
rect 49820 33686 49844 33738
rect 49684 33684 49740 33686
rect 49788 33684 49844 33686
rect 49892 33684 49948 33740
rect 48300 33068 48356 33124
rect 48188 32956 48244 33012
rect 50428 33122 50484 33124
rect 50428 33070 50430 33122
rect 50430 33070 50482 33122
rect 50482 33070 50484 33122
rect 50428 33068 50484 33070
rect 50092 32562 50148 32564
rect 50092 32510 50094 32562
rect 50094 32510 50146 32562
rect 50146 32510 50148 32562
rect 50092 32508 50148 32510
rect 50876 32508 50932 32564
rect 49268 32116 49324 32172
rect 49372 32170 49428 32172
rect 49476 32170 49532 32172
rect 49372 32118 49396 32170
rect 49396 32118 49428 32170
rect 49476 32118 49520 32170
rect 49520 32118 49532 32170
rect 49372 32116 49428 32118
rect 49476 32116 49532 32118
rect 49580 32116 49636 32172
rect 49684 32170 49740 32172
rect 49788 32170 49844 32172
rect 49684 32118 49696 32170
rect 49696 32118 49740 32170
rect 49788 32118 49820 32170
rect 49820 32118 49844 32170
rect 49684 32116 49740 32118
rect 49788 32116 49844 32118
rect 49892 32116 49948 32172
rect 46844 31948 46900 32004
rect 51212 32284 51268 32340
rect 52668 38892 52724 38948
rect 53004 36764 53060 36820
rect 52444 36540 52500 36596
rect 52780 36540 52836 36596
rect 52780 36316 52836 36372
rect 54012 40348 54068 40404
rect 54572 40236 54628 40292
rect 53768 39172 53824 39228
rect 53872 39226 53928 39228
rect 53976 39226 54032 39228
rect 53872 39174 53896 39226
rect 53896 39174 53928 39226
rect 53976 39174 54020 39226
rect 54020 39174 54032 39226
rect 53872 39172 53928 39174
rect 53976 39172 54032 39174
rect 54080 39172 54136 39228
rect 54184 39226 54240 39228
rect 54288 39226 54344 39228
rect 54184 39174 54196 39226
rect 54196 39174 54240 39226
rect 54288 39174 54320 39226
rect 54320 39174 54344 39226
rect 54184 39172 54240 39174
rect 54288 39172 54344 39174
rect 54392 39172 54448 39228
rect 53900 38946 53956 38948
rect 53900 38894 53902 38946
rect 53902 38894 53954 38946
rect 53954 38894 53956 38946
rect 53900 38892 53956 38894
rect 54796 40460 54852 40516
rect 54908 41804 54964 41860
rect 54572 37772 54628 37828
rect 53768 37604 53824 37660
rect 53872 37658 53928 37660
rect 53976 37658 54032 37660
rect 53872 37606 53896 37658
rect 53896 37606 53928 37658
rect 53976 37606 54020 37658
rect 54020 37606 54032 37658
rect 53872 37604 53928 37606
rect 53976 37604 54032 37606
rect 54080 37604 54136 37660
rect 54184 37658 54240 37660
rect 54288 37658 54344 37660
rect 54184 37606 54196 37658
rect 54196 37606 54240 37658
rect 54288 37606 54320 37658
rect 54320 37606 54344 37658
rect 54184 37604 54240 37606
rect 54288 37604 54344 37606
rect 54392 37604 54448 37660
rect 53228 37324 53284 37380
rect 54572 37378 54628 37380
rect 54572 37326 54574 37378
rect 54574 37326 54626 37378
rect 54626 37326 54628 37378
rect 54572 37324 54628 37326
rect 54012 37154 54068 37156
rect 54012 37102 54014 37154
rect 54014 37102 54066 37154
rect 54066 37102 54068 37154
rect 54012 37100 54068 37102
rect 53900 36988 53956 37044
rect 53900 36258 53956 36260
rect 53900 36206 53902 36258
rect 53902 36206 53954 36258
rect 53954 36206 53956 36258
rect 53900 36204 53956 36206
rect 53452 36092 53508 36148
rect 53768 36036 53824 36092
rect 53872 36090 53928 36092
rect 53976 36090 54032 36092
rect 53872 36038 53896 36090
rect 53896 36038 53928 36090
rect 53976 36038 54020 36090
rect 54020 36038 54032 36090
rect 53872 36036 53928 36038
rect 53976 36036 54032 36038
rect 54080 36036 54136 36092
rect 54184 36090 54240 36092
rect 54288 36090 54344 36092
rect 54184 36038 54196 36090
rect 54196 36038 54240 36090
rect 54288 36038 54320 36090
rect 54320 36038 54344 36090
rect 54184 36036 54240 36038
rect 54288 36036 54344 36038
rect 54392 36036 54448 36092
rect 53564 35868 53620 35924
rect 53788 35698 53844 35700
rect 53788 35646 53790 35698
rect 53790 35646 53842 35698
rect 53842 35646 53844 35698
rect 53788 35644 53844 35646
rect 53452 35532 53508 35588
rect 52668 34972 52724 35028
rect 52332 34130 52388 34132
rect 52332 34078 52334 34130
rect 52334 34078 52386 34130
rect 52386 34078 52388 34130
rect 52332 34076 52388 34078
rect 53228 34636 53284 34692
rect 53116 32508 53172 32564
rect 54124 34972 54180 35028
rect 54796 34748 54852 34804
rect 54684 34690 54740 34692
rect 54684 34638 54686 34690
rect 54686 34638 54738 34690
rect 54738 34638 54740 34690
rect 54684 34636 54740 34638
rect 53768 34468 53824 34524
rect 53872 34522 53928 34524
rect 53976 34522 54032 34524
rect 53872 34470 53896 34522
rect 53896 34470 53928 34522
rect 53976 34470 54020 34522
rect 54020 34470 54032 34522
rect 53872 34468 53928 34470
rect 53976 34468 54032 34470
rect 54080 34468 54136 34524
rect 54184 34522 54240 34524
rect 54288 34522 54344 34524
rect 54184 34470 54196 34522
rect 54196 34470 54240 34522
rect 54288 34470 54320 34522
rect 54320 34470 54344 34522
rect 54184 34468 54240 34470
rect 54288 34468 54344 34470
rect 54392 34468 54448 34524
rect 53768 32900 53824 32956
rect 53872 32954 53928 32956
rect 53976 32954 54032 32956
rect 53872 32902 53896 32954
rect 53896 32902 53928 32954
rect 53976 32902 54020 32954
rect 54020 32902 54032 32954
rect 53872 32900 53928 32902
rect 53976 32900 54032 32902
rect 54080 32900 54136 32956
rect 54184 32954 54240 32956
rect 54288 32954 54344 32956
rect 54184 32902 54196 32954
rect 54196 32902 54240 32954
rect 54288 32902 54320 32954
rect 54320 32902 54344 32954
rect 54184 32900 54240 32902
rect 54288 32900 54344 32902
rect 54392 32900 54448 32956
rect 54572 32732 54628 32788
rect 53788 32562 53844 32564
rect 53788 32510 53790 32562
rect 53790 32510 53842 32562
rect 53842 32510 53844 32562
rect 53788 32508 53844 32510
rect 53340 32396 53396 32452
rect 56364 48802 56420 48804
rect 56364 48750 56366 48802
rect 56366 48750 56418 48802
rect 56418 48750 56420 48802
rect 56364 48748 56420 48750
rect 57372 48748 57428 48804
rect 57036 47180 57092 47236
rect 55244 46674 55300 46676
rect 55244 46622 55246 46674
rect 55246 46622 55298 46674
rect 55298 46622 55300 46674
rect 55244 46620 55300 46622
rect 55356 46508 55412 46564
rect 55132 41916 55188 41972
rect 55244 46172 55300 46228
rect 55020 41692 55076 41748
rect 55580 46060 55636 46116
rect 57260 46508 57316 46564
rect 56588 46060 56644 46116
rect 56812 45778 56868 45780
rect 56812 45726 56814 45778
rect 56814 45726 56866 45778
rect 56866 45726 56868 45778
rect 56812 45724 56868 45726
rect 56028 45612 56084 45668
rect 56700 45612 56756 45668
rect 56924 45666 56980 45668
rect 56924 45614 56926 45666
rect 56926 45614 56978 45666
rect 56978 45614 56980 45666
rect 56924 45612 56980 45614
rect 55468 44322 55524 44324
rect 55468 44270 55470 44322
rect 55470 44270 55522 44322
rect 55522 44270 55524 44322
rect 55468 44268 55524 44270
rect 55692 44268 55748 44324
rect 55916 44156 55972 44212
rect 56700 44044 56756 44100
rect 56028 43650 56084 43652
rect 56028 43598 56030 43650
rect 56030 43598 56082 43650
rect 56082 43598 56084 43650
rect 56028 43596 56084 43598
rect 56812 43708 56868 43764
rect 56924 44210 56980 44212
rect 56924 44158 56926 44210
rect 56926 44158 56978 44210
rect 56978 44158 56980 44210
rect 56924 44156 56980 44158
rect 55356 41020 55412 41076
rect 55580 41970 55636 41972
rect 55580 41918 55582 41970
rect 55582 41918 55634 41970
rect 55634 41918 55636 41970
rect 55580 41916 55636 41918
rect 58044 52108 58100 52164
rect 58604 52274 58660 52276
rect 58604 52222 58606 52274
rect 58606 52222 58658 52274
rect 58658 52222 58660 52274
rect 58604 52220 58660 52222
rect 62768 54852 62824 54908
rect 62872 54906 62928 54908
rect 62976 54906 63032 54908
rect 62872 54854 62896 54906
rect 62896 54854 62928 54906
rect 62976 54854 63020 54906
rect 63020 54854 63032 54906
rect 62872 54852 62928 54854
rect 62976 54852 63032 54854
rect 63080 54852 63136 54908
rect 63184 54906 63240 54908
rect 63288 54906 63344 54908
rect 63184 54854 63196 54906
rect 63196 54854 63240 54906
rect 63288 54854 63320 54906
rect 63320 54854 63344 54906
rect 63184 54852 63240 54854
rect 63288 54852 63344 54854
rect 63392 54852 63448 54908
rect 60172 53788 60228 53844
rect 59052 52220 59108 52276
rect 60508 52274 60564 52276
rect 60508 52222 60510 52274
rect 60510 52222 60562 52274
rect 60562 52222 60564 52274
rect 60508 52220 60564 52222
rect 65324 53842 65380 53844
rect 65324 53790 65326 53842
rect 65326 53790 65378 53842
rect 65378 53790 65380 53842
rect 65324 53788 65380 53790
rect 61852 52108 61908 52164
rect 62076 53676 62132 53732
rect 65212 53730 65268 53732
rect 65212 53678 65214 53730
rect 65214 53678 65266 53730
rect 65266 53678 65268 53730
rect 65212 53676 65268 53678
rect 66780 54348 66836 54404
rect 66556 53900 66612 53956
rect 64876 53618 64932 53620
rect 64876 53566 64878 53618
rect 64878 53566 64930 53618
rect 64930 53566 64932 53618
rect 64876 53564 64932 53566
rect 62768 53284 62824 53340
rect 62872 53338 62928 53340
rect 62976 53338 63032 53340
rect 62872 53286 62896 53338
rect 62896 53286 62928 53338
rect 62976 53286 63020 53338
rect 63020 53286 63032 53338
rect 62872 53284 62928 53286
rect 62976 53284 63032 53286
rect 63080 53284 63136 53340
rect 63184 53338 63240 53340
rect 63288 53338 63344 53340
rect 63184 53286 63196 53338
rect 63196 53286 63240 53338
rect 63288 53286 63320 53338
rect 63320 53286 63344 53338
rect 63184 53284 63240 53286
rect 63288 53284 63344 53286
rect 63392 53284 63448 53340
rect 64540 53004 64596 53060
rect 66108 53676 66164 53732
rect 65436 53004 65492 53060
rect 62076 52780 62132 52836
rect 65212 52946 65268 52948
rect 65212 52894 65214 52946
rect 65214 52894 65266 52946
rect 65266 52894 65268 52946
rect 65212 52892 65268 52894
rect 62636 52668 62692 52724
rect 63420 52162 63476 52164
rect 63420 52110 63422 52162
rect 63422 52110 63474 52162
rect 63474 52110 63476 52162
rect 63420 52108 63476 52110
rect 63868 52162 63924 52164
rect 63868 52110 63870 52162
rect 63870 52110 63922 52162
rect 63922 52110 63924 52162
rect 63868 52108 63924 52110
rect 68460 56082 68516 56084
rect 68460 56030 68462 56082
rect 68462 56030 68514 56082
rect 68514 56030 68516 56082
rect 68460 56028 68516 56030
rect 67268 55636 67324 55692
rect 67372 55690 67428 55692
rect 67476 55690 67532 55692
rect 67372 55638 67396 55690
rect 67396 55638 67428 55690
rect 67476 55638 67520 55690
rect 67520 55638 67532 55690
rect 67372 55636 67428 55638
rect 67476 55636 67532 55638
rect 67580 55636 67636 55692
rect 67684 55690 67740 55692
rect 67788 55690 67844 55692
rect 67684 55638 67696 55690
rect 67696 55638 67740 55690
rect 67788 55638 67820 55690
rect 67820 55638 67844 55690
rect 67684 55636 67740 55638
rect 67788 55636 67844 55638
rect 67892 55636 67948 55692
rect 76268 55636 76324 55692
rect 76372 55690 76428 55692
rect 76476 55690 76532 55692
rect 76372 55638 76396 55690
rect 76396 55638 76428 55690
rect 76476 55638 76520 55690
rect 76520 55638 76532 55690
rect 76372 55636 76428 55638
rect 76476 55636 76532 55638
rect 76580 55636 76636 55692
rect 76684 55690 76740 55692
rect 76788 55690 76844 55692
rect 76684 55638 76696 55690
rect 76696 55638 76740 55690
rect 76788 55638 76820 55690
rect 76820 55638 76844 55690
rect 76684 55636 76740 55638
rect 76788 55636 76844 55638
rect 76892 55636 76948 55692
rect 67268 54068 67324 54124
rect 67372 54122 67428 54124
rect 67476 54122 67532 54124
rect 67372 54070 67396 54122
rect 67396 54070 67428 54122
rect 67476 54070 67520 54122
rect 67520 54070 67532 54122
rect 67372 54068 67428 54070
rect 67476 54068 67532 54070
rect 67580 54068 67636 54124
rect 67684 54122 67740 54124
rect 67788 54122 67844 54124
rect 67684 54070 67696 54122
rect 67696 54070 67740 54122
rect 67788 54070 67820 54122
rect 67820 54070 67844 54122
rect 67684 54068 67740 54070
rect 67788 54068 67844 54070
rect 67892 54068 67948 54124
rect 66892 53676 66948 53732
rect 67116 53900 67172 53956
rect 68684 55074 68740 55076
rect 68684 55022 68686 55074
rect 68686 55022 68738 55074
rect 68738 55022 68740 55074
rect 68684 55020 68740 55022
rect 81676 55020 81732 55076
rect 82124 56028 82180 56084
rect 71768 54852 71824 54908
rect 71872 54906 71928 54908
rect 71976 54906 72032 54908
rect 71872 54854 71896 54906
rect 71896 54854 71928 54906
rect 71976 54854 72020 54906
rect 72020 54854 72032 54906
rect 71872 54852 71928 54854
rect 71976 54852 72032 54854
rect 72080 54852 72136 54908
rect 72184 54906 72240 54908
rect 72288 54906 72344 54908
rect 72184 54854 72196 54906
rect 72196 54854 72240 54906
rect 72288 54854 72320 54906
rect 72320 54854 72344 54906
rect 72184 54852 72240 54854
rect 72288 54852 72344 54854
rect 72392 54852 72448 54908
rect 80768 54852 80824 54908
rect 80872 54906 80928 54908
rect 80976 54906 81032 54908
rect 80872 54854 80896 54906
rect 80896 54854 80928 54906
rect 80976 54854 81020 54906
rect 81020 54854 81032 54906
rect 80872 54852 80928 54854
rect 80976 54852 81032 54854
rect 81080 54852 81136 54908
rect 81184 54906 81240 54908
rect 81288 54906 81344 54908
rect 81184 54854 81196 54906
rect 81196 54854 81240 54906
rect 81288 54854 81320 54906
rect 81320 54854 81344 54906
rect 81184 54852 81240 54854
rect 81288 54852 81344 54854
rect 81392 54852 81448 54908
rect 97692 58492 97748 58548
rect 95900 56700 95956 56756
rect 89768 56420 89824 56476
rect 89872 56474 89928 56476
rect 89976 56474 90032 56476
rect 89872 56422 89896 56474
rect 89896 56422 89928 56474
rect 89976 56422 90020 56474
rect 90020 56422 90032 56474
rect 89872 56420 89928 56422
rect 89976 56420 90032 56422
rect 90080 56420 90136 56476
rect 90184 56474 90240 56476
rect 90288 56474 90344 56476
rect 90184 56422 90196 56474
rect 90196 56422 90240 56474
rect 90288 56422 90320 56474
rect 90320 56422 90344 56474
rect 90184 56420 90240 56422
rect 90288 56420 90344 56422
rect 90392 56420 90448 56476
rect 93212 56082 93268 56084
rect 93212 56030 93214 56082
rect 93214 56030 93266 56082
rect 93266 56030 93268 56082
rect 93212 56028 93268 56030
rect 96348 56082 96404 56084
rect 96348 56030 96350 56082
rect 96350 56030 96402 56082
rect 96402 56030 96404 56082
rect 96348 56028 96404 56030
rect 85268 55636 85324 55692
rect 85372 55690 85428 55692
rect 85476 55690 85532 55692
rect 85372 55638 85396 55690
rect 85396 55638 85428 55690
rect 85476 55638 85520 55690
rect 85520 55638 85532 55690
rect 85372 55636 85428 55638
rect 85476 55636 85532 55638
rect 85580 55636 85636 55692
rect 85684 55690 85740 55692
rect 85788 55690 85844 55692
rect 85684 55638 85696 55690
rect 85696 55638 85740 55690
rect 85788 55638 85820 55690
rect 85820 55638 85844 55690
rect 85684 55636 85740 55638
rect 85788 55636 85844 55638
rect 85892 55636 85948 55692
rect 94268 55636 94324 55692
rect 94372 55690 94428 55692
rect 94476 55690 94532 55692
rect 94372 55638 94396 55690
rect 94396 55638 94428 55690
rect 94476 55638 94520 55690
rect 94520 55638 94532 55690
rect 94372 55636 94428 55638
rect 94476 55636 94532 55638
rect 94580 55636 94636 55692
rect 94684 55690 94740 55692
rect 94788 55690 94844 55692
rect 94684 55638 94696 55690
rect 94696 55638 94740 55690
rect 94788 55638 94820 55690
rect 94820 55638 94844 55690
rect 94684 55636 94740 55638
rect 94788 55636 94844 55638
rect 94892 55636 94948 55692
rect 97244 56028 97300 56084
rect 89768 54852 89824 54908
rect 89872 54906 89928 54908
rect 89976 54906 90032 54908
rect 89872 54854 89896 54906
rect 89896 54854 89928 54906
rect 89976 54854 90020 54906
rect 90020 54854 90032 54906
rect 89872 54852 89928 54854
rect 89976 54852 90032 54854
rect 90080 54852 90136 54908
rect 90184 54906 90240 54908
rect 90288 54906 90344 54908
rect 90184 54854 90196 54906
rect 90196 54854 90240 54906
rect 90288 54854 90320 54906
rect 90320 54854 90344 54906
rect 90184 54852 90240 54854
rect 90288 54852 90344 54854
rect 90392 54852 90448 54908
rect 76268 54068 76324 54124
rect 76372 54122 76428 54124
rect 76476 54122 76532 54124
rect 76372 54070 76396 54122
rect 76396 54070 76428 54122
rect 76476 54070 76520 54122
rect 76520 54070 76532 54122
rect 76372 54068 76428 54070
rect 76476 54068 76532 54070
rect 76580 54068 76636 54124
rect 76684 54122 76740 54124
rect 76788 54122 76844 54124
rect 76684 54070 76696 54122
rect 76696 54070 76740 54122
rect 76788 54070 76820 54122
rect 76820 54070 76844 54122
rect 76684 54068 76740 54070
rect 76788 54068 76844 54070
rect 76892 54068 76948 54124
rect 68348 53900 68404 53956
rect 66668 53618 66724 53620
rect 66668 53566 66670 53618
rect 66670 53566 66722 53618
rect 66722 53566 66724 53618
rect 66668 53564 66724 53566
rect 66332 53452 66388 53508
rect 67676 53506 67732 53508
rect 67676 53454 67678 53506
rect 67678 53454 67730 53506
rect 67730 53454 67732 53506
rect 67676 53452 67732 53454
rect 70700 53618 70756 53620
rect 70700 53566 70702 53618
rect 70702 53566 70754 53618
rect 70754 53566 70756 53618
rect 70700 53564 70756 53566
rect 72828 53452 72884 53508
rect 67228 53116 67284 53172
rect 68796 52946 68852 52948
rect 68796 52894 68798 52946
rect 68798 52894 68850 52946
rect 68850 52894 68852 52946
rect 68796 52892 68852 52894
rect 75740 53452 75796 53508
rect 71768 53284 71824 53340
rect 71872 53338 71928 53340
rect 71976 53338 72032 53340
rect 71872 53286 71896 53338
rect 71896 53286 71928 53338
rect 71976 53286 72020 53338
rect 72020 53286 72032 53338
rect 71872 53284 71928 53286
rect 71976 53284 72032 53286
rect 72080 53284 72136 53340
rect 72184 53338 72240 53340
rect 72288 53338 72344 53340
rect 72184 53286 72196 53338
rect 72196 53286 72240 53338
rect 72288 53286 72320 53338
rect 72320 53286 72344 53338
rect 72184 53284 72240 53286
rect 72288 53284 72344 53286
rect 72392 53284 72448 53340
rect 69580 52892 69636 52948
rect 66556 52668 66612 52724
rect 68124 52668 68180 52724
rect 71260 52668 71316 52724
rect 67268 52500 67324 52556
rect 67372 52554 67428 52556
rect 67476 52554 67532 52556
rect 67372 52502 67396 52554
rect 67396 52502 67428 52554
rect 67476 52502 67520 52554
rect 67520 52502 67532 52554
rect 67372 52500 67428 52502
rect 67476 52500 67532 52502
rect 67580 52500 67636 52556
rect 67684 52554 67740 52556
rect 67788 52554 67844 52556
rect 67684 52502 67696 52554
rect 67696 52502 67740 52554
rect 67788 52502 67820 52554
rect 67820 52502 67844 52554
rect 67684 52500 67740 52502
rect 67788 52500 67844 52502
rect 67892 52500 67948 52556
rect 65100 52108 65156 52164
rect 62768 51716 62824 51772
rect 62872 51770 62928 51772
rect 62976 51770 63032 51772
rect 62872 51718 62896 51770
rect 62896 51718 62928 51770
rect 62976 51718 63020 51770
rect 63020 51718 63032 51770
rect 62872 51716 62928 51718
rect 62976 51716 63032 51718
rect 63080 51716 63136 51772
rect 63184 51770 63240 51772
rect 63288 51770 63344 51772
rect 63184 51718 63196 51770
rect 63196 51718 63240 51770
rect 63288 51718 63320 51770
rect 63320 51718 63344 51770
rect 63184 51716 63240 51718
rect 63288 51716 63344 51718
rect 63392 51716 63448 51772
rect 61740 51266 61796 51268
rect 61740 51214 61742 51266
rect 61742 51214 61794 51266
rect 61794 51214 61796 51266
rect 61740 51212 61796 51214
rect 62188 51212 62244 51268
rect 58268 50932 58324 50988
rect 58372 50986 58428 50988
rect 58476 50986 58532 50988
rect 58372 50934 58396 50986
rect 58396 50934 58428 50986
rect 58476 50934 58520 50986
rect 58520 50934 58532 50986
rect 58372 50932 58428 50934
rect 58476 50932 58532 50934
rect 58580 50932 58636 50988
rect 58684 50986 58740 50988
rect 58788 50986 58844 50988
rect 58684 50934 58696 50986
rect 58696 50934 58740 50986
rect 58788 50934 58820 50986
rect 58820 50934 58844 50986
rect 58684 50932 58740 50934
rect 58788 50932 58844 50934
rect 58892 50932 58948 50988
rect 63308 50482 63364 50484
rect 63308 50430 63310 50482
rect 63310 50430 63362 50482
rect 63362 50430 63364 50482
rect 63308 50428 63364 50430
rect 62768 50148 62824 50204
rect 62872 50202 62928 50204
rect 62976 50202 63032 50204
rect 62872 50150 62896 50202
rect 62896 50150 62928 50202
rect 62976 50150 63020 50202
rect 63020 50150 63032 50202
rect 62872 50148 62928 50150
rect 62976 50148 63032 50150
rect 63080 50148 63136 50204
rect 63184 50202 63240 50204
rect 63288 50202 63344 50204
rect 63184 50150 63196 50202
rect 63196 50150 63240 50202
rect 63288 50150 63320 50202
rect 63320 50150 63344 50202
rect 63184 50148 63240 50150
rect 63288 50148 63344 50150
rect 63392 50148 63448 50204
rect 60620 49698 60676 49700
rect 60620 49646 60622 49698
rect 60622 49646 60674 49698
rect 60674 49646 60676 49698
rect 60620 49644 60676 49646
rect 61964 49644 62020 49700
rect 61292 49532 61348 49588
rect 58268 49364 58324 49420
rect 58372 49418 58428 49420
rect 58476 49418 58532 49420
rect 58372 49366 58396 49418
rect 58396 49366 58428 49418
rect 58476 49366 58520 49418
rect 58520 49366 58532 49418
rect 58372 49364 58428 49366
rect 58476 49364 58532 49366
rect 58580 49364 58636 49420
rect 58684 49418 58740 49420
rect 58788 49418 58844 49420
rect 58684 49366 58696 49418
rect 58696 49366 58740 49418
rect 58788 49366 58820 49418
rect 58820 49366 58844 49418
rect 58684 49364 58740 49366
rect 58788 49364 58844 49366
rect 58892 49364 58948 49420
rect 57596 47346 57652 47348
rect 57596 47294 57598 47346
rect 57598 47294 57650 47346
rect 57650 47294 57652 47346
rect 57596 47292 57652 47294
rect 58268 47796 58324 47852
rect 58372 47850 58428 47852
rect 58476 47850 58532 47852
rect 58372 47798 58396 47850
rect 58396 47798 58428 47850
rect 58476 47798 58520 47850
rect 58520 47798 58532 47850
rect 58372 47796 58428 47798
rect 58476 47796 58532 47798
rect 58580 47796 58636 47852
rect 58684 47850 58740 47852
rect 58788 47850 58844 47852
rect 58684 47798 58696 47850
rect 58696 47798 58740 47850
rect 58788 47798 58820 47850
rect 58820 47798 58844 47850
rect 58684 47796 58740 47798
rect 58788 47796 58844 47798
rect 58892 47796 58948 47852
rect 58380 47234 58436 47236
rect 58380 47182 58382 47234
rect 58382 47182 58434 47234
rect 58434 47182 58436 47234
rect 58380 47180 58436 47182
rect 57820 46844 57876 46900
rect 57260 44156 57316 44212
rect 57484 44268 57540 44324
rect 58268 46562 58324 46564
rect 58268 46510 58270 46562
rect 58270 46510 58322 46562
rect 58322 46510 58324 46562
rect 58268 46508 58324 46510
rect 60060 46396 60116 46452
rect 60172 46620 60228 46676
rect 58268 46228 58324 46284
rect 58372 46282 58428 46284
rect 58476 46282 58532 46284
rect 58372 46230 58396 46282
rect 58396 46230 58428 46282
rect 58476 46230 58520 46282
rect 58520 46230 58532 46282
rect 58372 46228 58428 46230
rect 58476 46228 58532 46230
rect 58580 46228 58636 46284
rect 58684 46282 58740 46284
rect 58788 46282 58844 46284
rect 58684 46230 58696 46282
rect 58696 46230 58740 46282
rect 58788 46230 58820 46282
rect 58820 46230 58844 46282
rect 58684 46228 58740 46230
rect 58788 46228 58844 46230
rect 58892 46228 58948 46284
rect 58044 45724 58100 45780
rect 61292 45218 61348 45220
rect 61292 45166 61294 45218
rect 61294 45166 61346 45218
rect 61346 45166 61348 45218
rect 61292 45164 61348 45166
rect 61740 44994 61796 44996
rect 61740 44942 61742 44994
rect 61742 44942 61794 44994
rect 61794 44942 61796 44994
rect 61740 44940 61796 44942
rect 58492 44828 58548 44884
rect 58268 44660 58324 44716
rect 58372 44714 58428 44716
rect 58476 44714 58532 44716
rect 58372 44662 58396 44714
rect 58396 44662 58428 44714
rect 58476 44662 58520 44714
rect 58520 44662 58532 44714
rect 58372 44660 58428 44662
rect 58476 44660 58532 44662
rect 58580 44660 58636 44716
rect 58684 44714 58740 44716
rect 58788 44714 58844 44716
rect 58684 44662 58696 44714
rect 58696 44662 58740 44714
rect 58788 44662 58820 44714
rect 58820 44662 58844 44714
rect 58684 44660 58740 44662
rect 58788 44660 58844 44662
rect 58892 44660 58948 44716
rect 58492 44322 58548 44324
rect 58492 44270 58494 44322
rect 58494 44270 58546 44322
rect 58546 44270 58548 44322
rect 58492 44268 58548 44270
rect 57932 44098 57988 44100
rect 57932 44046 57934 44098
rect 57934 44046 57986 44098
rect 57986 44046 57988 44098
rect 57932 44044 57988 44046
rect 57708 43708 57764 43764
rect 60172 43762 60228 43764
rect 60172 43710 60174 43762
rect 60174 43710 60226 43762
rect 60226 43710 60228 43762
rect 60172 43708 60228 43710
rect 57820 43596 57876 43652
rect 56924 41916 56980 41972
rect 56028 41858 56084 41860
rect 56028 41806 56030 41858
rect 56030 41806 56082 41858
rect 56082 41806 56084 41858
rect 56028 41804 56084 41806
rect 57484 41804 57540 41860
rect 55468 41580 55524 41636
rect 56140 41692 56196 41748
rect 57596 41580 57652 41636
rect 57596 41244 57652 41300
rect 57036 41186 57092 41188
rect 57036 41134 57038 41186
rect 57038 41134 57090 41186
rect 57090 41134 57092 41186
rect 57036 41132 57092 41134
rect 57820 41074 57876 41076
rect 57820 41022 57822 41074
rect 57822 41022 57874 41074
rect 57874 41022 57876 41074
rect 57820 41020 57876 41022
rect 59388 43650 59444 43652
rect 59388 43598 59390 43650
rect 59390 43598 59442 43650
rect 59442 43598 59444 43650
rect 59388 43596 59444 43598
rect 60956 43596 61012 43652
rect 58268 43092 58324 43148
rect 58372 43146 58428 43148
rect 58476 43146 58532 43148
rect 58372 43094 58396 43146
rect 58396 43094 58428 43146
rect 58476 43094 58520 43146
rect 58520 43094 58532 43146
rect 58372 43092 58428 43094
rect 58476 43092 58532 43094
rect 58580 43092 58636 43148
rect 58684 43146 58740 43148
rect 58788 43146 58844 43148
rect 58684 43094 58696 43146
rect 58696 43094 58740 43146
rect 58788 43094 58820 43146
rect 58820 43094 58844 43146
rect 58684 43092 58740 43094
rect 58788 43092 58844 43094
rect 58892 43092 58948 43148
rect 60956 42812 61012 42868
rect 55692 40348 55748 40404
rect 57708 40348 57764 40404
rect 55356 40236 55412 40292
rect 55804 38556 55860 38612
rect 56700 38556 56756 38612
rect 58268 41524 58324 41580
rect 58372 41578 58428 41580
rect 58476 41578 58532 41580
rect 58372 41526 58396 41578
rect 58396 41526 58428 41578
rect 58476 41526 58520 41578
rect 58520 41526 58532 41578
rect 58372 41524 58428 41526
rect 58476 41524 58532 41526
rect 58580 41524 58636 41580
rect 58684 41578 58740 41580
rect 58788 41578 58844 41580
rect 58684 41526 58696 41578
rect 58696 41526 58740 41578
rect 58788 41526 58820 41578
rect 58820 41526 58844 41578
rect 58684 41524 58740 41526
rect 58788 41524 58844 41526
rect 58892 41524 58948 41580
rect 58716 41356 58772 41412
rect 59276 41356 59332 41412
rect 60508 41020 60564 41076
rect 58604 40402 58660 40404
rect 58604 40350 58606 40402
rect 58606 40350 58658 40402
rect 58658 40350 58660 40402
rect 58604 40348 58660 40350
rect 58268 39956 58324 40012
rect 58372 40010 58428 40012
rect 58476 40010 58532 40012
rect 58372 39958 58396 40010
rect 58396 39958 58428 40010
rect 58476 39958 58520 40010
rect 58520 39958 58532 40010
rect 58372 39956 58428 39958
rect 58476 39956 58532 39958
rect 58580 39956 58636 40012
rect 58684 40010 58740 40012
rect 58788 40010 58844 40012
rect 58684 39958 58696 40010
rect 58696 39958 58740 40010
rect 58788 39958 58820 40010
rect 58820 39958 58844 40010
rect 58684 39956 58740 39958
rect 58788 39956 58844 39958
rect 58892 39956 58948 40012
rect 58044 38892 58100 38948
rect 57820 38556 57876 38612
rect 56364 37826 56420 37828
rect 56364 37774 56366 37826
rect 56366 37774 56418 37826
rect 56418 37774 56420 37826
rect 56364 37772 56420 37774
rect 57932 37548 57988 37604
rect 55244 37100 55300 37156
rect 57484 37100 57540 37156
rect 56812 36876 56868 36932
rect 56028 36316 56084 36372
rect 57372 36316 57428 36372
rect 57148 35922 57204 35924
rect 57148 35870 57150 35922
rect 57150 35870 57202 35922
rect 57202 35870 57204 35922
rect 57148 35868 57204 35870
rect 56028 35698 56084 35700
rect 56028 35646 56030 35698
rect 56030 35646 56082 35698
rect 56082 35646 56084 35698
rect 56028 35644 56084 35646
rect 57148 35698 57204 35700
rect 57148 35646 57150 35698
rect 57150 35646 57202 35698
rect 57202 35646 57204 35698
rect 57148 35644 57204 35646
rect 56700 35586 56756 35588
rect 56700 35534 56702 35586
rect 56702 35534 56754 35586
rect 56754 35534 56756 35586
rect 56700 35532 56756 35534
rect 55356 34242 55412 34244
rect 55356 34190 55358 34242
rect 55358 34190 55410 34242
rect 55410 34190 55412 34242
rect 55356 34188 55412 34190
rect 60172 38834 60228 38836
rect 60172 38782 60174 38834
rect 60174 38782 60226 38834
rect 60226 38782 60228 38834
rect 60172 38780 60228 38782
rect 58268 38388 58324 38444
rect 58372 38442 58428 38444
rect 58476 38442 58532 38444
rect 58372 38390 58396 38442
rect 58396 38390 58428 38442
rect 58476 38390 58520 38442
rect 58520 38390 58532 38442
rect 58372 38388 58428 38390
rect 58476 38388 58532 38390
rect 58580 38388 58636 38444
rect 58684 38442 58740 38444
rect 58788 38442 58844 38444
rect 58684 38390 58696 38442
rect 58696 38390 58740 38442
rect 58788 38390 58820 38442
rect 58820 38390 58844 38442
rect 58684 38388 58740 38390
rect 58788 38388 58844 38390
rect 58892 38388 58948 38444
rect 59276 37938 59332 37940
rect 59276 37886 59278 37938
rect 59278 37886 59330 37938
rect 59330 37886 59332 37938
rect 59276 37884 59332 37886
rect 59948 37826 60004 37828
rect 59948 37774 59950 37826
rect 59950 37774 60002 37826
rect 60002 37774 60004 37826
rect 59948 37772 60004 37774
rect 61852 42866 61908 42868
rect 61852 42814 61854 42866
rect 61854 42814 61906 42866
rect 61906 42814 61908 42866
rect 61852 42812 61908 42814
rect 61740 41132 61796 41188
rect 62300 49644 62356 49700
rect 62076 49586 62132 49588
rect 62076 49534 62078 49586
rect 62078 49534 62130 49586
rect 62130 49534 62132 49586
rect 62076 49532 62132 49534
rect 62860 49532 62916 49588
rect 62768 48580 62824 48636
rect 62872 48634 62928 48636
rect 62976 48634 63032 48636
rect 62872 48582 62896 48634
rect 62896 48582 62928 48634
rect 62976 48582 63020 48634
rect 63020 48582 63032 48634
rect 62872 48580 62928 48582
rect 62976 48580 63032 48582
rect 63080 48580 63136 48636
rect 63184 48634 63240 48636
rect 63288 48634 63344 48636
rect 63184 48582 63196 48634
rect 63196 48582 63240 48634
rect 63288 48582 63320 48634
rect 63320 48582 63344 48634
rect 63184 48580 63240 48582
rect 63288 48580 63344 48582
rect 63392 48580 63448 48636
rect 62768 47012 62824 47068
rect 62872 47066 62928 47068
rect 62976 47066 63032 47068
rect 62872 47014 62896 47066
rect 62896 47014 62928 47066
rect 62976 47014 63020 47066
rect 63020 47014 63032 47066
rect 62872 47012 62928 47014
rect 62976 47012 63032 47014
rect 63080 47012 63136 47068
rect 63184 47066 63240 47068
rect 63288 47066 63344 47068
rect 63184 47014 63196 47066
rect 63196 47014 63240 47066
rect 63288 47014 63320 47066
rect 63320 47014 63344 47066
rect 63184 47012 63240 47014
rect 63288 47012 63344 47014
rect 63392 47012 63448 47068
rect 62636 45612 62692 45668
rect 62076 45164 62132 45220
rect 64540 50482 64596 50484
rect 64540 50430 64542 50482
rect 64542 50430 64594 50482
rect 64594 50430 64596 50482
rect 64540 50428 64596 50430
rect 64092 49532 64148 49588
rect 63644 49420 63700 49476
rect 64988 49756 65044 49812
rect 64876 49532 64932 49588
rect 63644 48972 63700 49028
rect 64204 48914 64260 48916
rect 64204 48862 64206 48914
rect 64206 48862 64258 48914
rect 64258 48862 64260 48914
rect 64204 48860 64260 48862
rect 63868 48466 63924 48468
rect 63868 48414 63870 48466
rect 63870 48414 63922 48466
rect 63922 48414 63924 48466
rect 63868 48412 63924 48414
rect 64540 48354 64596 48356
rect 64540 48302 64542 48354
rect 64542 48302 64594 48354
rect 64594 48302 64596 48354
rect 64540 48300 64596 48302
rect 67268 50932 67324 50988
rect 67372 50986 67428 50988
rect 67476 50986 67532 50988
rect 67372 50934 67396 50986
rect 67396 50934 67428 50986
rect 67476 50934 67520 50986
rect 67520 50934 67532 50986
rect 67372 50932 67428 50934
rect 67476 50932 67532 50934
rect 67580 50932 67636 50988
rect 67684 50986 67740 50988
rect 67788 50986 67844 50988
rect 67684 50934 67696 50986
rect 67696 50934 67740 50986
rect 67788 50934 67820 50986
rect 67820 50934 67844 50986
rect 67684 50932 67740 50934
rect 67788 50932 67844 50934
rect 67892 50932 67948 50988
rect 68124 50316 68180 50372
rect 69244 50316 69300 50372
rect 65772 49810 65828 49812
rect 65772 49758 65774 49810
rect 65774 49758 65826 49810
rect 65826 49758 65828 49810
rect 65772 49756 65828 49758
rect 71768 51716 71824 51772
rect 71872 51770 71928 51772
rect 71976 51770 72032 51772
rect 71872 51718 71896 51770
rect 71896 51718 71928 51770
rect 71976 51718 72020 51770
rect 72020 51718 72032 51770
rect 71872 51716 71928 51718
rect 71976 51716 72032 51718
rect 72080 51716 72136 51772
rect 72184 51770 72240 51772
rect 72288 51770 72344 51772
rect 72184 51718 72196 51770
rect 72196 51718 72240 51770
rect 72288 51718 72320 51770
rect 72320 51718 72344 51770
rect 72184 51716 72240 51718
rect 72288 51716 72344 51718
rect 72392 51716 72448 51772
rect 71372 51490 71428 51492
rect 71372 51438 71374 51490
rect 71374 51438 71426 51490
rect 71426 51438 71428 51490
rect 71372 51436 71428 51438
rect 72492 51436 72548 51492
rect 71768 50148 71824 50204
rect 71872 50202 71928 50204
rect 71976 50202 72032 50204
rect 71872 50150 71896 50202
rect 71896 50150 71928 50202
rect 71976 50150 72020 50202
rect 72020 50150 72032 50202
rect 71872 50148 71928 50150
rect 71976 50148 72032 50150
rect 72080 50148 72136 50204
rect 72184 50202 72240 50204
rect 72288 50202 72344 50204
rect 72184 50150 72196 50202
rect 72196 50150 72240 50202
rect 72288 50150 72320 50202
rect 72320 50150 72344 50202
rect 72184 50148 72240 50150
rect 72288 50148 72344 50150
rect 72392 50148 72448 50204
rect 74284 51212 74340 51268
rect 73164 50482 73220 50484
rect 73164 50430 73166 50482
rect 73166 50430 73218 50482
rect 73218 50430 73220 50482
rect 73164 50428 73220 50430
rect 65884 49532 65940 49588
rect 65100 49026 65156 49028
rect 65100 48974 65102 49026
rect 65102 48974 65154 49026
rect 65154 48974 65156 49026
rect 65100 48972 65156 48974
rect 68908 49586 68964 49588
rect 68908 49534 68910 49586
rect 68910 49534 68962 49586
rect 68962 49534 68964 49586
rect 68908 49532 68964 49534
rect 67268 49364 67324 49420
rect 67372 49418 67428 49420
rect 67476 49418 67532 49420
rect 67372 49366 67396 49418
rect 67396 49366 67428 49418
rect 67476 49366 67520 49418
rect 67520 49366 67532 49418
rect 67372 49364 67428 49366
rect 67476 49364 67532 49366
rect 67580 49364 67636 49420
rect 67684 49418 67740 49420
rect 67788 49418 67844 49420
rect 67684 49366 67696 49418
rect 67696 49366 67740 49418
rect 67788 49366 67820 49418
rect 67820 49366 67844 49418
rect 67684 49364 67740 49366
rect 67788 49364 67844 49366
rect 67892 49364 67948 49420
rect 65324 48914 65380 48916
rect 65324 48862 65326 48914
rect 65326 48862 65378 48914
rect 65378 48862 65380 48914
rect 65324 48860 65380 48862
rect 71708 49698 71764 49700
rect 71708 49646 71710 49698
rect 71710 49646 71762 49698
rect 71762 49646 71764 49698
rect 71708 49644 71764 49646
rect 72940 49644 72996 49700
rect 71260 48972 71316 49028
rect 65548 48412 65604 48468
rect 65100 48354 65156 48356
rect 65100 48302 65102 48354
rect 65102 48302 65154 48354
rect 65154 48302 65156 48354
rect 65100 48300 65156 48302
rect 64540 47516 64596 47572
rect 63868 47180 63924 47236
rect 64652 45836 64708 45892
rect 62768 45444 62824 45500
rect 62872 45498 62928 45500
rect 62976 45498 63032 45500
rect 62872 45446 62896 45498
rect 62896 45446 62928 45498
rect 62976 45446 63020 45498
rect 63020 45446 63032 45498
rect 62872 45444 62928 45446
rect 62976 45444 63032 45446
rect 63080 45444 63136 45500
rect 63184 45498 63240 45500
rect 63288 45498 63344 45500
rect 63184 45446 63196 45498
rect 63196 45446 63240 45498
rect 63288 45446 63320 45498
rect 63320 45446 63344 45498
rect 63184 45444 63240 45446
rect 63288 45444 63344 45446
rect 63392 45444 63448 45500
rect 64092 45666 64148 45668
rect 64092 45614 64094 45666
rect 64094 45614 64146 45666
rect 64146 45614 64148 45666
rect 64092 45612 64148 45614
rect 64652 45666 64708 45668
rect 64652 45614 64654 45666
rect 64654 45614 64706 45666
rect 64706 45614 64708 45666
rect 64652 45612 64708 45614
rect 63532 45388 63588 45444
rect 64540 45388 64596 45444
rect 63308 45218 63364 45220
rect 63308 45166 63310 45218
rect 63310 45166 63362 45218
rect 63362 45166 63364 45218
rect 63308 45164 63364 45166
rect 61964 41020 62020 41076
rect 62076 44940 62132 44996
rect 63532 44940 63588 44996
rect 63084 44492 63140 44548
rect 64428 44546 64484 44548
rect 64428 44494 64430 44546
rect 64430 44494 64482 44546
rect 64482 44494 64484 44546
rect 64428 44492 64484 44494
rect 63532 44098 63588 44100
rect 63532 44046 63534 44098
rect 63534 44046 63586 44098
rect 63586 44046 63588 44098
rect 63532 44044 63588 44046
rect 62768 43876 62824 43932
rect 62872 43930 62928 43932
rect 62976 43930 63032 43932
rect 62872 43878 62896 43930
rect 62896 43878 62928 43930
rect 62976 43878 63020 43930
rect 63020 43878 63032 43930
rect 62872 43876 62928 43878
rect 62976 43876 63032 43878
rect 63080 43876 63136 43932
rect 63184 43930 63240 43932
rect 63288 43930 63344 43932
rect 63184 43878 63196 43930
rect 63196 43878 63240 43930
rect 63288 43878 63320 43930
rect 63320 43878 63344 43930
rect 63184 43876 63240 43878
rect 63288 43876 63344 43878
rect 63392 43876 63448 43932
rect 63420 43708 63476 43764
rect 64092 43708 64148 43764
rect 64652 44044 64708 44100
rect 64540 43426 64596 43428
rect 64540 43374 64542 43426
rect 64542 43374 64594 43426
rect 64594 43374 64596 43426
rect 64540 43372 64596 43374
rect 62768 42308 62824 42364
rect 62872 42362 62928 42364
rect 62976 42362 63032 42364
rect 62872 42310 62896 42362
rect 62896 42310 62928 42362
rect 62976 42310 63020 42362
rect 63020 42310 63032 42362
rect 62872 42308 62928 42310
rect 62976 42308 63032 42310
rect 63080 42308 63136 42364
rect 63184 42362 63240 42364
rect 63288 42362 63344 42364
rect 63184 42310 63196 42362
rect 63196 42310 63240 42362
rect 63288 42310 63320 42362
rect 63320 42310 63344 42362
rect 63184 42308 63240 42310
rect 63288 42308 63344 42310
rect 63392 42308 63448 42364
rect 62076 40908 62132 40964
rect 60956 39004 61012 39060
rect 60956 38780 61012 38836
rect 60620 37938 60676 37940
rect 60620 37886 60622 37938
rect 60622 37886 60674 37938
rect 60674 37886 60676 37938
rect 60620 37884 60676 37886
rect 60508 37772 60564 37828
rect 61180 37772 61236 37828
rect 61740 37938 61796 37940
rect 61740 37886 61742 37938
rect 61742 37886 61794 37938
rect 61794 37886 61796 37938
rect 61740 37884 61796 37886
rect 60956 37548 61012 37604
rect 59948 36988 60004 37044
rect 58268 36820 58324 36876
rect 58372 36874 58428 36876
rect 58476 36874 58532 36876
rect 58372 36822 58396 36874
rect 58396 36822 58428 36874
rect 58476 36822 58520 36874
rect 58520 36822 58532 36874
rect 58372 36820 58428 36822
rect 58476 36820 58532 36822
rect 58580 36820 58636 36876
rect 58684 36874 58740 36876
rect 58788 36874 58844 36876
rect 58684 36822 58696 36874
rect 58696 36822 58740 36874
rect 58788 36822 58820 36874
rect 58820 36822 58844 36874
rect 58684 36820 58740 36822
rect 58788 36820 58844 36822
rect 58892 36820 58948 36876
rect 57372 34242 57428 34244
rect 57372 34190 57374 34242
rect 57374 34190 57426 34242
rect 57426 34190 57428 34242
rect 57372 34188 57428 34190
rect 57820 35532 57876 35588
rect 58268 35252 58324 35308
rect 58372 35306 58428 35308
rect 58476 35306 58532 35308
rect 58372 35254 58396 35306
rect 58396 35254 58428 35306
rect 58476 35254 58520 35306
rect 58520 35254 58532 35306
rect 58372 35252 58428 35254
rect 58476 35252 58532 35254
rect 58580 35252 58636 35308
rect 58684 35306 58740 35308
rect 58788 35306 58844 35308
rect 58684 35254 58696 35306
rect 58696 35254 58740 35306
rect 58788 35254 58820 35306
rect 58820 35254 58844 35306
rect 58684 35252 58740 35254
rect 58788 35252 58844 35254
rect 58892 35252 58948 35308
rect 57708 34860 57764 34916
rect 58940 34914 58996 34916
rect 58940 34862 58942 34914
rect 58942 34862 58994 34914
rect 58994 34862 58996 34914
rect 58940 34860 58996 34862
rect 61516 34748 61572 34804
rect 58156 34412 58212 34468
rect 60732 34524 60788 34580
rect 55244 32786 55300 32788
rect 55244 32734 55246 32786
rect 55246 32734 55298 32786
rect 55298 32734 55300 32786
rect 55244 32732 55300 32734
rect 55692 32786 55748 32788
rect 55692 32734 55694 32786
rect 55694 32734 55746 32786
rect 55746 32734 55748 32786
rect 55692 32732 55748 32734
rect 56364 32732 56420 32788
rect 58268 33684 58324 33740
rect 58372 33738 58428 33740
rect 58476 33738 58532 33740
rect 58372 33686 58396 33738
rect 58396 33686 58428 33738
rect 58476 33686 58520 33738
rect 58520 33686 58532 33738
rect 58372 33684 58428 33686
rect 58476 33684 58532 33686
rect 58580 33684 58636 33740
rect 58684 33738 58740 33740
rect 58788 33738 58844 33740
rect 58684 33686 58696 33738
rect 58696 33686 58740 33738
rect 58788 33686 58820 33738
rect 58820 33686 58844 33738
rect 58684 33684 58740 33686
rect 58788 33684 58844 33686
rect 58892 33684 58948 33740
rect 59836 33180 59892 33236
rect 57148 32732 57204 32788
rect 57820 32732 57876 32788
rect 56028 32674 56084 32676
rect 56028 32622 56030 32674
rect 56030 32622 56082 32674
rect 56082 32622 56084 32674
rect 56028 32620 56084 32622
rect 57260 32674 57316 32676
rect 57260 32622 57262 32674
rect 57262 32622 57314 32674
rect 57314 32622 57316 32674
rect 57260 32620 57316 32622
rect 59836 32620 59892 32676
rect 60284 33068 60340 33124
rect 57036 32562 57092 32564
rect 57036 32510 57038 32562
rect 57038 32510 57090 32562
rect 57090 32510 57092 32562
rect 57036 32508 57092 32510
rect 59164 32508 59220 32564
rect 53116 32060 53172 32116
rect 47180 30994 47236 30996
rect 47180 30942 47182 30994
rect 47182 30942 47234 30994
rect 47234 30942 47236 30994
rect 47180 30940 47236 30942
rect 46956 30882 47012 30884
rect 46956 30830 46958 30882
rect 46958 30830 47010 30882
rect 47010 30830 47012 30882
rect 46956 30828 47012 30830
rect 46844 30156 46900 30212
rect 47068 30210 47124 30212
rect 47068 30158 47070 30210
rect 47070 30158 47122 30210
rect 47122 30158 47124 30210
rect 47068 30156 47124 30158
rect 49268 30548 49324 30604
rect 49372 30602 49428 30604
rect 49476 30602 49532 30604
rect 49372 30550 49396 30602
rect 49396 30550 49428 30602
rect 49476 30550 49520 30602
rect 49520 30550 49532 30602
rect 49372 30548 49428 30550
rect 49476 30548 49532 30550
rect 49580 30548 49636 30604
rect 49684 30602 49740 30604
rect 49788 30602 49844 30604
rect 49684 30550 49696 30602
rect 49696 30550 49740 30602
rect 49788 30550 49820 30602
rect 49820 30550 49844 30602
rect 49684 30548 49740 30550
rect 49788 30548 49844 30550
rect 49892 30548 49948 30604
rect 49756 30210 49812 30212
rect 49756 30158 49758 30210
rect 49758 30158 49810 30210
rect 49810 30158 49812 30210
rect 49756 30156 49812 30158
rect 49196 30098 49252 30100
rect 49196 30046 49198 30098
rect 49198 30046 49250 30098
rect 49250 30046 49252 30098
rect 49196 30044 49252 30046
rect 49308 29708 49364 29764
rect 46956 29426 47012 29428
rect 46956 29374 46958 29426
rect 46958 29374 47010 29426
rect 47010 29374 47012 29426
rect 46956 29372 47012 29374
rect 50540 29708 50596 29764
rect 49756 29148 49812 29204
rect 49268 28980 49324 29036
rect 49372 29034 49428 29036
rect 49476 29034 49532 29036
rect 49372 28982 49396 29034
rect 49396 28982 49428 29034
rect 49476 28982 49520 29034
rect 49520 28982 49532 29034
rect 49372 28980 49428 28982
rect 49476 28980 49532 28982
rect 49580 28980 49636 29036
rect 49684 29034 49740 29036
rect 49788 29034 49844 29036
rect 49684 28982 49696 29034
rect 49696 28982 49740 29034
rect 49788 28982 49820 29034
rect 49820 28982 49844 29034
rect 49684 28980 49740 28982
rect 49788 28980 49844 28982
rect 49892 28980 49948 29036
rect 48076 27804 48132 27860
rect 51772 27916 51828 27972
rect 49196 27858 49252 27860
rect 49196 27806 49198 27858
rect 49198 27806 49250 27858
rect 49250 27806 49252 27858
rect 49196 27804 49252 27806
rect 46844 27746 46900 27748
rect 46844 27694 46846 27746
rect 46846 27694 46898 27746
rect 46898 27694 46900 27746
rect 46844 27692 46900 27694
rect 49268 27412 49324 27468
rect 49372 27466 49428 27468
rect 49476 27466 49532 27468
rect 49372 27414 49396 27466
rect 49396 27414 49428 27466
rect 49476 27414 49520 27466
rect 49520 27414 49532 27466
rect 49372 27412 49428 27414
rect 49476 27412 49532 27414
rect 49580 27412 49636 27468
rect 49684 27466 49740 27468
rect 49788 27466 49844 27468
rect 49684 27414 49696 27466
rect 49696 27414 49740 27466
rect 49788 27414 49820 27466
rect 49820 27414 49844 27466
rect 49684 27412 49740 27414
rect 49788 27412 49844 27414
rect 49892 27412 49948 27468
rect 48412 26236 48468 26292
rect 50428 26290 50484 26292
rect 50428 26238 50430 26290
rect 50430 26238 50482 26290
rect 50482 26238 50484 26290
rect 50428 26236 50484 26238
rect 49268 25844 49324 25900
rect 49372 25898 49428 25900
rect 49476 25898 49532 25900
rect 49372 25846 49396 25898
rect 49396 25846 49428 25898
rect 49476 25846 49520 25898
rect 49520 25846 49532 25898
rect 49372 25844 49428 25846
rect 49476 25844 49532 25846
rect 49580 25844 49636 25900
rect 49684 25898 49740 25900
rect 49788 25898 49844 25900
rect 49684 25846 49696 25898
rect 49696 25846 49740 25898
rect 49788 25846 49820 25898
rect 49820 25846 49844 25898
rect 49684 25844 49740 25846
rect 49788 25844 49844 25846
rect 49892 25844 49948 25900
rect 47628 25282 47684 25284
rect 47628 25230 47630 25282
rect 47630 25230 47682 25282
rect 47682 25230 47684 25282
rect 47628 25228 47684 25230
rect 49268 24276 49324 24332
rect 49372 24330 49428 24332
rect 49476 24330 49532 24332
rect 49372 24278 49396 24330
rect 49396 24278 49428 24330
rect 49476 24278 49520 24330
rect 49520 24278 49532 24330
rect 49372 24276 49428 24278
rect 49476 24276 49532 24278
rect 49580 24276 49636 24332
rect 49684 24330 49740 24332
rect 49788 24330 49844 24332
rect 49684 24278 49696 24330
rect 49696 24278 49740 24330
rect 49788 24278 49820 24330
rect 49820 24278 49844 24330
rect 49684 24276 49740 24278
rect 49788 24276 49844 24278
rect 49892 24276 49948 24332
rect 49268 22708 49324 22764
rect 49372 22762 49428 22764
rect 49476 22762 49532 22764
rect 49372 22710 49396 22762
rect 49396 22710 49428 22762
rect 49476 22710 49520 22762
rect 49520 22710 49532 22762
rect 49372 22708 49428 22710
rect 49476 22708 49532 22710
rect 49580 22708 49636 22764
rect 49684 22762 49740 22764
rect 49788 22762 49844 22764
rect 49684 22710 49696 22762
rect 49696 22710 49740 22762
rect 49788 22710 49820 22762
rect 49820 22710 49844 22762
rect 49684 22708 49740 22710
rect 49788 22708 49844 22710
rect 49892 22708 49948 22764
rect 46956 21420 47012 21476
rect 49268 21140 49324 21196
rect 49372 21194 49428 21196
rect 49476 21194 49532 21196
rect 49372 21142 49396 21194
rect 49396 21142 49428 21194
rect 49476 21142 49520 21194
rect 49520 21142 49532 21194
rect 49372 21140 49428 21142
rect 49476 21140 49532 21142
rect 49580 21140 49636 21196
rect 49684 21194 49740 21196
rect 49788 21194 49844 21196
rect 49684 21142 49696 21194
rect 49696 21142 49740 21194
rect 49788 21142 49820 21194
rect 49820 21142 49844 21194
rect 49684 21140 49740 21142
rect 49788 21140 49844 21142
rect 49892 21140 49948 21196
rect 46956 20636 47012 20692
rect 49268 19572 49324 19628
rect 49372 19626 49428 19628
rect 49476 19626 49532 19628
rect 49372 19574 49396 19626
rect 49396 19574 49428 19626
rect 49476 19574 49520 19626
rect 49520 19574 49532 19626
rect 49372 19572 49428 19574
rect 49476 19572 49532 19574
rect 49580 19572 49636 19628
rect 49684 19626 49740 19628
rect 49788 19626 49844 19628
rect 49684 19574 49696 19626
rect 49696 19574 49740 19626
rect 49788 19574 49820 19626
rect 49820 19574 49844 19626
rect 49684 19572 49740 19574
rect 49788 19572 49844 19574
rect 49892 19572 49948 19628
rect 49268 18004 49324 18060
rect 49372 18058 49428 18060
rect 49476 18058 49532 18060
rect 49372 18006 49396 18058
rect 49396 18006 49428 18058
rect 49476 18006 49520 18058
rect 49520 18006 49532 18058
rect 49372 18004 49428 18006
rect 49476 18004 49532 18006
rect 49580 18004 49636 18060
rect 49684 18058 49740 18060
rect 49788 18058 49844 18060
rect 49684 18006 49696 18058
rect 49696 18006 49740 18058
rect 49788 18006 49820 18058
rect 49820 18006 49844 18058
rect 49684 18004 49740 18006
rect 49788 18004 49844 18006
rect 49892 18004 49948 18060
rect 49268 16436 49324 16492
rect 49372 16490 49428 16492
rect 49476 16490 49532 16492
rect 49372 16438 49396 16490
rect 49396 16438 49428 16490
rect 49476 16438 49520 16490
rect 49520 16438 49532 16490
rect 49372 16436 49428 16438
rect 49476 16436 49532 16438
rect 49580 16436 49636 16492
rect 49684 16490 49740 16492
rect 49788 16490 49844 16492
rect 49684 16438 49696 16490
rect 49696 16438 49740 16490
rect 49788 16438 49820 16490
rect 49820 16438 49844 16490
rect 49684 16436 49740 16438
rect 49788 16436 49844 16438
rect 49892 16436 49948 16492
rect 49268 14868 49324 14924
rect 49372 14922 49428 14924
rect 49476 14922 49532 14924
rect 49372 14870 49396 14922
rect 49396 14870 49428 14922
rect 49476 14870 49520 14922
rect 49520 14870 49532 14922
rect 49372 14868 49428 14870
rect 49476 14868 49532 14870
rect 49580 14868 49636 14924
rect 49684 14922 49740 14924
rect 49788 14922 49844 14924
rect 49684 14870 49696 14922
rect 49696 14870 49740 14922
rect 49788 14870 49820 14922
rect 49820 14870 49844 14922
rect 49684 14868 49740 14870
rect 49788 14868 49844 14870
rect 49892 14868 49948 14924
rect 44768 14084 44824 14140
rect 44872 14138 44928 14140
rect 44976 14138 45032 14140
rect 44872 14086 44896 14138
rect 44896 14086 44928 14138
rect 44976 14086 45020 14138
rect 45020 14086 45032 14138
rect 44872 14084 44928 14086
rect 44976 14084 45032 14086
rect 45080 14084 45136 14140
rect 45184 14138 45240 14140
rect 45288 14138 45344 14140
rect 45184 14086 45196 14138
rect 45196 14086 45240 14138
rect 45288 14086 45320 14138
rect 45320 14086 45344 14138
rect 45184 14084 45240 14086
rect 45288 14084 45344 14086
rect 45392 14084 45448 14140
rect 45388 13692 45444 13748
rect 44768 12516 44824 12572
rect 44872 12570 44928 12572
rect 44976 12570 45032 12572
rect 44872 12518 44896 12570
rect 44896 12518 44928 12570
rect 44976 12518 45020 12570
rect 45020 12518 45032 12570
rect 44872 12516 44928 12518
rect 44976 12516 45032 12518
rect 45080 12516 45136 12572
rect 45184 12570 45240 12572
rect 45288 12570 45344 12572
rect 45184 12518 45196 12570
rect 45196 12518 45240 12570
rect 45288 12518 45320 12570
rect 45320 12518 45344 12570
rect 45184 12516 45240 12518
rect 45288 12516 45344 12518
rect 45392 12516 45448 12572
rect 44604 11452 44660 11508
rect 45948 14476 46004 14532
rect 45612 11452 45668 11508
rect 44768 10948 44824 11004
rect 44872 11002 44928 11004
rect 44976 11002 45032 11004
rect 44872 10950 44896 11002
rect 44896 10950 44928 11002
rect 44976 10950 45020 11002
rect 45020 10950 45032 11002
rect 44872 10948 44928 10950
rect 44976 10948 45032 10950
rect 45080 10948 45136 11004
rect 45184 11002 45240 11004
rect 45288 11002 45344 11004
rect 45184 10950 45196 11002
rect 45196 10950 45240 11002
rect 45288 10950 45320 11002
rect 45320 10950 45344 11002
rect 45184 10948 45240 10950
rect 45288 10948 45344 10950
rect 45392 10948 45448 11004
rect 45052 9938 45108 9940
rect 45052 9886 45054 9938
rect 45054 9886 45106 9938
rect 45106 9886 45108 9938
rect 45052 9884 45108 9886
rect 45164 9602 45220 9604
rect 45164 9550 45166 9602
rect 45166 9550 45218 9602
rect 45218 9550 45220 9602
rect 45164 9548 45220 9550
rect 44768 9380 44824 9436
rect 44872 9434 44928 9436
rect 44976 9434 45032 9436
rect 44872 9382 44896 9434
rect 44896 9382 44928 9434
rect 44976 9382 45020 9434
rect 45020 9382 45032 9434
rect 44872 9380 44928 9382
rect 44976 9380 45032 9382
rect 45080 9380 45136 9436
rect 45184 9434 45240 9436
rect 45288 9434 45344 9436
rect 45184 9382 45196 9434
rect 45196 9382 45240 9434
rect 45288 9382 45320 9434
rect 45320 9382 45344 9434
rect 45184 9380 45240 9382
rect 45288 9380 45344 9382
rect 45392 9380 45448 9436
rect 45388 9212 45444 9268
rect 44828 8146 44884 8148
rect 44828 8094 44830 8146
rect 44830 8094 44882 8146
rect 44882 8094 44884 8146
rect 44828 8092 44884 8094
rect 44768 7812 44824 7868
rect 44872 7866 44928 7868
rect 44976 7866 45032 7868
rect 44872 7814 44896 7866
rect 44896 7814 44928 7866
rect 44976 7814 45020 7866
rect 45020 7814 45032 7866
rect 44872 7812 44928 7814
rect 44976 7812 45032 7814
rect 45080 7812 45136 7868
rect 45184 7866 45240 7868
rect 45288 7866 45344 7868
rect 45184 7814 45196 7866
rect 45196 7814 45240 7866
rect 45288 7814 45320 7866
rect 45320 7814 45344 7866
rect 45184 7812 45240 7814
rect 45288 7812 45344 7814
rect 45392 7812 45448 7868
rect 44380 5180 44436 5236
rect 45388 6636 45444 6692
rect 46732 14530 46788 14532
rect 46732 14478 46734 14530
rect 46734 14478 46786 14530
rect 46786 14478 46788 14530
rect 46732 14476 46788 14478
rect 47068 14364 47124 14420
rect 52108 14252 52164 14308
rect 52444 27692 52500 27748
rect 48972 13916 49028 13972
rect 46172 13692 46228 13748
rect 46060 13580 46116 13636
rect 47180 12908 47236 12964
rect 47740 12796 47796 12852
rect 46844 12236 46900 12292
rect 46508 12124 46564 12180
rect 46172 9884 46228 9940
rect 45836 8876 45892 8932
rect 45388 6466 45444 6468
rect 45388 6414 45390 6466
rect 45390 6414 45442 6466
rect 45442 6414 45444 6466
rect 45388 6412 45444 6414
rect 44768 6244 44824 6300
rect 44872 6298 44928 6300
rect 44976 6298 45032 6300
rect 44872 6246 44896 6298
rect 44896 6246 44928 6298
rect 44976 6246 45020 6298
rect 45020 6246 45032 6298
rect 44872 6244 44928 6246
rect 44976 6244 45032 6246
rect 45080 6244 45136 6300
rect 45184 6298 45240 6300
rect 45288 6298 45344 6300
rect 45184 6246 45196 6298
rect 45196 6246 45240 6298
rect 45288 6246 45320 6298
rect 45320 6246 45344 6298
rect 45184 6244 45240 6246
rect 45288 6244 45344 6246
rect 45392 6244 45448 6300
rect 44940 6076 44996 6132
rect 44940 5234 44996 5236
rect 44940 5182 44942 5234
rect 44942 5182 44994 5234
rect 44994 5182 44996 5234
rect 44940 5180 44996 5182
rect 45276 4956 45332 5012
rect 45836 6636 45892 6692
rect 44604 4732 44660 4788
rect 44768 4676 44824 4732
rect 44872 4730 44928 4732
rect 44976 4730 45032 4732
rect 44872 4678 44896 4730
rect 44896 4678 44928 4730
rect 44976 4678 45020 4730
rect 45020 4678 45032 4730
rect 44872 4676 44928 4678
rect 44976 4676 45032 4678
rect 45080 4676 45136 4732
rect 45184 4730 45240 4732
rect 45288 4730 45344 4732
rect 45184 4678 45196 4730
rect 45196 4678 45240 4730
rect 45288 4678 45320 4730
rect 45320 4678 45344 4730
rect 45184 4676 45240 4678
rect 45288 4676 45344 4678
rect 45392 4676 45448 4732
rect 46284 8258 46340 8260
rect 46284 8206 46286 8258
rect 46286 8206 46338 8258
rect 46338 8206 46340 8258
rect 46284 8204 46340 8206
rect 46060 6412 46116 6468
rect 46172 8092 46228 8148
rect 46284 7980 46340 8036
rect 46396 5964 46452 6020
rect 46284 5628 46340 5684
rect 46620 4898 46676 4900
rect 46620 4846 46622 4898
rect 46622 4846 46674 4898
rect 46674 4846 46676 4898
rect 46620 4844 46676 4846
rect 45276 3778 45332 3780
rect 45276 3726 45278 3778
rect 45278 3726 45330 3778
rect 45330 3726 45332 3778
rect 45276 3724 45332 3726
rect 47180 12012 47236 12068
rect 47068 11282 47124 11284
rect 47068 11230 47070 11282
rect 47070 11230 47122 11282
rect 47122 11230 47124 11282
rect 47068 11228 47124 11230
rect 47068 6748 47124 6804
rect 48860 12290 48916 12292
rect 48860 12238 48862 12290
rect 48862 12238 48914 12290
rect 48914 12238 48916 12290
rect 48860 12236 48916 12238
rect 48748 12178 48804 12180
rect 48748 12126 48750 12178
rect 48750 12126 48802 12178
rect 48802 12126 48804 12178
rect 48748 12124 48804 12126
rect 48188 12066 48244 12068
rect 48188 12014 48190 12066
rect 48190 12014 48242 12066
rect 48242 12014 48244 12066
rect 48188 12012 48244 12014
rect 51660 13804 51716 13860
rect 53452 32338 53508 32340
rect 53452 32286 53454 32338
rect 53454 32286 53506 32338
rect 53506 32286 53508 32338
rect 53452 32284 53508 32286
rect 54460 32060 54516 32116
rect 58268 32116 58324 32172
rect 58372 32170 58428 32172
rect 58476 32170 58532 32172
rect 58372 32118 58396 32170
rect 58396 32118 58428 32170
rect 58476 32118 58520 32170
rect 58520 32118 58532 32170
rect 58372 32116 58428 32118
rect 58476 32116 58532 32118
rect 58580 32116 58636 32172
rect 58684 32170 58740 32172
rect 58788 32170 58844 32172
rect 58684 32118 58696 32170
rect 58696 32118 58740 32170
rect 58788 32118 58820 32170
rect 58820 32118 58844 32170
rect 58684 32116 58740 32118
rect 58788 32116 58844 32118
rect 58892 32116 58948 32172
rect 55356 31500 55412 31556
rect 53768 31332 53824 31388
rect 53872 31386 53928 31388
rect 53976 31386 54032 31388
rect 53872 31334 53896 31386
rect 53896 31334 53928 31386
rect 53976 31334 54020 31386
rect 54020 31334 54032 31386
rect 53872 31332 53928 31334
rect 53976 31332 54032 31334
rect 54080 31332 54136 31388
rect 54184 31386 54240 31388
rect 54288 31386 54344 31388
rect 54184 31334 54196 31386
rect 54196 31334 54240 31386
rect 54288 31334 54320 31386
rect 54320 31334 54344 31386
rect 54184 31332 54240 31334
rect 54288 31332 54344 31334
rect 54392 31332 54448 31388
rect 53768 29764 53824 29820
rect 53872 29818 53928 29820
rect 53976 29818 54032 29820
rect 53872 29766 53896 29818
rect 53896 29766 53928 29818
rect 53976 29766 54020 29818
rect 54020 29766 54032 29818
rect 53872 29764 53928 29766
rect 53976 29764 54032 29766
rect 54080 29764 54136 29820
rect 54184 29818 54240 29820
rect 54288 29818 54344 29820
rect 54184 29766 54196 29818
rect 54196 29766 54240 29818
rect 54288 29766 54320 29818
rect 54320 29766 54344 29818
rect 54184 29764 54240 29766
rect 54288 29764 54344 29766
rect 54392 29764 54448 29820
rect 53228 29484 53284 29540
rect 54236 29538 54292 29540
rect 54236 29486 54238 29538
rect 54238 29486 54290 29538
rect 54290 29486 54292 29538
rect 54236 29484 54292 29486
rect 55244 29484 55300 29540
rect 54908 29372 54964 29428
rect 53676 29202 53732 29204
rect 53676 29150 53678 29202
rect 53678 29150 53730 29202
rect 53730 29150 53732 29202
rect 53676 29148 53732 29150
rect 52892 27916 52948 27972
rect 52892 26348 52948 26404
rect 55020 28530 55076 28532
rect 55020 28478 55022 28530
rect 55022 28478 55074 28530
rect 55074 28478 55076 28530
rect 55020 28476 55076 28478
rect 53768 28196 53824 28252
rect 53872 28250 53928 28252
rect 53976 28250 54032 28252
rect 53872 28198 53896 28250
rect 53896 28198 53928 28250
rect 53976 28198 54020 28250
rect 54020 28198 54032 28250
rect 53872 28196 53928 28198
rect 53976 28196 54032 28198
rect 54080 28196 54136 28252
rect 54184 28250 54240 28252
rect 54288 28250 54344 28252
rect 54184 28198 54196 28250
rect 54196 28198 54240 28250
rect 54288 28198 54320 28250
rect 54320 28198 54344 28250
rect 54184 28196 54240 28198
rect 54288 28196 54344 28198
rect 54392 28196 54448 28252
rect 53676 27916 53732 27972
rect 56476 31554 56532 31556
rect 56476 31502 56478 31554
rect 56478 31502 56530 31554
rect 56530 31502 56532 31554
rect 56476 31500 56532 31502
rect 58268 30548 58324 30604
rect 58372 30602 58428 30604
rect 58476 30602 58532 30604
rect 58372 30550 58396 30602
rect 58396 30550 58428 30602
rect 58476 30550 58520 30602
rect 58520 30550 58532 30602
rect 58372 30548 58428 30550
rect 58476 30548 58532 30550
rect 58580 30548 58636 30604
rect 58684 30602 58740 30604
rect 58788 30602 58844 30604
rect 58684 30550 58696 30602
rect 58696 30550 58740 30602
rect 58788 30550 58820 30602
rect 58820 30550 58844 30602
rect 58684 30548 58740 30550
rect 58788 30548 58844 30550
rect 58892 30548 58948 30604
rect 59052 29986 59108 29988
rect 59052 29934 59054 29986
rect 59054 29934 59106 29986
rect 59106 29934 59108 29986
rect 59052 29932 59108 29934
rect 54572 27132 54628 27188
rect 53564 26796 53620 26852
rect 53768 26628 53824 26684
rect 53872 26682 53928 26684
rect 53976 26682 54032 26684
rect 53872 26630 53896 26682
rect 53896 26630 53928 26682
rect 53976 26630 54020 26682
rect 54020 26630 54032 26682
rect 53872 26628 53928 26630
rect 53976 26628 54032 26630
rect 54080 26628 54136 26684
rect 54184 26682 54240 26684
rect 54288 26682 54344 26684
rect 54184 26630 54196 26682
rect 54196 26630 54240 26682
rect 54288 26630 54320 26682
rect 54320 26630 54344 26682
rect 54184 26628 54240 26630
rect 54288 26628 54344 26630
rect 54392 26628 54448 26684
rect 53452 26348 53508 26404
rect 53788 26402 53844 26404
rect 53788 26350 53790 26402
rect 53790 26350 53842 26402
rect 53842 26350 53844 26402
rect 53788 26348 53844 26350
rect 56924 29538 56980 29540
rect 56924 29486 56926 29538
rect 56926 29486 56978 29538
rect 56978 29486 56980 29538
rect 56924 29484 56980 29486
rect 57596 29538 57652 29540
rect 57596 29486 57598 29538
rect 57598 29486 57650 29538
rect 57650 29486 57652 29538
rect 57596 29484 57652 29486
rect 56812 29426 56868 29428
rect 56812 29374 56814 29426
rect 56814 29374 56866 29426
rect 56866 29374 56868 29426
rect 56812 29372 56868 29374
rect 56924 28476 56980 28532
rect 58268 28980 58324 29036
rect 58372 29034 58428 29036
rect 58476 29034 58532 29036
rect 58372 28982 58396 29034
rect 58396 28982 58428 29034
rect 58476 28982 58520 29034
rect 58520 28982 58532 29034
rect 58372 28980 58428 28982
rect 58476 28980 58532 28982
rect 58580 28980 58636 29036
rect 58684 29034 58740 29036
rect 58788 29034 58844 29036
rect 58684 28982 58696 29034
rect 58696 28982 58740 29034
rect 58788 28982 58820 29034
rect 58820 28982 58844 29034
rect 58684 28980 58740 28982
rect 58788 28980 58844 28982
rect 58892 28980 58948 29036
rect 61628 34188 61684 34244
rect 61068 33516 61124 33572
rect 60844 33458 60900 33460
rect 60844 33406 60846 33458
rect 60846 33406 60898 33458
rect 60898 33406 60900 33458
rect 60844 33404 60900 33406
rect 61068 32732 61124 32788
rect 60284 32450 60340 32452
rect 60284 32398 60286 32450
rect 60286 32398 60338 32450
rect 60338 32398 60340 32450
rect 60284 32396 60340 32398
rect 62768 40740 62824 40796
rect 62872 40794 62928 40796
rect 62976 40794 63032 40796
rect 62872 40742 62896 40794
rect 62896 40742 62928 40794
rect 62976 40742 63020 40794
rect 63020 40742 63032 40794
rect 62872 40740 62928 40742
rect 62976 40740 63032 40742
rect 63080 40740 63136 40796
rect 63184 40794 63240 40796
rect 63288 40794 63344 40796
rect 63184 40742 63196 40794
rect 63196 40742 63240 40794
rect 63288 40742 63320 40794
rect 63320 40742 63344 40794
rect 63184 40740 63240 40742
rect 63288 40740 63344 40742
rect 63392 40740 63448 40796
rect 62768 39172 62824 39228
rect 62872 39226 62928 39228
rect 62976 39226 63032 39228
rect 62872 39174 62896 39226
rect 62896 39174 62928 39226
rect 62976 39174 63020 39226
rect 63020 39174 63032 39226
rect 62872 39172 62928 39174
rect 62976 39172 63032 39174
rect 63080 39172 63136 39228
rect 63184 39226 63240 39228
rect 63288 39226 63344 39228
rect 63184 39174 63196 39226
rect 63196 39174 63240 39226
rect 63288 39174 63320 39226
rect 63320 39174 63344 39226
rect 63184 39172 63240 39174
rect 63288 39172 63344 39174
rect 63392 39172 63448 39228
rect 63868 38332 63924 38388
rect 62768 37604 62824 37660
rect 62872 37658 62928 37660
rect 62976 37658 63032 37660
rect 62872 37606 62896 37658
rect 62896 37606 62928 37658
rect 62976 37606 63020 37658
rect 63020 37606 63032 37658
rect 62872 37604 62928 37606
rect 62976 37604 63032 37606
rect 63080 37604 63136 37660
rect 63184 37658 63240 37660
rect 63288 37658 63344 37660
rect 63184 37606 63196 37658
rect 63196 37606 63240 37658
rect 63288 37606 63320 37658
rect 63320 37606 63344 37658
rect 63184 37604 63240 37606
rect 63288 37604 63344 37606
rect 63392 37604 63448 37660
rect 64652 41186 64708 41188
rect 64652 41134 64654 41186
rect 64654 41134 64706 41186
rect 64706 41134 64708 41186
rect 64652 41132 64708 41134
rect 64652 39788 64708 39844
rect 64428 38332 64484 38388
rect 64540 38780 64596 38836
rect 63868 37100 63924 37156
rect 62768 36036 62824 36092
rect 62872 36090 62928 36092
rect 62976 36090 63032 36092
rect 62872 36038 62896 36090
rect 62896 36038 62928 36090
rect 62976 36038 63020 36090
rect 63020 36038 63032 36090
rect 62872 36036 62928 36038
rect 62976 36036 63032 36038
rect 63080 36036 63136 36092
rect 63184 36090 63240 36092
rect 63288 36090 63344 36092
rect 63184 36038 63196 36090
rect 63196 36038 63240 36090
rect 63288 36038 63320 36090
rect 63320 36038 63344 36090
rect 63184 36036 63240 36038
rect 63288 36036 63344 36038
rect 63392 36036 63448 36092
rect 64540 35644 64596 35700
rect 64988 46786 65044 46788
rect 64988 46734 64990 46786
rect 64990 46734 65042 46786
rect 65042 46734 65044 46786
rect 64988 46732 65044 46734
rect 64876 46620 64932 46676
rect 67268 47796 67324 47852
rect 67372 47850 67428 47852
rect 67476 47850 67532 47852
rect 67372 47798 67396 47850
rect 67396 47798 67428 47850
rect 67476 47798 67520 47850
rect 67520 47798 67532 47850
rect 67372 47796 67428 47798
rect 67476 47796 67532 47798
rect 67580 47796 67636 47852
rect 67684 47850 67740 47852
rect 67788 47850 67844 47852
rect 67684 47798 67696 47850
rect 67696 47798 67740 47850
rect 67788 47798 67820 47850
rect 67820 47798 67844 47850
rect 67684 47796 67740 47798
rect 67788 47796 67844 47798
rect 67892 47796 67948 47852
rect 65436 46786 65492 46788
rect 65436 46734 65438 46786
rect 65438 46734 65490 46786
rect 65490 46734 65492 46786
rect 65436 46732 65492 46734
rect 65772 46674 65828 46676
rect 65772 46622 65774 46674
rect 65774 46622 65826 46674
rect 65826 46622 65828 46674
rect 65772 46620 65828 46622
rect 65324 45836 65380 45892
rect 65212 44210 65268 44212
rect 65212 44158 65214 44210
rect 65214 44158 65266 44210
rect 65266 44158 65268 44210
rect 65212 44156 65268 44158
rect 64988 42812 65044 42868
rect 64988 42530 65044 42532
rect 64988 42478 64990 42530
rect 64990 42478 65042 42530
rect 65042 42478 65044 42530
rect 64988 42476 65044 42478
rect 65212 41132 65268 41188
rect 65884 44156 65940 44212
rect 65436 43538 65492 43540
rect 65436 43486 65438 43538
rect 65438 43486 65490 43538
rect 65490 43486 65492 43538
rect 65436 43484 65492 43486
rect 65548 43372 65604 43428
rect 66332 43372 66388 43428
rect 65660 42812 65716 42868
rect 66780 46450 66836 46452
rect 66780 46398 66782 46450
rect 66782 46398 66834 46450
rect 66834 46398 66836 46450
rect 66780 46396 66836 46398
rect 67268 46228 67324 46284
rect 67372 46282 67428 46284
rect 67476 46282 67532 46284
rect 67372 46230 67396 46282
rect 67396 46230 67428 46282
rect 67476 46230 67520 46282
rect 67520 46230 67532 46282
rect 67372 46228 67428 46230
rect 67476 46228 67532 46230
rect 67580 46228 67636 46284
rect 67684 46282 67740 46284
rect 67788 46282 67844 46284
rect 67684 46230 67696 46282
rect 67696 46230 67740 46282
rect 67788 46230 67820 46282
rect 67820 46230 67844 46282
rect 67684 46228 67740 46230
rect 67788 46228 67844 46230
rect 67892 46228 67948 46284
rect 67788 45388 67844 45444
rect 67268 44660 67324 44716
rect 67372 44714 67428 44716
rect 67476 44714 67532 44716
rect 67372 44662 67396 44714
rect 67396 44662 67428 44714
rect 67476 44662 67520 44714
rect 67520 44662 67532 44714
rect 67372 44660 67428 44662
rect 67476 44660 67532 44662
rect 67580 44660 67636 44716
rect 67684 44714 67740 44716
rect 67788 44714 67844 44716
rect 67684 44662 67696 44714
rect 67696 44662 67740 44714
rect 67788 44662 67820 44714
rect 67820 44662 67844 44714
rect 67684 44660 67740 44662
rect 67788 44660 67844 44662
rect 67892 44660 67948 44716
rect 67004 43538 67060 43540
rect 67004 43486 67006 43538
rect 67006 43486 67058 43538
rect 67058 43486 67060 43538
rect 67004 43484 67060 43486
rect 66668 42812 66724 42868
rect 66444 42700 66500 42756
rect 65324 39788 65380 39844
rect 64876 36594 64932 36596
rect 64876 36542 64878 36594
rect 64878 36542 64930 36594
rect 64930 36542 64932 36594
rect 64876 36540 64932 36542
rect 64316 34972 64372 35028
rect 62768 34468 62824 34524
rect 62872 34522 62928 34524
rect 62976 34522 63032 34524
rect 62872 34470 62896 34522
rect 62896 34470 62928 34522
rect 62976 34470 63020 34522
rect 63020 34470 63032 34522
rect 62872 34468 62928 34470
rect 62976 34468 63032 34470
rect 63080 34468 63136 34524
rect 63184 34522 63240 34524
rect 63288 34522 63344 34524
rect 63184 34470 63196 34522
rect 63196 34470 63240 34522
rect 63288 34470 63320 34522
rect 63320 34470 63344 34522
rect 63184 34468 63240 34470
rect 63288 34468 63344 34470
rect 63392 34468 63448 34524
rect 62972 34188 63028 34244
rect 62076 33404 62132 33460
rect 61852 33346 61908 33348
rect 61852 33294 61854 33346
rect 61854 33294 61906 33346
rect 61906 33294 61908 33346
rect 61852 33292 61908 33294
rect 62524 33516 62580 33572
rect 62412 33292 62468 33348
rect 61740 32562 61796 32564
rect 61740 32510 61742 32562
rect 61742 32510 61794 32562
rect 61794 32510 61796 32562
rect 61740 32508 61796 32510
rect 63644 33628 63700 33684
rect 63196 33068 63252 33124
rect 62768 32900 62824 32956
rect 62872 32954 62928 32956
rect 62976 32954 63032 32956
rect 62872 32902 62896 32954
rect 62896 32902 62928 32954
rect 62976 32902 63020 32954
rect 63020 32902 63032 32954
rect 62872 32900 62928 32902
rect 62976 32900 63032 32902
rect 63080 32900 63136 32956
rect 63184 32954 63240 32956
rect 63288 32954 63344 32956
rect 63184 32902 63196 32954
rect 63196 32902 63240 32954
rect 63288 32902 63320 32954
rect 63320 32902 63344 32954
rect 63184 32900 63240 32902
rect 63288 32900 63344 32902
rect 63392 32900 63448 32956
rect 63308 32674 63364 32676
rect 63308 32622 63310 32674
rect 63310 32622 63362 32674
rect 63362 32622 63364 32674
rect 63308 32620 63364 32622
rect 62972 32562 63028 32564
rect 62972 32510 62974 32562
rect 62974 32510 63026 32562
rect 63026 32510 63028 32562
rect 62972 32508 63028 32510
rect 63756 33068 63812 33124
rect 64652 34748 64708 34804
rect 65996 40908 66052 40964
rect 66108 40460 66164 40516
rect 65548 40402 65604 40404
rect 65548 40350 65550 40402
rect 65550 40350 65602 40402
rect 65602 40350 65604 40402
rect 65548 40348 65604 40350
rect 66556 40402 66612 40404
rect 66556 40350 66558 40402
rect 66558 40350 66610 40402
rect 66610 40350 66612 40402
rect 66556 40348 66612 40350
rect 65548 39004 65604 39060
rect 67268 43092 67324 43148
rect 67372 43146 67428 43148
rect 67476 43146 67532 43148
rect 67372 43094 67396 43146
rect 67396 43094 67428 43146
rect 67476 43094 67520 43146
rect 67520 43094 67532 43146
rect 67372 43092 67428 43094
rect 67476 43092 67532 43094
rect 67580 43092 67636 43148
rect 67684 43146 67740 43148
rect 67788 43146 67844 43148
rect 67684 43094 67696 43146
rect 67696 43094 67740 43146
rect 67788 43094 67820 43146
rect 67820 43094 67844 43146
rect 67684 43092 67740 43094
rect 67788 43092 67844 43094
rect 67892 43092 67948 43148
rect 70476 45612 70532 45668
rect 68908 45106 68964 45108
rect 68908 45054 68910 45106
rect 68910 45054 68962 45106
rect 68962 45054 68964 45106
rect 68908 45052 68964 45054
rect 70140 45106 70196 45108
rect 70140 45054 70142 45106
rect 70142 45054 70194 45106
rect 70194 45054 70196 45106
rect 70140 45052 70196 45054
rect 72156 49026 72212 49028
rect 72156 48974 72158 49026
rect 72158 48974 72210 49026
rect 72210 48974 72212 49026
rect 72156 48972 72212 48974
rect 72716 48972 72772 49028
rect 71820 48914 71876 48916
rect 71820 48862 71822 48914
rect 71822 48862 71874 48914
rect 71874 48862 71876 48914
rect 71820 48860 71876 48862
rect 71768 48580 71824 48636
rect 71872 48634 71928 48636
rect 71976 48634 72032 48636
rect 71872 48582 71896 48634
rect 71896 48582 71928 48634
rect 71976 48582 72020 48634
rect 72020 48582 72032 48634
rect 71872 48580 71928 48582
rect 71976 48580 72032 48582
rect 72080 48580 72136 48636
rect 72184 48634 72240 48636
rect 72288 48634 72344 48636
rect 72184 48582 72196 48634
rect 72196 48582 72240 48634
rect 72288 48582 72320 48634
rect 72320 48582 72344 48634
rect 72184 48580 72240 48582
rect 72288 48580 72344 48582
rect 72392 48580 72448 48636
rect 71708 48242 71764 48244
rect 71708 48190 71710 48242
rect 71710 48190 71762 48242
rect 71762 48190 71764 48242
rect 71708 48188 71764 48190
rect 72380 48242 72436 48244
rect 72380 48190 72382 48242
rect 72382 48190 72434 48242
rect 72434 48190 72436 48242
rect 72380 48188 72436 48190
rect 74284 50428 74340 50484
rect 74956 50428 75012 50484
rect 72940 48636 72996 48692
rect 73612 48300 73668 48356
rect 74060 48412 74116 48468
rect 74620 48412 74676 48468
rect 74172 48354 74228 48356
rect 74172 48302 74174 48354
rect 74174 48302 74226 48354
rect 74226 48302 74228 48354
rect 74172 48300 74228 48302
rect 73500 48188 73556 48244
rect 74396 48242 74452 48244
rect 74396 48190 74398 48242
rect 74398 48190 74450 48242
rect 74450 48190 74452 48242
rect 74396 48188 74452 48190
rect 72940 47964 72996 48020
rect 74060 47234 74116 47236
rect 74060 47182 74062 47234
rect 74062 47182 74114 47234
rect 74114 47182 74116 47234
rect 74060 47180 74116 47182
rect 71768 47012 71824 47068
rect 71872 47066 71928 47068
rect 71976 47066 72032 47068
rect 71872 47014 71896 47066
rect 71896 47014 71928 47066
rect 71976 47014 72020 47066
rect 72020 47014 72032 47066
rect 71872 47012 71928 47014
rect 71976 47012 72032 47014
rect 72080 47012 72136 47068
rect 72184 47066 72240 47068
rect 72288 47066 72344 47068
rect 72184 47014 72196 47066
rect 72196 47014 72240 47066
rect 72288 47014 72320 47066
rect 72320 47014 72344 47066
rect 72184 47012 72240 47014
rect 72288 47012 72344 47014
rect 72392 47012 72448 47068
rect 74620 48076 74676 48132
rect 80768 53284 80824 53340
rect 80872 53338 80928 53340
rect 80976 53338 81032 53340
rect 80872 53286 80896 53338
rect 80896 53286 80928 53338
rect 80976 53286 81020 53338
rect 81020 53286 81032 53338
rect 80872 53284 80928 53286
rect 80976 53284 81032 53286
rect 81080 53284 81136 53340
rect 81184 53338 81240 53340
rect 81288 53338 81344 53340
rect 81184 53286 81196 53338
rect 81196 53286 81240 53338
rect 81288 53286 81320 53338
rect 81320 53286 81344 53338
rect 81184 53284 81240 53286
rect 81288 53284 81344 53286
rect 81392 53284 81448 53340
rect 85268 54068 85324 54124
rect 85372 54122 85428 54124
rect 85476 54122 85532 54124
rect 85372 54070 85396 54122
rect 85396 54070 85428 54122
rect 85476 54070 85520 54122
rect 85520 54070 85532 54122
rect 85372 54068 85428 54070
rect 85476 54068 85532 54070
rect 85580 54068 85636 54124
rect 85684 54122 85740 54124
rect 85788 54122 85844 54124
rect 85684 54070 85696 54122
rect 85696 54070 85740 54122
rect 85788 54070 85820 54122
rect 85820 54070 85844 54122
rect 85684 54068 85740 54070
rect 85788 54068 85844 54070
rect 85892 54068 85948 54124
rect 94268 54068 94324 54124
rect 94372 54122 94428 54124
rect 94476 54122 94532 54124
rect 94372 54070 94396 54122
rect 94396 54070 94428 54122
rect 94476 54070 94520 54122
rect 94520 54070 94532 54122
rect 94372 54068 94428 54070
rect 94476 54068 94532 54070
rect 94580 54068 94636 54124
rect 94684 54122 94740 54124
rect 94788 54122 94844 54124
rect 94684 54070 94696 54122
rect 94696 54070 94740 54122
rect 94788 54070 94820 54122
rect 94820 54070 94844 54122
rect 94684 54068 94740 54070
rect 94788 54068 94844 54070
rect 94892 54068 94948 54124
rect 89768 53284 89824 53340
rect 89872 53338 89928 53340
rect 89976 53338 90032 53340
rect 89872 53286 89896 53338
rect 89896 53286 89928 53338
rect 89976 53286 90020 53338
rect 90020 53286 90032 53338
rect 89872 53284 89928 53286
rect 89976 53284 90032 53286
rect 90080 53284 90136 53340
rect 90184 53338 90240 53340
rect 90288 53338 90344 53340
rect 90184 53286 90196 53338
rect 90196 53286 90240 53338
rect 90288 53286 90320 53338
rect 90320 53286 90344 53338
rect 90184 53284 90240 53286
rect 90288 53284 90344 53286
rect 90392 53284 90448 53340
rect 81452 52780 81508 52836
rect 76268 52500 76324 52556
rect 76372 52554 76428 52556
rect 76476 52554 76532 52556
rect 76372 52502 76396 52554
rect 76396 52502 76428 52554
rect 76476 52502 76520 52554
rect 76520 52502 76532 52554
rect 76372 52500 76428 52502
rect 76476 52500 76532 52502
rect 76580 52500 76636 52556
rect 76684 52554 76740 52556
rect 76788 52554 76844 52556
rect 76684 52502 76696 52554
rect 76696 52502 76740 52554
rect 76788 52502 76820 52554
rect 76820 52502 76844 52554
rect 76684 52500 76740 52502
rect 76788 52500 76844 52502
rect 76892 52500 76948 52556
rect 85268 52500 85324 52556
rect 85372 52554 85428 52556
rect 85476 52554 85532 52556
rect 85372 52502 85396 52554
rect 85396 52502 85428 52554
rect 85476 52502 85520 52554
rect 85520 52502 85532 52554
rect 85372 52500 85428 52502
rect 85476 52500 85532 52502
rect 85580 52500 85636 52556
rect 85684 52554 85740 52556
rect 85788 52554 85844 52556
rect 85684 52502 85696 52554
rect 85696 52502 85740 52554
rect 85788 52502 85820 52554
rect 85820 52502 85844 52554
rect 85684 52500 85740 52502
rect 85788 52500 85844 52502
rect 85892 52500 85948 52556
rect 94268 52500 94324 52556
rect 94372 52554 94428 52556
rect 94476 52554 94532 52556
rect 94372 52502 94396 52554
rect 94396 52502 94428 52554
rect 94476 52502 94520 52554
rect 94520 52502 94532 52554
rect 94372 52500 94428 52502
rect 94476 52500 94532 52502
rect 94580 52500 94636 52556
rect 94684 52554 94740 52556
rect 94788 52554 94844 52556
rect 94684 52502 94696 52554
rect 94696 52502 94740 52554
rect 94788 52502 94820 52554
rect 94820 52502 94844 52554
rect 94684 52500 94740 52502
rect 94788 52500 94844 52502
rect 94892 52500 94948 52556
rect 80768 51716 80824 51772
rect 80872 51770 80928 51772
rect 80976 51770 81032 51772
rect 80872 51718 80896 51770
rect 80896 51718 80928 51770
rect 80976 51718 81020 51770
rect 81020 51718 81032 51770
rect 80872 51716 80928 51718
rect 80976 51716 81032 51718
rect 81080 51716 81136 51772
rect 81184 51770 81240 51772
rect 81288 51770 81344 51772
rect 81184 51718 81196 51770
rect 81196 51718 81240 51770
rect 81288 51718 81320 51770
rect 81320 51718 81344 51770
rect 81184 51716 81240 51718
rect 81288 51716 81344 51718
rect 81392 51716 81448 51772
rect 89768 51716 89824 51772
rect 89872 51770 89928 51772
rect 89976 51770 90032 51772
rect 89872 51718 89896 51770
rect 89896 51718 89928 51770
rect 89976 51718 90020 51770
rect 90020 51718 90032 51770
rect 89872 51716 89928 51718
rect 89976 51716 90032 51718
rect 90080 51716 90136 51772
rect 90184 51770 90240 51772
rect 90288 51770 90344 51772
rect 90184 51718 90196 51770
rect 90196 51718 90240 51770
rect 90288 51718 90320 51770
rect 90320 51718 90344 51770
rect 90184 51716 90240 51718
rect 90288 51716 90344 51718
rect 90392 51716 90448 51772
rect 90972 51602 91028 51604
rect 90972 51550 90974 51602
rect 90974 51550 91026 51602
rect 91026 51550 91028 51602
rect 90972 51548 91028 51550
rect 76636 51266 76692 51268
rect 76636 51214 76638 51266
rect 76638 51214 76690 51266
rect 76690 51214 76692 51266
rect 76636 51212 76692 51214
rect 76268 50932 76324 50988
rect 76372 50986 76428 50988
rect 76476 50986 76532 50988
rect 76372 50934 76396 50986
rect 76396 50934 76428 50986
rect 76476 50934 76520 50986
rect 76520 50934 76532 50986
rect 76372 50932 76428 50934
rect 76476 50932 76532 50934
rect 76580 50932 76636 50988
rect 76684 50986 76740 50988
rect 76788 50986 76844 50988
rect 76684 50934 76696 50986
rect 76696 50934 76740 50986
rect 76788 50934 76820 50986
rect 76820 50934 76844 50986
rect 76684 50932 76740 50934
rect 76788 50932 76844 50934
rect 76892 50932 76948 50988
rect 76524 50540 76580 50596
rect 79660 51212 79716 51268
rect 77308 50594 77364 50596
rect 77308 50542 77310 50594
rect 77310 50542 77362 50594
rect 77362 50542 77364 50594
rect 77308 50540 77364 50542
rect 77980 50428 78036 50484
rect 85268 50932 85324 50988
rect 85372 50986 85428 50988
rect 85476 50986 85532 50988
rect 85372 50934 85396 50986
rect 85396 50934 85428 50986
rect 85476 50934 85520 50986
rect 85520 50934 85532 50986
rect 85372 50932 85428 50934
rect 85476 50932 85532 50934
rect 85580 50932 85636 50988
rect 85684 50986 85740 50988
rect 85788 50986 85844 50988
rect 85684 50934 85696 50986
rect 85696 50934 85740 50986
rect 85788 50934 85820 50986
rect 85820 50934 85844 50986
rect 85684 50932 85740 50934
rect 85788 50932 85844 50934
rect 85892 50932 85948 50988
rect 80444 50482 80500 50484
rect 80444 50430 80446 50482
rect 80446 50430 80498 50482
rect 80498 50430 80500 50482
rect 80444 50428 80500 50430
rect 75740 49756 75796 49812
rect 77196 49810 77252 49812
rect 77196 49758 77198 49810
rect 77198 49758 77250 49810
rect 77250 49758 77252 49810
rect 77196 49756 77252 49758
rect 76188 49698 76244 49700
rect 76188 49646 76190 49698
rect 76190 49646 76242 49698
rect 76242 49646 76244 49698
rect 76188 49644 76244 49646
rect 77420 49644 77476 49700
rect 77644 49756 77700 49812
rect 76268 49364 76324 49420
rect 76372 49418 76428 49420
rect 76476 49418 76532 49420
rect 76372 49366 76396 49418
rect 76396 49366 76428 49418
rect 76476 49366 76520 49418
rect 76520 49366 76532 49418
rect 76372 49364 76428 49366
rect 76476 49364 76532 49366
rect 76580 49364 76636 49420
rect 76684 49418 76740 49420
rect 76788 49418 76844 49420
rect 76684 49366 76696 49418
rect 76696 49366 76740 49418
rect 76788 49366 76820 49418
rect 76820 49366 76844 49418
rect 76684 49364 76740 49366
rect 76788 49364 76844 49366
rect 76892 49364 76948 49420
rect 77644 49138 77700 49140
rect 77644 49086 77646 49138
rect 77646 49086 77698 49138
rect 77698 49086 77700 49138
rect 77644 49084 77700 49086
rect 77196 48354 77252 48356
rect 77196 48302 77198 48354
rect 77198 48302 77250 48354
rect 77250 48302 77252 48354
rect 77196 48300 77252 48302
rect 77980 49084 78036 49140
rect 76412 48242 76468 48244
rect 76412 48190 76414 48242
rect 76414 48190 76466 48242
rect 76466 48190 76468 48242
rect 76412 48188 76468 48190
rect 75964 48130 76020 48132
rect 75964 48078 75966 48130
rect 75966 48078 76018 48130
rect 76018 48078 76020 48130
rect 75964 48076 76020 48078
rect 75292 47628 75348 47684
rect 74956 47180 75012 47236
rect 73052 46620 73108 46676
rect 72940 45890 72996 45892
rect 72940 45838 72942 45890
rect 72942 45838 72994 45890
rect 72994 45838 72996 45890
rect 72940 45836 72996 45838
rect 73388 45724 73444 45780
rect 71932 45666 71988 45668
rect 71932 45614 71934 45666
rect 71934 45614 71986 45666
rect 71986 45614 71988 45666
rect 71932 45612 71988 45614
rect 73052 45666 73108 45668
rect 73052 45614 73054 45666
rect 73054 45614 73106 45666
rect 73106 45614 73108 45666
rect 73052 45612 73108 45614
rect 71372 45388 71428 45444
rect 71768 45444 71824 45500
rect 71872 45498 71928 45500
rect 71976 45498 72032 45500
rect 71872 45446 71896 45498
rect 71896 45446 71928 45498
rect 71976 45446 72020 45498
rect 72020 45446 72032 45498
rect 71872 45444 71928 45446
rect 71976 45444 72032 45446
rect 72080 45444 72136 45500
rect 72184 45498 72240 45500
rect 72288 45498 72344 45500
rect 72184 45446 72196 45498
rect 72196 45446 72240 45498
rect 72288 45446 72320 45498
rect 72320 45446 72344 45498
rect 72184 45444 72240 45446
rect 72288 45444 72344 45446
rect 72392 45444 72448 45500
rect 69468 44994 69524 44996
rect 69468 44942 69470 44994
rect 69470 44942 69522 44994
rect 69522 44942 69524 44994
rect 69468 44940 69524 44942
rect 69692 44322 69748 44324
rect 69692 44270 69694 44322
rect 69694 44270 69746 44322
rect 69746 44270 69748 44322
rect 69692 44268 69748 44270
rect 71260 45106 71316 45108
rect 71260 45054 71262 45106
rect 71262 45054 71314 45106
rect 71314 45054 71316 45106
rect 71260 45052 71316 45054
rect 73612 44994 73668 44996
rect 73612 44942 73614 44994
rect 73614 44942 73666 44994
rect 73666 44942 73668 44994
rect 73612 44940 73668 44942
rect 74508 46674 74564 46676
rect 74508 46622 74510 46674
rect 74510 46622 74562 46674
rect 74562 46622 74564 46674
rect 74508 46620 74564 46622
rect 74508 44940 74564 44996
rect 71260 44268 71316 44324
rect 73612 44322 73668 44324
rect 73612 44270 73614 44322
rect 73614 44270 73666 44322
rect 73666 44270 73668 44322
rect 73612 44268 73668 44270
rect 73052 44098 73108 44100
rect 73052 44046 73054 44098
rect 73054 44046 73106 44098
rect 73106 44046 73108 44098
rect 73052 44044 73108 44046
rect 73276 44044 73332 44100
rect 71768 43876 71824 43932
rect 71872 43930 71928 43932
rect 71976 43930 72032 43932
rect 71872 43878 71896 43930
rect 71896 43878 71928 43930
rect 71976 43878 72020 43930
rect 72020 43878 72032 43930
rect 71872 43876 71928 43878
rect 71976 43876 72032 43878
rect 72080 43876 72136 43932
rect 72184 43930 72240 43932
rect 72288 43930 72344 43932
rect 72184 43878 72196 43930
rect 72196 43878 72240 43930
rect 72288 43878 72320 43930
rect 72320 43878 72344 43930
rect 72184 43876 72240 43878
rect 72288 43876 72344 43878
rect 72392 43876 72448 43932
rect 67004 42140 67060 42196
rect 67004 41916 67060 41972
rect 67900 42700 67956 42756
rect 67788 41970 67844 41972
rect 67788 41918 67790 41970
rect 67790 41918 67842 41970
rect 67842 41918 67844 41970
rect 67788 41916 67844 41918
rect 67268 41524 67324 41580
rect 67372 41578 67428 41580
rect 67476 41578 67532 41580
rect 67372 41526 67396 41578
rect 67396 41526 67428 41578
rect 67476 41526 67520 41578
rect 67520 41526 67532 41578
rect 67372 41524 67428 41526
rect 67476 41524 67532 41526
rect 67580 41524 67636 41580
rect 67684 41578 67740 41580
rect 67788 41578 67844 41580
rect 67684 41526 67696 41578
rect 67696 41526 67740 41578
rect 67788 41526 67820 41578
rect 67820 41526 67844 41578
rect 67684 41524 67740 41526
rect 67788 41524 67844 41526
rect 67892 41524 67948 41580
rect 66892 40178 66948 40180
rect 66892 40126 66894 40178
rect 66894 40126 66946 40178
rect 66946 40126 66948 40178
rect 66892 40124 66948 40126
rect 67116 40908 67172 40964
rect 67452 40514 67508 40516
rect 67452 40462 67454 40514
rect 67454 40462 67506 40514
rect 67506 40462 67508 40514
rect 67452 40460 67508 40462
rect 67676 40124 67732 40180
rect 67268 39956 67324 40012
rect 67372 40010 67428 40012
rect 67476 40010 67532 40012
rect 67372 39958 67396 40010
rect 67396 39958 67428 40010
rect 67476 39958 67520 40010
rect 67520 39958 67532 40010
rect 67372 39956 67428 39958
rect 67476 39956 67532 39958
rect 67580 39956 67636 40012
rect 67684 40010 67740 40012
rect 67788 40010 67844 40012
rect 67684 39958 67696 40010
rect 67696 39958 67740 40010
rect 67788 39958 67820 40010
rect 67820 39958 67844 40010
rect 67684 39956 67740 39958
rect 67788 39956 67844 39958
rect 67892 39956 67948 40012
rect 70700 43538 70756 43540
rect 70700 43486 70702 43538
rect 70702 43486 70754 43538
rect 70754 43486 70756 43538
rect 70700 43484 70756 43486
rect 71708 43650 71764 43652
rect 71708 43598 71710 43650
rect 71710 43598 71762 43650
rect 71762 43598 71764 43650
rect 71708 43596 71764 43598
rect 73948 43932 74004 43988
rect 72492 43596 72548 43652
rect 72380 43538 72436 43540
rect 72380 43486 72382 43538
rect 72382 43486 72434 43538
rect 72434 43486 72436 43538
rect 72380 43484 72436 43486
rect 71260 43372 71316 43428
rect 69356 42530 69412 42532
rect 69356 42478 69358 42530
rect 69358 42478 69410 42530
rect 69410 42478 69412 42530
rect 69356 42476 69412 42478
rect 72492 42530 72548 42532
rect 72492 42478 72494 42530
rect 72494 42478 72546 42530
rect 72546 42478 72548 42530
rect 72492 42476 72548 42478
rect 71768 42308 71824 42364
rect 71872 42362 71928 42364
rect 71976 42362 72032 42364
rect 71872 42310 71896 42362
rect 71896 42310 71928 42362
rect 71976 42310 72020 42362
rect 72020 42310 72032 42362
rect 71872 42308 71928 42310
rect 71976 42308 72032 42310
rect 72080 42308 72136 42364
rect 72184 42362 72240 42364
rect 72288 42362 72344 42364
rect 72184 42310 72196 42362
rect 72196 42310 72240 42362
rect 72288 42310 72320 42362
rect 72320 42310 72344 42362
rect 72184 42308 72240 42310
rect 72288 42308 72344 42310
rect 72392 42308 72448 42364
rect 72268 41804 72324 41860
rect 72268 41244 72324 41300
rect 71372 41020 71428 41076
rect 68124 40572 68180 40628
rect 66892 39452 66948 39508
rect 66668 39058 66724 39060
rect 66668 39006 66670 39058
rect 66670 39006 66722 39058
rect 66722 39006 66724 39058
rect 66668 39004 66724 39006
rect 67004 38892 67060 38948
rect 66108 38332 66164 38388
rect 66444 37826 66500 37828
rect 66444 37774 66446 37826
rect 66446 37774 66498 37826
rect 66498 37774 66500 37826
rect 66444 37772 66500 37774
rect 66108 37660 66164 37716
rect 67228 38780 67284 38836
rect 68348 39788 68404 39844
rect 71768 40740 71824 40796
rect 71872 40794 71928 40796
rect 71976 40794 72032 40796
rect 71872 40742 71896 40794
rect 71896 40742 71928 40794
rect 71976 40742 72020 40794
rect 72020 40742 72032 40794
rect 71872 40740 71928 40742
rect 71976 40740 72032 40742
rect 72080 40740 72136 40796
rect 72184 40794 72240 40796
rect 72288 40794 72344 40796
rect 72184 40742 72196 40794
rect 72196 40742 72240 40794
rect 72288 40742 72320 40794
rect 72320 40742 72344 40794
rect 72184 40740 72240 40742
rect 72288 40740 72344 40742
rect 72392 40740 72448 40796
rect 71596 40572 71652 40628
rect 73164 43596 73220 43652
rect 72716 43426 72772 43428
rect 72716 43374 72718 43426
rect 72718 43374 72770 43426
rect 72770 43374 72772 43426
rect 72716 43372 72772 43374
rect 74508 42476 74564 42532
rect 74620 44268 74676 44324
rect 75068 44322 75124 44324
rect 75068 44270 75070 44322
rect 75070 44270 75122 44322
rect 75122 44270 75124 44322
rect 75068 44268 75124 44270
rect 74956 43932 75012 43988
rect 74620 42140 74676 42196
rect 72268 40626 72324 40628
rect 72268 40574 72270 40626
rect 72270 40574 72322 40626
rect 72322 40574 72324 40626
rect 72268 40572 72324 40574
rect 73500 41804 73556 41860
rect 71708 40402 71764 40404
rect 71708 40350 71710 40402
rect 71710 40350 71762 40402
rect 71762 40350 71764 40402
rect 71708 40348 71764 40350
rect 69692 40178 69748 40180
rect 69692 40126 69694 40178
rect 69694 40126 69746 40178
rect 69746 40126 69748 40178
rect 69692 40124 69748 40126
rect 68460 39506 68516 39508
rect 68460 39454 68462 39506
rect 68462 39454 68514 39506
rect 68514 39454 68516 39506
rect 68460 39452 68516 39454
rect 67788 39004 67844 39060
rect 68012 38946 68068 38948
rect 68012 38894 68014 38946
rect 68014 38894 68066 38946
rect 68066 38894 68068 38946
rect 68012 38892 68068 38894
rect 67268 38388 67324 38444
rect 67372 38442 67428 38444
rect 67476 38442 67532 38444
rect 67372 38390 67396 38442
rect 67396 38390 67428 38442
rect 67476 38390 67520 38442
rect 67520 38390 67532 38442
rect 67372 38388 67428 38390
rect 67476 38388 67532 38390
rect 67580 38388 67636 38444
rect 67684 38442 67740 38444
rect 67788 38442 67844 38444
rect 67684 38390 67696 38442
rect 67696 38390 67740 38442
rect 67788 38390 67820 38442
rect 67820 38390 67844 38442
rect 67684 38388 67740 38390
rect 67788 38388 67844 38390
rect 67892 38388 67948 38444
rect 67788 38220 67844 38276
rect 67116 37772 67172 37828
rect 67228 37996 67284 38052
rect 66892 36988 66948 37044
rect 67676 37772 67732 37828
rect 68572 38220 68628 38276
rect 69020 39788 69076 39844
rect 74172 41020 74228 41076
rect 73948 40402 74004 40404
rect 73948 40350 73950 40402
rect 73950 40350 74002 40402
rect 74002 40350 74004 40402
rect 73948 40348 74004 40350
rect 71768 39172 71824 39228
rect 71872 39226 71928 39228
rect 71976 39226 72032 39228
rect 71872 39174 71896 39226
rect 71896 39174 71928 39226
rect 71976 39174 72020 39226
rect 72020 39174 72032 39226
rect 71872 39172 71928 39174
rect 71976 39172 72032 39174
rect 72080 39172 72136 39228
rect 72184 39226 72240 39228
rect 72288 39226 72344 39228
rect 72184 39174 72196 39226
rect 72196 39174 72240 39226
rect 72288 39174 72320 39226
rect 72320 39174 72344 39226
rect 72184 39172 72240 39174
rect 72288 39172 72344 39174
rect 72392 39172 72448 39228
rect 75852 45836 75908 45892
rect 75404 44268 75460 44324
rect 75292 43314 75348 43316
rect 75292 43262 75294 43314
rect 75294 43262 75346 43314
rect 75346 43262 75348 43314
rect 75292 43260 75348 43262
rect 74732 41074 74788 41076
rect 74732 41022 74734 41074
rect 74734 41022 74786 41074
rect 74786 41022 74788 41074
rect 74732 41020 74788 41022
rect 74172 40236 74228 40292
rect 69020 38834 69076 38836
rect 69020 38782 69022 38834
rect 69022 38782 69074 38834
rect 69074 38782 69076 38834
rect 69020 38780 69076 38782
rect 68572 38050 68628 38052
rect 68572 37998 68574 38050
rect 68574 37998 68626 38050
rect 68626 37998 68628 38050
rect 68572 37996 68628 37998
rect 68348 37938 68404 37940
rect 68348 37886 68350 37938
rect 68350 37886 68402 37938
rect 68402 37886 68404 37938
rect 68348 37884 68404 37886
rect 74844 38834 74900 38836
rect 74844 38782 74846 38834
rect 74846 38782 74898 38834
rect 74898 38782 74900 38834
rect 74844 38780 74900 38782
rect 72380 37884 72436 37940
rect 68236 37548 68292 37604
rect 67228 36988 67284 37044
rect 68684 36988 68740 37044
rect 67268 36820 67324 36876
rect 67372 36874 67428 36876
rect 67476 36874 67532 36876
rect 67372 36822 67396 36874
rect 67396 36822 67428 36874
rect 67476 36822 67520 36874
rect 67520 36822 67532 36874
rect 67372 36820 67428 36822
rect 67476 36820 67532 36822
rect 67580 36820 67636 36876
rect 67684 36874 67740 36876
rect 67788 36874 67844 36876
rect 67684 36822 67696 36874
rect 67696 36822 67740 36874
rect 67788 36822 67820 36874
rect 67820 36822 67844 36874
rect 67684 36820 67740 36822
rect 67788 36820 67844 36822
rect 67892 36820 67948 36876
rect 65548 36540 65604 36596
rect 67452 36594 67508 36596
rect 67452 36542 67454 36594
rect 67454 36542 67506 36594
rect 67506 36542 67508 36594
rect 67452 36540 67508 36542
rect 65436 36316 65492 36372
rect 71932 37826 71988 37828
rect 71932 37774 71934 37826
rect 71934 37774 71986 37826
rect 71986 37774 71988 37826
rect 71932 37772 71988 37774
rect 72604 37772 72660 37828
rect 68908 37548 68964 37604
rect 71768 37604 71824 37660
rect 71872 37658 71928 37660
rect 71976 37658 72032 37660
rect 71872 37606 71896 37658
rect 71896 37606 71928 37658
rect 71976 37606 72020 37658
rect 72020 37606 72032 37658
rect 71872 37604 71928 37606
rect 71976 37604 72032 37606
rect 72080 37604 72136 37660
rect 72184 37658 72240 37660
rect 72288 37658 72344 37660
rect 72184 37606 72196 37658
rect 72196 37606 72240 37658
rect 72288 37606 72320 37658
rect 72320 37606 72344 37658
rect 72184 37604 72240 37606
rect 72288 37604 72344 37606
rect 72392 37604 72448 37660
rect 68796 36764 68852 36820
rect 69468 36876 69524 36932
rect 68796 36594 68852 36596
rect 68796 36542 68798 36594
rect 68798 36542 68850 36594
rect 68850 36542 68852 36594
rect 68796 36540 68852 36542
rect 67788 36370 67844 36372
rect 67788 36318 67790 36370
rect 67790 36318 67842 36370
rect 67842 36318 67844 36370
rect 67788 36316 67844 36318
rect 67268 35252 67324 35308
rect 67372 35306 67428 35308
rect 67476 35306 67532 35308
rect 67372 35254 67396 35306
rect 67396 35254 67428 35306
rect 67476 35254 67520 35306
rect 67520 35254 67532 35306
rect 67372 35252 67428 35254
rect 67476 35252 67532 35254
rect 67580 35252 67636 35308
rect 67684 35306 67740 35308
rect 67788 35306 67844 35308
rect 67684 35254 67696 35306
rect 67696 35254 67740 35306
rect 67788 35254 67820 35306
rect 67820 35254 67844 35306
rect 67684 35252 67740 35254
rect 67788 35252 67844 35254
rect 67892 35252 67948 35308
rect 67004 34636 67060 34692
rect 64652 33628 64708 33684
rect 64540 32508 64596 32564
rect 62524 31948 62580 32004
rect 64092 32002 64148 32004
rect 64092 31950 64094 32002
rect 64094 31950 64146 32002
rect 64146 31950 64148 32002
rect 64092 31948 64148 31950
rect 63532 31836 63588 31892
rect 64428 31890 64484 31892
rect 64428 31838 64430 31890
rect 64430 31838 64482 31890
rect 64482 31838 64484 31890
rect 64428 31836 64484 31838
rect 64652 31500 64708 31556
rect 62768 31332 62824 31388
rect 62872 31386 62928 31388
rect 62976 31386 63032 31388
rect 62872 31334 62896 31386
rect 62896 31334 62928 31386
rect 62976 31334 63020 31386
rect 63020 31334 63032 31386
rect 62872 31332 62928 31334
rect 62976 31332 63032 31334
rect 63080 31332 63136 31388
rect 63184 31386 63240 31388
rect 63288 31386 63344 31388
rect 63184 31334 63196 31386
rect 63196 31334 63240 31386
rect 63288 31334 63320 31386
rect 63320 31334 63344 31386
rect 63184 31332 63240 31334
rect 63288 31332 63344 31334
rect 63392 31332 63448 31388
rect 61628 29932 61684 29988
rect 60732 28812 60788 28868
rect 60732 28588 60788 28644
rect 61292 28588 61348 28644
rect 57260 27916 57316 27972
rect 57932 27692 57988 27748
rect 56924 27020 56980 27076
rect 57036 26850 57092 26852
rect 57036 26798 57038 26850
rect 57038 26798 57090 26850
rect 57090 26798 57092 26850
rect 57036 26796 57092 26798
rect 56028 26684 56084 26740
rect 57820 27074 57876 27076
rect 57820 27022 57822 27074
rect 57822 27022 57874 27074
rect 57874 27022 57876 27074
rect 57820 27020 57876 27022
rect 62768 29764 62824 29820
rect 62872 29818 62928 29820
rect 62976 29818 63032 29820
rect 62872 29766 62896 29818
rect 62896 29766 62928 29818
rect 62976 29766 63020 29818
rect 63020 29766 63032 29818
rect 62872 29764 62928 29766
rect 62976 29764 63032 29766
rect 63080 29764 63136 29820
rect 63184 29818 63240 29820
rect 63288 29818 63344 29820
rect 63184 29766 63196 29818
rect 63196 29766 63240 29818
rect 63288 29766 63320 29818
rect 63320 29766 63344 29818
rect 63184 29764 63240 29766
rect 63288 29764 63344 29766
rect 63392 29764 63448 29820
rect 61628 29596 61684 29652
rect 64652 29484 64708 29540
rect 61740 28866 61796 28868
rect 61740 28814 61742 28866
rect 61742 28814 61794 28866
rect 61794 28814 61796 28866
rect 61740 28812 61796 28814
rect 61180 28530 61236 28532
rect 61180 28478 61182 28530
rect 61182 28478 61234 28530
rect 61234 28478 61236 28530
rect 61180 28476 61236 28478
rect 62972 28588 63028 28644
rect 61068 28364 61124 28420
rect 58268 27412 58324 27468
rect 58372 27466 58428 27468
rect 58476 27466 58532 27468
rect 58372 27414 58396 27466
rect 58396 27414 58428 27466
rect 58476 27414 58520 27466
rect 58520 27414 58532 27466
rect 58372 27412 58428 27414
rect 58476 27412 58532 27414
rect 58580 27412 58636 27468
rect 58684 27466 58740 27468
rect 58788 27466 58844 27468
rect 58684 27414 58696 27466
rect 58696 27414 58740 27466
rect 58788 27414 58820 27466
rect 58820 27414 58844 27466
rect 58684 27412 58740 27414
rect 58788 27412 58844 27414
rect 58892 27412 58948 27468
rect 58044 26684 58100 26740
rect 57036 26290 57092 26292
rect 57036 26238 57038 26290
rect 57038 26238 57090 26290
rect 57090 26238 57092 26290
rect 57036 26236 57092 26238
rect 54572 25506 54628 25508
rect 54572 25454 54574 25506
rect 54574 25454 54626 25506
rect 54626 25454 54628 25506
rect 54572 25452 54628 25454
rect 53768 25060 53824 25116
rect 53872 25114 53928 25116
rect 53976 25114 54032 25116
rect 53872 25062 53896 25114
rect 53896 25062 53928 25114
rect 53976 25062 54020 25114
rect 54020 25062 54032 25114
rect 53872 25060 53928 25062
rect 53976 25060 54032 25062
rect 54080 25060 54136 25116
rect 54184 25114 54240 25116
rect 54288 25114 54344 25116
rect 54184 25062 54196 25114
rect 54196 25062 54240 25114
rect 54288 25062 54320 25114
rect 54320 25062 54344 25114
rect 54184 25060 54240 25062
rect 54288 25060 54344 25062
rect 54392 25060 54448 25116
rect 53768 23492 53824 23548
rect 53872 23546 53928 23548
rect 53976 23546 54032 23548
rect 53872 23494 53896 23546
rect 53896 23494 53928 23546
rect 53976 23494 54020 23546
rect 54020 23494 54032 23546
rect 53872 23492 53928 23494
rect 53976 23492 54032 23494
rect 54080 23492 54136 23548
rect 54184 23546 54240 23548
rect 54288 23546 54344 23548
rect 54184 23494 54196 23546
rect 54196 23494 54240 23546
rect 54288 23494 54320 23546
rect 54320 23494 54344 23546
rect 54184 23492 54240 23494
rect 54288 23492 54344 23494
rect 54392 23492 54448 23548
rect 53768 21924 53824 21980
rect 53872 21978 53928 21980
rect 53976 21978 54032 21980
rect 53872 21926 53896 21978
rect 53896 21926 53928 21978
rect 53976 21926 54020 21978
rect 54020 21926 54032 21978
rect 53872 21924 53928 21926
rect 53976 21924 54032 21926
rect 54080 21924 54136 21980
rect 54184 21978 54240 21980
rect 54288 21978 54344 21980
rect 54184 21926 54196 21978
rect 54196 21926 54240 21978
rect 54288 21926 54320 21978
rect 54320 21926 54344 21978
rect 54184 21924 54240 21926
rect 54288 21924 54344 21926
rect 54392 21924 54448 21980
rect 56028 20972 56084 21028
rect 55468 20914 55524 20916
rect 55468 20862 55470 20914
rect 55470 20862 55522 20914
rect 55522 20862 55524 20914
rect 55468 20860 55524 20862
rect 57932 26290 57988 26292
rect 57932 26238 57934 26290
rect 57934 26238 57986 26290
rect 57986 26238 57988 26290
rect 57932 26236 57988 26238
rect 57148 25564 57204 25620
rect 60172 27970 60228 27972
rect 60172 27918 60174 27970
rect 60174 27918 60226 27970
rect 60226 27918 60228 27970
rect 60172 27916 60228 27918
rect 59948 27244 60004 27300
rect 60620 27244 60676 27300
rect 60508 26962 60564 26964
rect 60508 26910 60510 26962
rect 60510 26910 60562 26962
rect 60562 26910 60564 26962
rect 60508 26908 60564 26910
rect 59612 26684 59668 26740
rect 59948 26796 60004 26852
rect 59612 26514 59668 26516
rect 59612 26462 59614 26514
rect 59614 26462 59666 26514
rect 59666 26462 59668 26514
rect 59612 26460 59668 26462
rect 58492 26402 58548 26404
rect 58492 26350 58494 26402
rect 58494 26350 58546 26402
rect 58546 26350 58548 26402
rect 58492 26348 58548 26350
rect 60060 26514 60116 26516
rect 60060 26462 60062 26514
rect 60062 26462 60114 26514
rect 60114 26462 60116 26514
rect 60060 26460 60116 26462
rect 59948 26402 60004 26404
rect 59948 26350 59950 26402
rect 59950 26350 60002 26402
rect 60002 26350 60004 26402
rect 59948 26348 60004 26350
rect 60060 26066 60116 26068
rect 60060 26014 60062 26066
rect 60062 26014 60114 26066
rect 60114 26014 60116 26066
rect 60060 26012 60116 26014
rect 58268 25844 58324 25900
rect 58372 25898 58428 25900
rect 58476 25898 58532 25900
rect 58372 25846 58396 25898
rect 58396 25846 58428 25898
rect 58476 25846 58520 25898
rect 58520 25846 58532 25898
rect 58372 25844 58428 25846
rect 58476 25844 58532 25846
rect 58580 25844 58636 25900
rect 58684 25898 58740 25900
rect 58788 25898 58844 25900
rect 58684 25846 58696 25898
rect 58696 25846 58740 25898
rect 58788 25846 58820 25898
rect 58820 25846 58844 25898
rect 58684 25844 58740 25846
rect 58788 25844 58844 25846
rect 58892 25844 58948 25900
rect 58044 25618 58100 25620
rect 58044 25566 58046 25618
rect 58046 25566 58098 25618
rect 58098 25566 58100 25618
rect 58044 25564 58100 25566
rect 60172 24946 60228 24948
rect 60172 24894 60174 24946
rect 60174 24894 60226 24946
rect 60226 24894 60228 24946
rect 60172 24892 60228 24894
rect 60844 27074 60900 27076
rect 60844 27022 60846 27074
rect 60846 27022 60898 27074
rect 60898 27022 60900 27074
rect 60844 27020 60900 27022
rect 63196 28642 63252 28644
rect 63196 28590 63198 28642
rect 63198 28590 63250 28642
rect 63250 28590 63252 28642
rect 63196 28588 63252 28590
rect 63532 28588 63588 28644
rect 61628 28364 61684 28420
rect 61068 26796 61124 26852
rect 61180 28028 61236 28084
rect 60620 24946 60676 24948
rect 60620 24894 60622 24946
rect 60622 24894 60674 24946
rect 60674 24894 60676 24946
rect 60620 24892 60676 24894
rect 59388 24668 59444 24724
rect 58268 24276 58324 24332
rect 58372 24330 58428 24332
rect 58476 24330 58532 24332
rect 58372 24278 58396 24330
rect 58396 24278 58428 24330
rect 58476 24278 58520 24330
rect 58520 24278 58532 24330
rect 58372 24276 58428 24278
rect 58476 24276 58532 24278
rect 58580 24276 58636 24332
rect 58684 24330 58740 24332
rect 58788 24330 58844 24332
rect 58684 24278 58696 24330
rect 58696 24278 58740 24330
rect 58788 24278 58820 24330
rect 58820 24278 58844 24330
rect 58684 24276 58740 24278
rect 58788 24276 58844 24278
rect 58892 24276 58948 24332
rect 59724 23826 59780 23828
rect 59724 23774 59726 23826
rect 59726 23774 59778 23826
rect 59778 23774 59780 23826
rect 59724 23772 59780 23774
rect 60620 24498 60676 24500
rect 60620 24446 60622 24498
rect 60622 24446 60674 24498
rect 60674 24446 60676 24498
rect 60620 24444 60676 24446
rect 61180 23996 61236 24052
rect 60508 23772 60564 23828
rect 61068 23826 61124 23828
rect 61068 23774 61070 23826
rect 61070 23774 61122 23826
rect 61122 23774 61124 23826
rect 61068 23772 61124 23774
rect 58268 22708 58324 22764
rect 58372 22762 58428 22764
rect 58476 22762 58532 22764
rect 58372 22710 58396 22762
rect 58396 22710 58428 22762
rect 58476 22710 58520 22762
rect 58520 22710 58532 22762
rect 58372 22708 58428 22710
rect 58476 22708 58532 22710
rect 58580 22708 58636 22764
rect 58684 22762 58740 22764
rect 58788 22762 58844 22764
rect 58684 22710 58696 22762
rect 58696 22710 58740 22762
rect 58788 22710 58820 22762
rect 58820 22710 58844 22762
rect 58684 22708 58740 22710
rect 58788 22708 58844 22710
rect 58892 22708 58948 22764
rect 60284 23660 60340 23716
rect 60732 23324 60788 23380
rect 60060 22316 60116 22372
rect 58268 21140 58324 21196
rect 58372 21194 58428 21196
rect 58476 21194 58532 21196
rect 58372 21142 58396 21194
rect 58396 21142 58428 21194
rect 58476 21142 58520 21194
rect 58520 21142 58532 21194
rect 58372 21140 58428 21142
rect 58476 21140 58532 21142
rect 58580 21140 58636 21196
rect 58684 21194 58740 21196
rect 58788 21194 58844 21196
rect 58684 21142 58696 21194
rect 58696 21142 58740 21194
rect 58788 21142 58820 21194
rect 58820 21142 58844 21194
rect 58684 21140 58740 21142
rect 58788 21140 58844 21142
rect 58892 21140 58948 21196
rect 56700 20972 56756 21028
rect 56028 20802 56084 20804
rect 56028 20750 56030 20802
rect 56030 20750 56082 20802
rect 56082 20750 56084 20802
rect 56028 20748 56084 20750
rect 56140 20860 56196 20916
rect 56364 20802 56420 20804
rect 56364 20750 56366 20802
rect 56366 20750 56418 20802
rect 56418 20750 56420 20802
rect 56364 20748 56420 20750
rect 53768 20356 53824 20412
rect 53872 20410 53928 20412
rect 53976 20410 54032 20412
rect 53872 20358 53896 20410
rect 53896 20358 53928 20410
rect 53976 20358 54020 20410
rect 54020 20358 54032 20410
rect 53872 20356 53928 20358
rect 53976 20356 54032 20358
rect 54080 20356 54136 20412
rect 54184 20410 54240 20412
rect 54288 20410 54344 20412
rect 54184 20358 54196 20410
rect 54196 20358 54240 20410
rect 54288 20358 54320 20410
rect 54320 20358 54344 20410
rect 54184 20356 54240 20358
rect 54288 20356 54344 20358
rect 54392 20356 54448 20412
rect 58268 19572 58324 19628
rect 58372 19626 58428 19628
rect 58476 19626 58532 19628
rect 58372 19574 58396 19626
rect 58396 19574 58428 19626
rect 58476 19574 58520 19626
rect 58520 19574 58532 19626
rect 58372 19572 58428 19574
rect 58476 19572 58532 19574
rect 58580 19572 58636 19628
rect 58684 19626 58740 19628
rect 58788 19626 58844 19628
rect 58684 19574 58696 19626
rect 58696 19574 58740 19626
rect 58788 19574 58820 19626
rect 58820 19574 58844 19626
rect 58684 19572 58740 19574
rect 58788 19572 58844 19574
rect 58892 19572 58948 19628
rect 53768 18788 53824 18844
rect 53872 18842 53928 18844
rect 53976 18842 54032 18844
rect 53872 18790 53896 18842
rect 53896 18790 53928 18842
rect 53976 18790 54020 18842
rect 54020 18790 54032 18842
rect 53872 18788 53928 18790
rect 53976 18788 54032 18790
rect 54080 18788 54136 18844
rect 54184 18842 54240 18844
rect 54288 18842 54344 18844
rect 54184 18790 54196 18842
rect 54196 18790 54240 18842
rect 54288 18790 54320 18842
rect 54320 18790 54344 18842
rect 54184 18788 54240 18790
rect 54288 18788 54344 18790
rect 54392 18788 54448 18844
rect 58268 18004 58324 18060
rect 58372 18058 58428 18060
rect 58476 18058 58532 18060
rect 58372 18006 58396 18058
rect 58396 18006 58428 18058
rect 58476 18006 58520 18058
rect 58520 18006 58532 18058
rect 58372 18004 58428 18006
rect 58476 18004 58532 18006
rect 58580 18004 58636 18060
rect 58684 18058 58740 18060
rect 58788 18058 58844 18060
rect 58684 18006 58696 18058
rect 58696 18006 58740 18058
rect 58788 18006 58820 18058
rect 58820 18006 58844 18058
rect 58684 18004 58740 18006
rect 58788 18004 58844 18006
rect 58892 18004 58948 18060
rect 53768 17220 53824 17276
rect 53872 17274 53928 17276
rect 53976 17274 54032 17276
rect 53872 17222 53896 17274
rect 53896 17222 53928 17274
rect 53976 17222 54020 17274
rect 54020 17222 54032 17274
rect 53872 17220 53928 17222
rect 53976 17220 54032 17222
rect 54080 17220 54136 17276
rect 54184 17274 54240 17276
rect 54288 17274 54344 17276
rect 54184 17222 54196 17274
rect 54196 17222 54240 17274
rect 54288 17222 54320 17274
rect 54320 17222 54344 17274
rect 54184 17220 54240 17222
rect 54288 17220 54344 17222
rect 54392 17220 54448 17276
rect 58268 16436 58324 16492
rect 58372 16490 58428 16492
rect 58476 16490 58532 16492
rect 58372 16438 58396 16490
rect 58396 16438 58428 16490
rect 58476 16438 58520 16490
rect 58520 16438 58532 16490
rect 58372 16436 58428 16438
rect 58476 16436 58532 16438
rect 58580 16436 58636 16492
rect 58684 16490 58740 16492
rect 58788 16490 58844 16492
rect 58684 16438 58696 16490
rect 58696 16438 58740 16490
rect 58788 16438 58820 16490
rect 58820 16438 58844 16490
rect 58684 16436 58740 16438
rect 58788 16436 58844 16438
rect 58892 16436 58948 16492
rect 53768 15652 53824 15708
rect 53872 15706 53928 15708
rect 53976 15706 54032 15708
rect 53872 15654 53896 15706
rect 53896 15654 53928 15706
rect 53976 15654 54020 15706
rect 54020 15654 54032 15706
rect 53872 15652 53928 15654
rect 53976 15652 54032 15654
rect 54080 15652 54136 15708
rect 54184 15706 54240 15708
rect 54288 15706 54344 15708
rect 54184 15654 54196 15706
rect 54196 15654 54240 15706
rect 54288 15654 54320 15706
rect 54320 15654 54344 15706
rect 54184 15652 54240 15654
rect 54288 15652 54344 15654
rect 54392 15652 54448 15708
rect 52444 13804 52500 13860
rect 58268 14868 58324 14924
rect 58372 14922 58428 14924
rect 58476 14922 58532 14924
rect 58372 14870 58396 14922
rect 58396 14870 58428 14922
rect 58476 14870 58520 14922
rect 58520 14870 58532 14922
rect 58372 14868 58428 14870
rect 58476 14868 58532 14870
rect 58580 14868 58636 14924
rect 58684 14922 58740 14924
rect 58788 14922 58844 14924
rect 58684 14870 58696 14922
rect 58696 14870 58740 14922
rect 58788 14870 58820 14922
rect 58820 14870 58844 14922
rect 58684 14868 58740 14870
rect 58788 14868 58844 14870
rect 58892 14868 58948 14924
rect 53768 14084 53824 14140
rect 53872 14138 53928 14140
rect 53976 14138 54032 14140
rect 53872 14086 53896 14138
rect 53896 14086 53928 14138
rect 53976 14086 54020 14138
rect 54020 14086 54032 14138
rect 53872 14084 53928 14086
rect 53976 14084 54032 14086
rect 54080 14084 54136 14140
rect 54184 14138 54240 14140
rect 54288 14138 54344 14140
rect 54184 14086 54196 14138
rect 54196 14086 54240 14138
rect 54288 14086 54320 14138
rect 54320 14086 54344 14138
rect 54184 14084 54240 14086
rect 54288 14084 54344 14086
rect 54392 14084 54448 14140
rect 53004 13916 53060 13972
rect 49268 13300 49324 13356
rect 49372 13354 49428 13356
rect 49476 13354 49532 13356
rect 49372 13302 49396 13354
rect 49396 13302 49428 13354
rect 49476 13302 49520 13354
rect 49520 13302 49532 13354
rect 49372 13300 49428 13302
rect 49476 13300 49532 13302
rect 49580 13300 49636 13356
rect 49684 13354 49740 13356
rect 49788 13354 49844 13356
rect 49684 13302 49696 13354
rect 49696 13302 49740 13354
rect 49788 13302 49820 13354
rect 49820 13302 49844 13354
rect 49684 13300 49740 13302
rect 49788 13300 49844 13302
rect 49892 13300 49948 13356
rect 49532 12850 49588 12852
rect 49532 12798 49534 12850
rect 49534 12798 49586 12850
rect 49586 12798 49588 12850
rect 49532 12796 49588 12798
rect 49268 11732 49324 11788
rect 49372 11786 49428 11788
rect 49476 11786 49532 11788
rect 49372 11734 49396 11786
rect 49396 11734 49428 11786
rect 49476 11734 49520 11786
rect 49520 11734 49532 11786
rect 49372 11732 49428 11734
rect 49476 11732 49532 11734
rect 49580 11732 49636 11788
rect 49684 11786 49740 11788
rect 49788 11786 49844 11788
rect 49684 11734 49696 11786
rect 49696 11734 49740 11786
rect 49788 11734 49820 11786
rect 49820 11734 49844 11786
rect 49684 11732 49740 11734
rect 49788 11732 49844 11734
rect 49892 11732 49948 11788
rect 49268 10164 49324 10220
rect 49372 10218 49428 10220
rect 49476 10218 49532 10220
rect 49372 10166 49396 10218
rect 49396 10166 49428 10218
rect 49476 10166 49520 10218
rect 49520 10166 49532 10218
rect 49372 10164 49428 10166
rect 49476 10164 49532 10166
rect 49580 10164 49636 10220
rect 49684 10218 49740 10220
rect 49788 10218 49844 10220
rect 49684 10166 49696 10218
rect 49696 10166 49740 10218
rect 49788 10166 49820 10218
rect 49820 10166 49844 10218
rect 49684 10164 49740 10166
rect 49788 10164 49844 10166
rect 49892 10164 49948 10220
rect 50428 12684 50484 12740
rect 50876 12738 50932 12740
rect 50876 12686 50878 12738
rect 50878 12686 50930 12738
rect 50930 12686 50932 12738
rect 50876 12684 50932 12686
rect 48748 8204 48804 8260
rect 48076 7308 48132 7364
rect 49268 8596 49324 8652
rect 49372 8650 49428 8652
rect 49476 8650 49532 8652
rect 49372 8598 49396 8650
rect 49396 8598 49428 8650
rect 49476 8598 49520 8650
rect 49520 8598 49532 8650
rect 49372 8596 49428 8598
rect 49476 8596 49532 8598
rect 49580 8596 49636 8652
rect 49684 8650 49740 8652
rect 49788 8650 49844 8652
rect 49684 8598 49696 8650
rect 49696 8598 49740 8650
rect 49788 8598 49820 8650
rect 49820 8598 49844 8650
rect 49684 8596 49740 8598
rect 49788 8596 49844 8598
rect 49892 8596 49948 8652
rect 48972 7980 49028 8036
rect 49868 8316 49924 8372
rect 49868 7698 49924 7700
rect 49868 7646 49870 7698
rect 49870 7646 49922 7698
rect 49922 7646 49924 7698
rect 49868 7644 49924 7646
rect 48636 6860 48692 6916
rect 48188 5906 48244 5908
rect 48188 5854 48190 5906
rect 48190 5854 48242 5906
rect 48242 5854 48244 5906
rect 48188 5852 48244 5854
rect 49268 7028 49324 7084
rect 49372 7082 49428 7084
rect 49476 7082 49532 7084
rect 49372 7030 49396 7082
rect 49396 7030 49428 7082
rect 49476 7030 49520 7082
rect 49520 7030 49532 7082
rect 49372 7028 49428 7030
rect 49476 7028 49532 7030
rect 49580 7028 49636 7084
rect 49684 7082 49740 7084
rect 49788 7082 49844 7084
rect 49684 7030 49696 7082
rect 49696 7030 49740 7082
rect 49788 7030 49820 7082
rect 49820 7030 49844 7082
rect 49684 7028 49740 7030
rect 49788 7028 49844 7030
rect 49892 7028 49948 7084
rect 49084 6860 49140 6916
rect 50316 8316 50372 8372
rect 50204 7756 50260 7812
rect 50092 6636 50148 6692
rect 49980 6524 50036 6580
rect 49308 6412 49364 6468
rect 48972 5682 49028 5684
rect 48972 5630 48974 5682
rect 48974 5630 49026 5682
rect 49026 5630 49028 5682
rect 48972 5628 49028 5630
rect 50092 6076 50148 6132
rect 49268 5460 49324 5516
rect 49372 5514 49428 5516
rect 49476 5514 49532 5516
rect 49372 5462 49396 5514
rect 49396 5462 49428 5514
rect 49476 5462 49520 5514
rect 49520 5462 49532 5514
rect 49372 5460 49428 5462
rect 49476 5460 49532 5462
rect 49580 5460 49636 5516
rect 49684 5514 49740 5516
rect 49788 5514 49844 5516
rect 49684 5462 49696 5514
rect 49696 5462 49740 5514
rect 49788 5462 49820 5514
rect 49820 5462 49844 5514
rect 49684 5460 49740 5462
rect 49788 5460 49844 5462
rect 49892 5460 49948 5516
rect 48300 5122 48356 5124
rect 48300 5070 48302 5122
rect 48302 5070 48354 5122
rect 48354 5070 48356 5122
rect 48300 5068 48356 5070
rect 48188 4338 48244 4340
rect 48188 4286 48190 4338
rect 48190 4286 48242 4338
rect 48242 4286 48244 4338
rect 48188 4284 48244 4286
rect 49868 5068 49924 5124
rect 49420 4956 49476 5012
rect 49756 4450 49812 4452
rect 49756 4398 49758 4450
rect 49758 4398 49810 4450
rect 49810 4398 49812 4450
rect 49756 4396 49812 4398
rect 49980 4450 50036 4452
rect 49980 4398 49982 4450
rect 49982 4398 50034 4450
rect 50034 4398 50036 4450
rect 49980 4396 50036 4398
rect 48524 4060 48580 4116
rect 49196 4114 49252 4116
rect 49196 4062 49198 4114
rect 49198 4062 49250 4114
rect 49250 4062 49252 4114
rect 49196 4060 49252 4062
rect 49268 3892 49324 3948
rect 49372 3946 49428 3948
rect 49476 3946 49532 3948
rect 49372 3894 49396 3946
rect 49396 3894 49428 3946
rect 49476 3894 49520 3946
rect 49520 3894 49532 3946
rect 49372 3892 49428 3894
rect 49476 3892 49532 3894
rect 49580 3892 49636 3948
rect 49684 3946 49740 3948
rect 49788 3946 49844 3948
rect 49684 3894 49696 3946
rect 49696 3894 49740 3946
rect 49788 3894 49820 3946
rect 49820 3894 49844 3946
rect 49684 3892 49740 3894
rect 49788 3892 49844 3894
rect 49892 3892 49948 3948
rect 51100 10108 51156 10164
rect 50428 6076 50484 6132
rect 51324 12738 51380 12740
rect 51324 12686 51326 12738
rect 51326 12686 51378 12738
rect 51378 12686 51380 12738
rect 51324 12684 51380 12686
rect 51212 7644 51268 7700
rect 50764 4844 50820 4900
rect 50204 4396 50260 4452
rect 44940 3554 44996 3556
rect 44940 3502 44942 3554
rect 44942 3502 44994 3554
rect 44994 3502 44996 3554
rect 44940 3500 44996 3502
rect 46396 3500 46452 3556
rect 43820 3442 43876 3444
rect 43820 3390 43822 3442
rect 43822 3390 43874 3442
rect 43874 3390 43876 3442
rect 43820 3388 43876 3390
rect 43932 3330 43988 3332
rect 43932 3278 43934 3330
rect 43934 3278 43986 3330
rect 43986 3278 43988 3330
rect 43932 3276 43988 3278
rect 50204 3724 50260 3780
rect 49308 3554 49364 3556
rect 49308 3502 49310 3554
rect 49310 3502 49362 3554
rect 49362 3502 49364 3554
rect 49308 3500 49364 3502
rect 46732 3442 46788 3444
rect 46732 3390 46734 3442
rect 46734 3390 46786 3442
rect 46786 3390 46788 3442
rect 46732 3388 46788 3390
rect 48860 3442 48916 3444
rect 48860 3390 48862 3442
rect 48862 3390 48914 3442
rect 48914 3390 48916 3442
rect 48860 3388 48916 3390
rect 49420 3388 49476 3444
rect 55580 13970 55636 13972
rect 55580 13918 55582 13970
rect 55582 13918 55634 13970
rect 55634 13918 55636 13970
rect 55580 13916 55636 13918
rect 55132 13858 55188 13860
rect 55132 13806 55134 13858
rect 55134 13806 55186 13858
rect 55186 13806 55188 13858
rect 55132 13804 55188 13806
rect 52332 13634 52388 13636
rect 52332 13582 52334 13634
rect 52334 13582 52386 13634
rect 52386 13582 52388 13634
rect 52332 13580 52388 13582
rect 52108 9996 52164 10052
rect 51884 7532 51940 7588
rect 51996 7474 52052 7476
rect 51996 7422 51998 7474
rect 51998 7422 52050 7474
rect 52050 7422 52052 7474
rect 51996 7420 52052 7422
rect 51772 5234 51828 5236
rect 51772 5182 51774 5234
rect 51774 5182 51826 5234
rect 51826 5182 51828 5234
rect 51772 5180 51828 5182
rect 52332 4508 52388 4564
rect 51436 4060 51492 4116
rect 52780 7420 52836 7476
rect 54572 13746 54628 13748
rect 54572 13694 54574 13746
rect 54574 13694 54626 13746
rect 54626 13694 54628 13746
rect 54572 13692 54628 13694
rect 58940 13468 58996 13524
rect 58268 13300 58324 13356
rect 58372 13354 58428 13356
rect 58476 13354 58532 13356
rect 58372 13302 58396 13354
rect 58396 13302 58428 13354
rect 58476 13302 58520 13354
rect 58520 13302 58532 13354
rect 58372 13300 58428 13302
rect 58476 13300 58532 13302
rect 58580 13300 58636 13356
rect 58684 13354 58740 13356
rect 58788 13354 58844 13356
rect 58684 13302 58696 13354
rect 58696 13302 58740 13354
rect 58788 13302 58820 13354
rect 58820 13302 58844 13354
rect 58684 13300 58740 13302
rect 58788 13300 58844 13302
rect 58892 13300 58948 13356
rect 53768 12516 53824 12572
rect 53872 12570 53928 12572
rect 53976 12570 54032 12572
rect 53872 12518 53896 12570
rect 53896 12518 53928 12570
rect 53976 12518 54020 12570
rect 54020 12518 54032 12570
rect 53872 12516 53928 12518
rect 53976 12516 54032 12518
rect 54080 12516 54136 12572
rect 54184 12570 54240 12572
rect 54288 12570 54344 12572
rect 54184 12518 54196 12570
rect 54196 12518 54240 12570
rect 54288 12518 54320 12570
rect 54320 12518 54344 12570
rect 54184 12516 54240 12518
rect 54288 12516 54344 12518
rect 54392 12516 54448 12572
rect 57820 12348 57876 12404
rect 53768 10948 53824 11004
rect 53872 11002 53928 11004
rect 53976 11002 54032 11004
rect 53872 10950 53896 11002
rect 53896 10950 53928 11002
rect 53976 10950 54020 11002
rect 54020 10950 54032 11002
rect 53872 10948 53928 10950
rect 53976 10948 54032 10950
rect 54080 10948 54136 11004
rect 54184 11002 54240 11004
rect 54288 11002 54344 11004
rect 54184 10950 54196 11002
rect 54196 10950 54240 11002
rect 54288 10950 54320 11002
rect 54320 10950 54344 11002
rect 54184 10948 54240 10950
rect 54288 10948 54344 10950
rect 54392 10948 54448 11004
rect 54684 10108 54740 10164
rect 53768 9380 53824 9436
rect 53872 9434 53928 9436
rect 53976 9434 54032 9436
rect 53872 9382 53896 9434
rect 53896 9382 53928 9434
rect 53976 9382 54020 9434
rect 54020 9382 54032 9434
rect 53872 9380 53928 9382
rect 53976 9380 54032 9382
rect 54080 9380 54136 9436
rect 54184 9434 54240 9436
rect 54288 9434 54344 9436
rect 54184 9382 54196 9434
rect 54196 9382 54240 9434
rect 54288 9382 54320 9434
rect 54320 9382 54344 9434
rect 54184 9380 54240 9382
rect 54288 9380 54344 9382
rect 54392 9380 54448 9436
rect 53768 7812 53824 7868
rect 53872 7866 53928 7868
rect 53976 7866 54032 7868
rect 53872 7814 53896 7866
rect 53896 7814 53928 7866
rect 53976 7814 54020 7866
rect 54020 7814 54032 7866
rect 53872 7812 53928 7814
rect 53976 7812 54032 7814
rect 54080 7812 54136 7868
rect 54184 7866 54240 7868
rect 54288 7866 54344 7868
rect 54184 7814 54196 7866
rect 54196 7814 54240 7866
rect 54288 7814 54320 7866
rect 54320 7814 54344 7866
rect 54184 7812 54240 7814
rect 54288 7812 54344 7814
rect 54392 7812 54448 7868
rect 56140 8316 56196 8372
rect 54684 8146 54740 8148
rect 54684 8094 54686 8146
rect 54686 8094 54738 8146
rect 54738 8094 54740 8146
rect 54684 8092 54740 8094
rect 53788 6412 53844 6468
rect 53768 6244 53824 6300
rect 53872 6298 53928 6300
rect 53976 6298 54032 6300
rect 53872 6246 53896 6298
rect 53896 6246 53928 6298
rect 53976 6246 54020 6298
rect 54020 6246 54032 6298
rect 53872 6244 53928 6246
rect 53976 6244 54032 6246
rect 54080 6244 54136 6300
rect 54184 6298 54240 6300
rect 54288 6298 54344 6300
rect 54184 6246 54196 6298
rect 54196 6246 54240 6298
rect 54288 6246 54320 6298
rect 54320 6246 54344 6298
rect 54184 6244 54240 6246
rect 54288 6244 54344 6246
rect 54392 6244 54448 6300
rect 54572 5852 54628 5908
rect 54684 7644 54740 7700
rect 53452 5292 53508 5348
rect 53228 5180 53284 5236
rect 55356 7420 55412 7476
rect 54908 6578 54964 6580
rect 54908 6526 54910 6578
rect 54910 6526 54962 6578
rect 54962 6526 54964 6578
rect 54908 6524 54964 6526
rect 56588 7474 56644 7476
rect 56588 7422 56590 7474
rect 56590 7422 56642 7474
rect 56642 7422 56644 7474
rect 56588 7420 56644 7422
rect 53768 4676 53824 4732
rect 53872 4730 53928 4732
rect 53976 4730 54032 4732
rect 53872 4678 53896 4730
rect 53896 4678 53928 4730
rect 53976 4678 54020 4730
rect 54020 4678 54032 4730
rect 53872 4676 53928 4678
rect 53976 4676 54032 4678
rect 54080 4676 54136 4732
rect 54184 4730 54240 4732
rect 54288 4730 54344 4732
rect 54184 4678 54196 4730
rect 54196 4678 54240 4730
rect 54288 4678 54320 4730
rect 54320 4678 54344 4730
rect 54184 4676 54240 4678
rect 54288 4676 54344 4678
rect 54392 4676 54448 4732
rect 52780 4450 52836 4452
rect 52780 4398 52782 4450
rect 52782 4398 52834 4450
rect 52834 4398 52836 4450
rect 52780 4396 52836 4398
rect 57148 5180 57204 5236
rect 56700 3724 56756 3780
rect 57484 4060 57540 4116
rect 52444 3612 52500 3668
rect 55468 3666 55524 3668
rect 55468 3614 55470 3666
rect 55470 3614 55522 3666
rect 55522 3614 55524 3666
rect 55468 3612 55524 3614
rect 59052 12348 59108 12404
rect 60284 13468 60340 13524
rect 58268 11732 58324 11788
rect 58372 11786 58428 11788
rect 58476 11786 58532 11788
rect 58372 11734 58396 11786
rect 58396 11734 58428 11786
rect 58476 11734 58520 11786
rect 58520 11734 58532 11786
rect 58372 11732 58428 11734
rect 58476 11732 58532 11734
rect 58580 11732 58636 11788
rect 58684 11786 58740 11788
rect 58788 11786 58844 11788
rect 58684 11734 58696 11786
rect 58696 11734 58740 11786
rect 58788 11734 58820 11786
rect 58820 11734 58844 11786
rect 58684 11732 58740 11734
rect 58788 11732 58844 11734
rect 58892 11732 58948 11788
rect 58156 11394 58212 11396
rect 58156 11342 58158 11394
rect 58158 11342 58210 11394
rect 58210 11342 58212 11394
rect 58156 11340 58212 11342
rect 57820 8316 57876 8372
rect 59388 11116 59444 11172
rect 58268 10164 58324 10220
rect 58372 10218 58428 10220
rect 58476 10218 58532 10220
rect 58372 10166 58396 10218
rect 58396 10166 58428 10218
rect 58476 10166 58520 10218
rect 58520 10166 58532 10218
rect 58372 10164 58428 10166
rect 58476 10164 58532 10166
rect 58580 10164 58636 10220
rect 58684 10218 58740 10220
rect 58788 10218 58844 10220
rect 58684 10166 58696 10218
rect 58696 10166 58740 10218
rect 58788 10166 58820 10218
rect 58820 10166 58844 10218
rect 58684 10164 58740 10166
rect 58788 10164 58844 10166
rect 58892 10164 58948 10220
rect 59276 9996 59332 10052
rect 58268 8596 58324 8652
rect 58372 8650 58428 8652
rect 58476 8650 58532 8652
rect 58372 8598 58396 8650
rect 58396 8598 58428 8650
rect 58476 8598 58520 8650
rect 58520 8598 58532 8650
rect 58372 8596 58428 8598
rect 58476 8596 58532 8598
rect 58580 8596 58636 8652
rect 58684 8650 58740 8652
rect 58788 8650 58844 8652
rect 58684 8598 58696 8650
rect 58696 8598 58740 8650
rect 58788 8598 58820 8650
rect 58820 8598 58844 8650
rect 58684 8596 58740 8598
rect 58788 8596 58844 8598
rect 58892 8596 58948 8652
rect 58828 8370 58884 8372
rect 58828 8318 58830 8370
rect 58830 8318 58882 8370
rect 58882 8318 58884 8370
rect 58828 8316 58884 8318
rect 59164 7532 59220 7588
rect 58268 7028 58324 7084
rect 58372 7082 58428 7084
rect 58476 7082 58532 7084
rect 58372 7030 58396 7082
rect 58396 7030 58428 7082
rect 58476 7030 58520 7082
rect 58520 7030 58532 7082
rect 58372 7028 58428 7030
rect 58476 7028 58532 7030
rect 58580 7028 58636 7084
rect 58684 7082 58740 7084
rect 58788 7082 58844 7084
rect 58684 7030 58696 7082
rect 58696 7030 58740 7082
rect 58788 7030 58820 7082
rect 58820 7030 58844 7082
rect 58684 7028 58740 7030
rect 58788 7028 58844 7030
rect 58892 7028 58948 7084
rect 58044 6636 58100 6692
rect 58828 6748 58884 6804
rect 59052 6524 59108 6580
rect 57932 5292 57988 5348
rect 58268 5460 58324 5516
rect 58372 5514 58428 5516
rect 58476 5514 58532 5516
rect 58372 5462 58396 5514
rect 58396 5462 58428 5514
rect 58476 5462 58520 5514
rect 58520 5462 58532 5514
rect 58372 5460 58428 5462
rect 58476 5460 58532 5462
rect 58580 5460 58636 5516
rect 58684 5514 58740 5516
rect 58788 5514 58844 5516
rect 58684 5462 58696 5514
rect 58696 5462 58740 5514
rect 58788 5462 58820 5514
rect 58820 5462 58844 5514
rect 58684 5460 58740 5462
rect 58788 5460 58844 5462
rect 58892 5460 58948 5516
rect 58716 5292 58772 5348
rect 59164 5122 59220 5124
rect 59164 5070 59166 5122
rect 59166 5070 59218 5122
rect 59218 5070 59220 5122
rect 59164 5068 59220 5070
rect 59836 6300 59892 6356
rect 59612 5010 59668 5012
rect 59612 4958 59614 5010
rect 59614 4958 59666 5010
rect 59666 4958 59668 5010
rect 59612 4956 59668 4958
rect 59276 4284 59332 4340
rect 59388 4844 59444 4900
rect 59388 4060 59444 4116
rect 58268 3892 58324 3948
rect 58372 3946 58428 3948
rect 58476 3946 58532 3948
rect 58372 3894 58396 3946
rect 58396 3894 58428 3946
rect 58476 3894 58520 3946
rect 58520 3894 58532 3946
rect 58372 3892 58428 3894
rect 58476 3892 58532 3894
rect 58580 3892 58636 3948
rect 58684 3946 58740 3948
rect 58788 3946 58844 3948
rect 58684 3894 58696 3946
rect 58696 3894 58740 3946
rect 58788 3894 58820 3946
rect 58820 3894 58844 3946
rect 58684 3892 58740 3894
rect 58788 3892 58844 3894
rect 58892 3892 58948 3948
rect 59052 3724 59108 3780
rect 50428 3500 50484 3556
rect 54572 3554 54628 3556
rect 54572 3502 54574 3554
rect 54574 3502 54626 3554
rect 54626 3502 54628 3554
rect 54572 3500 54628 3502
rect 55020 3554 55076 3556
rect 55020 3502 55022 3554
rect 55022 3502 55074 3554
rect 55074 3502 55076 3554
rect 55020 3500 55076 3502
rect 58156 3554 58212 3556
rect 58156 3502 58158 3554
rect 58158 3502 58210 3554
rect 58210 3502 58212 3554
rect 58156 3500 58212 3502
rect 59836 3612 59892 3668
rect 60620 11170 60676 11172
rect 60620 11118 60622 11170
rect 60622 11118 60674 11170
rect 60674 11118 60676 11170
rect 60620 11116 60676 11118
rect 60508 6690 60564 6692
rect 60508 6638 60510 6690
rect 60510 6638 60562 6690
rect 60562 6638 60564 6690
rect 60508 6636 60564 6638
rect 61068 11170 61124 11172
rect 61068 11118 61070 11170
rect 61070 11118 61122 11170
rect 61122 11118 61124 11170
rect 61068 11116 61124 11118
rect 62636 28364 62692 28420
rect 63084 28418 63140 28420
rect 63084 28366 63086 28418
rect 63086 28366 63138 28418
rect 63138 28366 63140 28418
rect 63084 28364 63140 28366
rect 62768 28196 62824 28252
rect 62872 28250 62928 28252
rect 62976 28250 63032 28252
rect 62872 28198 62896 28250
rect 62896 28198 62928 28250
rect 62976 28198 63020 28250
rect 63020 28198 63032 28250
rect 62872 28196 62928 28198
rect 62976 28196 63032 28198
rect 63080 28196 63136 28252
rect 63184 28250 63240 28252
rect 63288 28250 63344 28252
rect 63184 28198 63196 28250
rect 63196 28198 63240 28250
rect 63288 28198 63320 28250
rect 63320 28198 63344 28250
rect 63184 28196 63240 28198
rect 63288 28196 63344 28198
rect 63392 28196 63448 28252
rect 61740 27580 61796 27636
rect 62748 27074 62804 27076
rect 62748 27022 62750 27074
rect 62750 27022 62802 27074
rect 62802 27022 62804 27074
rect 62748 27020 62804 27022
rect 61740 26962 61796 26964
rect 61740 26910 61742 26962
rect 61742 26910 61794 26962
rect 61794 26910 61796 26962
rect 61740 26908 61796 26910
rect 61404 26850 61460 26852
rect 61404 26798 61406 26850
rect 61406 26798 61458 26850
rect 61458 26798 61460 26850
rect 61404 26796 61460 26798
rect 62300 26962 62356 26964
rect 62300 26910 62302 26962
rect 62302 26910 62354 26962
rect 62354 26910 62356 26962
rect 62300 26908 62356 26910
rect 62300 26684 62356 26740
rect 62768 26628 62824 26684
rect 62872 26682 62928 26684
rect 62976 26682 63032 26684
rect 62872 26630 62896 26682
rect 62896 26630 62928 26682
rect 62976 26630 63020 26682
rect 63020 26630 63032 26682
rect 62872 26628 62928 26630
rect 62976 26628 63032 26630
rect 63080 26628 63136 26684
rect 63184 26682 63240 26684
rect 63288 26682 63344 26684
rect 63184 26630 63196 26682
rect 63196 26630 63240 26682
rect 63288 26630 63320 26682
rect 63320 26630 63344 26682
rect 63184 26628 63240 26630
rect 63288 26628 63344 26630
rect 63392 26628 63448 26684
rect 62300 26290 62356 26292
rect 62300 26238 62302 26290
rect 62302 26238 62354 26290
rect 62354 26238 62356 26290
rect 62300 26236 62356 26238
rect 62972 25506 63028 25508
rect 62972 25454 62974 25506
rect 62974 25454 63026 25506
rect 63026 25454 63028 25506
rect 62972 25452 63028 25454
rect 62076 24444 62132 24500
rect 61404 23714 61460 23716
rect 61404 23662 61406 23714
rect 61406 23662 61458 23714
rect 61458 23662 61460 23714
rect 61404 23660 61460 23662
rect 62524 25282 62580 25284
rect 62524 25230 62526 25282
rect 62526 25230 62578 25282
rect 62578 25230 62580 25282
rect 62524 25228 62580 25230
rect 64428 28642 64484 28644
rect 64428 28590 64430 28642
rect 64430 28590 64482 28642
rect 64482 28590 64484 28642
rect 64428 28588 64484 28590
rect 65100 31666 65156 31668
rect 65100 31614 65102 31666
rect 65102 31614 65154 31666
rect 65154 31614 65156 31666
rect 65100 31612 65156 31614
rect 65100 31164 65156 31220
rect 65324 31554 65380 31556
rect 65324 31502 65326 31554
rect 65326 31502 65378 31554
rect 65378 31502 65380 31554
rect 65324 31500 65380 31502
rect 66108 33628 66164 33684
rect 67900 34690 67956 34692
rect 67900 34638 67902 34690
rect 67902 34638 67954 34690
rect 67954 34638 67956 34690
rect 67900 34636 67956 34638
rect 68124 35980 68180 36036
rect 68460 35980 68516 36036
rect 68236 35644 68292 35700
rect 68012 34188 68068 34244
rect 67004 33628 67060 33684
rect 67268 33684 67324 33740
rect 67372 33738 67428 33740
rect 67476 33738 67532 33740
rect 67372 33686 67396 33738
rect 67396 33686 67428 33738
rect 67476 33686 67520 33738
rect 67520 33686 67532 33738
rect 67372 33684 67428 33686
rect 67476 33684 67532 33686
rect 67580 33684 67636 33740
rect 67684 33738 67740 33740
rect 67788 33738 67844 33740
rect 67684 33686 67696 33738
rect 67696 33686 67740 33738
rect 67788 33686 67820 33738
rect 67820 33686 67844 33738
rect 67684 33684 67740 33686
rect 67788 33684 67844 33686
rect 67892 33684 67948 33740
rect 66668 33122 66724 33124
rect 66668 33070 66670 33122
rect 66670 33070 66722 33122
rect 66722 33070 66724 33122
rect 66668 33068 66724 33070
rect 68348 35308 68404 35364
rect 69468 36316 69524 36372
rect 69580 36764 69636 36820
rect 73948 37884 74004 37940
rect 74284 37938 74340 37940
rect 74284 37886 74286 37938
rect 74286 37886 74338 37938
rect 74338 37886 74340 37938
rect 74284 37884 74340 37886
rect 73500 36540 73556 36596
rect 71768 36036 71824 36092
rect 71872 36090 71928 36092
rect 71976 36090 72032 36092
rect 71872 36038 71896 36090
rect 71896 36038 71928 36090
rect 71976 36038 72020 36090
rect 72020 36038 72032 36090
rect 71872 36036 71928 36038
rect 71976 36036 72032 36038
rect 72080 36036 72136 36092
rect 72184 36090 72240 36092
rect 72288 36090 72344 36092
rect 72184 36038 72196 36090
rect 72196 36038 72240 36090
rect 72288 36038 72320 36090
rect 72320 36038 72344 36090
rect 72184 36036 72240 36038
rect 72288 36036 72344 36038
rect 72392 36036 72448 36092
rect 69580 35868 69636 35924
rect 71932 35868 71988 35924
rect 68908 35308 68964 35364
rect 73724 35868 73780 35924
rect 68236 32620 68292 32676
rect 71148 34690 71204 34692
rect 71148 34638 71150 34690
rect 71150 34638 71202 34690
rect 71202 34638 71204 34690
rect 71148 34636 71204 34638
rect 67268 32116 67324 32172
rect 67372 32170 67428 32172
rect 67476 32170 67532 32172
rect 67372 32118 67396 32170
rect 67396 32118 67428 32170
rect 67476 32118 67520 32170
rect 67520 32118 67532 32170
rect 67372 32116 67428 32118
rect 67476 32116 67532 32118
rect 67580 32116 67636 32172
rect 67684 32170 67740 32172
rect 67788 32170 67844 32172
rect 67684 32118 67696 32170
rect 67696 32118 67740 32170
rect 67788 32118 67820 32170
rect 67820 32118 67844 32170
rect 67684 32116 67740 32118
rect 67788 32116 67844 32118
rect 67892 32116 67948 32172
rect 67004 31836 67060 31892
rect 67900 31836 67956 31892
rect 65212 30940 65268 30996
rect 64764 28588 64820 28644
rect 63644 27580 63700 27636
rect 63868 27020 63924 27076
rect 63308 25282 63364 25284
rect 63308 25230 63310 25282
rect 63310 25230 63362 25282
rect 63362 25230 63364 25282
rect 63308 25228 63364 25230
rect 62768 25060 62824 25116
rect 62872 25114 62928 25116
rect 62976 25114 63032 25116
rect 62872 25062 62896 25114
rect 62896 25062 62928 25114
rect 62976 25062 63020 25114
rect 63020 25062 63032 25114
rect 62872 25060 62928 25062
rect 62976 25060 63032 25062
rect 63080 25060 63136 25116
rect 63184 25114 63240 25116
rect 63288 25114 63344 25116
rect 63184 25062 63196 25114
rect 63196 25062 63240 25114
rect 63288 25062 63320 25114
rect 63320 25062 63344 25114
rect 63184 25060 63240 25062
rect 63288 25060 63344 25062
rect 63392 25060 63448 25116
rect 62768 23492 62824 23548
rect 62872 23546 62928 23548
rect 62976 23546 63032 23548
rect 62872 23494 62896 23546
rect 62896 23494 62928 23546
rect 62976 23494 63020 23546
rect 63020 23494 63032 23546
rect 62872 23492 62928 23494
rect 62976 23492 63032 23494
rect 63080 23492 63136 23548
rect 63184 23546 63240 23548
rect 63288 23546 63344 23548
rect 63184 23494 63196 23546
rect 63196 23494 63240 23546
rect 63288 23494 63320 23546
rect 63320 23494 63344 23546
rect 63184 23492 63240 23494
rect 63288 23492 63344 23494
rect 63392 23492 63448 23548
rect 64540 26236 64596 26292
rect 62972 23154 63028 23156
rect 62972 23102 62974 23154
rect 62974 23102 63026 23154
rect 63026 23102 63028 23154
rect 62972 23100 63028 23102
rect 64204 23100 64260 23156
rect 62768 21924 62824 21980
rect 62872 21978 62928 21980
rect 62976 21978 63032 21980
rect 62872 21926 62896 21978
rect 62896 21926 62928 21978
rect 62976 21926 63020 21978
rect 63020 21926 63032 21978
rect 62872 21924 62928 21926
rect 62976 21924 63032 21926
rect 63080 21924 63136 21980
rect 63184 21978 63240 21980
rect 63288 21978 63344 21980
rect 63184 21926 63196 21978
rect 63196 21926 63240 21978
rect 63288 21926 63320 21978
rect 63320 21926 63344 21978
rect 63184 21924 63240 21926
rect 63288 21924 63344 21926
rect 63392 21924 63448 21980
rect 65996 31164 66052 31220
rect 65436 30994 65492 30996
rect 65436 30942 65438 30994
rect 65438 30942 65490 30994
rect 65490 30942 65492 30994
rect 65436 30940 65492 30942
rect 66556 31554 66612 31556
rect 66556 31502 66558 31554
rect 66558 31502 66610 31554
rect 66610 31502 66612 31554
rect 66556 31500 66612 31502
rect 67268 30548 67324 30604
rect 67372 30602 67428 30604
rect 67476 30602 67532 30604
rect 67372 30550 67396 30602
rect 67396 30550 67428 30602
rect 67476 30550 67520 30602
rect 67520 30550 67532 30602
rect 67372 30548 67428 30550
rect 67476 30548 67532 30550
rect 67580 30548 67636 30604
rect 67684 30602 67740 30604
rect 67788 30602 67844 30604
rect 67684 30550 67696 30602
rect 67696 30550 67740 30602
rect 67788 30550 67820 30602
rect 67820 30550 67844 30602
rect 67684 30548 67740 30550
rect 67788 30548 67844 30550
rect 67892 30548 67948 30604
rect 66668 30156 66724 30212
rect 67268 28980 67324 29036
rect 67372 29034 67428 29036
rect 67476 29034 67532 29036
rect 67372 28982 67396 29034
rect 67396 28982 67428 29034
rect 67476 28982 67520 29034
rect 67520 28982 67532 29034
rect 67372 28980 67428 28982
rect 67476 28980 67532 28982
rect 67580 28980 67636 29036
rect 67684 29034 67740 29036
rect 67788 29034 67844 29036
rect 67684 28982 67696 29034
rect 67696 28982 67740 29034
rect 67788 28982 67820 29034
rect 67820 28982 67844 29034
rect 67684 28980 67740 28982
rect 67788 28980 67844 28982
rect 67892 28980 67948 29036
rect 68348 29314 68404 29316
rect 68348 29262 68350 29314
rect 68350 29262 68402 29314
rect 68402 29262 68404 29314
rect 68348 29260 68404 29262
rect 65660 27970 65716 27972
rect 65660 27918 65662 27970
rect 65662 27918 65714 27970
rect 65714 27918 65716 27970
rect 65660 27916 65716 27918
rect 66332 27916 66388 27972
rect 65660 27634 65716 27636
rect 65660 27582 65662 27634
rect 65662 27582 65714 27634
rect 65714 27582 65716 27634
rect 65660 27580 65716 27582
rect 65436 26236 65492 26292
rect 65324 25564 65380 25620
rect 64988 25506 65044 25508
rect 64988 25454 64990 25506
rect 64990 25454 65042 25506
rect 65042 25454 65044 25506
rect 64988 25452 65044 25454
rect 64652 23772 64708 23828
rect 65212 23548 65268 23604
rect 64652 21698 64708 21700
rect 64652 21646 64654 21698
rect 64654 21646 64706 21698
rect 64706 21646 64708 21698
rect 64652 21644 64708 21646
rect 65100 21698 65156 21700
rect 65100 21646 65102 21698
rect 65102 21646 65154 21698
rect 65154 21646 65156 21698
rect 65100 21644 65156 21646
rect 64540 20972 64596 21028
rect 65212 21026 65268 21028
rect 65212 20974 65214 21026
rect 65214 20974 65266 21026
rect 65266 20974 65268 21026
rect 65212 20972 65268 20974
rect 64652 20860 64708 20916
rect 62768 20356 62824 20412
rect 62872 20410 62928 20412
rect 62976 20410 63032 20412
rect 62872 20358 62896 20410
rect 62896 20358 62928 20410
rect 62976 20358 63020 20410
rect 63020 20358 63032 20410
rect 62872 20356 62928 20358
rect 62976 20356 63032 20358
rect 63080 20356 63136 20412
rect 63184 20410 63240 20412
rect 63288 20410 63344 20412
rect 63184 20358 63196 20410
rect 63196 20358 63240 20410
rect 63288 20358 63320 20410
rect 63320 20358 63344 20410
rect 63184 20356 63240 20358
rect 63288 20356 63344 20358
rect 63392 20356 63448 20412
rect 62768 18788 62824 18844
rect 62872 18842 62928 18844
rect 62976 18842 63032 18844
rect 62872 18790 62896 18842
rect 62896 18790 62928 18842
rect 62976 18790 63020 18842
rect 63020 18790 63032 18842
rect 62872 18788 62928 18790
rect 62976 18788 63032 18790
rect 63080 18788 63136 18844
rect 63184 18842 63240 18844
rect 63288 18842 63344 18844
rect 63184 18790 63196 18842
rect 63196 18790 63240 18842
rect 63288 18790 63320 18842
rect 63320 18790 63344 18842
rect 63184 18788 63240 18790
rect 63288 18788 63344 18790
rect 63392 18788 63448 18844
rect 62768 17220 62824 17276
rect 62872 17274 62928 17276
rect 62976 17274 63032 17276
rect 62872 17222 62896 17274
rect 62896 17222 62928 17274
rect 62976 17222 63020 17274
rect 63020 17222 63032 17274
rect 62872 17220 62928 17222
rect 62976 17220 63032 17222
rect 63080 17220 63136 17276
rect 63184 17274 63240 17276
rect 63288 17274 63344 17276
rect 63184 17222 63196 17274
rect 63196 17222 63240 17274
rect 63288 17222 63320 17274
rect 63320 17222 63344 17274
rect 63184 17220 63240 17222
rect 63288 17220 63344 17222
rect 63392 17220 63448 17276
rect 62768 15652 62824 15708
rect 62872 15706 62928 15708
rect 62976 15706 63032 15708
rect 62872 15654 62896 15706
rect 62896 15654 62928 15706
rect 62976 15654 63020 15706
rect 63020 15654 63032 15706
rect 62872 15652 62928 15654
rect 62976 15652 63032 15654
rect 63080 15652 63136 15708
rect 63184 15706 63240 15708
rect 63288 15706 63344 15708
rect 63184 15654 63196 15706
rect 63196 15654 63240 15706
rect 63288 15654 63320 15706
rect 63320 15654 63344 15706
rect 63184 15652 63240 15654
rect 63288 15652 63344 15654
rect 63392 15652 63448 15708
rect 66332 27244 66388 27300
rect 68348 28700 68404 28756
rect 66780 26684 66836 26740
rect 65772 25618 65828 25620
rect 65772 25566 65774 25618
rect 65774 25566 65826 25618
rect 65826 25566 65828 25618
rect 65772 25564 65828 25566
rect 66332 24946 66388 24948
rect 66332 24894 66334 24946
rect 66334 24894 66386 24946
rect 66386 24894 66388 24946
rect 66332 24892 66388 24894
rect 67268 27412 67324 27468
rect 67372 27466 67428 27468
rect 67476 27466 67532 27468
rect 67372 27414 67396 27466
rect 67396 27414 67428 27466
rect 67476 27414 67520 27466
rect 67520 27414 67532 27466
rect 67372 27412 67428 27414
rect 67476 27412 67532 27414
rect 67580 27412 67636 27468
rect 67684 27466 67740 27468
rect 67788 27466 67844 27468
rect 67684 27414 67696 27466
rect 67696 27414 67740 27466
rect 67788 27414 67820 27466
rect 67820 27414 67844 27466
rect 67684 27412 67740 27414
rect 67788 27412 67844 27414
rect 67892 27412 67948 27468
rect 67228 27244 67284 27300
rect 67564 27244 67620 27300
rect 71768 34468 71824 34524
rect 71872 34522 71928 34524
rect 71976 34522 72032 34524
rect 71872 34470 71896 34522
rect 71896 34470 71928 34522
rect 71976 34470 72020 34522
rect 72020 34470 72032 34522
rect 71872 34468 71928 34470
rect 71976 34468 72032 34470
rect 72080 34468 72136 34524
rect 72184 34522 72240 34524
rect 72288 34522 72344 34524
rect 72184 34470 72196 34522
rect 72196 34470 72240 34522
rect 72288 34470 72320 34522
rect 72320 34470 72344 34522
rect 72184 34468 72240 34470
rect 72288 34468 72344 34470
rect 72392 34468 72448 34524
rect 72492 34354 72548 34356
rect 72492 34302 72494 34354
rect 72494 34302 72546 34354
rect 72546 34302 72548 34354
rect 72492 34300 72548 34302
rect 73388 34130 73444 34132
rect 73388 34078 73390 34130
rect 73390 34078 73442 34130
rect 73442 34078 73444 34130
rect 73388 34076 73444 34078
rect 74732 35420 74788 35476
rect 74508 34354 74564 34356
rect 74508 34302 74510 34354
rect 74510 34302 74562 34354
rect 74562 34302 74564 34354
rect 74508 34300 74564 34302
rect 74284 34130 74340 34132
rect 74284 34078 74286 34130
rect 74286 34078 74338 34130
rect 74338 34078 74340 34130
rect 74284 34076 74340 34078
rect 75068 40236 75124 40292
rect 75404 42530 75460 42532
rect 75404 42478 75406 42530
rect 75406 42478 75458 42530
rect 75458 42478 75460 42530
rect 75404 42476 75460 42478
rect 75740 41916 75796 41972
rect 75628 40962 75684 40964
rect 75628 40910 75630 40962
rect 75630 40910 75682 40962
rect 75682 40910 75684 40962
rect 75628 40908 75684 40910
rect 75404 39004 75460 39060
rect 74956 37826 75012 37828
rect 74956 37774 74958 37826
rect 74958 37774 75010 37826
rect 75010 37774 75012 37826
rect 74956 37772 75012 37774
rect 75404 38220 75460 38276
rect 75628 37996 75684 38052
rect 75292 37100 75348 37156
rect 77420 48242 77476 48244
rect 77420 48190 77422 48242
rect 77422 48190 77474 48242
rect 77474 48190 77476 48242
rect 77420 48188 77476 48190
rect 76972 48076 77028 48132
rect 76268 47796 76324 47852
rect 76372 47850 76428 47852
rect 76476 47850 76532 47852
rect 76372 47798 76396 47850
rect 76396 47798 76428 47850
rect 76476 47798 76520 47850
rect 76520 47798 76532 47850
rect 76372 47796 76428 47798
rect 76476 47796 76532 47798
rect 76580 47796 76636 47852
rect 76684 47850 76740 47852
rect 76788 47850 76844 47852
rect 76684 47798 76696 47850
rect 76696 47798 76740 47850
rect 76788 47798 76820 47850
rect 76820 47798 76844 47850
rect 76684 47796 76740 47798
rect 76788 47796 76844 47798
rect 76892 47796 76948 47852
rect 77420 47964 77476 48020
rect 77308 47292 77364 47348
rect 76636 46562 76692 46564
rect 76636 46510 76638 46562
rect 76638 46510 76690 46562
rect 76690 46510 76692 46562
rect 76636 46508 76692 46510
rect 76268 46228 76324 46284
rect 76372 46282 76428 46284
rect 76476 46282 76532 46284
rect 76372 46230 76396 46282
rect 76396 46230 76428 46282
rect 76476 46230 76520 46282
rect 76520 46230 76532 46282
rect 76372 46228 76428 46230
rect 76476 46228 76532 46230
rect 76580 46228 76636 46284
rect 76684 46282 76740 46284
rect 76788 46282 76844 46284
rect 76684 46230 76696 46282
rect 76696 46230 76740 46282
rect 76788 46230 76820 46282
rect 76820 46230 76844 46282
rect 76684 46228 76740 46230
rect 76788 46228 76844 46230
rect 76892 46228 76948 46284
rect 77084 45890 77140 45892
rect 77084 45838 77086 45890
rect 77086 45838 77138 45890
rect 77138 45838 77140 45890
rect 77084 45836 77140 45838
rect 77308 45890 77364 45892
rect 77308 45838 77310 45890
rect 77310 45838 77362 45890
rect 77362 45838 77364 45890
rect 77308 45836 77364 45838
rect 78876 49084 78932 49140
rect 78428 48860 78484 48916
rect 78316 48354 78372 48356
rect 78316 48302 78318 48354
rect 78318 48302 78370 48354
rect 78370 48302 78372 48354
rect 78316 48300 78372 48302
rect 78092 47964 78148 48020
rect 78092 47292 78148 47348
rect 77420 45666 77476 45668
rect 77420 45614 77422 45666
rect 77422 45614 77474 45666
rect 77474 45614 77476 45666
rect 77420 45612 77476 45614
rect 76748 45218 76804 45220
rect 76748 45166 76750 45218
rect 76750 45166 76802 45218
rect 76802 45166 76804 45218
rect 76748 45164 76804 45166
rect 76300 44994 76356 44996
rect 76300 44942 76302 44994
rect 76302 44942 76354 44994
rect 76354 44942 76356 44994
rect 76300 44940 76356 44942
rect 76268 44660 76324 44716
rect 76372 44714 76428 44716
rect 76476 44714 76532 44716
rect 76372 44662 76396 44714
rect 76396 44662 76428 44714
rect 76476 44662 76520 44714
rect 76520 44662 76532 44714
rect 76372 44660 76428 44662
rect 76476 44660 76532 44662
rect 76580 44660 76636 44716
rect 76684 44714 76740 44716
rect 76788 44714 76844 44716
rect 76684 44662 76696 44714
rect 76696 44662 76740 44714
rect 76788 44662 76820 44714
rect 76820 44662 76844 44714
rect 76684 44660 76740 44662
rect 76788 44660 76844 44662
rect 76892 44660 76948 44716
rect 76636 44098 76692 44100
rect 76636 44046 76638 44098
rect 76638 44046 76690 44098
rect 76690 44046 76692 44098
rect 76636 44044 76692 44046
rect 77756 45218 77812 45220
rect 77756 45166 77758 45218
rect 77758 45166 77810 45218
rect 77810 45166 77812 45218
rect 77756 45164 77812 45166
rect 77532 44940 77588 44996
rect 77308 44044 77364 44100
rect 76972 43650 77028 43652
rect 76972 43598 76974 43650
rect 76974 43598 77026 43650
rect 77026 43598 77028 43650
rect 76972 43596 77028 43598
rect 77420 43596 77476 43652
rect 76268 43092 76324 43148
rect 76372 43146 76428 43148
rect 76476 43146 76532 43148
rect 76372 43094 76396 43146
rect 76396 43094 76428 43146
rect 76476 43094 76520 43146
rect 76520 43094 76532 43146
rect 76372 43092 76428 43094
rect 76476 43092 76532 43094
rect 76580 43092 76636 43148
rect 76684 43146 76740 43148
rect 76788 43146 76844 43148
rect 76684 43094 76696 43146
rect 76696 43094 76740 43146
rect 76788 43094 76820 43146
rect 76820 43094 76844 43146
rect 76684 43092 76740 43094
rect 76788 43092 76844 43094
rect 76892 43092 76948 43148
rect 77196 43260 77252 43316
rect 77084 42476 77140 42532
rect 76860 41970 76916 41972
rect 76860 41918 76862 41970
rect 76862 41918 76914 41970
rect 76914 41918 76916 41970
rect 76860 41916 76916 41918
rect 76412 41858 76468 41860
rect 76412 41806 76414 41858
rect 76414 41806 76466 41858
rect 76466 41806 76468 41858
rect 76412 41804 76468 41806
rect 76268 41524 76324 41580
rect 76372 41578 76428 41580
rect 76476 41578 76532 41580
rect 76372 41526 76396 41578
rect 76396 41526 76428 41578
rect 76476 41526 76520 41578
rect 76520 41526 76532 41578
rect 76372 41524 76428 41526
rect 76476 41524 76532 41526
rect 76580 41524 76636 41580
rect 76684 41578 76740 41580
rect 76788 41578 76844 41580
rect 76684 41526 76696 41578
rect 76696 41526 76740 41578
rect 76788 41526 76820 41578
rect 76820 41526 76844 41578
rect 76684 41524 76740 41526
rect 76788 41524 76844 41526
rect 76892 41524 76948 41580
rect 76748 41356 76804 41412
rect 76188 41132 76244 41188
rect 76300 41074 76356 41076
rect 76300 41022 76302 41074
rect 76302 41022 76354 41074
rect 76354 41022 76356 41074
rect 76300 41020 76356 41022
rect 76860 41074 76916 41076
rect 76860 41022 76862 41074
rect 76862 41022 76914 41074
rect 76914 41022 76916 41074
rect 76860 41020 76916 41022
rect 76412 40908 76468 40964
rect 76300 40796 76356 40852
rect 76972 40348 77028 40404
rect 75964 39788 76020 39844
rect 76268 39956 76324 40012
rect 76372 40010 76428 40012
rect 76476 40010 76532 40012
rect 76372 39958 76396 40010
rect 76396 39958 76428 40010
rect 76476 39958 76520 40010
rect 76520 39958 76532 40010
rect 76372 39956 76428 39958
rect 76476 39956 76532 39958
rect 76580 39956 76636 40012
rect 76684 40010 76740 40012
rect 76788 40010 76844 40012
rect 76684 39958 76696 40010
rect 76696 39958 76740 40010
rect 76788 39958 76820 40010
rect 76820 39958 76844 40010
rect 76684 39956 76740 39958
rect 76788 39956 76844 39958
rect 76892 39956 76948 40012
rect 77980 42028 78036 42084
rect 77868 41858 77924 41860
rect 77868 41806 77870 41858
rect 77870 41806 77922 41858
rect 77922 41806 77924 41858
rect 77868 41804 77924 41806
rect 80768 50148 80824 50204
rect 80872 50202 80928 50204
rect 80976 50202 81032 50204
rect 80872 50150 80896 50202
rect 80896 50150 80928 50202
rect 80976 50150 81020 50202
rect 81020 50150 81032 50202
rect 80872 50148 80928 50150
rect 80976 50148 81032 50150
rect 81080 50148 81136 50204
rect 81184 50202 81240 50204
rect 81288 50202 81344 50204
rect 81184 50150 81196 50202
rect 81196 50150 81240 50202
rect 81288 50150 81320 50202
rect 81320 50150 81344 50202
rect 81184 50148 81240 50150
rect 81288 50148 81344 50150
rect 81392 50148 81448 50204
rect 85268 49364 85324 49420
rect 85372 49418 85428 49420
rect 85476 49418 85532 49420
rect 85372 49366 85396 49418
rect 85396 49366 85428 49418
rect 85476 49366 85520 49418
rect 85520 49366 85532 49418
rect 85372 49364 85428 49366
rect 85476 49364 85532 49366
rect 85580 49364 85636 49420
rect 85684 49418 85740 49420
rect 85788 49418 85844 49420
rect 85684 49366 85696 49418
rect 85696 49366 85740 49418
rect 85788 49366 85820 49418
rect 85820 49366 85844 49418
rect 85684 49364 85740 49366
rect 85788 49364 85844 49366
rect 85892 49364 85948 49420
rect 85036 48914 85092 48916
rect 85036 48862 85038 48914
rect 85038 48862 85090 48914
rect 85090 48862 85092 48914
rect 85036 48860 85092 48862
rect 79548 48188 79604 48244
rect 85820 49026 85876 49028
rect 85820 48974 85822 49026
rect 85822 48974 85874 49026
rect 85874 48974 85876 49026
rect 85820 48972 85876 48974
rect 89768 50148 89824 50204
rect 89872 50202 89928 50204
rect 89976 50202 90032 50204
rect 89872 50150 89896 50202
rect 89896 50150 89928 50202
rect 89976 50150 90020 50202
rect 90020 50150 90032 50202
rect 89872 50148 89928 50150
rect 89976 50148 90032 50150
rect 90080 50148 90136 50204
rect 90184 50202 90240 50204
rect 90288 50202 90344 50204
rect 90184 50150 90196 50202
rect 90196 50150 90240 50202
rect 90288 50150 90320 50202
rect 90320 50150 90344 50202
rect 90184 50148 90240 50150
rect 90288 50148 90344 50150
rect 90392 50148 90448 50204
rect 90524 49644 90580 49700
rect 94268 50932 94324 50988
rect 94372 50986 94428 50988
rect 94476 50986 94532 50988
rect 94372 50934 94396 50986
rect 94396 50934 94428 50986
rect 94476 50934 94520 50986
rect 94520 50934 94532 50986
rect 94372 50932 94428 50934
rect 94476 50932 94532 50934
rect 94580 50932 94636 50988
rect 94684 50986 94740 50988
rect 94788 50986 94844 50988
rect 94684 50934 94696 50986
rect 94696 50934 94740 50986
rect 94788 50934 94820 50986
rect 94820 50934 94844 50986
rect 94684 50932 94740 50934
rect 94788 50932 94844 50934
rect 94892 50932 94948 50988
rect 92428 49698 92484 49700
rect 92428 49646 92430 49698
rect 92430 49646 92482 49698
rect 92482 49646 92484 49698
rect 92428 49644 92484 49646
rect 95452 49644 95508 49700
rect 94268 49364 94324 49420
rect 94372 49418 94428 49420
rect 94476 49418 94532 49420
rect 94372 49366 94396 49418
rect 94396 49366 94428 49418
rect 94476 49366 94520 49418
rect 94520 49366 94532 49418
rect 94372 49364 94428 49366
rect 94476 49364 94532 49366
rect 94580 49364 94636 49420
rect 94684 49418 94740 49420
rect 94788 49418 94844 49420
rect 94684 49366 94696 49418
rect 94696 49366 94740 49418
rect 94788 49366 94820 49418
rect 94820 49366 94844 49418
rect 94684 49364 94740 49366
rect 94788 49364 94844 49366
rect 94892 49364 94948 49420
rect 90748 49196 90804 49252
rect 90188 49026 90244 49028
rect 90188 48974 90190 49026
rect 90190 48974 90242 49026
rect 90242 48974 90244 49026
rect 90188 48972 90244 48974
rect 89628 48860 89684 48916
rect 90524 48860 90580 48916
rect 80768 48580 80824 48636
rect 80872 48634 80928 48636
rect 80976 48634 81032 48636
rect 80872 48582 80896 48634
rect 80896 48582 80928 48634
rect 80976 48582 81020 48634
rect 81020 48582 81032 48634
rect 80872 48580 80928 48582
rect 80976 48580 81032 48582
rect 81080 48580 81136 48636
rect 81184 48634 81240 48636
rect 81288 48634 81344 48636
rect 81184 48582 81196 48634
rect 81196 48582 81240 48634
rect 81288 48582 81320 48634
rect 81320 48582 81344 48634
rect 81184 48580 81240 48582
rect 81288 48580 81344 48582
rect 81392 48580 81448 48636
rect 80556 48242 80612 48244
rect 80556 48190 80558 48242
rect 80558 48190 80610 48242
rect 80610 48190 80612 48242
rect 80556 48188 80612 48190
rect 80768 47012 80824 47068
rect 80872 47066 80928 47068
rect 80976 47066 81032 47068
rect 80872 47014 80896 47066
rect 80896 47014 80928 47066
rect 80976 47014 81020 47066
rect 81020 47014 81032 47066
rect 80872 47012 80928 47014
rect 80976 47012 81032 47014
rect 81080 47012 81136 47068
rect 81184 47066 81240 47068
rect 81288 47066 81344 47068
rect 81184 47014 81196 47066
rect 81196 47014 81240 47066
rect 81288 47014 81320 47066
rect 81320 47014 81344 47066
rect 81184 47012 81240 47014
rect 81288 47012 81344 47014
rect 81392 47012 81448 47068
rect 79100 46002 79156 46004
rect 79100 45950 79102 46002
rect 79102 45950 79154 46002
rect 79154 45950 79156 46002
rect 79100 45948 79156 45950
rect 79548 45948 79604 46004
rect 78652 45724 78708 45780
rect 78316 45612 78372 45668
rect 79324 45778 79380 45780
rect 79324 45726 79326 45778
rect 79326 45726 79378 45778
rect 79378 45726 79380 45778
rect 79324 45724 79380 45726
rect 78316 44210 78372 44212
rect 78316 44158 78318 44210
rect 78318 44158 78370 44210
rect 78370 44158 78372 44210
rect 78316 44156 78372 44158
rect 78204 41916 78260 41972
rect 79100 42082 79156 42084
rect 79100 42030 79102 42082
rect 79102 42030 79154 42082
rect 79154 42030 79156 42082
rect 79100 42028 79156 42030
rect 78652 41356 78708 41412
rect 77644 40962 77700 40964
rect 77644 40910 77646 40962
rect 77646 40910 77698 40962
rect 77698 40910 77700 40962
rect 77644 40908 77700 40910
rect 78540 40908 78596 40964
rect 77196 39004 77252 39060
rect 76860 38722 76916 38724
rect 76860 38670 76862 38722
rect 76862 38670 76914 38722
rect 76914 38670 76916 38722
rect 76860 38668 76916 38670
rect 77196 38668 77252 38724
rect 76268 38388 76324 38444
rect 76372 38442 76428 38444
rect 76476 38442 76532 38444
rect 76372 38390 76396 38442
rect 76396 38390 76428 38442
rect 76476 38390 76520 38442
rect 76520 38390 76532 38442
rect 76372 38388 76428 38390
rect 76476 38388 76532 38390
rect 76580 38388 76636 38444
rect 76684 38442 76740 38444
rect 76788 38442 76844 38444
rect 76684 38390 76696 38442
rect 76696 38390 76740 38442
rect 76788 38390 76820 38442
rect 76820 38390 76844 38442
rect 76684 38388 76740 38390
rect 76788 38388 76844 38390
rect 76892 38388 76948 38444
rect 77196 38220 77252 38276
rect 77420 38892 77476 38948
rect 77756 40402 77812 40404
rect 77756 40350 77758 40402
rect 77758 40350 77810 40402
rect 77810 40350 77812 40402
rect 77756 40348 77812 40350
rect 78092 40290 78148 40292
rect 78092 40238 78094 40290
rect 78094 40238 78146 40290
rect 78146 40238 78148 40290
rect 78092 40236 78148 40238
rect 77756 39788 77812 39844
rect 77756 39004 77812 39060
rect 76188 37772 76244 37828
rect 76300 37938 76356 37940
rect 76300 37886 76302 37938
rect 76302 37886 76354 37938
rect 76354 37886 76356 37938
rect 76300 37884 76356 37886
rect 77532 37772 77588 37828
rect 76860 37490 76916 37492
rect 76860 37438 76862 37490
rect 76862 37438 76914 37490
rect 76914 37438 76916 37490
rect 76860 37436 76916 37438
rect 77532 37436 77588 37492
rect 76188 37154 76244 37156
rect 76188 37102 76190 37154
rect 76190 37102 76242 37154
rect 76242 37102 76244 37154
rect 76188 37100 76244 37102
rect 75740 36876 75796 36932
rect 78540 39058 78596 39060
rect 78540 39006 78542 39058
rect 78542 39006 78594 39058
rect 78594 39006 78596 39058
rect 78540 39004 78596 39006
rect 77868 38668 77924 38724
rect 82796 45948 82852 46004
rect 79884 45890 79940 45892
rect 79884 45838 79886 45890
rect 79886 45838 79938 45890
rect 79938 45838 79940 45890
rect 79884 45836 79940 45838
rect 80556 45836 80612 45892
rect 80768 45444 80824 45500
rect 80872 45498 80928 45500
rect 80976 45498 81032 45500
rect 80872 45446 80896 45498
rect 80896 45446 80928 45498
rect 80976 45446 81020 45498
rect 81020 45446 81032 45498
rect 80872 45444 80928 45446
rect 80976 45444 81032 45446
rect 81080 45444 81136 45500
rect 81184 45498 81240 45500
rect 81288 45498 81344 45500
rect 81184 45446 81196 45498
rect 81196 45446 81240 45498
rect 81288 45446 81320 45498
rect 81320 45446 81344 45498
rect 81184 45444 81240 45446
rect 81288 45444 81344 45446
rect 81392 45444 81448 45500
rect 79772 44210 79828 44212
rect 79772 44158 79774 44210
rect 79774 44158 79826 44210
rect 79826 44158 79828 44210
rect 79772 44156 79828 44158
rect 80108 43708 80164 43764
rect 80768 43876 80824 43932
rect 80872 43930 80928 43932
rect 80976 43930 81032 43932
rect 80872 43878 80896 43930
rect 80896 43878 80928 43930
rect 80976 43878 81020 43930
rect 81020 43878 81032 43930
rect 80872 43876 80928 43878
rect 80976 43876 81032 43878
rect 81080 43876 81136 43932
rect 81184 43930 81240 43932
rect 81288 43930 81344 43932
rect 81184 43878 81196 43930
rect 81196 43878 81240 43930
rect 81288 43878 81320 43930
rect 81320 43878 81344 43930
rect 81184 43876 81240 43878
rect 81288 43876 81344 43878
rect 81392 43876 81448 43932
rect 81340 43708 81396 43764
rect 83692 48354 83748 48356
rect 83692 48302 83694 48354
rect 83694 48302 83746 48354
rect 83746 48302 83748 48354
rect 83692 48300 83748 48302
rect 85148 48188 85204 48244
rect 85268 47796 85324 47852
rect 85372 47850 85428 47852
rect 85476 47850 85532 47852
rect 85372 47798 85396 47850
rect 85396 47798 85428 47850
rect 85476 47798 85520 47850
rect 85520 47798 85532 47850
rect 85372 47796 85428 47798
rect 85476 47796 85532 47798
rect 85580 47796 85636 47852
rect 85684 47850 85740 47852
rect 85788 47850 85844 47852
rect 85684 47798 85696 47850
rect 85696 47798 85740 47850
rect 85788 47798 85820 47850
rect 85820 47798 85844 47850
rect 85684 47796 85740 47798
rect 85788 47796 85844 47798
rect 85892 47796 85948 47852
rect 85484 46396 85540 46452
rect 85268 46228 85324 46284
rect 85372 46282 85428 46284
rect 85476 46282 85532 46284
rect 85372 46230 85396 46282
rect 85396 46230 85428 46282
rect 85476 46230 85520 46282
rect 85520 46230 85532 46282
rect 85372 46228 85428 46230
rect 85476 46228 85532 46230
rect 85580 46228 85636 46284
rect 85684 46282 85740 46284
rect 85788 46282 85844 46284
rect 85684 46230 85696 46282
rect 85696 46230 85740 46282
rect 85788 46230 85820 46282
rect 85820 46230 85844 46282
rect 85684 46228 85740 46230
rect 85788 46228 85844 46230
rect 85892 46228 85948 46284
rect 86380 46396 86436 46452
rect 89768 48580 89824 48636
rect 89872 48634 89928 48636
rect 89976 48634 90032 48636
rect 89872 48582 89896 48634
rect 89896 48582 89928 48634
rect 89976 48582 90020 48634
rect 90020 48582 90032 48634
rect 89872 48580 89928 48582
rect 89976 48580 90032 48582
rect 90080 48580 90136 48636
rect 90184 48634 90240 48636
rect 90288 48634 90344 48636
rect 90184 48582 90196 48634
rect 90196 48582 90240 48634
rect 90288 48582 90320 48634
rect 90320 48582 90344 48634
rect 90184 48580 90240 48582
rect 90288 48580 90344 48582
rect 90392 48580 90448 48636
rect 91196 48242 91252 48244
rect 91196 48190 91198 48242
rect 91198 48190 91250 48242
rect 91250 48190 91252 48242
rect 91196 48188 91252 48190
rect 89768 47012 89824 47068
rect 89872 47066 89928 47068
rect 89976 47066 90032 47068
rect 89872 47014 89896 47066
rect 89896 47014 89928 47066
rect 89976 47014 90020 47066
rect 90020 47014 90032 47066
rect 89872 47012 89928 47014
rect 89976 47012 90032 47014
rect 90080 47012 90136 47068
rect 90184 47066 90240 47068
rect 90288 47066 90344 47068
rect 90184 47014 90196 47066
rect 90196 47014 90240 47066
rect 90288 47014 90320 47066
rect 90320 47014 90344 47066
rect 90184 47012 90240 47014
rect 90288 47012 90344 47014
rect 90392 47012 90448 47068
rect 83580 45666 83636 45668
rect 83580 45614 83582 45666
rect 83582 45614 83634 45666
rect 83634 45614 83636 45666
rect 83580 45612 83636 45614
rect 86940 46450 86996 46452
rect 86940 46398 86942 46450
rect 86942 46398 86994 46450
rect 86994 46398 86996 46450
rect 86940 46396 86996 46398
rect 89628 46396 89684 46452
rect 89628 45724 89684 45780
rect 89068 45666 89124 45668
rect 89068 45614 89070 45666
rect 89070 45614 89122 45666
rect 89122 45614 89124 45666
rect 89068 45612 89124 45614
rect 89964 45612 90020 45668
rect 89768 45444 89824 45500
rect 89872 45498 89928 45500
rect 89976 45498 90032 45500
rect 89872 45446 89896 45498
rect 89896 45446 89928 45498
rect 89976 45446 90020 45498
rect 90020 45446 90032 45498
rect 89872 45444 89928 45446
rect 89976 45444 90032 45446
rect 90080 45444 90136 45500
rect 90184 45498 90240 45500
rect 90288 45498 90344 45500
rect 90184 45446 90196 45498
rect 90196 45446 90240 45498
rect 90288 45446 90320 45498
rect 90320 45446 90344 45498
rect 90184 45444 90240 45446
rect 90288 45444 90344 45446
rect 90392 45444 90448 45500
rect 86716 45164 86772 45220
rect 92316 48242 92372 48244
rect 92316 48190 92318 48242
rect 92318 48190 92370 48242
rect 92370 48190 92372 48242
rect 92316 48188 92372 48190
rect 91644 47628 91700 47684
rect 92540 47628 92596 47684
rect 92652 47458 92708 47460
rect 92652 47406 92654 47458
rect 92654 47406 92706 47458
rect 92706 47406 92708 47458
rect 92652 47404 92708 47406
rect 93100 48636 93156 48692
rect 96236 48636 96292 48692
rect 94268 47796 94324 47852
rect 94372 47850 94428 47852
rect 94476 47850 94532 47852
rect 94372 47798 94396 47850
rect 94396 47798 94428 47850
rect 94476 47798 94520 47850
rect 94520 47798 94532 47850
rect 94372 47796 94428 47798
rect 94476 47796 94532 47798
rect 94580 47796 94636 47852
rect 94684 47850 94740 47852
rect 94788 47850 94844 47852
rect 94684 47798 94696 47850
rect 94696 47798 94740 47850
rect 94788 47798 94820 47850
rect 94820 47798 94844 47850
rect 94684 47796 94740 47798
rect 94788 47796 94844 47798
rect 94892 47796 94948 47852
rect 93436 47404 93492 47460
rect 91980 46732 92036 46788
rect 91868 46674 91924 46676
rect 91868 46622 91870 46674
rect 91870 46622 91922 46674
rect 91922 46622 91924 46674
rect 91868 46620 91924 46622
rect 92540 46786 92596 46788
rect 92540 46734 92542 46786
rect 92542 46734 92594 46786
rect 92594 46734 92596 46786
rect 92540 46732 92596 46734
rect 92876 46620 92932 46676
rect 91308 45500 91364 45556
rect 92540 45612 92596 45668
rect 91196 45330 91252 45332
rect 91196 45278 91198 45330
rect 91198 45278 91250 45330
rect 91250 45278 91252 45330
rect 91196 45276 91252 45278
rect 91980 45276 92036 45332
rect 90636 45218 90692 45220
rect 90636 45166 90638 45218
rect 90638 45166 90690 45218
rect 90690 45166 90692 45218
rect 90636 45164 90692 45166
rect 85268 44660 85324 44716
rect 85372 44714 85428 44716
rect 85476 44714 85532 44716
rect 85372 44662 85396 44714
rect 85396 44662 85428 44714
rect 85476 44662 85520 44714
rect 85520 44662 85532 44714
rect 85372 44660 85428 44662
rect 85476 44660 85532 44662
rect 85580 44660 85636 44716
rect 85684 44714 85740 44716
rect 85788 44714 85844 44716
rect 85684 44662 85696 44714
rect 85696 44662 85740 44714
rect 85788 44662 85820 44714
rect 85820 44662 85844 44714
rect 85684 44660 85740 44662
rect 85788 44660 85844 44662
rect 85892 44660 85948 44716
rect 89768 43876 89824 43932
rect 89872 43930 89928 43932
rect 89976 43930 90032 43932
rect 89872 43878 89896 43930
rect 89896 43878 89928 43930
rect 89976 43878 90020 43930
rect 90020 43878 90032 43930
rect 89872 43876 89928 43878
rect 89976 43876 90032 43878
rect 90080 43876 90136 43932
rect 90184 43930 90240 43932
rect 90288 43930 90344 43932
rect 90184 43878 90196 43930
rect 90196 43878 90240 43930
rect 90288 43878 90320 43930
rect 90320 43878 90344 43930
rect 90184 43876 90240 43878
rect 90288 43876 90344 43878
rect 90392 43876 90448 43932
rect 88396 43708 88452 43764
rect 80768 42308 80824 42364
rect 80872 42362 80928 42364
rect 80976 42362 81032 42364
rect 80872 42310 80896 42362
rect 80896 42310 80928 42362
rect 80976 42310 81020 42362
rect 81020 42310 81032 42362
rect 80872 42308 80928 42310
rect 80976 42308 81032 42310
rect 81080 42308 81136 42364
rect 81184 42362 81240 42364
rect 81288 42362 81344 42364
rect 81184 42310 81196 42362
rect 81196 42310 81240 42362
rect 81288 42310 81320 42362
rect 81320 42310 81344 42362
rect 81184 42308 81240 42310
rect 81288 42308 81344 42310
rect 81392 42308 81448 42364
rect 80556 41916 80612 41972
rect 80892 41916 80948 41972
rect 81676 41916 81732 41972
rect 81564 41410 81620 41412
rect 81564 41358 81566 41410
rect 81566 41358 81618 41410
rect 81618 41358 81620 41410
rect 81564 41356 81620 41358
rect 80892 40962 80948 40964
rect 80892 40910 80894 40962
rect 80894 40910 80946 40962
rect 80946 40910 80948 40962
rect 80892 40908 80948 40910
rect 80768 40740 80824 40796
rect 80872 40794 80928 40796
rect 80976 40794 81032 40796
rect 80872 40742 80896 40794
rect 80896 40742 80928 40794
rect 80976 40742 81020 40794
rect 81020 40742 81032 40794
rect 80872 40740 80928 40742
rect 80976 40740 81032 40742
rect 81080 40740 81136 40796
rect 81184 40794 81240 40796
rect 81288 40794 81344 40796
rect 81184 40742 81196 40794
rect 81196 40742 81240 40794
rect 81288 40742 81320 40794
rect 81320 40742 81344 40794
rect 81184 40740 81240 40742
rect 81288 40740 81344 40742
rect 81392 40740 81448 40796
rect 80768 39172 80824 39228
rect 80872 39226 80928 39228
rect 80976 39226 81032 39228
rect 80872 39174 80896 39226
rect 80896 39174 80928 39226
rect 80976 39174 81020 39226
rect 81020 39174 81032 39226
rect 80872 39172 80928 39174
rect 80976 39172 81032 39174
rect 81080 39172 81136 39228
rect 81184 39226 81240 39228
rect 81288 39226 81344 39228
rect 81184 39174 81196 39226
rect 81196 39174 81240 39226
rect 81288 39174 81320 39226
rect 81320 39174 81344 39226
rect 81184 39172 81240 39174
rect 81288 39172 81344 39174
rect 81392 39172 81448 39228
rect 79548 38668 79604 38724
rect 78316 37772 78372 37828
rect 78540 37996 78596 38052
rect 79324 38050 79380 38052
rect 79324 37998 79326 38050
rect 79326 37998 79378 38050
rect 79378 37998 79380 38050
rect 79324 37996 79380 37998
rect 84476 43650 84532 43652
rect 84476 43598 84478 43650
rect 84478 43598 84530 43650
rect 84530 43598 84532 43650
rect 84476 43596 84532 43598
rect 85268 43092 85324 43148
rect 85372 43146 85428 43148
rect 85476 43146 85532 43148
rect 85372 43094 85396 43146
rect 85396 43094 85428 43146
rect 85476 43094 85520 43146
rect 85520 43094 85532 43146
rect 85372 43092 85428 43094
rect 85476 43092 85532 43094
rect 85580 43092 85636 43148
rect 85684 43146 85740 43148
rect 85788 43146 85844 43148
rect 85684 43094 85696 43146
rect 85696 43094 85740 43146
rect 85788 43094 85820 43146
rect 85820 43094 85844 43146
rect 85684 43092 85740 43094
rect 85788 43092 85844 43094
rect 85892 43092 85948 43148
rect 83468 41916 83524 41972
rect 87164 41970 87220 41972
rect 87164 41918 87166 41970
rect 87166 41918 87218 41970
rect 87218 41918 87220 41970
rect 87164 41916 87220 41918
rect 85268 41524 85324 41580
rect 85372 41578 85428 41580
rect 85476 41578 85532 41580
rect 85372 41526 85396 41578
rect 85396 41526 85428 41578
rect 85476 41526 85520 41578
rect 85520 41526 85532 41578
rect 85372 41524 85428 41526
rect 85476 41524 85532 41526
rect 85580 41524 85636 41580
rect 85684 41578 85740 41580
rect 85788 41578 85844 41580
rect 85684 41526 85696 41578
rect 85696 41526 85740 41578
rect 85788 41526 85820 41578
rect 85820 41526 85844 41578
rect 85684 41524 85740 41526
rect 85788 41524 85844 41526
rect 85892 41524 85948 41580
rect 84140 40684 84196 40740
rect 82124 39730 82180 39732
rect 82124 39678 82126 39730
rect 82126 39678 82178 39730
rect 82178 39678 82180 39730
rect 82124 39676 82180 39678
rect 83020 39618 83076 39620
rect 83020 39566 83022 39618
rect 83022 39566 83074 39618
rect 83074 39566 83076 39618
rect 83020 39564 83076 39566
rect 83916 39618 83972 39620
rect 83916 39566 83918 39618
rect 83918 39566 83970 39618
rect 83970 39566 83972 39618
rect 83916 39564 83972 39566
rect 84924 39618 84980 39620
rect 84924 39566 84926 39618
rect 84926 39566 84978 39618
rect 84978 39566 84980 39618
rect 84924 39564 84980 39566
rect 85372 40626 85428 40628
rect 85372 40574 85374 40626
rect 85374 40574 85426 40626
rect 85426 40574 85428 40626
rect 85372 40572 85428 40574
rect 85932 40626 85988 40628
rect 85932 40574 85934 40626
rect 85934 40574 85986 40626
rect 85986 40574 85988 40626
rect 85932 40572 85988 40574
rect 86268 40514 86324 40516
rect 86268 40462 86270 40514
rect 86270 40462 86322 40514
rect 86322 40462 86324 40514
rect 86268 40460 86324 40462
rect 86828 40460 86884 40516
rect 85268 39956 85324 40012
rect 85372 40010 85428 40012
rect 85476 40010 85532 40012
rect 85372 39958 85396 40010
rect 85396 39958 85428 40010
rect 85476 39958 85520 40010
rect 85520 39958 85532 40010
rect 85372 39956 85428 39958
rect 85476 39956 85532 39958
rect 85580 39956 85636 40012
rect 85684 40010 85740 40012
rect 85788 40010 85844 40012
rect 85684 39958 85696 40010
rect 85696 39958 85740 40010
rect 85788 39958 85820 40010
rect 85820 39958 85844 40010
rect 85684 39956 85740 39958
rect 85788 39956 85844 39958
rect 85892 39956 85948 40012
rect 82684 39004 82740 39060
rect 83468 39004 83524 39060
rect 83916 38892 83972 38948
rect 82460 37826 82516 37828
rect 82460 37774 82462 37826
rect 82462 37774 82514 37826
rect 82514 37774 82516 37826
rect 82460 37772 82516 37774
rect 83468 37826 83524 37828
rect 83468 37774 83470 37826
rect 83470 37774 83522 37826
rect 83522 37774 83524 37826
rect 83468 37772 83524 37774
rect 80768 37604 80824 37660
rect 80872 37658 80928 37660
rect 80976 37658 81032 37660
rect 80872 37606 80896 37658
rect 80896 37606 80928 37658
rect 80976 37606 81020 37658
rect 81020 37606 81032 37658
rect 80872 37604 80928 37606
rect 80976 37604 81032 37606
rect 81080 37604 81136 37660
rect 81184 37658 81240 37660
rect 81288 37658 81344 37660
rect 81184 37606 81196 37658
rect 81196 37606 81240 37658
rect 81288 37606 81320 37658
rect 81320 37606 81344 37658
rect 81184 37604 81240 37606
rect 81288 37604 81344 37606
rect 81392 37604 81448 37660
rect 83468 37324 83524 37380
rect 84364 39452 84420 39508
rect 84812 39506 84868 39508
rect 84812 39454 84814 39506
rect 84814 39454 84866 39506
rect 84866 39454 84868 39506
rect 84812 39452 84868 39454
rect 84476 39004 84532 39060
rect 84140 37884 84196 37940
rect 84252 37826 84308 37828
rect 84252 37774 84254 37826
rect 84254 37774 84306 37826
rect 84306 37774 84308 37826
rect 84252 37772 84308 37774
rect 85820 39394 85876 39396
rect 85820 39342 85822 39394
rect 85822 39342 85874 39394
rect 85874 39342 85876 39394
rect 85820 39340 85876 39342
rect 85260 39058 85316 39060
rect 85260 39006 85262 39058
rect 85262 39006 85314 39058
rect 85314 39006 85316 39058
rect 85260 39004 85316 39006
rect 84700 38946 84756 38948
rect 84700 38894 84702 38946
rect 84702 38894 84754 38946
rect 84754 38894 84756 38946
rect 84700 38892 84756 38894
rect 85268 38388 85324 38444
rect 85372 38442 85428 38444
rect 85476 38442 85532 38444
rect 85372 38390 85396 38442
rect 85396 38390 85428 38442
rect 85476 38390 85520 38442
rect 85520 38390 85532 38442
rect 85372 38388 85428 38390
rect 85476 38388 85532 38390
rect 85580 38388 85636 38444
rect 85684 38442 85740 38444
rect 85788 38442 85844 38444
rect 85684 38390 85696 38442
rect 85696 38390 85740 38442
rect 85788 38390 85820 38442
rect 85820 38390 85844 38442
rect 85684 38388 85740 38390
rect 85788 38388 85844 38390
rect 85892 38388 85948 38444
rect 77756 37100 77812 37156
rect 76268 36820 76324 36876
rect 76372 36874 76428 36876
rect 76476 36874 76532 36876
rect 76372 36822 76396 36874
rect 76396 36822 76428 36874
rect 76476 36822 76520 36874
rect 76520 36822 76532 36874
rect 76372 36820 76428 36822
rect 76476 36820 76532 36822
rect 76580 36820 76636 36876
rect 76684 36874 76740 36876
rect 76788 36874 76844 36876
rect 76684 36822 76696 36874
rect 76696 36822 76740 36874
rect 76788 36822 76820 36874
rect 76820 36822 76844 36874
rect 76684 36820 76740 36822
rect 76788 36820 76844 36822
rect 76892 36820 76948 36876
rect 77196 36594 77252 36596
rect 77196 36542 77198 36594
rect 77198 36542 77250 36594
rect 77250 36542 77252 36594
rect 77196 36540 77252 36542
rect 76268 35252 76324 35308
rect 76372 35306 76428 35308
rect 76476 35306 76532 35308
rect 76372 35254 76396 35306
rect 76396 35254 76428 35306
rect 76476 35254 76520 35306
rect 76520 35254 76532 35306
rect 76372 35252 76428 35254
rect 76476 35252 76532 35254
rect 76580 35252 76636 35308
rect 76684 35306 76740 35308
rect 76788 35306 76844 35308
rect 76684 35254 76696 35306
rect 76696 35254 76740 35306
rect 76788 35254 76820 35306
rect 76820 35254 76844 35306
rect 76684 35252 76740 35254
rect 76788 35252 76844 35254
rect 76892 35252 76948 35308
rect 84252 36652 84308 36708
rect 77980 36428 78036 36484
rect 81564 36316 81620 36372
rect 78428 36204 78484 36260
rect 78988 36258 79044 36260
rect 78988 36206 78990 36258
rect 78990 36206 79042 36258
rect 79042 36206 79044 36258
rect 78988 36204 79044 36206
rect 80768 36036 80824 36092
rect 80872 36090 80928 36092
rect 80976 36090 81032 36092
rect 80872 36038 80896 36090
rect 80896 36038 80928 36090
rect 80976 36038 81020 36090
rect 81020 36038 81032 36090
rect 80872 36036 80928 36038
rect 80976 36036 81032 36038
rect 81080 36036 81136 36092
rect 81184 36090 81240 36092
rect 81288 36090 81344 36092
rect 81184 36038 81196 36090
rect 81196 36038 81240 36090
rect 81288 36038 81320 36090
rect 81320 36038 81344 36090
rect 81184 36036 81240 36038
rect 81288 36036 81344 36038
rect 81392 36036 81448 36092
rect 78428 35922 78484 35924
rect 78428 35870 78430 35922
rect 78430 35870 78482 35922
rect 78482 35870 78484 35922
rect 78428 35868 78484 35870
rect 78876 35698 78932 35700
rect 78876 35646 78878 35698
rect 78878 35646 78930 35698
rect 78930 35646 78932 35698
rect 78876 35644 78932 35646
rect 78092 35308 78148 35364
rect 80220 35810 80276 35812
rect 80220 35758 80222 35810
rect 80222 35758 80274 35810
rect 80274 35758 80276 35810
rect 80220 35756 80276 35758
rect 84812 36204 84868 36260
rect 81564 35756 81620 35812
rect 79996 35698 80052 35700
rect 79996 35646 79998 35698
rect 79998 35646 80050 35698
rect 80050 35646 80052 35698
rect 79996 35644 80052 35646
rect 80332 35420 80388 35476
rect 79100 35308 79156 35364
rect 80780 35308 80836 35364
rect 84588 35644 84644 35700
rect 84924 37772 84980 37828
rect 85484 37772 85540 37828
rect 85932 37826 85988 37828
rect 85932 37774 85934 37826
rect 85934 37774 85986 37826
rect 85986 37774 85988 37826
rect 85932 37772 85988 37774
rect 91084 45164 91140 45220
rect 91756 45164 91812 45220
rect 96012 46620 96068 46676
rect 94268 46228 94324 46284
rect 94372 46282 94428 46284
rect 94476 46282 94532 46284
rect 94372 46230 94396 46282
rect 94396 46230 94428 46282
rect 94476 46230 94520 46282
rect 94520 46230 94532 46282
rect 94372 46228 94428 46230
rect 94476 46228 94532 46230
rect 94580 46228 94636 46284
rect 94684 46282 94740 46284
rect 94788 46282 94844 46284
rect 94684 46230 94696 46282
rect 94696 46230 94740 46282
rect 94788 46230 94820 46282
rect 94820 46230 94844 46282
rect 94684 46228 94740 46230
rect 94788 46228 94844 46230
rect 94892 46228 94948 46284
rect 95676 45666 95732 45668
rect 95676 45614 95678 45666
rect 95678 45614 95730 45666
rect 95730 45614 95732 45666
rect 95676 45612 95732 45614
rect 95004 45500 95060 45556
rect 94268 44660 94324 44716
rect 94372 44714 94428 44716
rect 94476 44714 94532 44716
rect 94372 44662 94396 44714
rect 94396 44662 94428 44714
rect 94476 44662 94520 44714
rect 94520 44662 94532 44714
rect 94372 44660 94428 44662
rect 94476 44660 94532 44662
rect 94580 44660 94636 44716
rect 94684 44714 94740 44716
rect 94788 44714 94844 44716
rect 94684 44662 94696 44714
rect 94696 44662 94740 44714
rect 94788 44662 94820 44714
rect 94820 44662 94844 44714
rect 94684 44660 94740 44662
rect 94788 44660 94844 44662
rect 94892 44660 94948 44716
rect 90860 43708 90916 43764
rect 88844 42476 88900 42532
rect 90076 42530 90132 42532
rect 90076 42478 90078 42530
rect 90078 42478 90130 42530
rect 90130 42478 90132 42530
rect 90076 42476 90132 42478
rect 89768 42308 89824 42364
rect 89872 42362 89928 42364
rect 89976 42362 90032 42364
rect 89872 42310 89896 42362
rect 89896 42310 89928 42362
rect 89976 42310 90020 42362
rect 90020 42310 90032 42362
rect 89872 42308 89928 42310
rect 89976 42308 90032 42310
rect 90080 42308 90136 42364
rect 90184 42362 90240 42364
rect 90288 42362 90344 42364
rect 90184 42310 90196 42362
rect 90196 42310 90240 42362
rect 90288 42310 90320 42362
rect 90320 42310 90344 42362
rect 90184 42308 90240 42310
rect 90288 42308 90344 42310
rect 90392 42308 90448 42364
rect 89180 41970 89236 41972
rect 89180 41918 89182 41970
rect 89182 41918 89234 41970
rect 89234 41918 89236 41970
rect 89180 41916 89236 41918
rect 89768 40740 89824 40796
rect 89872 40794 89928 40796
rect 89976 40794 90032 40796
rect 89872 40742 89896 40794
rect 89896 40742 89928 40794
rect 89976 40742 90020 40794
rect 90020 40742 90032 40794
rect 89872 40740 89928 40742
rect 89976 40740 90032 40742
rect 90080 40740 90136 40796
rect 90184 40794 90240 40796
rect 90288 40794 90344 40796
rect 90184 40742 90196 40794
rect 90196 40742 90240 40794
rect 90288 40742 90320 40794
rect 90320 40742 90344 40794
rect 90184 40740 90240 40742
rect 90288 40740 90344 40742
rect 90392 40740 90448 40796
rect 92316 43708 92372 43764
rect 87500 40236 87556 40292
rect 89516 40460 89572 40516
rect 87164 39618 87220 39620
rect 87164 39566 87166 39618
rect 87166 39566 87218 39618
rect 87218 39566 87220 39618
rect 87164 39564 87220 39566
rect 90748 40460 90804 40516
rect 89068 38892 89124 38948
rect 87164 38556 87220 38612
rect 89068 38108 89124 38164
rect 87500 38050 87556 38052
rect 87500 37998 87502 38050
rect 87502 37998 87554 38050
rect 87554 37998 87556 38050
rect 87500 37996 87556 37998
rect 86828 37490 86884 37492
rect 86828 37438 86830 37490
rect 86830 37438 86882 37490
rect 86882 37438 86884 37490
rect 86828 37436 86884 37438
rect 88060 37490 88116 37492
rect 88060 37438 88062 37490
rect 88062 37438 88114 37490
rect 88114 37438 88116 37490
rect 88060 37436 88116 37438
rect 90300 39394 90356 39396
rect 90300 39342 90302 39394
rect 90302 39342 90354 39394
rect 90354 39342 90356 39394
rect 90300 39340 90356 39342
rect 89768 39172 89824 39228
rect 89872 39226 89928 39228
rect 89976 39226 90032 39228
rect 89872 39174 89896 39226
rect 89896 39174 89928 39226
rect 89976 39174 90020 39226
rect 90020 39174 90032 39226
rect 89872 39172 89928 39174
rect 89976 39172 90032 39174
rect 90080 39172 90136 39228
rect 90184 39226 90240 39228
rect 90288 39226 90344 39228
rect 90184 39174 90196 39226
rect 90196 39174 90240 39226
rect 90288 39174 90320 39226
rect 90320 39174 90344 39226
rect 90184 39172 90240 39174
rect 90288 39172 90344 39174
rect 90392 39172 90448 39228
rect 89740 39058 89796 39060
rect 89740 39006 89742 39058
rect 89742 39006 89794 39058
rect 89794 39006 89796 39058
rect 89740 39004 89796 39006
rect 90972 43426 91028 43428
rect 90972 43374 90974 43426
rect 90974 43374 91026 43426
rect 91026 43374 91028 43426
rect 90972 43372 91028 43374
rect 94556 43372 94612 43428
rect 94268 43092 94324 43148
rect 94372 43146 94428 43148
rect 94476 43146 94532 43148
rect 94372 43094 94396 43146
rect 94396 43094 94428 43146
rect 94476 43094 94520 43146
rect 94520 43094 94532 43146
rect 94372 43092 94428 43094
rect 94476 43092 94532 43094
rect 94580 43092 94636 43148
rect 94684 43146 94740 43148
rect 94788 43146 94844 43148
rect 94684 43094 94696 43146
rect 94696 43094 94740 43146
rect 94788 43094 94820 43146
rect 94820 43094 94844 43146
rect 94684 43092 94740 43094
rect 94788 43092 94844 43094
rect 94892 43092 94948 43148
rect 92764 42978 92820 42980
rect 92764 42926 92766 42978
rect 92766 42926 92818 42978
rect 92818 42926 92820 42978
rect 92764 42924 92820 42926
rect 92316 42476 92372 42532
rect 93100 42530 93156 42532
rect 93100 42478 93102 42530
rect 93102 42478 93154 42530
rect 93154 42478 93156 42530
rect 93100 42476 93156 42478
rect 94268 41524 94324 41580
rect 94372 41578 94428 41580
rect 94476 41578 94532 41580
rect 94372 41526 94396 41578
rect 94396 41526 94428 41578
rect 94476 41526 94520 41578
rect 94520 41526 94532 41578
rect 94372 41524 94428 41526
rect 94476 41524 94532 41526
rect 94580 41524 94636 41580
rect 94684 41578 94740 41580
rect 94788 41578 94844 41580
rect 94684 41526 94696 41578
rect 94696 41526 94740 41578
rect 94788 41526 94820 41578
rect 94820 41526 94844 41578
rect 94684 41524 94740 41526
rect 94788 41524 94844 41526
rect 94892 41524 94948 41580
rect 96124 45724 96180 45780
rect 96236 45612 96292 45668
rect 95340 42924 95396 42980
rect 97020 51548 97076 51604
rect 96908 46674 96964 46676
rect 96908 46622 96910 46674
rect 96910 46622 96962 46674
rect 96962 46622 96964 46674
rect 96908 46620 96964 46622
rect 98140 56082 98196 56084
rect 98140 56030 98142 56082
rect 98142 56030 98194 56082
rect 98194 56030 98196 56082
rect 98140 56028 98196 56030
rect 98028 54908 98084 54964
rect 98028 53116 98084 53172
rect 97692 51324 97748 51380
rect 98028 49532 98084 49588
rect 98028 47740 98084 47796
rect 98028 45948 98084 46004
rect 98028 44210 98084 44212
rect 98028 44158 98030 44210
rect 98030 44158 98082 44210
rect 98082 44158 98084 44210
rect 98028 44156 98084 44158
rect 96236 42812 96292 42868
rect 91084 40124 91140 40180
rect 91644 40124 91700 40180
rect 90860 39004 90916 39060
rect 90188 38946 90244 38948
rect 90188 38894 90190 38946
rect 90190 38894 90242 38946
rect 90242 38894 90244 38946
rect 90188 38892 90244 38894
rect 90972 38946 91028 38948
rect 90972 38894 90974 38946
rect 90974 38894 91026 38946
rect 91026 38894 91028 38946
rect 90972 38892 91028 38894
rect 90972 37996 91028 38052
rect 91308 38946 91364 38948
rect 91308 38894 91310 38946
rect 91310 38894 91362 38946
rect 91362 38894 91364 38946
rect 91308 38892 91364 38894
rect 89768 37604 89824 37660
rect 89872 37658 89928 37660
rect 89976 37658 90032 37660
rect 89872 37606 89896 37658
rect 89896 37606 89928 37658
rect 89976 37606 90020 37658
rect 90020 37606 90032 37658
rect 89872 37604 89928 37606
rect 89976 37604 90032 37606
rect 90080 37604 90136 37660
rect 90184 37658 90240 37660
rect 90288 37658 90344 37660
rect 90184 37606 90196 37658
rect 90196 37606 90240 37658
rect 90288 37606 90320 37658
rect 90320 37606 90344 37658
rect 90184 37604 90240 37606
rect 90288 37604 90344 37606
rect 90392 37604 90448 37660
rect 89516 37436 89572 37492
rect 85372 36988 85428 37044
rect 87500 37042 87556 37044
rect 87500 36990 87502 37042
rect 87502 36990 87554 37042
rect 87554 36990 87556 37042
rect 87500 36988 87556 36990
rect 85268 36820 85324 36876
rect 85372 36874 85428 36876
rect 85476 36874 85532 36876
rect 85372 36822 85396 36874
rect 85396 36822 85428 36874
rect 85476 36822 85520 36874
rect 85520 36822 85532 36874
rect 85372 36820 85428 36822
rect 85476 36820 85532 36822
rect 85580 36820 85636 36876
rect 85684 36874 85740 36876
rect 85788 36874 85844 36876
rect 85684 36822 85696 36874
rect 85696 36822 85740 36874
rect 85788 36822 85820 36874
rect 85820 36822 85844 36874
rect 85684 36820 85740 36822
rect 85788 36820 85844 36822
rect 85892 36820 85948 36876
rect 89292 36204 89348 36260
rect 85484 35810 85540 35812
rect 85484 35758 85486 35810
rect 85486 35758 85538 35810
rect 85538 35758 85540 35810
rect 85484 35756 85540 35758
rect 89768 36036 89824 36092
rect 89872 36090 89928 36092
rect 89976 36090 90032 36092
rect 89872 36038 89896 36090
rect 89896 36038 89928 36090
rect 89976 36038 90020 36090
rect 90020 36038 90032 36090
rect 89872 36036 89928 36038
rect 89976 36036 90032 36038
rect 90080 36036 90136 36092
rect 90184 36090 90240 36092
rect 90288 36090 90344 36092
rect 90184 36038 90196 36090
rect 90196 36038 90240 36090
rect 90288 36038 90320 36090
rect 90320 36038 90344 36090
rect 90184 36036 90240 36038
rect 90288 36036 90344 36038
rect 90392 36036 90448 36092
rect 89516 35868 89572 35924
rect 85260 35698 85316 35700
rect 85260 35646 85262 35698
rect 85262 35646 85314 35698
rect 85314 35646 85316 35698
rect 85260 35644 85316 35646
rect 84924 35532 84980 35588
rect 85148 35420 85204 35476
rect 86044 35420 86100 35476
rect 86156 35644 86212 35700
rect 77644 34802 77700 34804
rect 77644 34750 77646 34802
rect 77646 34750 77698 34802
rect 77698 34750 77700 34802
rect 77644 34748 77700 34750
rect 80780 34802 80836 34804
rect 80780 34750 80782 34802
rect 80782 34750 80834 34802
rect 80834 34750 80836 34802
rect 80780 34748 80836 34750
rect 75180 34690 75236 34692
rect 75180 34638 75182 34690
rect 75182 34638 75234 34690
rect 75234 34638 75236 34690
rect 75180 34636 75236 34638
rect 75740 34300 75796 34356
rect 75852 34636 75908 34692
rect 71768 32900 71824 32956
rect 71872 32954 71928 32956
rect 71976 32954 72032 32956
rect 71872 32902 71896 32954
rect 71896 32902 71928 32954
rect 71976 32902 72020 32954
rect 72020 32902 72032 32954
rect 71872 32900 71928 32902
rect 71976 32900 72032 32902
rect 72080 32900 72136 32956
rect 72184 32954 72240 32956
rect 72288 32954 72344 32956
rect 72184 32902 72196 32954
rect 72196 32902 72240 32954
rect 72288 32902 72320 32954
rect 72320 32902 72344 32954
rect 72184 32900 72240 32902
rect 72288 32900 72344 32902
rect 72392 32900 72448 32956
rect 68572 31890 68628 31892
rect 68572 31838 68574 31890
rect 68574 31838 68626 31890
rect 68626 31838 68628 31890
rect 68572 31836 68628 31838
rect 70700 31836 70756 31892
rect 68908 31500 68964 31556
rect 69020 31388 69076 31444
rect 68572 30156 68628 30212
rect 69916 31388 69972 31444
rect 72940 31836 72996 31892
rect 73052 33292 73108 33348
rect 72940 31666 72996 31668
rect 72940 31614 72942 31666
rect 72942 31614 72994 31666
rect 72994 31614 72996 31666
rect 72940 31612 72996 31614
rect 70700 31388 70756 31444
rect 71148 31500 71204 31556
rect 69468 31106 69524 31108
rect 69468 31054 69470 31106
rect 69470 31054 69522 31106
rect 69522 31054 69524 31106
rect 69468 31052 69524 31054
rect 70364 30994 70420 30996
rect 70364 30942 70366 30994
rect 70366 30942 70418 30994
rect 70418 30942 70420 30994
rect 70364 30940 70420 30942
rect 69020 29596 69076 29652
rect 69692 29650 69748 29652
rect 69692 29598 69694 29650
rect 69694 29598 69746 29650
rect 69746 29598 69748 29650
rect 69692 29596 69748 29598
rect 69244 29426 69300 29428
rect 69244 29374 69246 29426
rect 69246 29374 69298 29426
rect 69298 29374 69300 29426
rect 69244 29372 69300 29374
rect 70476 29372 70532 29428
rect 68572 29260 68628 29316
rect 70700 28588 70756 28644
rect 72156 31554 72212 31556
rect 72156 31502 72158 31554
rect 72158 31502 72210 31554
rect 72210 31502 72212 31554
rect 72156 31500 72212 31502
rect 71768 31332 71824 31388
rect 71872 31386 71928 31388
rect 71976 31386 72032 31388
rect 71872 31334 71896 31386
rect 71896 31334 71928 31386
rect 71976 31334 72020 31386
rect 72020 31334 72032 31386
rect 71872 31332 71928 31334
rect 71976 31332 72032 31334
rect 72080 31332 72136 31388
rect 72184 31386 72240 31388
rect 72288 31386 72344 31388
rect 72184 31334 72196 31386
rect 72196 31334 72240 31386
rect 72288 31334 72320 31386
rect 72320 31334 72344 31386
rect 72184 31332 72240 31334
rect 72288 31332 72344 31334
rect 72392 31332 72448 31388
rect 74508 33292 74564 33348
rect 74060 31666 74116 31668
rect 74060 31614 74062 31666
rect 74062 31614 74114 31666
rect 74114 31614 74116 31666
rect 74060 31612 74116 31614
rect 74396 31554 74452 31556
rect 74396 31502 74398 31554
rect 74398 31502 74450 31554
rect 74450 31502 74452 31554
rect 74396 31500 74452 31502
rect 72268 30940 72324 30996
rect 72492 30210 72548 30212
rect 72492 30158 72494 30210
rect 72494 30158 72546 30210
rect 72546 30158 72548 30210
rect 72492 30156 72548 30158
rect 72828 30098 72884 30100
rect 72828 30046 72830 30098
rect 72830 30046 72882 30098
rect 72882 30046 72884 30098
rect 72828 30044 72884 30046
rect 71768 29764 71824 29820
rect 71872 29818 71928 29820
rect 71976 29818 72032 29820
rect 71872 29766 71896 29818
rect 71896 29766 71928 29818
rect 71976 29766 72020 29818
rect 72020 29766 72032 29818
rect 71872 29764 71928 29766
rect 71976 29764 72032 29766
rect 72080 29764 72136 29820
rect 72184 29818 72240 29820
rect 72288 29818 72344 29820
rect 72184 29766 72196 29818
rect 72196 29766 72240 29818
rect 72288 29766 72320 29818
rect 72320 29766 72344 29818
rect 72184 29764 72240 29766
rect 72288 29764 72344 29766
rect 72392 29764 72448 29820
rect 71932 28642 71988 28644
rect 71932 28590 71934 28642
rect 71934 28590 71986 28642
rect 71986 28590 71988 28642
rect 71932 28588 71988 28590
rect 72380 28642 72436 28644
rect 72380 28590 72382 28642
rect 72382 28590 72434 28642
rect 72434 28590 72436 28642
rect 72380 28588 72436 28590
rect 72716 28588 72772 28644
rect 71768 28196 71824 28252
rect 71872 28250 71928 28252
rect 71976 28250 72032 28252
rect 71872 28198 71896 28250
rect 71896 28198 71928 28250
rect 71976 28198 72020 28250
rect 72020 28198 72032 28250
rect 71872 28196 71928 28198
rect 71976 28196 72032 28198
rect 72080 28196 72136 28252
rect 72184 28250 72240 28252
rect 72288 28250 72344 28252
rect 72184 28198 72196 28250
rect 72196 28198 72240 28250
rect 72288 28198 72320 28250
rect 72320 28198 72344 28250
rect 72184 28196 72240 28198
rect 72288 28196 72344 28198
rect 72392 28196 72448 28252
rect 70812 27970 70868 27972
rect 70812 27918 70814 27970
rect 70814 27918 70866 27970
rect 70866 27918 70868 27970
rect 70812 27916 70868 27918
rect 71260 27970 71316 27972
rect 71260 27918 71262 27970
rect 71262 27918 71314 27970
rect 71314 27918 71316 27970
rect 71260 27916 71316 27918
rect 73052 27916 73108 27972
rect 67116 26796 67172 26852
rect 67340 26402 67396 26404
rect 67340 26350 67342 26402
rect 67342 26350 67394 26402
rect 67394 26350 67396 26402
rect 67340 26348 67396 26350
rect 68124 26402 68180 26404
rect 68124 26350 68126 26402
rect 68126 26350 68178 26402
rect 68178 26350 68180 26402
rect 68124 26348 68180 26350
rect 67268 25844 67324 25900
rect 67372 25898 67428 25900
rect 67476 25898 67532 25900
rect 67372 25846 67396 25898
rect 67396 25846 67428 25898
rect 67476 25846 67520 25898
rect 67520 25846 67532 25898
rect 67372 25844 67428 25846
rect 67476 25844 67532 25846
rect 67580 25844 67636 25900
rect 67684 25898 67740 25900
rect 67788 25898 67844 25900
rect 67684 25846 67696 25898
rect 67696 25846 67740 25898
rect 67788 25846 67820 25898
rect 67820 25846 67844 25898
rect 67684 25844 67740 25846
rect 67788 25844 67844 25846
rect 67892 25844 67948 25900
rect 72604 27132 72660 27188
rect 68908 26684 68964 26740
rect 67004 24892 67060 24948
rect 65548 23772 65604 23828
rect 66332 23548 66388 23604
rect 65996 23378 66052 23380
rect 65996 23326 65998 23378
rect 65998 23326 66050 23378
rect 66050 23326 66052 23378
rect 65996 23324 66052 23326
rect 67268 24276 67324 24332
rect 67372 24330 67428 24332
rect 67476 24330 67532 24332
rect 67372 24278 67396 24330
rect 67396 24278 67428 24330
rect 67476 24278 67520 24330
rect 67520 24278 67532 24330
rect 67372 24276 67428 24278
rect 67476 24276 67532 24278
rect 67580 24276 67636 24332
rect 67684 24330 67740 24332
rect 67788 24330 67844 24332
rect 67684 24278 67696 24330
rect 67696 24278 67740 24330
rect 67788 24278 67820 24330
rect 67820 24278 67844 24330
rect 67684 24276 67740 24278
rect 67788 24276 67844 24278
rect 67892 24276 67948 24332
rect 67004 23324 67060 23380
rect 67268 22708 67324 22764
rect 67372 22762 67428 22764
rect 67476 22762 67532 22764
rect 67372 22710 67396 22762
rect 67396 22710 67428 22762
rect 67476 22710 67520 22762
rect 67520 22710 67532 22762
rect 67372 22708 67428 22710
rect 67476 22708 67532 22710
rect 67580 22708 67636 22764
rect 67684 22762 67740 22764
rect 67788 22762 67844 22764
rect 67684 22710 67696 22762
rect 67696 22710 67740 22762
rect 67788 22710 67820 22762
rect 67820 22710 67844 22762
rect 67684 22708 67740 22710
rect 67788 22708 67844 22710
rect 67892 22708 67948 22764
rect 68572 22428 68628 22484
rect 68348 22370 68404 22372
rect 68348 22318 68350 22370
rect 68350 22318 68402 22370
rect 68402 22318 68404 22370
rect 68348 22316 68404 22318
rect 66668 21756 66724 21812
rect 67268 21140 67324 21196
rect 67372 21194 67428 21196
rect 67476 21194 67532 21196
rect 67372 21142 67396 21194
rect 67396 21142 67428 21194
rect 67476 21142 67520 21194
rect 67520 21142 67532 21194
rect 67372 21140 67428 21142
rect 67476 21140 67532 21142
rect 67580 21140 67636 21196
rect 67684 21194 67740 21196
rect 67788 21194 67844 21196
rect 67684 21142 67696 21194
rect 67696 21142 67740 21194
rect 67788 21142 67820 21194
rect 67820 21142 67844 21194
rect 67684 21140 67740 21142
rect 67788 21140 67844 21142
rect 67892 21140 67948 21196
rect 65548 20914 65604 20916
rect 65548 20862 65550 20914
rect 65550 20862 65602 20914
rect 65602 20862 65604 20914
rect 65548 20860 65604 20862
rect 65884 20972 65940 21028
rect 70476 26684 70532 26740
rect 71768 26628 71824 26684
rect 71872 26682 71928 26684
rect 71976 26682 72032 26684
rect 71872 26630 71896 26682
rect 71896 26630 71928 26682
rect 71976 26630 72020 26682
rect 72020 26630 72032 26682
rect 71872 26628 71928 26630
rect 71976 26628 72032 26630
rect 72080 26628 72136 26684
rect 72184 26682 72240 26684
rect 72288 26682 72344 26684
rect 72184 26630 72196 26682
rect 72196 26630 72240 26682
rect 72288 26630 72320 26682
rect 72320 26630 72344 26682
rect 72184 26628 72240 26630
rect 72288 26628 72344 26630
rect 72392 26628 72448 26684
rect 73164 27746 73220 27748
rect 73164 27694 73166 27746
rect 73166 27694 73218 27746
rect 73218 27694 73220 27746
rect 73164 27692 73220 27694
rect 73612 27692 73668 27748
rect 75068 33292 75124 33348
rect 76412 34690 76468 34692
rect 76412 34638 76414 34690
rect 76414 34638 76466 34690
rect 76466 34638 76468 34690
rect 76412 34636 76468 34638
rect 76188 34300 76244 34356
rect 80768 34468 80824 34524
rect 80872 34522 80928 34524
rect 80976 34522 81032 34524
rect 80872 34470 80896 34522
rect 80896 34470 80928 34522
rect 80976 34470 81020 34522
rect 81020 34470 81032 34522
rect 80872 34468 80928 34470
rect 80976 34468 81032 34470
rect 81080 34468 81136 34524
rect 81184 34522 81240 34524
rect 81288 34522 81344 34524
rect 81184 34470 81196 34522
rect 81196 34470 81240 34522
rect 81288 34470 81320 34522
rect 81320 34470 81344 34522
rect 81184 34468 81240 34470
rect 81288 34468 81344 34470
rect 81392 34468 81448 34524
rect 76412 34300 76468 34356
rect 84364 34300 84420 34356
rect 76524 34242 76580 34244
rect 76524 34190 76526 34242
rect 76526 34190 76578 34242
rect 76578 34190 76580 34242
rect 76524 34188 76580 34190
rect 76268 33684 76324 33740
rect 76372 33738 76428 33740
rect 76476 33738 76532 33740
rect 76372 33686 76396 33738
rect 76396 33686 76428 33738
rect 76476 33686 76520 33738
rect 76520 33686 76532 33738
rect 76372 33684 76428 33686
rect 76476 33684 76532 33686
rect 76580 33684 76636 33740
rect 76684 33738 76740 33740
rect 76788 33738 76844 33740
rect 76684 33686 76696 33738
rect 76696 33686 76740 33738
rect 76788 33686 76820 33738
rect 76820 33686 76844 33738
rect 76684 33684 76740 33686
rect 76788 33684 76844 33686
rect 76892 33684 76948 33740
rect 80768 32900 80824 32956
rect 80872 32954 80928 32956
rect 80976 32954 81032 32956
rect 80872 32902 80896 32954
rect 80896 32902 80928 32954
rect 80976 32902 81020 32954
rect 81020 32902 81032 32954
rect 80872 32900 80928 32902
rect 80976 32900 81032 32902
rect 81080 32900 81136 32956
rect 81184 32954 81240 32956
rect 81288 32954 81344 32956
rect 81184 32902 81196 32954
rect 81196 32902 81240 32954
rect 81288 32902 81320 32954
rect 81320 32902 81344 32954
rect 81184 32900 81240 32902
rect 81288 32900 81344 32902
rect 81392 32900 81448 32956
rect 75404 29372 75460 29428
rect 73052 26908 73108 26964
rect 74508 26796 74564 26852
rect 72716 26402 72772 26404
rect 72716 26350 72718 26402
rect 72718 26350 72770 26402
rect 72770 26350 72772 26402
rect 72716 26348 72772 26350
rect 73500 26402 73556 26404
rect 73500 26350 73502 26402
rect 73502 26350 73554 26402
rect 73554 26350 73556 26402
rect 73500 26348 73556 26350
rect 73164 26290 73220 26292
rect 73164 26238 73166 26290
rect 73166 26238 73218 26290
rect 73218 26238 73220 26290
rect 73164 26236 73220 26238
rect 74172 26236 74228 26292
rect 71768 25060 71824 25116
rect 71872 25114 71928 25116
rect 71976 25114 72032 25116
rect 71872 25062 71896 25114
rect 71896 25062 71928 25114
rect 71976 25062 72020 25114
rect 72020 25062 72032 25114
rect 71872 25060 71928 25062
rect 71976 25060 72032 25062
rect 72080 25060 72136 25116
rect 72184 25114 72240 25116
rect 72288 25114 72344 25116
rect 72184 25062 72196 25114
rect 72196 25062 72240 25114
rect 72288 25062 72320 25114
rect 72320 25062 72344 25114
rect 72184 25060 72240 25062
rect 72288 25060 72344 25062
rect 72392 25060 72448 25116
rect 68796 24892 68852 24948
rect 70252 24946 70308 24948
rect 70252 24894 70254 24946
rect 70254 24894 70306 24946
rect 70306 24894 70308 24946
rect 70252 24892 70308 24894
rect 71148 24892 71204 24948
rect 74508 26124 74564 26180
rect 75068 25340 75124 25396
rect 74508 25228 74564 25284
rect 74396 24834 74452 24836
rect 74396 24782 74398 24834
rect 74398 24782 74450 24834
rect 74450 24782 74452 24834
rect 74396 24780 74452 24782
rect 74956 25228 75012 25284
rect 69468 23324 69524 23380
rect 69804 23378 69860 23380
rect 69804 23326 69806 23378
rect 69806 23326 69858 23378
rect 69858 23326 69860 23378
rect 69804 23324 69860 23326
rect 69356 22876 69412 22932
rect 70588 22930 70644 22932
rect 70588 22878 70590 22930
rect 70590 22878 70642 22930
rect 70642 22878 70644 22930
rect 70588 22876 70644 22878
rect 69916 22482 69972 22484
rect 69916 22430 69918 22482
rect 69918 22430 69970 22482
rect 69970 22430 69972 22482
rect 69916 22428 69972 22430
rect 69468 21644 69524 21700
rect 70364 21644 70420 21700
rect 68684 20860 68740 20916
rect 67268 19572 67324 19628
rect 67372 19626 67428 19628
rect 67476 19626 67532 19628
rect 67372 19574 67396 19626
rect 67396 19574 67428 19626
rect 67476 19574 67520 19626
rect 67520 19574 67532 19626
rect 67372 19572 67428 19574
rect 67476 19572 67532 19574
rect 67580 19572 67636 19628
rect 67684 19626 67740 19628
rect 67788 19626 67844 19628
rect 67684 19574 67696 19626
rect 67696 19574 67740 19626
rect 67788 19574 67820 19626
rect 67820 19574 67844 19626
rect 67684 19572 67740 19574
rect 67788 19572 67844 19574
rect 67892 19572 67948 19628
rect 67268 18004 67324 18060
rect 67372 18058 67428 18060
rect 67476 18058 67532 18060
rect 67372 18006 67396 18058
rect 67396 18006 67428 18058
rect 67476 18006 67520 18058
rect 67520 18006 67532 18058
rect 67372 18004 67428 18006
rect 67476 18004 67532 18006
rect 67580 18004 67636 18060
rect 67684 18058 67740 18060
rect 67788 18058 67844 18060
rect 67684 18006 67696 18058
rect 67696 18006 67740 18058
rect 67788 18006 67820 18058
rect 67820 18006 67844 18058
rect 67684 18004 67740 18006
rect 67788 18004 67844 18006
rect 67892 18004 67948 18060
rect 67268 16436 67324 16492
rect 67372 16490 67428 16492
rect 67476 16490 67532 16492
rect 67372 16438 67396 16490
rect 67396 16438 67428 16490
rect 67476 16438 67520 16490
rect 67520 16438 67532 16490
rect 67372 16436 67428 16438
rect 67476 16436 67532 16438
rect 67580 16436 67636 16492
rect 67684 16490 67740 16492
rect 67788 16490 67844 16492
rect 67684 16438 67696 16490
rect 67696 16438 67740 16490
rect 67788 16438 67820 16490
rect 67820 16438 67844 16490
rect 67684 16436 67740 16438
rect 67788 16436 67844 16438
rect 67892 16436 67948 16492
rect 66220 16044 66276 16100
rect 62768 14084 62824 14140
rect 62872 14138 62928 14140
rect 62976 14138 63032 14140
rect 62872 14086 62896 14138
rect 62896 14086 62928 14138
rect 62976 14086 63020 14138
rect 63020 14086 63032 14138
rect 62872 14084 62928 14086
rect 62976 14084 63032 14086
rect 63080 14084 63136 14140
rect 63184 14138 63240 14140
rect 63288 14138 63344 14140
rect 63184 14086 63196 14138
rect 63196 14086 63240 14138
rect 63288 14086 63320 14138
rect 63320 14086 63344 14138
rect 63184 14084 63240 14086
rect 63288 14084 63344 14086
rect 63392 14084 63448 14140
rect 61292 11452 61348 11508
rect 61180 7084 61236 7140
rect 60284 4172 60340 4228
rect 60172 3836 60228 3892
rect 52668 3442 52724 3444
rect 52668 3390 52670 3442
rect 52670 3390 52722 3442
rect 52722 3390 52724 3442
rect 52668 3388 52724 3390
rect 42700 3164 42756 3220
rect 44768 3108 44824 3164
rect 44872 3162 44928 3164
rect 44976 3162 45032 3164
rect 44872 3110 44896 3162
rect 44896 3110 44928 3162
rect 44976 3110 45020 3162
rect 45020 3110 45032 3162
rect 44872 3108 44928 3110
rect 44976 3108 45032 3110
rect 45080 3108 45136 3164
rect 45184 3162 45240 3164
rect 45288 3162 45344 3164
rect 45184 3110 45196 3162
rect 45196 3110 45240 3162
rect 45288 3110 45320 3162
rect 45320 3110 45344 3162
rect 45184 3108 45240 3110
rect 45288 3108 45344 3110
rect 45392 3108 45448 3164
rect 60732 5234 60788 5236
rect 60732 5182 60734 5234
rect 60734 5182 60786 5234
rect 60786 5182 60788 5234
rect 60732 5180 60788 5182
rect 62768 12516 62824 12572
rect 62872 12570 62928 12572
rect 62976 12570 63032 12572
rect 62872 12518 62896 12570
rect 62896 12518 62928 12570
rect 62976 12518 63020 12570
rect 63020 12518 63032 12570
rect 62872 12516 62928 12518
rect 62976 12516 63032 12518
rect 63080 12516 63136 12572
rect 63184 12570 63240 12572
rect 63288 12570 63344 12572
rect 63184 12518 63196 12570
rect 63196 12518 63240 12570
rect 63288 12518 63320 12570
rect 63320 12518 63344 12570
rect 63184 12516 63240 12518
rect 63288 12516 63344 12518
rect 63392 12516 63448 12572
rect 62188 11506 62244 11508
rect 62188 11454 62190 11506
rect 62190 11454 62242 11506
rect 62242 11454 62244 11506
rect 62188 11452 62244 11454
rect 63644 11452 63700 11508
rect 62768 10948 62824 11004
rect 62872 11002 62928 11004
rect 62976 11002 63032 11004
rect 62872 10950 62896 11002
rect 62896 10950 62928 11002
rect 62976 10950 63020 11002
rect 63020 10950 63032 11002
rect 62872 10948 62928 10950
rect 62976 10948 63032 10950
rect 63080 10948 63136 11004
rect 63184 11002 63240 11004
rect 63288 11002 63344 11004
rect 63184 10950 63196 11002
rect 63196 10950 63240 11002
rect 63288 10950 63320 11002
rect 63320 10950 63344 11002
rect 63184 10948 63240 10950
rect 63288 10948 63344 10950
rect 63392 10948 63448 11004
rect 62768 9380 62824 9436
rect 62872 9434 62928 9436
rect 62976 9434 63032 9436
rect 62872 9382 62896 9434
rect 62896 9382 62928 9434
rect 62976 9382 63020 9434
rect 63020 9382 63032 9434
rect 62872 9380 62928 9382
rect 62976 9380 63032 9382
rect 63080 9380 63136 9436
rect 63184 9434 63240 9436
rect 63288 9434 63344 9436
rect 63184 9382 63196 9434
rect 63196 9382 63240 9434
rect 63288 9382 63320 9434
rect 63320 9382 63344 9434
rect 63184 9380 63240 9382
rect 63288 9380 63344 9382
rect 63392 9380 63448 9436
rect 62412 8316 62468 8372
rect 63644 10108 63700 10164
rect 61964 8258 62020 8260
rect 61964 8206 61966 8258
rect 61966 8206 62018 8258
rect 62018 8206 62020 8258
rect 61964 8204 62020 8206
rect 63084 7980 63140 8036
rect 62768 7812 62824 7868
rect 62872 7866 62928 7868
rect 62976 7866 63032 7868
rect 62872 7814 62896 7866
rect 62896 7814 62928 7866
rect 62976 7814 63020 7866
rect 63020 7814 63032 7866
rect 62872 7812 62928 7814
rect 62976 7812 63032 7814
rect 63080 7812 63136 7868
rect 63184 7866 63240 7868
rect 63288 7866 63344 7868
rect 63184 7814 63196 7866
rect 63196 7814 63240 7866
rect 63288 7814 63320 7866
rect 63320 7814 63344 7866
rect 63184 7812 63240 7814
rect 63288 7812 63344 7814
rect 63392 7812 63448 7868
rect 62188 6300 62244 6356
rect 62412 6636 62468 6692
rect 62636 6636 62692 6692
rect 62768 6244 62824 6300
rect 62872 6298 62928 6300
rect 62976 6298 63032 6300
rect 62872 6246 62896 6298
rect 62896 6246 62928 6298
rect 62976 6246 63020 6298
rect 63020 6246 63032 6298
rect 62872 6244 62928 6246
rect 62976 6244 63032 6246
rect 63080 6244 63136 6300
rect 63184 6298 63240 6300
rect 63288 6298 63344 6300
rect 63184 6246 63196 6298
rect 63196 6246 63240 6298
rect 63288 6246 63320 6298
rect 63320 6246 63344 6298
rect 63184 6244 63240 6246
rect 63288 6244 63344 6246
rect 63392 6244 63448 6300
rect 64428 7084 64484 7140
rect 64652 5292 64708 5348
rect 62768 4676 62824 4732
rect 62872 4730 62928 4732
rect 62976 4730 63032 4732
rect 62872 4678 62896 4730
rect 62896 4678 62928 4730
rect 62976 4678 63020 4730
rect 63020 4678 63032 4730
rect 62872 4676 62928 4678
rect 62976 4676 63032 4678
rect 63080 4676 63136 4732
rect 63184 4730 63240 4732
rect 63288 4730 63344 4732
rect 63184 4678 63196 4730
rect 63196 4678 63240 4730
rect 63288 4678 63320 4730
rect 63320 4678 63344 4730
rect 63184 4676 63240 4678
rect 63288 4676 63344 4678
rect 63392 4676 63448 4732
rect 63196 4562 63252 4564
rect 63196 4510 63198 4562
rect 63198 4510 63250 4562
rect 63250 4510 63252 4562
rect 63196 4508 63252 4510
rect 62748 4450 62804 4452
rect 62748 4398 62750 4450
rect 62750 4398 62802 4450
rect 62802 4398 62804 4450
rect 62748 4396 62804 4398
rect 62188 4226 62244 4228
rect 62188 4174 62190 4226
rect 62190 4174 62242 4226
rect 62242 4174 62244 4226
rect 62188 4172 62244 4174
rect 61740 3836 61796 3892
rect 60844 3778 60900 3780
rect 60844 3726 60846 3778
rect 60846 3726 60898 3778
rect 60898 3726 60900 3778
rect 60844 3724 60900 3726
rect 60732 3666 60788 3668
rect 60732 3614 60734 3666
rect 60734 3614 60786 3666
rect 60786 3614 60788 3666
rect 60732 3612 60788 3614
rect 67268 14868 67324 14924
rect 67372 14922 67428 14924
rect 67476 14922 67532 14924
rect 67372 14870 67396 14922
rect 67396 14870 67428 14922
rect 67476 14870 67520 14922
rect 67520 14870 67532 14922
rect 67372 14868 67428 14870
rect 67476 14868 67532 14870
rect 67580 14868 67636 14924
rect 67684 14922 67740 14924
rect 67788 14922 67844 14924
rect 67684 14870 67696 14922
rect 67696 14870 67740 14922
rect 67788 14870 67820 14922
rect 67820 14870 67844 14922
rect 67684 14868 67740 14870
rect 67788 14868 67844 14870
rect 67892 14868 67948 14924
rect 68348 14476 68404 14532
rect 65548 13692 65604 13748
rect 67268 13300 67324 13356
rect 67372 13354 67428 13356
rect 67476 13354 67532 13356
rect 67372 13302 67396 13354
rect 67396 13302 67428 13354
rect 67476 13302 67520 13354
rect 67520 13302 67532 13354
rect 67372 13300 67428 13302
rect 67476 13300 67532 13302
rect 67580 13300 67636 13356
rect 67684 13354 67740 13356
rect 67788 13354 67844 13356
rect 67684 13302 67696 13354
rect 67696 13302 67740 13354
rect 67788 13302 67820 13354
rect 67820 13302 67844 13354
rect 67684 13300 67740 13302
rect 67788 13300 67844 13302
rect 67892 13300 67948 13356
rect 65772 11340 65828 11396
rect 65548 6636 65604 6692
rect 65436 6524 65492 6580
rect 65324 4508 65380 4564
rect 65996 10108 66052 10164
rect 63532 3724 63588 3780
rect 62748 3666 62804 3668
rect 62748 3614 62750 3666
rect 62750 3614 62802 3666
rect 62802 3614 62804 3666
rect 62748 3612 62804 3614
rect 61292 3554 61348 3556
rect 61292 3502 61294 3554
rect 61294 3502 61346 3554
rect 61346 3502 61348 3554
rect 61292 3500 61348 3502
rect 63196 3554 63252 3556
rect 63196 3502 63198 3554
rect 63198 3502 63250 3554
rect 63250 3502 63252 3554
rect 63196 3500 63252 3502
rect 67268 11732 67324 11788
rect 67372 11786 67428 11788
rect 67476 11786 67532 11788
rect 67372 11734 67396 11786
rect 67396 11734 67428 11786
rect 67476 11734 67520 11786
rect 67520 11734 67532 11786
rect 67372 11732 67428 11734
rect 67476 11732 67532 11734
rect 67580 11732 67636 11788
rect 67684 11786 67740 11788
rect 67788 11786 67844 11788
rect 67684 11734 67696 11786
rect 67696 11734 67740 11786
rect 67788 11734 67820 11786
rect 67820 11734 67844 11786
rect 67684 11732 67740 11734
rect 67788 11732 67844 11734
rect 67892 11732 67948 11788
rect 67564 11618 67620 11620
rect 67564 11566 67566 11618
rect 67566 11566 67618 11618
rect 67618 11566 67620 11618
rect 67564 11564 67620 11566
rect 67268 10164 67324 10220
rect 67372 10218 67428 10220
rect 67476 10218 67532 10220
rect 67372 10166 67396 10218
rect 67396 10166 67428 10218
rect 67476 10166 67520 10218
rect 67520 10166 67532 10218
rect 67372 10164 67428 10166
rect 67476 10164 67532 10166
rect 67580 10164 67636 10220
rect 67684 10218 67740 10220
rect 67788 10218 67844 10220
rect 67684 10166 67696 10218
rect 67696 10166 67740 10218
rect 67788 10166 67820 10218
rect 67820 10166 67844 10218
rect 67684 10164 67740 10166
rect 67788 10164 67844 10166
rect 67892 10164 67948 10220
rect 67268 8596 67324 8652
rect 67372 8650 67428 8652
rect 67476 8650 67532 8652
rect 67372 8598 67396 8650
rect 67396 8598 67428 8650
rect 67476 8598 67520 8650
rect 67520 8598 67532 8650
rect 67372 8596 67428 8598
rect 67476 8596 67532 8598
rect 67580 8596 67636 8652
rect 67684 8650 67740 8652
rect 67788 8650 67844 8652
rect 67684 8598 67696 8650
rect 67696 8598 67740 8650
rect 67788 8598 67820 8650
rect 67820 8598 67844 8650
rect 67684 8596 67740 8598
rect 67788 8596 67844 8598
rect 67892 8596 67948 8652
rect 66220 8204 66276 8260
rect 66220 7868 66276 7924
rect 66444 7586 66500 7588
rect 66444 7534 66446 7586
rect 66446 7534 66498 7586
rect 66498 7534 66500 7586
rect 66444 7532 66500 7534
rect 67268 7028 67324 7084
rect 67372 7082 67428 7084
rect 67476 7082 67532 7084
rect 67372 7030 67396 7082
rect 67396 7030 67428 7082
rect 67476 7030 67520 7082
rect 67520 7030 67532 7082
rect 67372 7028 67428 7030
rect 67476 7028 67532 7030
rect 67580 7028 67636 7084
rect 67684 7082 67740 7084
rect 67788 7082 67844 7084
rect 67684 7030 67696 7082
rect 67696 7030 67740 7082
rect 67788 7030 67820 7082
rect 67820 7030 67844 7082
rect 67684 7028 67740 7030
rect 67788 7028 67844 7030
rect 67892 7028 67948 7084
rect 68124 7084 68180 7140
rect 67268 5460 67324 5516
rect 67372 5514 67428 5516
rect 67476 5514 67532 5516
rect 67372 5462 67396 5514
rect 67396 5462 67428 5514
rect 67476 5462 67520 5514
rect 67520 5462 67532 5514
rect 67372 5460 67428 5462
rect 67476 5460 67532 5462
rect 67580 5460 67636 5516
rect 67684 5514 67740 5516
rect 67788 5514 67844 5516
rect 67684 5462 67696 5514
rect 67696 5462 67740 5514
rect 67788 5462 67820 5514
rect 67820 5462 67844 5514
rect 67684 5460 67740 5462
rect 67788 5460 67844 5462
rect 67892 5460 67948 5516
rect 70028 14530 70084 14532
rect 70028 14478 70030 14530
rect 70030 14478 70082 14530
rect 70082 14478 70084 14530
rect 70028 14476 70084 14478
rect 68348 13692 68404 13748
rect 68348 11564 68404 11620
rect 67340 4956 67396 5012
rect 68348 5122 68404 5124
rect 68348 5070 68350 5122
rect 68350 5070 68402 5122
rect 68402 5070 68404 5122
rect 68348 5068 68404 5070
rect 68236 4956 68292 5012
rect 67268 3892 67324 3948
rect 67372 3946 67428 3948
rect 67476 3946 67532 3948
rect 67372 3894 67396 3946
rect 67396 3894 67428 3946
rect 67476 3894 67520 3946
rect 67520 3894 67532 3946
rect 67372 3892 67428 3894
rect 67476 3892 67532 3894
rect 67580 3892 67636 3948
rect 67684 3946 67740 3948
rect 67788 3946 67844 3948
rect 67684 3894 67696 3946
rect 67696 3894 67740 3946
rect 67788 3894 67820 3946
rect 67820 3894 67844 3946
rect 67684 3892 67740 3894
rect 67788 3892 67844 3894
rect 67892 3892 67948 3948
rect 69020 6578 69076 6580
rect 69020 6526 69022 6578
rect 69022 6526 69074 6578
rect 69074 6526 69076 6578
rect 69020 6524 69076 6526
rect 70140 6972 70196 7028
rect 69692 5964 69748 6020
rect 68460 3724 68516 3780
rect 69580 3778 69636 3780
rect 69580 3726 69582 3778
rect 69582 3726 69634 3778
rect 69634 3726 69636 3778
rect 69580 3724 69636 3726
rect 67452 3388 67508 3444
rect 71372 20524 71428 20580
rect 73500 23660 73556 23716
rect 71768 23492 71824 23548
rect 71872 23546 71928 23548
rect 71976 23546 72032 23548
rect 71872 23494 71896 23546
rect 71896 23494 71928 23546
rect 71976 23494 72020 23546
rect 72020 23494 72032 23546
rect 71872 23492 71928 23494
rect 71976 23492 72032 23494
rect 72080 23492 72136 23548
rect 72184 23546 72240 23548
rect 72288 23546 72344 23548
rect 72184 23494 72196 23546
rect 72196 23494 72240 23546
rect 72288 23494 72320 23546
rect 72320 23494 72344 23546
rect 72184 23492 72240 23494
rect 72288 23492 72344 23494
rect 72392 23492 72448 23548
rect 72156 23212 72212 23268
rect 72940 23266 72996 23268
rect 72940 23214 72942 23266
rect 72942 23214 72994 23266
rect 72994 23214 72996 23266
rect 72940 23212 72996 23214
rect 73724 23266 73780 23268
rect 73724 23214 73726 23266
rect 73726 23214 73778 23266
rect 73778 23214 73780 23266
rect 73724 23212 73780 23214
rect 74508 23266 74564 23268
rect 74508 23214 74510 23266
rect 74510 23214 74562 23266
rect 74562 23214 74564 23266
rect 74508 23212 74564 23214
rect 73724 22428 73780 22484
rect 75068 22428 75124 22484
rect 71768 21924 71824 21980
rect 71872 21978 71928 21980
rect 71976 21978 72032 21980
rect 71872 21926 71896 21978
rect 71896 21926 71928 21978
rect 71976 21926 72020 21978
rect 72020 21926 72032 21978
rect 71872 21924 71928 21926
rect 71976 21924 72032 21926
rect 72080 21924 72136 21980
rect 72184 21978 72240 21980
rect 72288 21978 72344 21980
rect 72184 21926 72196 21978
rect 72196 21926 72240 21978
rect 72288 21926 72320 21978
rect 72320 21926 72344 21978
rect 72184 21924 72240 21926
rect 72288 21924 72344 21926
rect 72392 21924 72448 21980
rect 74844 21980 74900 22036
rect 73500 21532 73556 21588
rect 72044 20802 72100 20804
rect 72044 20750 72046 20802
rect 72046 20750 72098 20802
rect 72098 20750 72100 20802
rect 72044 20748 72100 20750
rect 72156 20578 72212 20580
rect 72156 20526 72158 20578
rect 72158 20526 72210 20578
rect 72210 20526 72212 20578
rect 72156 20524 72212 20526
rect 72492 20524 72548 20580
rect 73052 20578 73108 20580
rect 73052 20526 73054 20578
rect 73054 20526 73106 20578
rect 73106 20526 73108 20578
rect 73052 20524 73108 20526
rect 71768 20356 71824 20412
rect 71872 20410 71928 20412
rect 71976 20410 72032 20412
rect 71872 20358 71896 20410
rect 71896 20358 71928 20410
rect 71976 20358 72020 20410
rect 72020 20358 72032 20410
rect 71872 20356 71928 20358
rect 71976 20356 72032 20358
rect 72080 20356 72136 20412
rect 72184 20410 72240 20412
rect 72288 20410 72344 20412
rect 72184 20358 72196 20410
rect 72196 20358 72240 20410
rect 72288 20358 72320 20410
rect 72320 20358 72344 20410
rect 72184 20356 72240 20358
rect 72288 20356 72344 20358
rect 72392 20356 72448 20412
rect 73388 20130 73444 20132
rect 73388 20078 73390 20130
rect 73390 20078 73442 20130
rect 73442 20078 73444 20130
rect 73388 20076 73444 20078
rect 75180 21698 75236 21700
rect 75180 21646 75182 21698
rect 75182 21646 75234 21698
rect 75234 21646 75236 21698
rect 75180 21644 75236 21646
rect 76268 32116 76324 32172
rect 76372 32170 76428 32172
rect 76476 32170 76532 32172
rect 76372 32118 76396 32170
rect 76396 32118 76428 32170
rect 76476 32118 76520 32170
rect 76520 32118 76532 32170
rect 76372 32116 76428 32118
rect 76476 32116 76532 32118
rect 76580 32116 76636 32172
rect 76684 32170 76740 32172
rect 76788 32170 76844 32172
rect 76684 32118 76696 32170
rect 76696 32118 76740 32170
rect 76788 32118 76820 32170
rect 76820 32118 76844 32170
rect 76684 32116 76740 32118
rect 76788 32116 76844 32118
rect 76892 32116 76948 32172
rect 80768 31332 80824 31388
rect 80872 31386 80928 31388
rect 80976 31386 81032 31388
rect 80872 31334 80896 31386
rect 80896 31334 80928 31386
rect 80976 31334 81020 31386
rect 81020 31334 81032 31386
rect 80872 31332 80928 31334
rect 80976 31332 81032 31334
rect 81080 31332 81136 31388
rect 81184 31386 81240 31388
rect 81288 31386 81344 31388
rect 81184 31334 81196 31386
rect 81196 31334 81240 31386
rect 81288 31334 81320 31386
rect 81320 31334 81344 31386
rect 81184 31332 81240 31334
rect 81288 31332 81344 31334
rect 81392 31332 81448 31388
rect 76268 30548 76324 30604
rect 76372 30602 76428 30604
rect 76476 30602 76532 30604
rect 76372 30550 76396 30602
rect 76396 30550 76428 30602
rect 76476 30550 76520 30602
rect 76520 30550 76532 30602
rect 76372 30548 76428 30550
rect 76476 30548 76532 30550
rect 76580 30548 76636 30604
rect 76684 30602 76740 30604
rect 76788 30602 76844 30604
rect 76684 30550 76696 30602
rect 76696 30550 76740 30602
rect 76788 30550 76820 30602
rect 76820 30550 76844 30602
rect 76684 30548 76740 30550
rect 76788 30548 76844 30550
rect 76892 30548 76948 30604
rect 85268 35252 85324 35308
rect 85372 35306 85428 35308
rect 85476 35306 85532 35308
rect 85372 35254 85396 35306
rect 85396 35254 85428 35306
rect 85476 35254 85520 35306
rect 85520 35254 85532 35306
rect 85372 35252 85428 35254
rect 85476 35252 85532 35254
rect 85580 35252 85636 35308
rect 85684 35306 85740 35308
rect 85788 35306 85844 35308
rect 85684 35254 85696 35306
rect 85696 35254 85740 35306
rect 85788 35254 85820 35306
rect 85820 35254 85844 35306
rect 85684 35252 85740 35254
rect 85788 35252 85844 35254
rect 85892 35252 85948 35308
rect 85372 35084 85428 35140
rect 85820 34748 85876 34804
rect 85372 34188 85428 34244
rect 85932 34242 85988 34244
rect 85932 34190 85934 34242
rect 85934 34190 85986 34242
rect 85986 34190 85988 34242
rect 85932 34188 85988 34190
rect 89964 35644 90020 35700
rect 94780 40460 94836 40516
rect 95340 40402 95396 40404
rect 95340 40350 95342 40402
rect 95342 40350 95394 40402
rect 95394 40350 95396 40402
rect 95340 40348 95396 40350
rect 96236 40572 96292 40628
rect 96124 40348 96180 40404
rect 94268 39956 94324 40012
rect 94372 40010 94428 40012
rect 94476 40010 94532 40012
rect 94372 39958 94396 40010
rect 94396 39958 94428 40010
rect 94476 39958 94520 40010
rect 94520 39958 94532 40010
rect 94372 39956 94428 39958
rect 94476 39956 94532 39958
rect 94580 39956 94636 40012
rect 94684 40010 94740 40012
rect 94788 40010 94844 40012
rect 94684 39958 94696 40010
rect 94696 39958 94740 40010
rect 94788 39958 94820 40010
rect 94820 39958 94844 40010
rect 94684 39956 94740 39958
rect 94788 39956 94844 39958
rect 94892 39956 94948 40012
rect 96236 39340 96292 39396
rect 94268 38388 94324 38444
rect 94372 38442 94428 38444
rect 94476 38442 94532 38444
rect 94372 38390 94396 38442
rect 94396 38390 94428 38442
rect 94476 38390 94520 38442
rect 94520 38390 94532 38442
rect 94372 38388 94428 38390
rect 94476 38388 94532 38390
rect 94580 38388 94636 38444
rect 94684 38442 94740 38444
rect 94788 38442 94844 38444
rect 94684 38390 94696 38442
rect 94696 38390 94740 38442
rect 94788 38390 94820 38442
rect 94820 38390 94844 38442
rect 94684 38388 94740 38390
rect 94788 38388 94844 38390
rect 94892 38388 94948 38444
rect 94268 36820 94324 36876
rect 94372 36874 94428 36876
rect 94476 36874 94532 36876
rect 94372 36822 94396 36874
rect 94396 36822 94428 36874
rect 94476 36822 94520 36874
rect 94520 36822 94532 36874
rect 94372 36820 94428 36822
rect 94476 36820 94532 36822
rect 94580 36820 94636 36876
rect 94684 36874 94740 36876
rect 94788 36874 94844 36876
rect 94684 36822 94696 36874
rect 94696 36822 94740 36874
rect 94788 36822 94820 36874
rect 94820 36822 94844 36874
rect 94684 36820 94740 36822
rect 94788 36820 94844 36822
rect 94892 36820 94948 36876
rect 91868 36258 91924 36260
rect 91868 36206 91870 36258
rect 91870 36206 91922 36258
rect 91922 36206 91924 36258
rect 91868 36204 91924 36206
rect 89068 34860 89124 34916
rect 88172 34802 88228 34804
rect 88172 34750 88174 34802
rect 88174 34750 88226 34802
rect 88226 34750 88228 34802
rect 88172 34748 88228 34750
rect 89768 34468 89824 34524
rect 89872 34522 89928 34524
rect 89976 34522 90032 34524
rect 89872 34470 89896 34522
rect 89896 34470 89928 34522
rect 89976 34470 90020 34522
rect 90020 34470 90032 34522
rect 89872 34468 89928 34470
rect 89976 34468 90032 34470
rect 90080 34468 90136 34524
rect 90184 34522 90240 34524
rect 90288 34522 90344 34524
rect 90184 34470 90196 34522
rect 90196 34470 90240 34522
rect 90288 34470 90320 34522
rect 90320 34470 90344 34522
rect 90184 34468 90240 34470
rect 90288 34468 90344 34470
rect 90392 34468 90448 34524
rect 87388 34300 87444 34356
rect 85268 33684 85324 33740
rect 85372 33738 85428 33740
rect 85476 33738 85532 33740
rect 85372 33686 85396 33738
rect 85396 33686 85428 33738
rect 85476 33686 85520 33738
rect 85520 33686 85532 33738
rect 85372 33684 85428 33686
rect 85476 33684 85532 33686
rect 85580 33684 85636 33740
rect 85684 33738 85740 33740
rect 85788 33738 85844 33740
rect 85684 33686 85696 33738
rect 85696 33686 85740 33738
rect 85788 33686 85820 33738
rect 85820 33686 85844 33738
rect 85684 33684 85740 33686
rect 85788 33684 85844 33686
rect 85892 33684 85948 33740
rect 89768 32900 89824 32956
rect 89872 32954 89928 32956
rect 89976 32954 90032 32956
rect 89872 32902 89896 32954
rect 89896 32902 89928 32954
rect 89976 32902 90020 32954
rect 90020 32902 90032 32954
rect 89872 32900 89928 32902
rect 89976 32900 90032 32902
rect 90080 32900 90136 32956
rect 90184 32954 90240 32956
rect 90288 32954 90344 32956
rect 90184 32902 90196 32954
rect 90196 32902 90240 32954
rect 90288 32902 90320 32954
rect 90320 32902 90344 32954
rect 90184 32900 90240 32902
rect 90288 32900 90344 32902
rect 90392 32900 90448 32956
rect 85268 32116 85324 32172
rect 85372 32170 85428 32172
rect 85476 32170 85532 32172
rect 85372 32118 85396 32170
rect 85396 32118 85428 32170
rect 85476 32118 85520 32170
rect 85520 32118 85532 32170
rect 85372 32116 85428 32118
rect 85476 32116 85532 32118
rect 85580 32116 85636 32172
rect 85684 32170 85740 32172
rect 85788 32170 85844 32172
rect 85684 32118 85696 32170
rect 85696 32118 85740 32170
rect 85788 32118 85820 32170
rect 85820 32118 85844 32170
rect 85684 32116 85740 32118
rect 85788 32116 85844 32118
rect 85892 32116 85948 32172
rect 89768 31332 89824 31388
rect 89872 31386 89928 31388
rect 89976 31386 90032 31388
rect 89872 31334 89896 31386
rect 89896 31334 89928 31386
rect 89976 31334 90020 31386
rect 90020 31334 90032 31386
rect 89872 31332 89928 31334
rect 89976 31332 90032 31334
rect 90080 31332 90136 31388
rect 90184 31386 90240 31388
rect 90288 31386 90344 31388
rect 90184 31334 90196 31386
rect 90196 31334 90240 31386
rect 90288 31334 90320 31386
rect 90320 31334 90344 31386
rect 90184 31332 90240 31334
rect 90288 31332 90344 31334
rect 90392 31332 90448 31388
rect 85268 30548 85324 30604
rect 85372 30602 85428 30604
rect 85476 30602 85532 30604
rect 85372 30550 85396 30602
rect 85396 30550 85428 30602
rect 85476 30550 85520 30602
rect 85520 30550 85532 30602
rect 85372 30548 85428 30550
rect 85476 30548 85532 30550
rect 85580 30548 85636 30604
rect 85684 30602 85740 30604
rect 85788 30602 85844 30604
rect 85684 30550 85696 30602
rect 85696 30550 85740 30602
rect 85788 30550 85820 30602
rect 85820 30550 85844 30602
rect 85684 30548 85740 30550
rect 85788 30548 85844 30550
rect 85892 30548 85948 30604
rect 77420 30156 77476 30212
rect 75852 29426 75908 29428
rect 75852 29374 75854 29426
rect 75854 29374 75906 29426
rect 75906 29374 75908 29426
rect 75852 29372 75908 29374
rect 83468 30210 83524 30212
rect 83468 30158 83470 30210
rect 83470 30158 83522 30210
rect 83522 30158 83524 30210
rect 83468 30156 83524 30158
rect 84476 30210 84532 30212
rect 84476 30158 84478 30210
rect 84478 30158 84530 30210
rect 84530 30158 84532 30210
rect 84476 30156 84532 30158
rect 92428 35980 92484 36036
rect 92988 35922 93044 35924
rect 92988 35870 92990 35922
rect 92990 35870 93042 35922
rect 93042 35870 93044 35922
rect 92988 35868 93044 35870
rect 93772 35922 93828 35924
rect 93772 35870 93774 35922
rect 93774 35870 93826 35922
rect 93826 35870 93828 35922
rect 93772 35868 93828 35870
rect 96236 36988 96292 37044
rect 96236 36370 96292 36372
rect 96236 36318 96238 36370
rect 96238 36318 96290 36370
rect 96290 36318 96292 36370
rect 96236 36316 96292 36318
rect 96124 35868 96180 35924
rect 94268 35252 94324 35308
rect 94372 35306 94428 35308
rect 94476 35306 94532 35308
rect 94372 35254 94396 35306
rect 94396 35254 94428 35306
rect 94476 35254 94520 35306
rect 94520 35254 94532 35306
rect 94372 35252 94428 35254
rect 94476 35252 94532 35254
rect 94580 35252 94636 35308
rect 94684 35306 94740 35308
rect 94788 35306 94844 35308
rect 94684 35254 94696 35306
rect 94696 35254 94740 35306
rect 94788 35254 94820 35306
rect 94820 35254 94844 35306
rect 94684 35252 94740 35254
rect 94788 35252 94844 35254
rect 94892 35252 94948 35308
rect 96236 34802 96292 34804
rect 96236 34750 96238 34802
rect 96238 34750 96290 34802
rect 96290 34750 96292 34802
rect 96236 34748 96292 34750
rect 94268 33684 94324 33740
rect 94372 33738 94428 33740
rect 94476 33738 94532 33740
rect 94372 33686 94396 33738
rect 94396 33686 94428 33738
rect 94476 33686 94520 33738
rect 94520 33686 94532 33738
rect 94372 33684 94428 33686
rect 94476 33684 94532 33686
rect 94580 33684 94636 33740
rect 94684 33738 94740 33740
rect 94788 33738 94844 33740
rect 94684 33686 94696 33738
rect 94696 33686 94740 33738
rect 94788 33686 94820 33738
rect 94820 33686 94844 33738
rect 94684 33684 94740 33686
rect 94788 33684 94844 33686
rect 94892 33684 94948 33740
rect 94268 32116 94324 32172
rect 94372 32170 94428 32172
rect 94476 32170 94532 32172
rect 94372 32118 94396 32170
rect 94396 32118 94428 32170
rect 94476 32118 94520 32170
rect 94520 32118 94532 32170
rect 94372 32116 94428 32118
rect 94476 32116 94532 32118
rect 94580 32116 94636 32172
rect 94684 32170 94740 32172
rect 94788 32170 94844 32172
rect 94684 32118 94696 32170
rect 94696 32118 94740 32170
rect 94788 32118 94820 32170
rect 94820 32118 94844 32170
rect 94684 32116 94740 32118
rect 94788 32116 94844 32118
rect 94892 32116 94948 32172
rect 94268 30548 94324 30604
rect 94372 30602 94428 30604
rect 94476 30602 94532 30604
rect 94372 30550 94396 30602
rect 94396 30550 94428 30602
rect 94476 30550 94520 30602
rect 94520 30550 94532 30602
rect 94372 30548 94428 30550
rect 94476 30548 94532 30550
rect 94580 30548 94636 30604
rect 94684 30602 94740 30604
rect 94788 30602 94844 30604
rect 94684 30550 94696 30602
rect 94696 30550 94740 30602
rect 94788 30550 94820 30602
rect 94820 30550 94844 30602
rect 94684 30548 94740 30550
rect 94788 30548 94844 30550
rect 94892 30548 94948 30604
rect 91308 30156 91364 30212
rect 80768 29764 80824 29820
rect 80872 29818 80928 29820
rect 80976 29818 81032 29820
rect 80872 29766 80896 29818
rect 80896 29766 80928 29818
rect 80976 29766 81020 29818
rect 81020 29766 81032 29818
rect 80872 29764 80928 29766
rect 80976 29764 81032 29766
rect 81080 29764 81136 29820
rect 81184 29818 81240 29820
rect 81288 29818 81344 29820
rect 81184 29766 81196 29818
rect 81196 29766 81240 29818
rect 81288 29766 81320 29818
rect 81320 29766 81344 29818
rect 81184 29764 81240 29766
rect 81288 29764 81344 29766
rect 81392 29764 81448 29820
rect 89768 29764 89824 29820
rect 89872 29818 89928 29820
rect 89976 29818 90032 29820
rect 89872 29766 89896 29818
rect 89896 29766 89928 29818
rect 89976 29766 90020 29818
rect 90020 29766 90032 29818
rect 89872 29764 89928 29766
rect 89976 29764 90032 29766
rect 90080 29764 90136 29820
rect 90184 29818 90240 29820
rect 90288 29818 90344 29820
rect 90184 29766 90196 29818
rect 90196 29766 90240 29818
rect 90288 29766 90320 29818
rect 90320 29766 90344 29818
rect 90184 29764 90240 29766
rect 90288 29764 90344 29766
rect 90392 29764 90448 29820
rect 77420 29372 77476 29428
rect 76268 28980 76324 29036
rect 76372 29034 76428 29036
rect 76476 29034 76532 29036
rect 76372 28982 76396 29034
rect 76396 28982 76428 29034
rect 76476 28982 76520 29034
rect 76520 28982 76532 29034
rect 76372 28980 76428 28982
rect 76476 28980 76532 28982
rect 76580 28980 76636 29036
rect 76684 29034 76740 29036
rect 76788 29034 76844 29036
rect 76684 28982 76696 29034
rect 76696 28982 76740 29034
rect 76788 28982 76820 29034
rect 76820 28982 76844 29034
rect 76684 28980 76740 28982
rect 76788 28980 76844 28982
rect 76892 28980 76948 29036
rect 76076 28812 76132 28868
rect 75964 27804 76020 27860
rect 75964 27132 76020 27188
rect 76188 28364 76244 28420
rect 76524 27858 76580 27860
rect 76524 27806 76526 27858
rect 76526 27806 76578 27858
rect 76578 27806 76580 27858
rect 76524 27804 76580 27806
rect 76268 27412 76324 27468
rect 76372 27466 76428 27468
rect 76476 27466 76532 27468
rect 76372 27414 76396 27466
rect 76396 27414 76428 27466
rect 76476 27414 76520 27466
rect 76520 27414 76532 27466
rect 76372 27412 76428 27414
rect 76476 27412 76532 27414
rect 76580 27412 76636 27468
rect 76684 27466 76740 27468
rect 76788 27466 76844 27468
rect 76684 27414 76696 27466
rect 76696 27414 76740 27466
rect 76788 27414 76820 27466
rect 76820 27414 76844 27466
rect 76684 27412 76740 27414
rect 76788 27412 76844 27414
rect 76892 27412 76948 27468
rect 85268 28980 85324 29036
rect 85372 29034 85428 29036
rect 85476 29034 85532 29036
rect 85372 28982 85396 29034
rect 85396 28982 85428 29034
rect 85476 28982 85520 29034
rect 85520 28982 85532 29034
rect 85372 28980 85428 28982
rect 85476 28980 85532 28982
rect 85580 28980 85636 29036
rect 85684 29034 85740 29036
rect 85788 29034 85844 29036
rect 85684 28982 85696 29034
rect 85696 28982 85740 29034
rect 85788 28982 85820 29034
rect 85820 28982 85844 29034
rect 85684 28980 85740 28982
rect 85788 28980 85844 28982
rect 85892 28980 85948 29036
rect 94268 28980 94324 29036
rect 94372 29034 94428 29036
rect 94476 29034 94532 29036
rect 94372 28982 94396 29034
rect 94396 28982 94428 29034
rect 94476 28982 94520 29034
rect 94520 28982 94532 29034
rect 94372 28980 94428 28982
rect 94476 28980 94532 28982
rect 94580 28980 94636 29036
rect 94684 29034 94740 29036
rect 94788 29034 94844 29036
rect 94684 28982 94696 29034
rect 94696 28982 94740 29034
rect 94788 28982 94820 29034
rect 94820 28982 94844 29034
rect 94684 28980 94740 28982
rect 94788 28980 94844 28982
rect 94892 28980 94948 29036
rect 77756 28418 77812 28420
rect 77756 28366 77758 28418
rect 77758 28366 77810 28418
rect 77810 28366 77812 28418
rect 77756 28364 77812 28366
rect 80768 28196 80824 28252
rect 80872 28250 80928 28252
rect 80976 28250 81032 28252
rect 80872 28198 80896 28250
rect 80896 28198 80928 28250
rect 80976 28198 81020 28250
rect 81020 28198 81032 28250
rect 80872 28196 80928 28198
rect 80976 28196 81032 28198
rect 81080 28196 81136 28252
rect 81184 28250 81240 28252
rect 81288 28250 81344 28252
rect 81184 28198 81196 28250
rect 81196 28198 81240 28250
rect 81288 28198 81320 28250
rect 81320 28198 81344 28250
rect 81184 28196 81240 28198
rect 81288 28196 81344 28198
rect 81392 28196 81448 28252
rect 89768 28196 89824 28252
rect 89872 28250 89928 28252
rect 89976 28250 90032 28252
rect 89872 28198 89896 28250
rect 89896 28198 89928 28250
rect 89976 28198 90020 28250
rect 90020 28198 90032 28250
rect 89872 28196 89928 28198
rect 89976 28196 90032 28198
rect 90080 28196 90136 28252
rect 90184 28250 90240 28252
rect 90288 28250 90344 28252
rect 90184 28198 90196 28250
rect 90196 28198 90240 28250
rect 90288 28198 90320 28250
rect 90320 28198 90344 28250
rect 90184 28196 90240 28198
rect 90288 28196 90344 28198
rect 90392 28196 90448 28252
rect 98028 42364 98084 42420
rect 98028 40572 98084 40628
rect 98028 38780 98084 38836
rect 98028 36988 98084 37044
rect 97692 35196 97748 35252
rect 96572 34130 96628 34132
rect 96572 34078 96574 34130
rect 96574 34078 96626 34130
rect 96626 34078 96628 34130
rect 96572 34076 96628 34078
rect 97020 34130 97076 34132
rect 97020 34078 97022 34130
rect 97022 34078 97074 34130
rect 97074 34078 97076 34130
rect 97020 34076 97076 34078
rect 97692 33404 97748 33460
rect 98028 31666 98084 31668
rect 98028 31614 98030 31666
rect 98030 31614 98082 31666
rect 98082 31614 98084 31666
rect 98028 31612 98084 31614
rect 96684 31554 96740 31556
rect 96684 31502 96686 31554
rect 96686 31502 96738 31554
rect 96738 31502 96740 31554
rect 96684 31500 96740 31502
rect 96684 30098 96740 30100
rect 96684 30046 96686 30098
rect 96686 30046 96738 30098
rect 96738 30046 96740 30098
rect 96684 30044 96740 30046
rect 98028 29820 98084 29876
rect 96572 28642 96628 28644
rect 96572 28590 96574 28642
rect 96574 28590 96626 28642
rect 96626 28590 96628 28642
rect 96572 28588 96628 28590
rect 97020 28642 97076 28644
rect 97020 28590 97022 28642
rect 97022 28590 97074 28642
rect 97074 28590 97076 28642
rect 97020 28588 97076 28590
rect 96348 28028 96404 28084
rect 97692 28028 97748 28084
rect 77532 27580 77588 27636
rect 76412 27186 76468 27188
rect 76412 27134 76414 27186
rect 76414 27134 76466 27186
rect 76466 27134 76468 27186
rect 76412 27132 76468 27134
rect 75740 26178 75796 26180
rect 75740 26126 75742 26178
rect 75742 26126 75794 26178
rect 75794 26126 75796 26178
rect 75740 26124 75796 26126
rect 76524 26348 76580 26404
rect 77084 26402 77140 26404
rect 77084 26350 77086 26402
rect 77086 26350 77138 26402
rect 77138 26350 77140 26402
rect 77084 26348 77140 26350
rect 75964 26124 76020 26180
rect 76076 26012 76132 26068
rect 76268 25844 76324 25900
rect 76372 25898 76428 25900
rect 76476 25898 76532 25900
rect 76372 25846 76396 25898
rect 76396 25846 76428 25898
rect 76476 25846 76520 25898
rect 76520 25846 76532 25898
rect 76372 25844 76428 25846
rect 76476 25844 76532 25846
rect 76580 25844 76636 25900
rect 76684 25898 76740 25900
rect 76788 25898 76844 25900
rect 76684 25846 76696 25898
rect 76696 25846 76740 25898
rect 76788 25846 76820 25898
rect 76820 25846 76844 25898
rect 76684 25844 76740 25846
rect 76788 25844 76844 25846
rect 76892 25844 76948 25900
rect 77420 25506 77476 25508
rect 77420 25454 77422 25506
rect 77422 25454 77474 25506
rect 77474 25454 77476 25506
rect 77420 25452 77476 25454
rect 77644 26236 77700 26292
rect 75964 25340 76020 25396
rect 75740 24780 75796 24836
rect 75740 23884 75796 23940
rect 76268 24276 76324 24332
rect 76372 24330 76428 24332
rect 76476 24330 76532 24332
rect 76372 24278 76396 24330
rect 76396 24278 76428 24330
rect 76476 24278 76520 24330
rect 76520 24278 76532 24330
rect 76372 24276 76428 24278
rect 76476 24276 76532 24278
rect 76580 24276 76636 24332
rect 76684 24330 76740 24332
rect 76788 24330 76844 24332
rect 76684 24278 76696 24330
rect 76696 24278 76740 24330
rect 76788 24278 76820 24330
rect 76820 24278 76844 24330
rect 76684 24276 76740 24278
rect 76788 24276 76844 24278
rect 76892 24276 76948 24332
rect 76300 23938 76356 23940
rect 76300 23886 76302 23938
rect 76302 23886 76354 23938
rect 76354 23886 76356 23938
rect 76300 23884 76356 23886
rect 76636 23324 76692 23380
rect 77980 26178 78036 26180
rect 77980 26126 77982 26178
rect 77982 26126 78034 26178
rect 78034 26126 78036 26178
rect 77980 26124 78036 26126
rect 79660 27634 79716 27636
rect 79660 27582 79662 27634
rect 79662 27582 79714 27634
rect 79714 27582 79716 27634
rect 79660 27580 79716 27582
rect 84028 27580 84084 27636
rect 80768 26628 80824 26684
rect 80872 26682 80928 26684
rect 80976 26682 81032 26684
rect 80872 26630 80896 26682
rect 80896 26630 80928 26682
rect 80976 26630 81020 26682
rect 81020 26630 81032 26682
rect 80872 26628 80928 26630
rect 80976 26628 81032 26630
rect 81080 26628 81136 26684
rect 81184 26682 81240 26684
rect 81288 26682 81344 26684
rect 81184 26630 81196 26682
rect 81196 26630 81240 26682
rect 81288 26630 81320 26682
rect 81320 26630 81344 26682
rect 81184 26628 81240 26630
rect 81288 26628 81344 26630
rect 81392 26628 81448 26684
rect 85268 27412 85324 27468
rect 85372 27466 85428 27468
rect 85476 27466 85532 27468
rect 85372 27414 85396 27466
rect 85396 27414 85428 27466
rect 85476 27414 85520 27466
rect 85520 27414 85532 27466
rect 85372 27412 85428 27414
rect 85476 27412 85532 27414
rect 85580 27412 85636 27468
rect 85684 27466 85740 27468
rect 85788 27466 85844 27468
rect 85684 27414 85696 27466
rect 85696 27414 85740 27466
rect 85788 27414 85820 27466
rect 85820 27414 85844 27466
rect 85684 27412 85740 27414
rect 85788 27412 85844 27414
rect 85892 27412 85948 27468
rect 94268 27412 94324 27468
rect 94372 27466 94428 27468
rect 94476 27466 94532 27468
rect 94372 27414 94396 27466
rect 94396 27414 94428 27466
rect 94476 27414 94520 27466
rect 94520 27414 94532 27466
rect 94372 27412 94428 27414
rect 94476 27412 94532 27414
rect 94580 27412 94636 27468
rect 94684 27466 94740 27468
rect 94788 27466 94844 27468
rect 94684 27414 94696 27466
rect 94696 27414 94740 27466
rect 94788 27414 94820 27466
rect 94820 27414 94844 27466
rect 94684 27412 94740 27414
rect 94788 27412 94844 27414
rect 94892 27412 94948 27468
rect 96572 27244 96628 27300
rect 89768 26628 89824 26684
rect 89872 26682 89928 26684
rect 89976 26682 90032 26684
rect 89872 26630 89896 26682
rect 89896 26630 89928 26682
rect 89976 26630 90020 26682
rect 90020 26630 90032 26682
rect 89872 26628 89928 26630
rect 89976 26628 90032 26630
rect 90080 26628 90136 26684
rect 90184 26682 90240 26684
rect 90288 26682 90344 26684
rect 90184 26630 90196 26682
rect 90196 26630 90240 26682
rect 90288 26630 90320 26682
rect 90320 26630 90344 26682
rect 90184 26628 90240 26630
rect 90288 26628 90344 26630
rect 90392 26628 90448 26684
rect 84252 26402 84308 26404
rect 84252 26350 84254 26402
rect 84254 26350 84306 26402
rect 84306 26350 84308 26402
rect 84252 26348 84308 26350
rect 96908 26348 96964 26404
rect 78876 26124 78932 26180
rect 85268 25844 85324 25900
rect 85372 25898 85428 25900
rect 85476 25898 85532 25900
rect 85372 25846 85396 25898
rect 85396 25846 85428 25898
rect 85476 25846 85520 25898
rect 85520 25846 85532 25898
rect 85372 25844 85428 25846
rect 85476 25844 85532 25846
rect 85580 25844 85636 25900
rect 85684 25898 85740 25900
rect 85788 25898 85844 25900
rect 85684 25846 85696 25898
rect 85696 25846 85740 25898
rect 85788 25846 85820 25898
rect 85820 25846 85844 25898
rect 85684 25844 85740 25846
rect 85788 25844 85844 25846
rect 85892 25844 85948 25900
rect 94268 25844 94324 25900
rect 94372 25898 94428 25900
rect 94476 25898 94532 25900
rect 94372 25846 94396 25898
rect 94396 25846 94428 25898
rect 94476 25846 94520 25898
rect 94520 25846 94532 25898
rect 94372 25844 94428 25846
rect 94476 25844 94532 25846
rect 94580 25844 94636 25900
rect 94684 25898 94740 25900
rect 94788 25898 94844 25900
rect 94684 25846 94696 25898
rect 94696 25846 94740 25898
rect 94788 25846 94820 25898
rect 94820 25846 94844 25898
rect 94684 25844 94740 25846
rect 94788 25844 94844 25846
rect 94892 25844 94948 25900
rect 78876 25564 78932 25620
rect 78092 24946 78148 24948
rect 78092 24894 78094 24946
rect 78094 24894 78146 24946
rect 78146 24894 78148 24946
rect 78092 24892 78148 24894
rect 78764 25506 78820 25508
rect 78764 25454 78766 25506
rect 78766 25454 78818 25506
rect 78818 25454 78820 25506
rect 78764 25452 78820 25454
rect 81116 25394 81172 25396
rect 81116 25342 81118 25394
rect 81118 25342 81170 25394
rect 81170 25342 81172 25394
rect 81116 25340 81172 25342
rect 80768 25060 80824 25116
rect 80872 25114 80928 25116
rect 80976 25114 81032 25116
rect 80872 25062 80896 25114
rect 80896 25062 80928 25114
rect 80976 25062 81020 25114
rect 81020 25062 81032 25114
rect 80872 25060 80928 25062
rect 80976 25060 81032 25062
rect 81080 25060 81136 25116
rect 81184 25114 81240 25116
rect 81288 25114 81344 25116
rect 81184 25062 81196 25114
rect 81196 25062 81240 25114
rect 81288 25062 81320 25114
rect 81320 25062 81344 25114
rect 81184 25060 81240 25062
rect 81288 25060 81344 25062
rect 81392 25060 81448 25116
rect 89768 25060 89824 25116
rect 89872 25114 89928 25116
rect 89976 25114 90032 25116
rect 89872 25062 89896 25114
rect 89896 25062 89928 25114
rect 89976 25062 90020 25114
rect 90020 25062 90032 25114
rect 89872 25060 89928 25062
rect 89976 25060 90032 25062
rect 90080 25060 90136 25116
rect 90184 25114 90240 25116
rect 90288 25114 90344 25116
rect 90184 25062 90196 25114
rect 90196 25062 90240 25114
rect 90288 25062 90320 25114
rect 90320 25062 90344 25114
rect 90184 25060 90240 25062
rect 90288 25060 90344 25062
rect 90392 25060 90448 25116
rect 81900 24892 81956 24948
rect 83132 24892 83188 24948
rect 80768 23492 80824 23548
rect 80872 23546 80928 23548
rect 80976 23546 81032 23548
rect 80872 23494 80896 23546
rect 80896 23494 80928 23546
rect 80976 23494 81020 23546
rect 81020 23494 81032 23546
rect 80872 23492 80928 23494
rect 80976 23492 81032 23494
rect 81080 23492 81136 23548
rect 81184 23546 81240 23548
rect 81288 23546 81344 23548
rect 81184 23494 81196 23546
rect 81196 23494 81240 23546
rect 81288 23494 81320 23546
rect 81320 23494 81344 23546
rect 81184 23492 81240 23494
rect 81288 23492 81344 23494
rect 81392 23492 81448 23548
rect 77756 23266 77812 23268
rect 77756 23214 77758 23266
rect 77758 23214 77810 23266
rect 77810 23214 77812 23266
rect 77756 23212 77812 23214
rect 78428 23154 78484 23156
rect 78428 23102 78430 23154
rect 78430 23102 78482 23154
rect 78482 23102 78484 23154
rect 78428 23100 78484 23102
rect 76268 22708 76324 22764
rect 76372 22762 76428 22764
rect 76476 22762 76532 22764
rect 76372 22710 76396 22762
rect 76396 22710 76428 22762
rect 76476 22710 76520 22762
rect 76520 22710 76532 22762
rect 76372 22708 76428 22710
rect 76476 22708 76532 22710
rect 76580 22708 76636 22764
rect 76684 22762 76740 22764
rect 76788 22762 76844 22764
rect 76684 22710 76696 22762
rect 76696 22710 76740 22762
rect 76788 22710 76820 22762
rect 76820 22710 76844 22762
rect 76684 22708 76740 22710
rect 76788 22708 76844 22710
rect 76892 22708 76948 22764
rect 75404 22316 75460 22372
rect 75628 22428 75684 22484
rect 75404 21980 75460 22036
rect 75292 21586 75348 21588
rect 75292 21534 75294 21586
rect 75294 21534 75346 21586
rect 75346 21534 75348 21586
rect 75292 21532 75348 21534
rect 73724 20914 73780 20916
rect 73724 20862 73726 20914
rect 73726 20862 73778 20914
rect 73778 20862 73780 20914
rect 73724 20860 73780 20862
rect 74172 20860 74228 20916
rect 74956 20524 75012 20580
rect 74396 20076 74452 20132
rect 74956 19852 75012 19908
rect 74396 19458 74452 19460
rect 74396 19406 74398 19458
rect 74398 19406 74450 19458
rect 74450 19406 74452 19458
rect 74396 19404 74452 19406
rect 71484 19068 71540 19124
rect 73836 19292 73892 19348
rect 75180 19404 75236 19460
rect 74732 19346 74788 19348
rect 74732 19294 74734 19346
rect 74734 19294 74786 19346
rect 74786 19294 74788 19346
rect 74732 19292 74788 19294
rect 71768 18788 71824 18844
rect 71872 18842 71928 18844
rect 71976 18842 72032 18844
rect 71872 18790 71896 18842
rect 71896 18790 71928 18842
rect 71976 18790 72020 18842
rect 72020 18790 72032 18842
rect 71872 18788 71928 18790
rect 71976 18788 72032 18790
rect 72080 18788 72136 18844
rect 72184 18842 72240 18844
rect 72288 18842 72344 18844
rect 72184 18790 72196 18842
rect 72196 18790 72240 18842
rect 72288 18790 72320 18842
rect 72320 18790 72344 18842
rect 72184 18788 72240 18790
rect 72288 18788 72344 18790
rect 72392 18788 72448 18844
rect 76300 22482 76356 22484
rect 76300 22430 76302 22482
rect 76302 22430 76354 22482
rect 76354 22430 76356 22482
rect 76300 22428 76356 22430
rect 77756 22482 77812 22484
rect 77756 22430 77758 22482
rect 77758 22430 77810 22482
rect 77810 22430 77812 22482
rect 77756 22428 77812 22430
rect 77756 22092 77812 22148
rect 80220 23100 80276 23156
rect 82572 23212 82628 23268
rect 82124 23154 82180 23156
rect 82124 23102 82126 23154
rect 82126 23102 82178 23154
rect 82178 23102 82180 23154
rect 82124 23100 82180 23102
rect 81452 22540 81508 22596
rect 82572 22370 82628 22372
rect 82572 22318 82574 22370
rect 82574 22318 82626 22370
rect 82626 22318 82628 22370
rect 82572 22316 82628 22318
rect 82684 22204 82740 22260
rect 83356 23154 83412 23156
rect 83356 23102 83358 23154
rect 83358 23102 83410 23154
rect 83410 23102 83412 23154
rect 83356 23100 83412 23102
rect 80892 22146 80948 22148
rect 80892 22094 80894 22146
rect 80894 22094 80946 22146
rect 80946 22094 80948 22146
rect 80892 22092 80948 22094
rect 80768 21924 80824 21980
rect 80872 21978 80928 21980
rect 80976 21978 81032 21980
rect 80872 21926 80896 21978
rect 80896 21926 80928 21978
rect 80976 21926 81020 21978
rect 81020 21926 81032 21978
rect 80872 21924 80928 21926
rect 80976 21924 81032 21926
rect 81080 21924 81136 21980
rect 81184 21978 81240 21980
rect 81288 21978 81344 21980
rect 81184 21926 81196 21978
rect 81196 21926 81240 21978
rect 81288 21926 81320 21978
rect 81320 21926 81344 21978
rect 81184 21924 81240 21926
rect 81288 21924 81344 21926
rect 81392 21924 81448 21980
rect 75740 21644 75796 21700
rect 77756 21644 77812 21700
rect 75852 21532 75908 21588
rect 76268 21140 76324 21196
rect 76372 21194 76428 21196
rect 76476 21194 76532 21196
rect 76372 21142 76396 21194
rect 76396 21142 76428 21194
rect 76476 21142 76520 21194
rect 76520 21142 76532 21194
rect 76372 21140 76428 21142
rect 76476 21140 76532 21142
rect 76580 21140 76636 21196
rect 76684 21194 76740 21196
rect 76788 21194 76844 21196
rect 76684 21142 76696 21194
rect 76696 21142 76740 21194
rect 76788 21142 76820 21194
rect 76820 21142 76844 21194
rect 76684 21140 76740 21142
rect 76788 21140 76844 21142
rect 76892 21140 76948 21196
rect 76300 20242 76356 20244
rect 76300 20190 76302 20242
rect 76302 20190 76354 20242
rect 76354 20190 76356 20242
rect 76300 20188 76356 20190
rect 78764 21532 78820 21588
rect 75628 19346 75684 19348
rect 75628 19294 75630 19346
rect 75630 19294 75682 19346
rect 75682 19294 75684 19346
rect 75628 19292 75684 19294
rect 76972 20018 77028 20020
rect 76972 19966 76974 20018
rect 76974 19966 77026 20018
rect 77026 19966 77028 20018
rect 76972 19964 77028 19966
rect 76524 19852 76580 19908
rect 77420 19906 77476 19908
rect 77420 19854 77422 19906
rect 77422 19854 77474 19906
rect 77474 19854 77476 19906
rect 77420 19852 77476 19854
rect 76268 19572 76324 19628
rect 76372 19626 76428 19628
rect 76476 19626 76532 19628
rect 76372 19574 76396 19626
rect 76396 19574 76428 19626
rect 76476 19574 76520 19626
rect 76520 19574 76532 19626
rect 76372 19572 76428 19574
rect 76476 19572 76532 19574
rect 76580 19572 76636 19628
rect 76684 19626 76740 19628
rect 76788 19626 76844 19628
rect 76684 19574 76696 19626
rect 76696 19574 76740 19626
rect 76788 19574 76820 19626
rect 76820 19574 76844 19626
rect 76684 19572 76740 19574
rect 76788 19572 76844 19574
rect 76892 19572 76948 19628
rect 71768 17220 71824 17276
rect 71872 17274 71928 17276
rect 71976 17274 72032 17276
rect 71872 17222 71896 17274
rect 71896 17222 71928 17274
rect 71976 17222 72020 17274
rect 72020 17222 72032 17274
rect 71872 17220 71928 17222
rect 71976 17220 72032 17222
rect 72080 17220 72136 17276
rect 72184 17274 72240 17276
rect 72288 17274 72344 17276
rect 72184 17222 72196 17274
rect 72196 17222 72240 17274
rect 72288 17222 72320 17274
rect 72320 17222 72344 17274
rect 72184 17220 72240 17222
rect 72288 17220 72344 17222
rect 72392 17220 72448 17276
rect 71768 15652 71824 15708
rect 71872 15706 71928 15708
rect 71976 15706 72032 15708
rect 71872 15654 71896 15706
rect 71896 15654 71928 15706
rect 71976 15654 72020 15706
rect 72020 15654 72032 15706
rect 71872 15652 71928 15654
rect 71976 15652 72032 15654
rect 72080 15652 72136 15708
rect 72184 15706 72240 15708
rect 72288 15706 72344 15708
rect 72184 15654 72196 15706
rect 72196 15654 72240 15706
rect 72288 15654 72320 15706
rect 72320 15654 72344 15706
rect 72184 15652 72240 15654
rect 72288 15652 72344 15654
rect 72392 15652 72448 15708
rect 70812 13804 70868 13860
rect 71768 14084 71824 14140
rect 71872 14138 71928 14140
rect 71976 14138 72032 14140
rect 71872 14086 71896 14138
rect 71896 14086 71928 14138
rect 71976 14086 72020 14138
rect 72020 14086 72032 14138
rect 71872 14084 71928 14086
rect 71976 14084 72032 14086
rect 72080 14084 72136 14140
rect 72184 14138 72240 14140
rect 72288 14138 72344 14140
rect 72184 14086 72196 14138
rect 72196 14086 72240 14138
rect 72288 14086 72320 14138
rect 72320 14086 72344 14138
rect 72184 14084 72240 14086
rect 72288 14084 72344 14086
rect 72392 14084 72448 14140
rect 72268 13858 72324 13860
rect 72268 13806 72270 13858
rect 72270 13806 72322 13858
rect 72322 13806 72324 13858
rect 72268 13804 72324 13806
rect 71768 12516 71824 12572
rect 71872 12570 71928 12572
rect 71976 12570 72032 12572
rect 71872 12518 71896 12570
rect 71896 12518 71928 12570
rect 71976 12518 72020 12570
rect 72020 12518 72032 12570
rect 71872 12516 71928 12518
rect 71976 12516 72032 12518
rect 72080 12516 72136 12572
rect 72184 12570 72240 12572
rect 72288 12570 72344 12572
rect 72184 12518 72196 12570
rect 72196 12518 72240 12570
rect 72288 12518 72320 12570
rect 72320 12518 72344 12570
rect 72184 12516 72240 12518
rect 72288 12516 72344 12518
rect 72392 12516 72448 12572
rect 72828 12236 72884 12292
rect 71372 12012 71428 12068
rect 70028 4956 70084 5012
rect 70924 8876 70980 8932
rect 70812 7868 70868 7924
rect 70028 4060 70084 4116
rect 70812 6188 70868 6244
rect 71036 8092 71092 8148
rect 71148 6636 71204 6692
rect 70812 5794 70868 5796
rect 70812 5742 70814 5794
rect 70814 5742 70866 5794
rect 70866 5742 70868 5794
rect 70812 5740 70868 5742
rect 70924 5628 70980 5684
rect 70700 4844 70756 4900
rect 70364 3612 70420 3668
rect 71036 3666 71092 3668
rect 71036 3614 71038 3666
rect 71038 3614 71090 3666
rect 71090 3614 71092 3666
rect 71036 3612 71092 3614
rect 72492 12066 72548 12068
rect 72492 12014 72494 12066
rect 72494 12014 72546 12066
rect 72546 12014 72548 12066
rect 72492 12012 72548 12014
rect 71768 10948 71824 11004
rect 71872 11002 71928 11004
rect 71976 11002 72032 11004
rect 71872 10950 71896 11002
rect 71896 10950 71928 11002
rect 71976 10950 72020 11002
rect 72020 10950 72032 11002
rect 71872 10948 71928 10950
rect 71976 10948 72032 10950
rect 72080 10948 72136 11004
rect 72184 11002 72240 11004
rect 72288 11002 72344 11004
rect 72184 10950 72196 11002
rect 72196 10950 72240 11002
rect 72288 10950 72320 11002
rect 72320 10950 72344 11002
rect 72184 10948 72240 10950
rect 72288 10948 72344 10950
rect 72392 10948 72448 11004
rect 71768 9380 71824 9436
rect 71872 9434 71928 9436
rect 71976 9434 72032 9436
rect 71872 9382 71896 9434
rect 71896 9382 71928 9434
rect 71976 9382 72020 9434
rect 72020 9382 72032 9434
rect 71872 9380 71928 9382
rect 71976 9380 72032 9382
rect 72080 9380 72136 9436
rect 72184 9434 72240 9436
rect 72288 9434 72344 9436
rect 72184 9382 72196 9434
rect 72196 9382 72240 9434
rect 72288 9382 72320 9434
rect 72320 9382 72344 9434
rect 72184 9380 72240 9382
rect 72288 9380 72344 9382
rect 72392 9380 72448 9436
rect 71372 5292 71428 5348
rect 72492 8930 72548 8932
rect 72492 8878 72494 8930
rect 72494 8878 72546 8930
rect 72546 8878 72548 8930
rect 72492 8876 72548 8878
rect 71768 7812 71824 7868
rect 71872 7866 71928 7868
rect 71976 7866 72032 7868
rect 71872 7814 71896 7866
rect 71896 7814 71928 7866
rect 71976 7814 72020 7866
rect 72020 7814 72032 7866
rect 71872 7812 71928 7814
rect 71976 7812 72032 7814
rect 72080 7812 72136 7868
rect 72184 7866 72240 7868
rect 72288 7866 72344 7868
rect 72184 7814 72196 7866
rect 72196 7814 72240 7866
rect 72288 7814 72320 7866
rect 72320 7814 72344 7866
rect 72184 7812 72240 7814
rect 72288 7812 72344 7814
rect 72392 7812 72448 7868
rect 71596 6412 71652 6468
rect 71768 6244 71824 6300
rect 71872 6298 71928 6300
rect 71976 6298 72032 6300
rect 71872 6246 71896 6298
rect 71896 6246 71928 6298
rect 71976 6246 72020 6298
rect 72020 6246 72032 6298
rect 71872 6244 71928 6246
rect 71976 6244 72032 6246
rect 72080 6244 72136 6300
rect 72184 6298 72240 6300
rect 72288 6298 72344 6300
rect 72184 6246 72196 6298
rect 72196 6246 72240 6298
rect 72288 6246 72320 6298
rect 72320 6246 72344 6298
rect 72184 6244 72240 6246
rect 72288 6244 72344 6246
rect 72392 6244 72448 6300
rect 71708 6076 71764 6132
rect 72492 6018 72548 6020
rect 72492 5966 72494 6018
rect 72494 5966 72546 6018
rect 72546 5966 72548 6018
rect 72492 5964 72548 5966
rect 73612 8988 73668 9044
rect 72828 7980 72884 8036
rect 72604 5628 72660 5684
rect 71768 4676 71824 4732
rect 71872 4730 71928 4732
rect 71976 4730 72032 4732
rect 71872 4678 71896 4730
rect 71896 4678 71928 4730
rect 71976 4678 72020 4730
rect 72020 4678 72032 4730
rect 71872 4676 71928 4678
rect 71976 4676 72032 4678
rect 72080 4676 72136 4732
rect 72184 4730 72240 4732
rect 72288 4730 72344 4732
rect 72184 4678 72196 4730
rect 72196 4678 72240 4730
rect 72288 4678 72320 4730
rect 72320 4678 72344 4730
rect 72184 4676 72240 4678
rect 72288 4676 72344 4678
rect 72392 4676 72448 4732
rect 71708 4226 71764 4228
rect 71708 4174 71710 4226
rect 71710 4174 71762 4226
rect 71762 4174 71764 4226
rect 71708 4172 71764 4174
rect 71596 4114 71652 4116
rect 71596 4062 71598 4114
rect 71598 4062 71650 4114
rect 71650 4062 71652 4114
rect 71596 4060 71652 4062
rect 71596 3500 71652 3556
rect 69692 3442 69748 3444
rect 69692 3390 69694 3442
rect 69694 3390 69746 3442
rect 69746 3390 69748 3442
rect 69692 3388 69748 3390
rect 53768 3108 53824 3164
rect 53872 3162 53928 3164
rect 53976 3162 54032 3164
rect 53872 3110 53896 3162
rect 53896 3110 53928 3162
rect 53976 3110 54020 3162
rect 54020 3110 54032 3162
rect 53872 3108 53928 3110
rect 53976 3108 54032 3110
rect 54080 3108 54136 3164
rect 54184 3162 54240 3164
rect 54288 3162 54344 3164
rect 54184 3110 54196 3162
rect 54196 3110 54240 3162
rect 54288 3110 54320 3162
rect 54320 3110 54344 3162
rect 54184 3108 54240 3110
rect 54288 3108 54344 3110
rect 54392 3108 54448 3164
rect 62768 3108 62824 3164
rect 62872 3162 62928 3164
rect 62976 3162 63032 3164
rect 62872 3110 62896 3162
rect 62896 3110 62928 3162
rect 62976 3110 63020 3162
rect 63020 3110 63032 3162
rect 62872 3108 62928 3110
rect 62976 3108 63032 3110
rect 63080 3108 63136 3164
rect 63184 3162 63240 3164
rect 63288 3162 63344 3164
rect 63184 3110 63196 3162
rect 63196 3110 63240 3162
rect 63288 3110 63320 3162
rect 63320 3110 63344 3162
rect 63184 3108 63240 3110
rect 63288 3108 63344 3110
rect 63392 3108 63448 3164
rect 71932 3388 71988 3444
rect 74060 13746 74116 13748
rect 74060 13694 74062 13746
rect 74062 13694 74114 13746
rect 74114 13694 74116 13746
rect 74060 13692 74116 13694
rect 76268 18004 76324 18060
rect 76372 18058 76428 18060
rect 76476 18058 76532 18060
rect 76372 18006 76396 18058
rect 76396 18006 76428 18058
rect 76476 18006 76520 18058
rect 76520 18006 76532 18058
rect 76372 18004 76428 18006
rect 76476 18004 76532 18006
rect 76580 18004 76636 18060
rect 76684 18058 76740 18060
rect 76788 18058 76844 18060
rect 76684 18006 76696 18058
rect 76696 18006 76740 18058
rect 76788 18006 76820 18058
rect 76820 18006 76844 18058
rect 76684 18004 76740 18006
rect 76788 18004 76844 18006
rect 76892 18004 76948 18060
rect 76268 16436 76324 16492
rect 76372 16490 76428 16492
rect 76476 16490 76532 16492
rect 76372 16438 76396 16490
rect 76396 16438 76428 16490
rect 76476 16438 76520 16490
rect 76520 16438 76532 16490
rect 76372 16436 76428 16438
rect 76476 16436 76532 16438
rect 76580 16436 76636 16492
rect 76684 16490 76740 16492
rect 76788 16490 76844 16492
rect 76684 16438 76696 16490
rect 76696 16438 76740 16490
rect 76788 16438 76820 16490
rect 76820 16438 76844 16490
rect 76684 16436 76740 16438
rect 76788 16436 76844 16438
rect 76892 16436 76948 16492
rect 76268 14868 76324 14924
rect 76372 14922 76428 14924
rect 76476 14922 76532 14924
rect 76372 14870 76396 14922
rect 76396 14870 76428 14922
rect 76476 14870 76520 14922
rect 76520 14870 76532 14922
rect 76372 14868 76428 14870
rect 76476 14868 76532 14870
rect 76580 14868 76636 14924
rect 76684 14922 76740 14924
rect 76788 14922 76844 14924
rect 76684 14870 76696 14922
rect 76696 14870 76740 14922
rect 76788 14870 76820 14922
rect 76820 14870 76844 14922
rect 76684 14868 76740 14870
rect 76788 14868 76844 14870
rect 76892 14868 76948 14924
rect 74844 13580 74900 13636
rect 77756 14028 77812 14084
rect 73836 12684 73892 12740
rect 74284 12738 74340 12740
rect 74284 12686 74286 12738
rect 74286 12686 74338 12738
rect 74338 12686 74340 12738
rect 74284 12684 74340 12686
rect 73948 6690 74004 6692
rect 73948 6638 73950 6690
rect 73950 6638 74002 6690
rect 74002 6638 74004 6690
rect 73948 6636 74004 6638
rect 74620 6860 74676 6916
rect 73948 6412 74004 6468
rect 74508 6466 74564 6468
rect 74508 6414 74510 6466
rect 74510 6414 74562 6466
rect 74562 6414 74564 6466
rect 74508 6412 74564 6414
rect 74508 5404 74564 5460
rect 74844 6076 74900 6132
rect 74508 5180 74564 5236
rect 73724 5068 73780 5124
rect 73276 4284 73332 4340
rect 74396 4060 74452 4116
rect 74284 3666 74340 3668
rect 74284 3614 74286 3666
rect 74286 3614 74338 3666
rect 74338 3614 74340 3666
rect 74284 3612 74340 3614
rect 73276 3442 73332 3444
rect 73276 3390 73278 3442
rect 73278 3390 73330 3442
rect 73330 3390 73332 3442
rect 73276 3388 73332 3390
rect 75516 13580 75572 13636
rect 76268 13300 76324 13356
rect 76372 13354 76428 13356
rect 76476 13354 76532 13356
rect 76372 13302 76396 13354
rect 76396 13302 76428 13354
rect 76476 13302 76520 13354
rect 76520 13302 76532 13354
rect 76372 13300 76428 13302
rect 76476 13300 76532 13302
rect 76580 13300 76636 13356
rect 76684 13354 76740 13356
rect 76788 13354 76844 13356
rect 76684 13302 76696 13354
rect 76696 13302 76740 13354
rect 76788 13302 76820 13354
rect 76820 13302 76844 13354
rect 76684 13300 76740 13302
rect 76788 13300 76844 13302
rect 76892 13300 76948 13356
rect 75068 10668 75124 10724
rect 76268 11732 76324 11788
rect 76372 11786 76428 11788
rect 76476 11786 76532 11788
rect 76372 11734 76396 11786
rect 76396 11734 76428 11786
rect 76476 11734 76520 11786
rect 76520 11734 76532 11786
rect 76372 11732 76428 11734
rect 76476 11732 76532 11734
rect 76580 11732 76636 11788
rect 76684 11786 76740 11788
rect 76788 11786 76844 11788
rect 76684 11734 76696 11786
rect 76696 11734 76740 11786
rect 76788 11734 76820 11786
rect 76820 11734 76844 11786
rect 76684 11732 76740 11734
rect 76788 11732 76844 11734
rect 76892 11732 76948 11788
rect 76076 10722 76132 10724
rect 76076 10670 76078 10722
rect 76078 10670 76130 10722
rect 76130 10670 76132 10722
rect 76076 10668 76132 10670
rect 76268 10164 76324 10220
rect 76372 10218 76428 10220
rect 76476 10218 76532 10220
rect 76372 10166 76396 10218
rect 76396 10166 76428 10218
rect 76476 10166 76520 10218
rect 76520 10166 76532 10218
rect 76372 10164 76428 10166
rect 76476 10164 76532 10166
rect 76580 10164 76636 10220
rect 76684 10218 76740 10220
rect 76788 10218 76844 10220
rect 76684 10166 76696 10218
rect 76696 10166 76740 10218
rect 76788 10166 76820 10218
rect 76820 10166 76844 10218
rect 76684 10164 76740 10166
rect 76788 10164 76844 10166
rect 76892 10164 76948 10220
rect 77308 13746 77364 13748
rect 77308 13694 77310 13746
rect 77310 13694 77362 13746
rect 77362 13694 77364 13746
rect 77308 13692 77364 13694
rect 77196 9100 77252 9156
rect 76076 9042 76132 9044
rect 76076 8990 76078 9042
rect 76078 8990 76130 9042
rect 76130 8990 76132 9042
rect 76076 8988 76132 8990
rect 76268 8596 76324 8652
rect 76372 8650 76428 8652
rect 76476 8650 76532 8652
rect 76372 8598 76396 8650
rect 76396 8598 76428 8650
rect 76476 8598 76520 8650
rect 76520 8598 76532 8650
rect 76372 8596 76428 8598
rect 76476 8596 76532 8598
rect 76580 8596 76636 8652
rect 76684 8650 76740 8652
rect 76788 8650 76844 8652
rect 76684 8598 76696 8650
rect 76696 8598 76740 8650
rect 76788 8598 76820 8650
rect 76820 8598 76844 8650
rect 76684 8596 76740 8598
rect 76788 8596 76844 8598
rect 76892 8596 76948 8652
rect 76412 8146 76468 8148
rect 76412 8094 76414 8146
rect 76414 8094 76466 8146
rect 76466 8094 76468 8146
rect 76412 8092 76468 8094
rect 77196 7474 77252 7476
rect 77196 7422 77198 7474
rect 77198 7422 77250 7474
rect 77250 7422 77252 7474
rect 77196 7420 77252 7422
rect 76268 7028 76324 7084
rect 76372 7082 76428 7084
rect 76476 7082 76532 7084
rect 76372 7030 76396 7082
rect 76396 7030 76428 7082
rect 76476 7030 76520 7082
rect 76520 7030 76532 7082
rect 76372 7028 76428 7030
rect 76476 7028 76532 7030
rect 76580 7028 76636 7084
rect 76684 7082 76740 7084
rect 76788 7082 76844 7084
rect 76684 7030 76696 7082
rect 76696 7030 76740 7082
rect 76788 7030 76820 7082
rect 76820 7030 76844 7082
rect 76684 7028 76740 7030
rect 76788 7028 76844 7030
rect 76892 7028 76948 7084
rect 77084 6748 77140 6804
rect 75516 6524 75572 6580
rect 75404 6466 75460 6468
rect 75404 6414 75406 6466
rect 75406 6414 75458 6466
rect 75458 6414 75460 6466
rect 75404 6412 75460 6414
rect 75292 4172 75348 4228
rect 74956 3724 75012 3780
rect 76188 5964 76244 6020
rect 75628 4450 75684 4452
rect 75628 4398 75630 4450
rect 75630 4398 75682 4450
rect 75682 4398 75684 4450
rect 75628 4396 75684 4398
rect 74396 3388 74452 3444
rect 75852 3388 75908 3444
rect 76268 5460 76324 5516
rect 76372 5514 76428 5516
rect 76476 5514 76532 5516
rect 76372 5462 76396 5514
rect 76396 5462 76428 5514
rect 76476 5462 76520 5514
rect 76520 5462 76532 5514
rect 76372 5460 76428 5462
rect 76476 5460 76532 5462
rect 76580 5460 76636 5516
rect 76684 5514 76740 5516
rect 76788 5514 76844 5516
rect 76684 5462 76696 5514
rect 76696 5462 76740 5514
rect 76788 5462 76820 5514
rect 76820 5462 76844 5514
rect 76684 5460 76740 5462
rect 76788 5460 76844 5462
rect 76892 5460 76948 5516
rect 76268 3892 76324 3948
rect 76372 3946 76428 3948
rect 76476 3946 76532 3948
rect 76372 3894 76396 3946
rect 76396 3894 76428 3946
rect 76476 3894 76520 3946
rect 76520 3894 76532 3946
rect 76372 3892 76428 3894
rect 76476 3892 76532 3894
rect 76580 3892 76636 3948
rect 76684 3946 76740 3948
rect 76788 3946 76844 3948
rect 76684 3894 76696 3946
rect 76696 3894 76740 3946
rect 76788 3894 76820 3946
rect 76820 3894 76844 3946
rect 76684 3892 76740 3894
rect 76788 3892 76844 3894
rect 76892 3892 76948 3948
rect 77308 5404 77364 5460
rect 77644 4172 77700 4228
rect 77756 13804 77812 13860
rect 78092 20130 78148 20132
rect 78092 20078 78094 20130
rect 78094 20078 78146 20130
rect 78146 20078 78148 20130
rect 78092 20076 78148 20078
rect 80556 21586 80612 21588
rect 80556 21534 80558 21586
rect 80558 21534 80610 21586
rect 80610 21534 80612 21586
rect 80556 21532 80612 21534
rect 80444 21196 80500 21252
rect 81004 21586 81060 21588
rect 81004 21534 81006 21586
rect 81006 21534 81058 21586
rect 81058 21534 81060 21586
rect 81004 21532 81060 21534
rect 81564 21532 81620 21588
rect 80108 20188 80164 20244
rect 80768 20356 80824 20412
rect 80872 20410 80928 20412
rect 80976 20410 81032 20412
rect 80872 20358 80896 20410
rect 80896 20358 80928 20410
rect 80976 20358 81020 20410
rect 81020 20358 81032 20410
rect 80872 20356 80928 20358
rect 80976 20356 81032 20358
rect 81080 20356 81136 20412
rect 81184 20410 81240 20412
rect 81288 20410 81344 20412
rect 81184 20358 81196 20410
rect 81196 20358 81240 20410
rect 81288 20358 81320 20410
rect 81320 20358 81344 20410
rect 81184 20356 81240 20358
rect 81288 20356 81344 20358
rect 81392 20356 81448 20412
rect 79772 20076 79828 20132
rect 77980 19964 78036 20020
rect 79212 19292 79268 19348
rect 79212 19010 79268 19012
rect 79212 18958 79214 19010
rect 79214 18958 79266 19010
rect 79266 18958 79268 19010
rect 79212 18956 79268 18958
rect 79660 18956 79716 19012
rect 81676 21196 81732 21252
rect 82684 21196 82740 21252
rect 81900 20242 81956 20244
rect 81900 20190 81902 20242
rect 81902 20190 81954 20242
rect 81954 20190 81956 20242
rect 81900 20188 81956 20190
rect 81564 20076 81620 20132
rect 80668 19852 80724 19908
rect 80444 19740 80500 19796
rect 81676 20018 81732 20020
rect 81676 19966 81678 20018
rect 81678 19966 81730 20018
rect 81730 19966 81732 20018
rect 81676 19964 81732 19966
rect 81004 19740 81060 19796
rect 80768 18788 80824 18844
rect 80872 18842 80928 18844
rect 80976 18842 81032 18844
rect 80872 18790 80896 18842
rect 80896 18790 80928 18842
rect 80976 18790 81020 18842
rect 81020 18790 81032 18842
rect 80872 18788 80928 18790
rect 80976 18788 81032 18790
rect 81080 18788 81136 18844
rect 81184 18842 81240 18844
rect 81288 18842 81344 18844
rect 81184 18790 81196 18842
rect 81196 18790 81240 18842
rect 81288 18790 81320 18842
rect 81320 18790 81344 18842
rect 81184 18788 81240 18790
rect 81288 18788 81344 18790
rect 81392 18788 81448 18844
rect 78428 14028 78484 14084
rect 78652 13692 78708 13748
rect 78204 10722 78260 10724
rect 78204 10670 78206 10722
rect 78206 10670 78258 10722
rect 78258 10670 78260 10722
rect 78204 10668 78260 10670
rect 78204 6578 78260 6580
rect 78204 6526 78206 6578
rect 78206 6526 78258 6578
rect 78258 6526 78260 6578
rect 78204 6524 78260 6526
rect 77980 5404 78036 5460
rect 78540 6130 78596 6132
rect 78540 6078 78542 6130
rect 78542 6078 78594 6130
rect 78594 6078 78596 6130
rect 78540 6076 78596 6078
rect 78876 12572 78932 12628
rect 80768 17220 80824 17276
rect 80872 17274 80928 17276
rect 80976 17274 81032 17276
rect 80872 17222 80896 17274
rect 80896 17222 80928 17274
rect 80976 17222 81020 17274
rect 81020 17222 81032 17274
rect 80872 17220 80928 17222
rect 80976 17220 81032 17222
rect 81080 17220 81136 17276
rect 81184 17274 81240 17276
rect 81288 17274 81344 17276
rect 81184 17222 81196 17274
rect 81196 17222 81240 17274
rect 81288 17222 81320 17274
rect 81320 17222 81344 17274
rect 81184 17220 81240 17222
rect 81288 17220 81344 17222
rect 81392 17220 81448 17276
rect 80768 15652 80824 15708
rect 80872 15706 80928 15708
rect 80976 15706 81032 15708
rect 80872 15654 80896 15706
rect 80896 15654 80928 15706
rect 80976 15654 81020 15706
rect 81020 15654 81032 15706
rect 80872 15652 80928 15654
rect 80976 15652 81032 15654
rect 81080 15652 81136 15708
rect 81184 15706 81240 15708
rect 81288 15706 81344 15708
rect 81184 15654 81196 15706
rect 81196 15654 81240 15706
rect 81288 15654 81320 15706
rect 81320 15654 81344 15706
rect 81184 15652 81240 15654
rect 81288 15652 81344 15654
rect 81392 15652 81448 15708
rect 80220 13858 80276 13860
rect 80220 13806 80222 13858
rect 80222 13806 80274 13858
rect 80274 13806 80276 13858
rect 80220 13804 80276 13806
rect 80108 13746 80164 13748
rect 80108 13694 80110 13746
rect 80110 13694 80162 13746
rect 80162 13694 80164 13746
rect 80108 13692 80164 13694
rect 79324 13634 79380 13636
rect 79324 13582 79326 13634
rect 79326 13582 79378 13634
rect 79378 13582 79380 13634
rect 79324 13580 79380 13582
rect 78316 4450 78372 4452
rect 78316 4398 78318 4450
rect 78318 4398 78370 4450
rect 78370 4398 78372 4450
rect 78316 4396 78372 4398
rect 78876 12066 78932 12068
rect 78876 12014 78878 12066
rect 78878 12014 78930 12066
rect 78930 12014 78932 12066
rect 78876 12012 78932 12014
rect 80108 12178 80164 12180
rect 80108 12126 80110 12178
rect 80110 12126 80162 12178
rect 80162 12126 80164 12178
rect 80108 12124 80164 12126
rect 79100 8988 79156 9044
rect 80556 14530 80612 14532
rect 80556 14478 80558 14530
rect 80558 14478 80610 14530
rect 80610 14478 80612 14530
rect 80556 14476 80612 14478
rect 97692 26236 97748 26292
rect 98028 24444 98084 24500
rect 85268 24276 85324 24332
rect 85372 24330 85428 24332
rect 85476 24330 85532 24332
rect 85372 24278 85396 24330
rect 85396 24278 85428 24330
rect 85476 24278 85520 24330
rect 85520 24278 85532 24330
rect 85372 24276 85428 24278
rect 85476 24276 85532 24278
rect 85580 24276 85636 24332
rect 85684 24330 85740 24332
rect 85788 24330 85844 24332
rect 85684 24278 85696 24330
rect 85696 24278 85740 24330
rect 85788 24278 85820 24330
rect 85820 24278 85844 24330
rect 85684 24276 85740 24278
rect 85788 24276 85844 24278
rect 85892 24276 85948 24332
rect 94268 24276 94324 24332
rect 94372 24330 94428 24332
rect 94476 24330 94532 24332
rect 94372 24278 94396 24330
rect 94396 24278 94428 24330
rect 94476 24278 94520 24330
rect 94520 24278 94532 24330
rect 94372 24276 94428 24278
rect 94476 24276 94532 24278
rect 94580 24276 94636 24332
rect 94684 24330 94740 24332
rect 94788 24330 94844 24332
rect 94684 24278 94696 24330
rect 94696 24278 94740 24330
rect 94788 24278 94820 24330
rect 94820 24278 94844 24330
rect 94684 24276 94740 24278
rect 94788 24276 94844 24278
rect 94892 24276 94948 24332
rect 89768 23492 89824 23548
rect 89872 23546 89928 23548
rect 89976 23546 90032 23548
rect 89872 23494 89896 23546
rect 89896 23494 89928 23546
rect 89976 23494 90020 23546
rect 90020 23494 90032 23546
rect 89872 23492 89928 23494
rect 89976 23492 90032 23494
rect 90080 23492 90136 23548
rect 90184 23546 90240 23548
rect 90288 23546 90344 23548
rect 90184 23494 90196 23546
rect 90196 23494 90240 23546
rect 90288 23494 90320 23546
rect 90320 23494 90344 23546
rect 90184 23492 90240 23494
rect 90288 23492 90344 23494
rect 90392 23492 90448 23548
rect 96572 23378 96628 23380
rect 96572 23326 96574 23378
rect 96574 23326 96626 23378
rect 96626 23326 96628 23378
rect 96572 23324 96628 23326
rect 85036 23212 85092 23268
rect 84588 22258 84644 22260
rect 84588 22206 84590 22258
rect 84590 22206 84642 22258
rect 84642 22206 84644 22258
rect 84588 22204 84644 22206
rect 84812 22258 84868 22260
rect 84812 22206 84814 22258
rect 84814 22206 84866 22258
rect 84866 22206 84868 22258
rect 84812 22204 84868 22206
rect 82908 20130 82964 20132
rect 82908 20078 82910 20130
rect 82910 20078 82962 20130
rect 82962 20078 82964 20130
rect 82908 20076 82964 20078
rect 83020 20018 83076 20020
rect 83020 19966 83022 20018
rect 83022 19966 83074 20018
rect 83074 19966 83076 20018
rect 83020 19964 83076 19966
rect 82796 19010 82852 19012
rect 82796 18958 82798 19010
rect 82798 18958 82850 19010
rect 82850 18958 82852 19010
rect 82796 18956 82852 18958
rect 83356 20130 83412 20132
rect 83356 20078 83358 20130
rect 83358 20078 83410 20130
rect 83410 20078 83412 20130
rect 83356 20076 83412 20078
rect 83580 17612 83636 17668
rect 84364 21308 84420 21364
rect 85708 23266 85764 23268
rect 85708 23214 85710 23266
rect 85710 23214 85762 23266
rect 85762 23214 85764 23266
rect 85708 23212 85764 23214
rect 85268 22708 85324 22764
rect 85372 22762 85428 22764
rect 85476 22762 85532 22764
rect 85372 22710 85396 22762
rect 85396 22710 85428 22762
rect 85476 22710 85520 22762
rect 85520 22710 85532 22762
rect 85372 22708 85428 22710
rect 85476 22708 85532 22710
rect 85580 22708 85636 22764
rect 85684 22762 85740 22764
rect 85788 22762 85844 22764
rect 85684 22710 85696 22762
rect 85696 22710 85740 22762
rect 85788 22710 85820 22762
rect 85820 22710 85844 22762
rect 85684 22708 85740 22710
rect 85788 22708 85844 22710
rect 85892 22708 85948 22764
rect 94268 22708 94324 22764
rect 94372 22762 94428 22764
rect 94476 22762 94532 22764
rect 94372 22710 94396 22762
rect 94396 22710 94428 22762
rect 94476 22710 94520 22762
rect 94520 22710 94532 22762
rect 94372 22708 94428 22710
rect 94476 22708 94532 22710
rect 94580 22708 94636 22764
rect 94684 22762 94740 22764
rect 94788 22762 94844 22764
rect 94684 22710 94696 22762
rect 94696 22710 94740 22762
rect 94788 22710 94820 22762
rect 94820 22710 94844 22762
rect 94684 22708 94740 22710
rect 94788 22708 94844 22710
rect 94892 22708 94948 22764
rect 98028 22652 98084 22708
rect 86492 22204 86548 22260
rect 89768 21924 89824 21980
rect 89872 21978 89928 21980
rect 89976 21978 90032 21980
rect 89872 21926 89896 21978
rect 89896 21926 89928 21978
rect 89976 21926 90020 21978
rect 90020 21926 90032 21978
rect 89872 21924 89928 21926
rect 89976 21924 90032 21926
rect 90080 21924 90136 21980
rect 90184 21978 90240 21980
rect 90288 21978 90344 21980
rect 90184 21926 90196 21978
rect 90196 21926 90240 21978
rect 90288 21926 90320 21978
rect 90320 21926 90344 21978
rect 90184 21924 90240 21926
rect 90288 21924 90344 21926
rect 90392 21924 90448 21980
rect 96572 21810 96628 21812
rect 96572 21758 96574 21810
rect 96574 21758 96626 21810
rect 96626 21758 96628 21810
rect 96572 21756 96628 21758
rect 85268 21140 85324 21196
rect 85372 21194 85428 21196
rect 85476 21194 85532 21196
rect 85372 21142 85396 21194
rect 85396 21142 85428 21194
rect 85476 21142 85520 21194
rect 85520 21142 85532 21194
rect 85372 21140 85428 21142
rect 85476 21140 85532 21142
rect 85580 21140 85636 21196
rect 85684 21194 85740 21196
rect 85788 21194 85844 21196
rect 85684 21142 85696 21194
rect 85696 21142 85740 21194
rect 85788 21142 85820 21194
rect 85820 21142 85844 21194
rect 85684 21140 85740 21142
rect 85788 21140 85844 21142
rect 85892 21140 85948 21196
rect 85036 20578 85092 20580
rect 85036 20526 85038 20578
rect 85038 20526 85090 20578
rect 85090 20526 85092 20578
rect 85036 20524 85092 20526
rect 84252 20076 84308 20132
rect 84700 19906 84756 19908
rect 84700 19854 84702 19906
rect 84702 19854 84754 19906
rect 84754 19854 84756 19906
rect 84700 19852 84756 19854
rect 85036 19852 85092 19908
rect 85372 20076 85428 20132
rect 85596 20130 85652 20132
rect 85596 20078 85598 20130
rect 85598 20078 85650 20130
rect 85650 20078 85652 20130
rect 85596 20076 85652 20078
rect 86156 20524 86212 20580
rect 85268 19572 85324 19628
rect 85372 19626 85428 19628
rect 85476 19626 85532 19628
rect 85372 19574 85396 19626
rect 85396 19574 85428 19626
rect 85476 19574 85520 19626
rect 85520 19574 85532 19626
rect 85372 19572 85428 19574
rect 85476 19572 85532 19574
rect 85580 19572 85636 19628
rect 85684 19626 85740 19628
rect 85788 19626 85844 19628
rect 85684 19574 85696 19626
rect 85696 19574 85740 19626
rect 85788 19574 85820 19626
rect 85820 19574 85844 19626
rect 85684 19572 85740 19574
rect 85788 19572 85844 19574
rect 85892 19572 85948 19628
rect 85148 19010 85204 19012
rect 85148 18958 85150 19010
rect 85150 18958 85202 19010
rect 85202 18958 85204 19010
rect 85148 18956 85204 18958
rect 85268 18004 85324 18060
rect 85372 18058 85428 18060
rect 85476 18058 85532 18060
rect 85372 18006 85396 18058
rect 85396 18006 85428 18058
rect 85476 18006 85520 18058
rect 85520 18006 85532 18058
rect 85372 18004 85428 18006
rect 85476 18004 85532 18006
rect 85580 18004 85636 18060
rect 85684 18058 85740 18060
rect 85788 18058 85844 18060
rect 85684 18006 85696 18058
rect 85696 18006 85740 18058
rect 85788 18006 85820 18058
rect 85820 18006 85844 18058
rect 85684 18004 85740 18006
rect 85788 18004 85844 18006
rect 85892 18004 85948 18060
rect 85708 17666 85764 17668
rect 85708 17614 85710 17666
rect 85710 17614 85762 17666
rect 85762 17614 85764 17666
rect 85708 17612 85764 17614
rect 83692 17388 83748 17444
rect 85268 16436 85324 16492
rect 85372 16490 85428 16492
rect 85476 16490 85532 16492
rect 85372 16438 85396 16490
rect 85396 16438 85428 16490
rect 85476 16438 85520 16490
rect 85520 16438 85532 16490
rect 85372 16436 85428 16438
rect 85476 16436 85532 16438
rect 85580 16436 85636 16492
rect 85684 16490 85740 16492
rect 85788 16490 85844 16492
rect 85684 16438 85696 16490
rect 85696 16438 85740 16490
rect 85788 16438 85820 16490
rect 85820 16438 85844 16490
rect 85684 16436 85740 16438
rect 85788 16436 85844 16438
rect 85892 16436 85948 16492
rect 85268 14868 85324 14924
rect 85372 14922 85428 14924
rect 85476 14922 85532 14924
rect 85372 14870 85396 14922
rect 85396 14870 85428 14922
rect 85476 14870 85520 14922
rect 85520 14870 85532 14922
rect 85372 14868 85428 14870
rect 85476 14868 85532 14870
rect 85580 14868 85636 14924
rect 85684 14922 85740 14924
rect 85788 14922 85844 14924
rect 85684 14870 85696 14922
rect 85696 14870 85740 14922
rect 85788 14870 85820 14922
rect 85820 14870 85844 14922
rect 85684 14868 85740 14870
rect 85788 14868 85844 14870
rect 85892 14868 85948 14924
rect 83020 14476 83076 14532
rect 80768 14084 80824 14140
rect 80872 14138 80928 14140
rect 80976 14138 81032 14140
rect 80872 14086 80896 14138
rect 80896 14086 80928 14138
rect 80976 14086 81020 14138
rect 81020 14086 81032 14138
rect 80872 14084 80928 14086
rect 80976 14084 81032 14086
rect 81080 14084 81136 14140
rect 81184 14138 81240 14140
rect 81288 14138 81344 14140
rect 81184 14086 81196 14138
rect 81196 14086 81240 14138
rect 81288 14086 81320 14138
rect 81320 14086 81344 14138
rect 81184 14084 81240 14086
rect 81288 14084 81344 14086
rect 81392 14084 81448 14140
rect 80444 13692 80500 13748
rect 81788 13746 81844 13748
rect 81788 13694 81790 13746
rect 81790 13694 81842 13746
rect 81842 13694 81844 13746
rect 81788 13692 81844 13694
rect 81788 12684 81844 12740
rect 80768 12516 80824 12572
rect 80872 12570 80928 12572
rect 80976 12570 81032 12572
rect 80872 12518 80896 12570
rect 80896 12518 80928 12570
rect 80976 12518 81020 12570
rect 81020 12518 81032 12570
rect 80872 12516 80928 12518
rect 80976 12516 81032 12518
rect 81080 12516 81136 12572
rect 81184 12570 81240 12572
rect 81288 12570 81344 12572
rect 81184 12518 81196 12570
rect 81196 12518 81240 12570
rect 81288 12518 81320 12570
rect 81320 12518 81344 12570
rect 81184 12516 81240 12518
rect 81288 12516 81344 12518
rect 81392 12516 81448 12572
rect 81564 12236 81620 12292
rect 81452 11116 81508 11172
rect 80768 10948 80824 11004
rect 80872 11002 80928 11004
rect 80976 11002 81032 11004
rect 80872 10950 80896 11002
rect 80896 10950 80928 11002
rect 80976 10950 81020 11002
rect 81020 10950 81032 11002
rect 80872 10948 80928 10950
rect 80976 10948 81032 10950
rect 81080 10948 81136 11004
rect 81184 11002 81240 11004
rect 81288 11002 81344 11004
rect 81184 10950 81196 11002
rect 81196 10950 81240 11002
rect 81288 10950 81320 11002
rect 81320 10950 81344 11002
rect 81184 10948 81240 10950
rect 81288 10948 81344 10950
rect 81392 10948 81448 11004
rect 80768 9380 80824 9436
rect 80872 9434 80928 9436
rect 80976 9434 81032 9436
rect 80872 9382 80896 9434
rect 80896 9382 80928 9434
rect 80976 9382 81020 9434
rect 81020 9382 81032 9434
rect 80872 9380 80928 9382
rect 80976 9380 81032 9382
rect 81080 9380 81136 9436
rect 81184 9434 81240 9436
rect 81288 9434 81344 9436
rect 81184 9382 81196 9434
rect 81196 9382 81240 9434
rect 81288 9382 81320 9434
rect 81320 9382 81344 9434
rect 81184 9380 81240 9382
rect 81288 9380 81344 9382
rect 81392 9380 81448 9436
rect 80668 9154 80724 9156
rect 80668 9102 80670 9154
rect 80670 9102 80722 9154
rect 80722 9102 80724 9154
rect 80668 9100 80724 9102
rect 83132 14418 83188 14420
rect 83132 14366 83134 14418
rect 83134 14366 83186 14418
rect 83186 14366 83188 14418
rect 83132 14364 83188 14366
rect 82236 14306 82292 14308
rect 82236 14254 82238 14306
rect 82238 14254 82290 14306
rect 82290 14254 82292 14306
rect 82236 14252 82292 14254
rect 81900 12012 81956 12068
rect 81900 8988 81956 9044
rect 82124 11116 82180 11172
rect 78876 4396 78932 4452
rect 77868 4284 77924 4340
rect 79436 4284 79492 4340
rect 80108 5906 80164 5908
rect 80108 5854 80110 5906
rect 80110 5854 80162 5906
rect 80162 5854 80164 5906
rect 80108 5852 80164 5854
rect 80768 7812 80824 7868
rect 80872 7866 80928 7868
rect 80976 7866 81032 7868
rect 80872 7814 80896 7866
rect 80896 7814 80928 7866
rect 80976 7814 81020 7866
rect 81020 7814 81032 7866
rect 80872 7812 80928 7814
rect 80976 7812 81032 7814
rect 81080 7812 81136 7868
rect 81184 7866 81240 7868
rect 81288 7866 81344 7868
rect 81184 7814 81196 7866
rect 81196 7814 81240 7866
rect 81288 7814 81320 7866
rect 81320 7814 81344 7866
rect 81184 7812 81240 7814
rect 81288 7812 81344 7814
rect 81392 7812 81448 7868
rect 80768 6244 80824 6300
rect 80872 6298 80928 6300
rect 80976 6298 81032 6300
rect 80872 6246 80896 6298
rect 80896 6246 80928 6298
rect 80976 6246 81020 6298
rect 81020 6246 81032 6298
rect 80872 6244 80928 6246
rect 80976 6244 81032 6246
rect 81080 6244 81136 6300
rect 81184 6298 81240 6300
rect 81288 6298 81344 6300
rect 81184 6246 81196 6298
rect 81196 6246 81240 6298
rect 81288 6246 81320 6298
rect 81320 6246 81344 6298
rect 81184 6244 81240 6246
rect 81288 6244 81344 6246
rect 81392 6244 81448 6300
rect 80444 5404 80500 5460
rect 81676 6748 81732 6804
rect 81788 6578 81844 6580
rect 81788 6526 81790 6578
rect 81790 6526 81842 6578
rect 81842 6526 81844 6578
rect 81788 6524 81844 6526
rect 81564 5292 81620 5348
rect 81676 6412 81732 6468
rect 80668 5180 80724 5236
rect 79996 4508 80052 4564
rect 81676 5068 81732 5124
rect 80768 4676 80824 4732
rect 80872 4730 80928 4732
rect 80976 4730 81032 4732
rect 80872 4678 80896 4730
rect 80896 4678 80928 4730
rect 80976 4678 81020 4730
rect 81020 4678 81032 4730
rect 80872 4676 80928 4678
rect 80976 4676 81032 4678
rect 81080 4676 81136 4732
rect 81184 4730 81240 4732
rect 81288 4730 81344 4732
rect 81184 4678 81196 4730
rect 81196 4678 81240 4730
rect 81288 4678 81320 4730
rect 81320 4678 81344 4730
rect 81184 4676 81240 4678
rect 81288 4676 81344 4678
rect 81392 4676 81448 4732
rect 79212 4172 79268 4228
rect 78876 4060 78932 4116
rect 78092 3612 78148 3668
rect 81900 5068 81956 5124
rect 82572 12178 82628 12180
rect 82572 12126 82574 12178
rect 82574 12126 82626 12178
rect 82626 12126 82628 12178
rect 82572 12124 82628 12126
rect 82236 10332 82292 10388
rect 82124 6636 82180 6692
rect 82796 13580 82852 13636
rect 83580 13580 83636 13636
rect 85268 13300 85324 13356
rect 85372 13354 85428 13356
rect 85476 13354 85532 13356
rect 85372 13302 85396 13354
rect 85396 13302 85428 13354
rect 85476 13302 85520 13354
rect 85520 13302 85532 13354
rect 85372 13300 85428 13302
rect 85476 13300 85532 13302
rect 85580 13300 85636 13356
rect 85684 13354 85740 13356
rect 85788 13354 85844 13356
rect 85684 13302 85696 13354
rect 85696 13302 85740 13354
rect 85788 13302 85820 13354
rect 85820 13302 85844 13354
rect 85684 13300 85740 13302
rect 85788 13300 85844 13302
rect 85892 13300 85948 13356
rect 83804 12066 83860 12068
rect 83804 12014 83806 12066
rect 83806 12014 83858 12066
rect 83858 12014 83860 12066
rect 83804 12012 83860 12014
rect 86044 12012 86100 12068
rect 85268 11732 85324 11788
rect 85372 11786 85428 11788
rect 85476 11786 85532 11788
rect 85372 11734 85396 11786
rect 85396 11734 85428 11786
rect 85476 11734 85520 11786
rect 85520 11734 85532 11786
rect 85372 11732 85428 11734
rect 85476 11732 85532 11734
rect 85580 11732 85636 11788
rect 85684 11786 85740 11788
rect 85788 11786 85844 11788
rect 85684 11734 85696 11786
rect 85696 11734 85740 11786
rect 85788 11734 85820 11786
rect 85820 11734 85844 11786
rect 85684 11732 85740 11734
rect 85788 11732 85844 11734
rect 85892 11732 85948 11788
rect 85268 10164 85324 10220
rect 85372 10218 85428 10220
rect 85476 10218 85532 10220
rect 85372 10166 85396 10218
rect 85396 10166 85428 10218
rect 85476 10166 85520 10218
rect 85520 10166 85532 10218
rect 85372 10164 85428 10166
rect 85476 10164 85532 10166
rect 85580 10164 85636 10220
rect 85684 10218 85740 10220
rect 85788 10218 85844 10220
rect 85684 10166 85696 10218
rect 85696 10166 85740 10218
rect 85788 10166 85820 10218
rect 85820 10166 85844 10218
rect 85684 10164 85740 10166
rect 85788 10164 85844 10166
rect 85892 10164 85948 10220
rect 82684 6636 82740 6692
rect 82796 9660 82852 9716
rect 82348 6466 82404 6468
rect 82348 6414 82350 6466
rect 82350 6414 82402 6466
rect 82402 6414 82404 6466
rect 82348 6412 82404 6414
rect 82124 5180 82180 5236
rect 82460 5068 82516 5124
rect 84028 9042 84084 9044
rect 84028 8990 84030 9042
rect 84030 8990 84082 9042
rect 84082 8990 84084 9042
rect 84028 8988 84084 8990
rect 83916 7420 83972 7476
rect 84028 6690 84084 6692
rect 84028 6638 84030 6690
rect 84030 6638 84082 6690
rect 84082 6638 84084 6690
rect 84028 6636 84084 6638
rect 85148 9996 85204 10052
rect 84364 9714 84420 9716
rect 84364 9662 84366 9714
rect 84366 9662 84418 9714
rect 84418 9662 84420 9714
rect 84364 9660 84420 9662
rect 85268 8596 85324 8652
rect 85372 8650 85428 8652
rect 85476 8650 85532 8652
rect 85372 8598 85396 8650
rect 85396 8598 85428 8650
rect 85476 8598 85520 8650
rect 85520 8598 85532 8650
rect 85372 8596 85428 8598
rect 85476 8596 85532 8598
rect 85580 8596 85636 8652
rect 85684 8650 85740 8652
rect 85788 8650 85844 8652
rect 85684 8598 85696 8650
rect 85696 8598 85740 8650
rect 85788 8598 85820 8650
rect 85820 8598 85844 8650
rect 85684 8596 85740 8598
rect 85788 8596 85844 8598
rect 85892 8596 85948 8652
rect 85268 7028 85324 7084
rect 85372 7082 85428 7084
rect 85476 7082 85532 7084
rect 85372 7030 85396 7082
rect 85396 7030 85428 7082
rect 85476 7030 85520 7082
rect 85520 7030 85532 7082
rect 85372 7028 85428 7030
rect 85476 7028 85532 7030
rect 85580 7028 85636 7084
rect 85684 7082 85740 7084
rect 85788 7082 85844 7084
rect 85684 7030 85696 7082
rect 85696 7030 85740 7082
rect 85788 7030 85820 7082
rect 85820 7030 85844 7082
rect 85684 7028 85740 7030
rect 85788 7028 85844 7030
rect 85892 7028 85948 7084
rect 85268 5460 85324 5516
rect 85372 5514 85428 5516
rect 85476 5514 85532 5516
rect 85372 5462 85396 5514
rect 85396 5462 85428 5514
rect 85476 5462 85520 5514
rect 85520 5462 85532 5514
rect 85372 5460 85428 5462
rect 85476 5460 85532 5462
rect 85580 5460 85636 5516
rect 85684 5514 85740 5516
rect 85788 5514 85844 5516
rect 85684 5462 85696 5514
rect 85696 5462 85740 5514
rect 85788 5462 85820 5514
rect 85820 5462 85844 5514
rect 85684 5460 85740 5462
rect 85788 5460 85844 5462
rect 85892 5460 85948 5516
rect 84700 5180 84756 5236
rect 83244 3612 83300 3668
rect 85932 4226 85988 4228
rect 85932 4174 85934 4226
rect 85934 4174 85986 4226
rect 85986 4174 85988 4226
rect 85932 4172 85988 4174
rect 85268 3892 85324 3948
rect 85372 3946 85428 3948
rect 85476 3946 85532 3948
rect 85372 3894 85396 3946
rect 85396 3894 85428 3946
rect 85476 3894 85520 3946
rect 85520 3894 85532 3946
rect 85372 3892 85428 3894
rect 85476 3892 85532 3894
rect 85580 3892 85636 3948
rect 85684 3946 85740 3948
rect 85788 3946 85844 3948
rect 85684 3894 85696 3946
rect 85696 3894 85740 3946
rect 85788 3894 85820 3946
rect 85820 3894 85844 3946
rect 85684 3892 85740 3894
rect 85788 3892 85844 3894
rect 85892 3892 85948 3948
rect 86156 6524 86212 6580
rect 94268 21140 94324 21196
rect 94372 21194 94428 21196
rect 94476 21194 94532 21196
rect 94372 21142 94396 21194
rect 94396 21142 94428 21194
rect 94476 21142 94520 21194
rect 94520 21142 94532 21194
rect 94372 21140 94428 21142
rect 94476 21140 94532 21142
rect 94580 21140 94636 21196
rect 94684 21194 94740 21196
rect 94788 21194 94844 21196
rect 94684 21142 94696 21194
rect 94696 21142 94740 21194
rect 94788 21142 94820 21194
rect 94820 21142 94844 21194
rect 94684 21140 94740 21142
rect 94788 21140 94844 21142
rect 94892 21140 94948 21196
rect 98028 20860 98084 20916
rect 89768 20356 89824 20412
rect 89872 20410 89928 20412
rect 89976 20410 90032 20412
rect 89872 20358 89896 20410
rect 89896 20358 89928 20410
rect 89976 20358 90020 20410
rect 90020 20358 90032 20410
rect 89872 20356 89928 20358
rect 89976 20356 90032 20358
rect 90080 20356 90136 20412
rect 90184 20410 90240 20412
rect 90288 20410 90344 20412
rect 90184 20358 90196 20410
rect 90196 20358 90240 20410
rect 90288 20358 90320 20410
rect 90320 20358 90344 20410
rect 90184 20356 90240 20358
rect 90288 20356 90344 20358
rect 90392 20356 90448 20412
rect 89068 20076 89124 20132
rect 94268 19572 94324 19628
rect 94372 19626 94428 19628
rect 94476 19626 94532 19628
rect 94372 19574 94396 19626
rect 94396 19574 94428 19626
rect 94476 19574 94520 19626
rect 94520 19574 94532 19626
rect 94372 19572 94428 19574
rect 94476 19572 94532 19574
rect 94580 19572 94636 19628
rect 94684 19626 94740 19628
rect 94788 19626 94844 19628
rect 94684 19574 94696 19626
rect 94696 19574 94740 19626
rect 94788 19574 94820 19626
rect 94820 19574 94844 19626
rect 94684 19572 94740 19574
rect 94788 19572 94844 19574
rect 94892 19572 94948 19628
rect 88284 19010 88340 19012
rect 88284 18958 88286 19010
rect 88286 18958 88338 19010
rect 88338 18958 88340 19010
rect 88284 18956 88340 18958
rect 96684 19122 96740 19124
rect 96684 19070 96686 19122
rect 96686 19070 96738 19122
rect 96738 19070 96740 19122
rect 96684 19068 96740 19070
rect 98028 19122 98084 19124
rect 98028 19070 98030 19122
rect 98030 19070 98082 19122
rect 98082 19070 98084 19122
rect 98028 19068 98084 19070
rect 89768 18788 89824 18844
rect 89872 18842 89928 18844
rect 89976 18842 90032 18844
rect 89872 18790 89896 18842
rect 89896 18790 89928 18842
rect 89976 18790 90020 18842
rect 90020 18790 90032 18842
rect 89872 18788 89928 18790
rect 89976 18788 90032 18790
rect 90080 18788 90136 18844
rect 90184 18842 90240 18844
rect 90288 18842 90344 18844
rect 90184 18790 90196 18842
rect 90196 18790 90240 18842
rect 90288 18790 90320 18842
rect 90320 18790 90344 18842
rect 90184 18788 90240 18790
rect 90288 18788 90344 18790
rect 90392 18788 90448 18844
rect 89068 18508 89124 18564
rect 89964 18562 90020 18564
rect 89964 18510 89966 18562
rect 89966 18510 90018 18562
rect 90018 18510 90020 18562
rect 89964 18508 90020 18510
rect 94268 18004 94324 18060
rect 94372 18058 94428 18060
rect 94476 18058 94532 18060
rect 94372 18006 94396 18058
rect 94396 18006 94428 18058
rect 94476 18006 94520 18058
rect 94520 18006 94532 18058
rect 94372 18004 94428 18006
rect 94476 18004 94532 18006
rect 94580 18004 94636 18060
rect 94684 18058 94740 18060
rect 94788 18058 94844 18060
rect 94684 18006 94696 18058
rect 94696 18006 94740 18058
rect 94788 18006 94820 18058
rect 94820 18006 94844 18058
rect 94684 18004 94740 18006
rect 94788 18004 94844 18006
rect 94892 18004 94948 18060
rect 89768 17220 89824 17276
rect 89872 17274 89928 17276
rect 89976 17274 90032 17276
rect 89872 17222 89896 17274
rect 89896 17222 89928 17274
rect 89976 17222 90020 17274
rect 90020 17222 90032 17274
rect 89872 17220 89928 17222
rect 89976 17220 90032 17222
rect 90080 17220 90136 17276
rect 90184 17274 90240 17276
rect 90288 17274 90344 17276
rect 90184 17222 90196 17274
rect 90196 17222 90240 17274
rect 90288 17222 90320 17274
rect 90320 17222 90344 17274
rect 90184 17220 90240 17222
rect 90288 17220 90344 17222
rect 90392 17220 90448 17276
rect 89768 15652 89824 15708
rect 89872 15706 89928 15708
rect 89976 15706 90032 15708
rect 89872 15654 89896 15706
rect 89896 15654 89928 15706
rect 89976 15654 90020 15706
rect 90020 15654 90032 15706
rect 89872 15652 89928 15654
rect 89976 15652 90032 15654
rect 90080 15652 90136 15708
rect 90184 15706 90240 15708
rect 90288 15706 90344 15708
rect 90184 15654 90196 15706
rect 90196 15654 90240 15706
rect 90288 15654 90320 15706
rect 90320 15654 90344 15706
rect 90184 15652 90240 15654
rect 90288 15652 90344 15654
rect 90392 15652 90448 15708
rect 88172 14252 88228 14308
rect 87388 9212 87444 9268
rect 88060 9996 88116 10052
rect 87500 8988 87556 9044
rect 87948 6802 88004 6804
rect 87948 6750 87950 6802
rect 87950 6750 88002 6802
rect 88002 6750 88004 6802
rect 87948 6748 88004 6750
rect 86268 4508 86324 4564
rect 89768 14084 89824 14140
rect 89872 14138 89928 14140
rect 89976 14138 90032 14140
rect 89872 14086 89896 14138
rect 89896 14086 89928 14138
rect 89976 14086 90020 14138
rect 90020 14086 90032 14138
rect 89872 14084 89928 14086
rect 89976 14084 90032 14086
rect 90080 14084 90136 14140
rect 90184 14138 90240 14140
rect 90288 14138 90344 14140
rect 90184 14086 90196 14138
rect 90196 14086 90240 14138
rect 90288 14086 90320 14138
rect 90320 14086 90344 14138
rect 90184 14084 90240 14086
rect 90288 14084 90344 14086
rect 90392 14084 90448 14140
rect 89768 12516 89824 12572
rect 89872 12570 89928 12572
rect 89976 12570 90032 12572
rect 89872 12518 89896 12570
rect 89896 12518 89928 12570
rect 89976 12518 90020 12570
rect 90020 12518 90032 12570
rect 89872 12516 89928 12518
rect 89976 12516 90032 12518
rect 90080 12516 90136 12572
rect 90184 12570 90240 12572
rect 90288 12570 90344 12572
rect 90184 12518 90196 12570
rect 90196 12518 90240 12570
rect 90288 12518 90320 12570
rect 90320 12518 90344 12570
rect 90184 12516 90240 12518
rect 90288 12516 90344 12518
rect 90392 12516 90448 12572
rect 89768 10948 89824 11004
rect 89872 11002 89928 11004
rect 89976 11002 90032 11004
rect 89872 10950 89896 11002
rect 89896 10950 89928 11002
rect 89976 10950 90020 11002
rect 90020 10950 90032 11002
rect 89872 10948 89928 10950
rect 89976 10948 90032 10950
rect 90080 10948 90136 11004
rect 90184 11002 90240 11004
rect 90288 11002 90344 11004
rect 90184 10950 90196 11002
rect 90196 10950 90240 11002
rect 90288 10950 90320 11002
rect 90320 10950 90344 11002
rect 90184 10948 90240 10950
rect 90288 10948 90344 10950
rect 90392 10948 90448 11004
rect 88956 10332 89012 10388
rect 89768 9380 89824 9436
rect 89872 9434 89928 9436
rect 89976 9434 90032 9436
rect 89872 9382 89896 9434
rect 89896 9382 89928 9434
rect 89976 9382 90020 9434
rect 90020 9382 90032 9434
rect 89872 9380 89928 9382
rect 89976 9380 90032 9382
rect 90080 9380 90136 9436
rect 90184 9434 90240 9436
rect 90288 9434 90344 9436
rect 90184 9382 90196 9434
rect 90196 9382 90240 9434
rect 90288 9382 90320 9434
rect 90320 9382 90344 9434
rect 90184 9380 90240 9382
rect 90288 9380 90344 9382
rect 90392 9380 90448 9436
rect 88956 8316 89012 8372
rect 89768 7812 89824 7868
rect 89872 7866 89928 7868
rect 89976 7866 90032 7868
rect 89872 7814 89896 7866
rect 89896 7814 89928 7866
rect 89976 7814 90020 7866
rect 90020 7814 90032 7866
rect 89872 7812 89928 7814
rect 89976 7812 90032 7814
rect 90080 7812 90136 7868
rect 90184 7866 90240 7868
rect 90288 7866 90344 7868
rect 90184 7814 90196 7866
rect 90196 7814 90240 7866
rect 90288 7814 90320 7866
rect 90320 7814 90344 7866
rect 90184 7812 90240 7814
rect 90288 7812 90344 7814
rect 90392 7812 90448 7868
rect 96684 17442 96740 17444
rect 96684 17390 96686 17442
rect 96686 17390 96738 17442
rect 96738 17390 96740 17442
rect 96684 17388 96740 17390
rect 98028 17276 98084 17332
rect 94268 16436 94324 16492
rect 94372 16490 94428 16492
rect 94476 16490 94532 16492
rect 94372 16438 94396 16490
rect 94396 16438 94428 16490
rect 94476 16438 94520 16490
rect 94520 16438 94532 16490
rect 94372 16436 94428 16438
rect 94476 16436 94532 16438
rect 94580 16436 94636 16492
rect 94684 16490 94740 16492
rect 94788 16490 94844 16492
rect 94684 16438 94696 16490
rect 94696 16438 94740 16490
rect 94788 16438 94820 16490
rect 94820 16438 94844 16490
rect 94684 16436 94740 16438
rect 94788 16436 94844 16438
rect 94892 16436 94948 16492
rect 96684 16098 96740 16100
rect 96684 16046 96686 16098
rect 96686 16046 96738 16098
rect 96738 16046 96740 16098
rect 96684 16044 96740 16046
rect 98028 15484 98084 15540
rect 94268 14868 94324 14924
rect 94372 14922 94428 14924
rect 94476 14922 94532 14924
rect 94372 14870 94396 14922
rect 94396 14870 94428 14922
rect 94476 14870 94520 14922
rect 94520 14870 94532 14922
rect 94372 14868 94428 14870
rect 94476 14868 94532 14870
rect 94580 14868 94636 14924
rect 94684 14922 94740 14924
rect 94788 14922 94844 14924
rect 94684 14870 94696 14922
rect 94696 14870 94740 14922
rect 94788 14870 94820 14922
rect 94820 14870 94844 14922
rect 94684 14868 94740 14870
rect 94788 14868 94844 14870
rect 94892 14868 94948 14924
rect 90860 14476 90916 14532
rect 90524 6636 90580 6692
rect 90748 8316 90804 8372
rect 89768 6244 89824 6300
rect 89872 6298 89928 6300
rect 89976 6298 90032 6300
rect 89872 6246 89896 6298
rect 89896 6246 89928 6298
rect 89976 6246 90020 6298
rect 90020 6246 90032 6298
rect 89872 6244 89928 6246
rect 89976 6244 90032 6246
rect 90080 6244 90136 6300
rect 90184 6298 90240 6300
rect 90288 6298 90344 6300
rect 90184 6246 90196 6298
rect 90196 6246 90240 6298
rect 90288 6246 90320 6298
rect 90320 6246 90344 6298
rect 90184 6244 90240 6246
rect 90288 6244 90344 6246
rect 90392 6244 90448 6300
rect 96908 14530 96964 14532
rect 96908 14478 96910 14530
rect 96910 14478 96962 14530
rect 96962 14478 96964 14530
rect 96908 14476 96964 14478
rect 98028 13692 98084 13748
rect 94268 13300 94324 13356
rect 94372 13354 94428 13356
rect 94476 13354 94532 13356
rect 94372 13302 94396 13354
rect 94396 13302 94428 13354
rect 94476 13302 94520 13354
rect 94520 13302 94532 13354
rect 94372 13300 94428 13302
rect 94476 13300 94532 13302
rect 94580 13300 94636 13356
rect 94684 13354 94740 13356
rect 94788 13354 94844 13356
rect 94684 13302 94696 13354
rect 94696 13302 94740 13354
rect 94788 13302 94820 13354
rect 94820 13302 94844 13354
rect 94684 13300 94740 13302
rect 94788 13300 94844 13302
rect 94892 13300 94948 13356
rect 96572 12290 96628 12292
rect 96572 12238 96574 12290
rect 96574 12238 96626 12290
rect 96626 12238 96628 12290
rect 96572 12236 96628 12238
rect 91196 12124 91252 12180
rect 89768 4676 89824 4732
rect 89872 4730 89928 4732
rect 89976 4730 90032 4732
rect 89872 4678 89896 4730
rect 89896 4678 89928 4730
rect 89976 4678 90020 4730
rect 90020 4678 90032 4730
rect 89872 4676 89928 4678
rect 89976 4676 90032 4678
rect 90080 4676 90136 4732
rect 90184 4730 90240 4732
rect 90288 4730 90344 4732
rect 90184 4678 90196 4730
rect 90196 4678 90240 4730
rect 90288 4678 90320 4730
rect 90320 4678 90344 4730
rect 90184 4676 90240 4678
rect 90288 4676 90344 4678
rect 90392 4676 90448 4732
rect 98028 11900 98084 11956
rect 94268 11732 94324 11788
rect 94372 11786 94428 11788
rect 94476 11786 94532 11788
rect 94372 11734 94396 11786
rect 94396 11734 94428 11786
rect 94476 11734 94520 11786
rect 94520 11734 94532 11786
rect 94372 11732 94428 11734
rect 94476 11732 94532 11734
rect 94580 11732 94636 11788
rect 94684 11786 94740 11788
rect 94788 11786 94844 11788
rect 94684 11734 94696 11786
rect 94696 11734 94740 11786
rect 94788 11734 94820 11786
rect 94820 11734 94844 11786
rect 94684 11732 94740 11734
rect 94788 11732 94844 11734
rect 94892 11732 94948 11788
rect 96684 10722 96740 10724
rect 96684 10670 96686 10722
rect 96686 10670 96738 10722
rect 96738 10670 96740 10722
rect 96684 10668 96740 10670
rect 94268 10164 94324 10220
rect 94372 10218 94428 10220
rect 94476 10218 94532 10220
rect 94372 10166 94396 10218
rect 94396 10166 94428 10218
rect 94476 10166 94520 10218
rect 94520 10166 94532 10218
rect 94372 10164 94428 10166
rect 94476 10164 94532 10166
rect 94580 10164 94636 10220
rect 94684 10218 94740 10220
rect 94788 10218 94844 10220
rect 94684 10166 94696 10218
rect 94696 10166 94740 10218
rect 94788 10166 94820 10218
rect 94820 10166 94844 10218
rect 94684 10164 94740 10166
rect 94788 10164 94844 10166
rect 94892 10164 94948 10220
rect 98028 10108 98084 10164
rect 96684 9266 96740 9268
rect 96684 9214 96686 9266
rect 96686 9214 96738 9266
rect 96738 9214 96740 9266
rect 96684 9212 96740 9214
rect 94268 8596 94324 8652
rect 94372 8650 94428 8652
rect 94476 8650 94532 8652
rect 94372 8598 94396 8650
rect 94396 8598 94428 8650
rect 94476 8598 94520 8650
rect 94520 8598 94532 8650
rect 94372 8596 94428 8598
rect 94476 8596 94532 8598
rect 94580 8596 94636 8652
rect 94684 8650 94740 8652
rect 94788 8650 94844 8652
rect 94684 8598 94696 8650
rect 94696 8598 94740 8650
rect 94788 8598 94820 8650
rect 94820 8598 94844 8650
rect 94684 8596 94740 8598
rect 94788 8596 94844 8598
rect 94892 8596 94948 8652
rect 97692 8316 97748 8372
rect 94268 7028 94324 7084
rect 94372 7082 94428 7084
rect 94476 7082 94532 7084
rect 94372 7030 94396 7082
rect 94396 7030 94428 7082
rect 94476 7030 94520 7082
rect 94520 7030 94532 7082
rect 94372 7028 94428 7030
rect 94476 7028 94532 7030
rect 94580 7028 94636 7084
rect 94684 7082 94740 7084
rect 94788 7082 94844 7084
rect 94684 7030 94696 7082
rect 94696 7030 94740 7082
rect 94788 7030 94820 7082
rect 94820 7030 94844 7082
rect 94684 7028 94740 7030
rect 94788 7028 94844 7030
rect 94892 7028 94948 7084
rect 96684 6690 96740 6692
rect 96684 6638 96686 6690
rect 96686 6638 96738 6690
rect 96738 6638 96740 6690
rect 96684 6636 96740 6638
rect 98028 6578 98084 6580
rect 98028 6526 98030 6578
rect 98030 6526 98082 6578
rect 98082 6526 98084 6578
rect 98028 6524 98084 6526
rect 94268 5460 94324 5516
rect 94372 5514 94428 5516
rect 94476 5514 94532 5516
rect 94372 5462 94396 5514
rect 94396 5462 94428 5514
rect 94476 5462 94520 5514
rect 94520 5462 94532 5514
rect 94372 5460 94428 5462
rect 94476 5460 94532 5462
rect 94580 5460 94636 5516
rect 94684 5514 94740 5516
rect 94788 5514 94844 5516
rect 94684 5462 94696 5514
rect 94696 5462 94740 5514
rect 94788 5462 94820 5514
rect 94820 5462 94844 5514
rect 94684 5460 94740 5462
rect 94788 5460 94844 5462
rect 94892 5460 94948 5516
rect 96572 5292 96628 5348
rect 97692 4732 97748 4788
rect 96684 4562 96740 4564
rect 96684 4510 96686 4562
rect 96686 4510 96738 4562
rect 96738 4510 96740 4562
rect 96684 4508 96740 4510
rect 86156 4172 86212 4228
rect 82908 3500 82964 3556
rect 76188 3276 76244 3332
rect 81900 3330 81956 3332
rect 81900 3278 81902 3330
rect 81902 3278 81954 3330
rect 81954 3278 81956 3330
rect 81900 3276 81956 3278
rect 71768 3108 71824 3164
rect 71872 3162 71928 3164
rect 71976 3162 72032 3164
rect 71872 3110 71896 3162
rect 71896 3110 71928 3162
rect 71976 3110 72020 3162
rect 72020 3110 72032 3162
rect 71872 3108 71928 3110
rect 71976 3108 72032 3110
rect 72080 3108 72136 3164
rect 72184 3162 72240 3164
rect 72288 3162 72344 3164
rect 72184 3110 72196 3162
rect 72196 3110 72240 3162
rect 72288 3110 72320 3162
rect 72320 3110 72344 3162
rect 72184 3108 72240 3110
rect 72288 3108 72344 3110
rect 72392 3108 72448 3164
rect 80768 3108 80824 3164
rect 80872 3162 80928 3164
rect 80976 3162 81032 3164
rect 80872 3110 80896 3162
rect 80896 3110 80928 3162
rect 80976 3110 81020 3162
rect 81020 3110 81032 3162
rect 80872 3108 80928 3110
rect 80976 3108 81032 3110
rect 81080 3108 81136 3164
rect 81184 3162 81240 3164
rect 81288 3162 81344 3164
rect 81184 3110 81196 3162
rect 81196 3110 81240 3162
rect 81288 3110 81320 3162
rect 81320 3110 81344 3162
rect 81184 3108 81240 3110
rect 81288 3108 81344 3110
rect 81392 3108 81448 3164
rect 94268 3892 94324 3948
rect 94372 3946 94428 3948
rect 94476 3946 94532 3948
rect 94372 3894 94396 3946
rect 94396 3894 94428 3946
rect 94476 3894 94520 3946
rect 94520 3894 94532 3946
rect 94372 3892 94428 3894
rect 94476 3892 94532 3894
rect 94580 3892 94636 3948
rect 94684 3946 94740 3948
rect 94788 3946 94844 3948
rect 94684 3894 94696 3946
rect 94696 3894 94740 3946
rect 94788 3894 94820 3946
rect 94820 3894 94844 3946
rect 94684 3892 94740 3894
rect 94788 3892 94844 3894
rect 94892 3892 94948 3948
rect 96348 3724 96404 3780
rect 86156 3554 86212 3556
rect 86156 3502 86158 3554
rect 86158 3502 86210 3554
rect 86210 3502 86212 3554
rect 86156 3500 86212 3502
rect 83244 3442 83300 3444
rect 83244 3390 83246 3442
rect 83246 3390 83298 3442
rect 83298 3390 83300 3442
rect 83244 3388 83300 3390
rect 96908 3724 96964 3780
rect 89768 3108 89824 3164
rect 89872 3162 89928 3164
rect 89976 3162 90032 3164
rect 89872 3110 89896 3162
rect 89896 3110 89928 3162
rect 89976 3110 90020 3162
rect 90020 3110 90032 3162
rect 89872 3108 89928 3110
rect 89976 3108 90032 3110
rect 90080 3108 90136 3164
rect 90184 3162 90240 3164
rect 90288 3162 90344 3164
rect 90184 3110 90196 3162
rect 90196 3110 90240 3162
rect 90288 3110 90320 3162
rect 90320 3110 90344 3162
rect 90184 3108 90240 3110
rect 90288 3108 90344 3110
rect 90392 3108 90448 3164
rect 94108 3442 94164 3444
rect 94108 3390 94110 3442
rect 94110 3390 94162 3442
rect 94162 3390 94164 3442
rect 94108 3388 94164 3390
rect 97692 2940 97748 2996
rect 97804 1148 97860 1204
<< metal3 >>
rect 99200 58548 100000 58576
rect 97682 58492 97692 58548
rect 97748 58492 100000 58548
rect 99200 58464 100000 58492
rect 99200 56756 100000 56784
rect 95890 56700 95900 56756
rect 95956 56700 100000 56756
rect 99200 56672 100000 56700
rect 8758 56420 8768 56476
rect 8824 56420 8872 56476
rect 8928 56420 8976 56476
rect 9032 56420 9080 56476
rect 9136 56420 9184 56476
rect 9240 56420 9288 56476
rect 9344 56420 9392 56476
rect 9448 56420 9458 56476
rect 17758 56420 17768 56476
rect 17824 56420 17872 56476
rect 17928 56420 17976 56476
rect 18032 56420 18080 56476
rect 18136 56420 18184 56476
rect 18240 56420 18288 56476
rect 18344 56420 18392 56476
rect 18448 56420 18458 56476
rect 26758 56420 26768 56476
rect 26824 56420 26872 56476
rect 26928 56420 26976 56476
rect 27032 56420 27080 56476
rect 27136 56420 27184 56476
rect 27240 56420 27288 56476
rect 27344 56420 27392 56476
rect 27448 56420 27458 56476
rect 35758 56420 35768 56476
rect 35824 56420 35872 56476
rect 35928 56420 35976 56476
rect 36032 56420 36080 56476
rect 36136 56420 36184 56476
rect 36240 56420 36288 56476
rect 36344 56420 36392 56476
rect 36448 56420 36458 56476
rect 44758 56420 44768 56476
rect 44824 56420 44872 56476
rect 44928 56420 44976 56476
rect 45032 56420 45080 56476
rect 45136 56420 45184 56476
rect 45240 56420 45288 56476
rect 45344 56420 45392 56476
rect 45448 56420 45458 56476
rect 53758 56420 53768 56476
rect 53824 56420 53872 56476
rect 53928 56420 53976 56476
rect 54032 56420 54080 56476
rect 54136 56420 54184 56476
rect 54240 56420 54288 56476
rect 54344 56420 54392 56476
rect 54448 56420 54458 56476
rect 62758 56420 62768 56476
rect 62824 56420 62872 56476
rect 62928 56420 62976 56476
rect 63032 56420 63080 56476
rect 63136 56420 63184 56476
rect 63240 56420 63288 56476
rect 63344 56420 63392 56476
rect 63448 56420 63458 56476
rect 71758 56420 71768 56476
rect 71824 56420 71872 56476
rect 71928 56420 71976 56476
rect 72032 56420 72080 56476
rect 72136 56420 72184 56476
rect 72240 56420 72288 56476
rect 72344 56420 72392 56476
rect 72448 56420 72458 56476
rect 80758 56420 80768 56476
rect 80824 56420 80872 56476
rect 80928 56420 80976 56476
rect 81032 56420 81080 56476
rect 81136 56420 81184 56476
rect 81240 56420 81288 56476
rect 81344 56420 81392 56476
rect 81448 56420 81458 56476
rect 89758 56420 89768 56476
rect 89824 56420 89872 56476
rect 89928 56420 89976 56476
rect 90032 56420 90080 56476
rect 90136 56420 90184 56476
rect 90240 56420 90288 56476
rect 90344 56420 90392 56476
rect 90448 56420 90458 56476
rect 31378 56252 31388 56308
rect 31444 56252 32172 56308
rect 32228 56252 32238 56308
rect 68338 56252 68348 56308
rect 68404 56252 69020 56308
rect 69076 56252 69086 56308
rect 2034 56140 2044 56196
rect 2100 56140 12124 56196
rect 12180 56140 12190 56196
rect 20066 56028 20076 56084
rect 20132 56028 25452 56084
rect 25508 56028 25518 56084
rect 67106 56028 67116 56084
rect 67172 56028 68460 56084
rect 68516 56028 68526 56084
rect 82114 56028 82124 56084
rect 82180 56028 93212 56084
rect 93268 56028 93278 56084
rect 96338 56028 96348 56084
rect 96404 56028 97244 56084
rect 97300 56028 98140 56084
rect 98196 56028 98206 56084
rect 8194 55916 8204 55972
rect 8260 55916 8764 55972
rect 8820 55916 26124 55972
rect 26180 55916 26190 55972
rect 0 55636 800 55664
rect 4258 55636 4268 55692
rect 4324 55636 4372 55692
rect 4428 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4788 55692
rect 4844 55636 4892 55692
rect 4948 55636 4958 55692
rect 13258 55636 13268 55692
rect 13324 55636 13372 55692
rect 13428 55636 13476 55692
rect 13532 55636 13580 55692
rect 13636 55636 13684 55692
rect 13740 55636 13788 55692
rect 13844 55636 13892 55692
rect 13948 55636 13958 55692
rect 22258 55636 22268 55692
rect 22324 55636 22372 55692
rect 22428 55636 22476 55692
rect 22532 55636 22580 55692
rect 22636 55636 22684 55692
rect 22740 55636 22788 55692
rect 22844 55636 22892 55692
rect 22948 55636 22958 55692
rect 31258 55636 31268 55692
rect 31324 55636 31372 55692
rect 31428 55636 31476 55692
rect 31532 55636 31580 55692
rect 31636 55636 31684 55692
rect 31740 55636 31788 55692
rect 31844 55636 31892 55692
rect 31948 55636 31958 55692
rect 40258 55636 40268 55692
rect 40324 55636 40372 55692
rect 40428 55636 40476 55692
rect 40532 55636 40580 55692
rect 40636 55636 40684 55692
rect 40740 55636 40788 55692
rect 40844 55636 40892 55692
rect 40948 55636 40958 55692
rect 49258 55636 49268 55692
rect 49324 55636 49372 55692
rect 49428 55636 49476 55692
rect 49532 55636 49580 55692
rect 49636 55636 49684 55692
rect 49740 55636 49788 55692
rect 49844 55636 49892 55692
rect 49948 55636 49958 55692
rect 58258 55636 58268 55692
rect 58324 55636 58372 55692
rect 58428 55636 58476 55692
rect 58532 55636 58580 55692
rect 58636 55636 58684 55692
rect 58740 55636 58788 55692
rect 58844 55636 58892 55692
rect 58948 55636 58958 55692
rect 67258 55636 67268 55692
rect 67324 55636 67372 55692
rect 67428 55636 67476 55692
rect 67532 55636 67580 55692
rect 67636 55636 67684 55692
rect 67740 55636 67788 55692
rect 67844 55636 67892 55692
rect 67948 55636 67958 55692
rect 76258 55636 76268 55692
rect 76324 55636 76372 55692
rect 76428 55636 76476 55692
rect 76532 55636 76580 55692
rect 76636 55636 76684 55692
rect 76740 55636 76788 55692
rect 76844 55636 76892 55692
rect 76948 55636 76958 55692
rect 85258 55636 85268 55692
rect 85324 55636 85372 55692
rect 85428 55636 85476 55692
rect 85532 55636 85580 55692
rect 85636 55636 85684 55692
rect 85740 55636 85788 55692
rect 85844 55636 85892 55692
rect 85948 55636 85958 55692
rect 94258 55636 94268 55692
rect 94324 55636 94372 55692
rect 94428 55636 94476 55692
rect 94532 55636 94580 55692
rect 94636 55636 94684 55692
rect 94740 55636 94788 55692
rect 94844 55636 94892 55692
rect 94948 55636 94958 55692
rect 0 55580 1708 55636
rect 1764 55580 2492 55636
rect 2548 55580 2558 55636
rect 0 55552 800 55580
rect 29250 55244 29260 55300
rect 29316 55244 33180 55300
rect 33236 55244 33628 55300
rect 33684 55244 37100 55300
rect 37156 55244 39788 55300
rect 39844 55244 43596 55300
rect 43652 55244 43708 55300
rect 43764 55244 44268 55300
rect 44324 55244 45164 55300
rect 45220 55244 45230 55300
rect 45938 55132 45948 55188
rect 46004 55132 48860 55188
rect 48916 55132 48926 55188
rect 1698 55020 1708 55076
rect 1764 55020 2492 55076
rect 2548 55020 2558 55076
rect 51762 55020 51772 55076
rect 51828 55020 52780 55076
rect 52836 55020 52846 55076
rect 53106 55020 53116 55076
rect 53172 55020 55468 55076
rect 57586 55020 57596 55076
rect 57652 55020 60508 55076
rect 60564 55020 60574 55076
rect 68674 55020 68684 55076
rect 68740 55020 81676 55076
rect 81732 55020 81742 55076
rect 8758 54852 8768 54908
rect 8824 54852 8872 54908
rect 8928 54852 8976 54908
rect 9032 54852 9080 54908
rect 9136 54852 9184 54908
rect 9240 54852 9288 54908
rect 9344 54852 9392 54908
rect 9448 54852 9458 54908
rect 17758 54852 17768 54908
rect 17824 54852 17872 54908
rect 17928 54852 17976 54908
rect 18032 54852 18080 54908
rect 18136 54852 18184 54908
rect 18240 54852 18288 54908
rect 18344 54852 18392 54908
rect 18448 54852 18458 54908
rect 26758 54852 26768 54908
rect 26824 54852 26872 54908
rect 26928 54852 26976 54908
rect 27032 54852 27080 54908
rect 27136 54852 27184 54908
rect 27240 54852 27288 54908
rect 27344 54852 27392 54908
rect 27448 54852 27458 54908
rect 35758 54852 35768 54908
rect 35824 54852 35872 54908
rect 35928 54852 35976 54908
rect 36032 54852 36080 54908
rect 36136 54852 36184 54908
rect 36240 54852 36288 54908
rect 36344 54852 36392 54908
rect 36448 54852 36458 54908
rect 44758 54852 44768 54908
rect 44824 54852 44872 54908
rect 44928 54852 44976 54908
rect 45032 54852 45080 54908
rect 45136 54852 45184 54908
rect 45240 54852 45288 54908
rect 45344 54852 45392 54908
rect 45448 54852 45458 54908
rect 53758 54852 53768 54908
rect 53824 54852 53872 54908
rect 53928 54852 53976 54908
rect 54032 54852 54080 54908
rect 54136 54852 54184 54908
rect 54240 54852 54288 54908
rect 54344 54852 54392 54908
rect 54448 54852 54458 54908
rect 55412 54852 55468 55020
rect 99200 54964 100000 54992
rect 98018 54908 98028 54964
rect 98084 54908 100000 54964
rect 62758 54852 62768 54908
rect 62824 54852 62872 54908
rect 62928 54852 62976 54908
rect 63032 54852 63080 54908
rect 63136 54852 63184 54908
rect 63240 54852 63288 54908
rect 63344 54852 63392 54908
rect 63448 54852 63458 54908
rect 71758 54852 71768 54908
rect 71824 54852 71872 54908
rect 71928 54852 71976 54908
rect 72032 54852 72080 54908
rect 72136 54852 72184 54908
rect 72240 54852 72288 54908
rect 72344 54852 72392 54908
rect 72448 54852 72458 54908
rect 80758 54852 80768 54908
rect 80824 54852 80872 54908
rect 80928 54852 80976 54908
rect 81032 54852 81080 54908
rect 81136 54852 81184 54908
rect 81240 54852 81288 54908
rect 81344 54852 81392 54908
rect 81448 54852 81458 54908
rect 89758 54852 89768 54908
rect 89824 54852 89872 54908
rect 89928 54852 89976 54908
rect 90032 54852 90080 54908
rect 90136 54852 90184 54908
rect 90240 54852 90288 54908
rect 90344 54852 90392 54908
rect 90448 54852 90458 54908
rect 99200 54880 100000 54908
rect 55412 54796 57820 54852
rect 57876 54796 57886 54852
rect 47730 54684 47740 54740
rect 47796 54684 59164 54740
rect 59220 54684 59230 54740
rect 41906 54572 41916 54628
rect 41972 54572 44156 54628
rect 44212 54572 44222 54628
rect 44594 54572 44604 54628
rect 44660 54572 44670 54628
rect 47954 54572 47964 54628
rect 48020 54572 49756 54628
rect 49812 54572 49822 54628
rect 57698 54572 57708 54628
rect 57764 54572 58380 54628
rect 58436 54572 59500 54628
rect 59556 54572 59566 54628
rect 0 54516 800 54544
rect 44604 54516 44660 54572
rect 0 54460 1708 54516
rect 1764 54460 1774 54516
rect 38882 54460 38892 54516
rect 38948 54460 40236 54516
rect 40292 54460 42588 54516
rect 42644 54460 44660 54516
rect 47852 54460 48748 54516
rect 48804 54460 52668 54516
rect 52724 54460 55580 54516
rect 55636 54460 56812 54516
rect 56868 54460 56878 54516
rect 0 54432 800 54460
rect 47852 54404 47908 54460
rect 39890 54348 39900 54404
rect 39956 54348 43260 54404
rect 43316 54348 43326 54404
rect 44146 54348 44156 54404
rect 44212 54348 47908 54404
rect 48066 54348 48076 54404
rect 48132 54348 52892 54404
rect 52948 54348 52958 54404
rect 57810 54348 57820 54404
rect 57876 54348 66780 54404
rect 66836 54348 66846 54404
rect 44930 54236 44940 54292
rect 44996 54236 56140 54292
rect 56196 54236 56812 54292
rect 56868 54236 56878 54292
rect 57474 54236 57484 54292
rect 57540 54236 58380 54292
rect 58436 54236 59276 54292
rect 59332 54236 59342 54292
rect 43250 54124 43260 54180
rect 43316 54124 44828 54180
rect 44884 54124 44894 54180
rect 52882 54124 52892 54180
rect 52948 54124 54236 54180
rect 54292 54124 54302 54180
rect 4258 54068 4268 54124
rect 4324 54068 4372 54124
rect 4428 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4788 54124
rect 4844 54068 4892 54124
rect 4948 54068 4958 54124
rect 13258 54068 13268 54124
rect 13324 54068 13372 54124
rect 13428 54068 13476 54124
rect 13532 54068 13580 54124
rect 13636 54068 13684 54124
rect 13740 54068 13788 54124
rect 13844 54068 13892 54124
rect 13948 54068 13958 54124
rect 22258 54068 22268 54124
rect 22324 54068 22372 54124
rect 22428 54068 22476 54124
rect 22532 54068 22580 54124
rect 22636 54068 22684 54124
rect 22740 54068 22788 54124
rect 22844 54068 22892 54124
rect 22948 54068 22958 54124
rect 31258 54068 31268 54124
rect 31324 54068 31372 54124
rect 31428 54068 31476 54124
rect 31532 54068 31580 54124
rect 31636 54068 31684 54124
rect 31740 54068 31788 54124
rect 31844 54068 31892 54124
rect 31948 54068 31958 54124
rect 40258 54068 40268 54124
rect 40324 54068 40372 54124
rect 40428 54068 40476 54124
rect 40532 54068 40580 54124
rect 40636 54068 40684 54124
rect 40740 54068 40788 54124
rect 40844 54068 40892 54124
rect 40948 54068 40958 54124
rect 49258 54068 49268 54124
rect 49324 54068 49372 54124
rect 49428 54068 49476 54124
rect 49532 54068 49580 54124
rect 49636 54068 49684 54124
rect 49740 54068 49788 54124
rect 49844 54068 49892 54124
rect 49948 54068 49958 54124
rect 58258 54068 58268 54124
rect 58324 54068 58372 54124
rect 58428 54068 58476 54124
rect 58532 54068 58580 54124
rect 58636 54068 58684 54124
rect 58740 54068 58788 54124
rect 58844 54068 58892 54124
rect 58948 54068 58958 54124
rect 67258 54068 67268 54124
rect 67324 54068 67372 54124
rect 67428 54068 67476 54124
rect 67532 54068 67580 54124
rect 67636 54068 67684 54124
rect 67740 54068 67788 54124
rect 67844 54068 67892 54124
rect 67948 54068 67958 54124
rect 76258 54068 76268 54124
rect 76324 54068 76372 54124
rect 76428 54068 76476 54124
rect 76532 54068 76580 54124
rect 76636 54068 76684 54124
rect 76740 54068 76788 54124
rect 76844 54068 76892 54124
rect 76948 54068 76958 54124
rect 85258 54068 85268 54124
rect 85324 54068 85372 54124
rect 85428 54068 85476 54124
rect 85532 54068 85580 54124
rect 85636 54068 85684 54124
rect 85740 54068 85788 54124
rect 85844 54068 85892 54124
rect 85948 54068 85958 54124
rect 94258 54068 94268 54124
rect 94324 54068 94372 54124
rect 94428 54068 94476 54124
rect 94532 54068 94580 54124
rect 94636 54068 94684 54124
rect 94740 54068 94788 54124
rect 94844 54068 94892 54124
rect 94948 54068 94958 54124
rect 28466 53900 28476 53956
rect 28532 53900 46732 53956
rect 46788 53900 46798 53956
rect 66546 53900 66556 53956
rect 66612 53900 67116 53956
rect 67172 53900 68348 53956
rect 68404 53900 68414 53956
rect 33954 53788 33964 53844
rect 34020 53788 35084 53844
rect 35140 53788 35150 53844
rect 35634 53788 35644 53844
rect 35700 53788 36764 53844
rect 36820 53788 36830 53844
rect 40114 53788 40124 53844
rect 40180 53788 41468 53844
rect 41524 53788 41534 53844
rect 57362 53788 57372 53844
rect 57428 53788 58044 53844
rect 58100 53788 58110 53844
rect 60162 53788 60172 53844
rect 60228 53788 65324 53844
rect 65380 53788 65390 53844
rect 36530 53676 36540 53732
rect 36596 53676 38220 53732
rect 38276 53676 39228 53732
rect 39284 53676 39294 53732
rect 44930 53676 44940 53732
rect 44996 53676 45948 53732
rect 46004 53676 50092 53732
rect 50148 53676 50158 53732
rect 51202 53676 51212 53732
rect 51268 53676 53900 53732
rect 53956 53676 53966 53732
rect 55412 53676 62076 53732
rect 62132 53676 62142 53732
rect 65202 53676 65212 53732
rect 65268 53676 66108 53732
rect 66164 53676 66892 53732
rect 66948 53676 66958 53732
rect 55412 53620 55468 53676
rect 30818 53564 30828 53620
rect 30884 53564 32060 53620
rect 32116 53564 35420 53620
rect 35476 53564 35486 53620
rect 35858 53564 35868 53620
rect 35924 53564 36596 53620
rect 50418 53564 50428 53620
rect 50484 53564 51660 53620
rect 51716 53564 55468 53620
rect 57810 53564 57820 53620
rect 57876 53564 64876 53620
rect 64932 53564 64942 53620
rect 66658 53564 66668 53620
rect 66724 53564 70700 53620
rect 70756 53564 70766 53620
rect 36540 53508 36596 53564
rect 29922 53452 29932 53508
rect 29988 53452 30716 53508
rect 30772 53452 30782 53508
rect 31266 53452 31276 53508
rect 31332 53452 34412 53508
rect 34468 53452 34478 53508
rect 34626 53452 34636 53508
rect 34692 53452 35196 53508
rect 35252 53452 36204 53508
rect 36260 53452 36270 53508
rect 36530 53452 36540 53508
rect 36596 53452 36606 53508
rect 47730 53452 47740 53508
rect 47796 53452 50764 53508
rect 50820 53452 51100 53508
rect 51156 53452 56028 53508
rect 56084 53452 56094 53508
rect 56354 53452 56364 53508
rect 56420 53452 66332 53508
rect 66388 53452 66398 53508
rect 67666 53452 67676 53508
rect 67732 53452 72828 53508
rect 72884 53452 75740 53508
rect 75796 53452 75806 53508
rect 0 53396 800 53424
rect 31276 53396 31332 53452
rect 56028 53396 56084 53452
rect 0 53340 1708 53396
rect 1764 53340 2492 53396
rect 2548 53340 2558 53396
rect 29250 53340 29260 53396
rect 29316 53340 30156 53396
rect 30212 53340 31332 53396
rect 36978 53340 36988 53396
rect 37044 53340 39452 53396
rect 39508 53340 39518 53396
rect 56028 53340 57484 53396
rect 57540 53340 57550 53396
rect 0 53312 800 53340
rect 8758 53284 8768 53340
rect 8824 53284 8872 53340
rect 8928 53284 8976 53340
rect 9032 53284 9080 53340
rect 9136 53284 9184 53340
rect 9240 53284 9288 53340
rect 9344 53284 9392 53340
rect 9448 53284 9458 53340
rect 17758 53284 17768 53340
rect 17824 53284 17872 53340
rect 17928 53284 17976 53340
rect 18032 53284 18080 53340
rect 18136 53284 18184 53340
rect 18240 53284 18288 53340
rect 18344 53284 18392 53340
rect 18448 53284 18458 53340
rect 26758 53284 26768 53340
rect 26824 53284 26872 53340
rect 26928 53284 26976 53340
rect 27032 53284 27080 53340
rect 27136 53284 27184 53340
rect 27240 53284 27288 53340
rect 27344 53284 27392 53340
rect 27448 53284 27458 53340
rect 35758 53284 35768 53340
rect 35824 53284 35872 53340
rect 35928 53284 35976 53340
rect 36032 53284 36080 53340
rect 36136 53284 36184 53340
rect 36240 53284 36288 53340
rect 36344 53284 36392 53340
rect 36448 53284 36458 53340
rect 44758 53284 44768 53340
rect 44824 53284 44872 53340
rect 44928 53284 44976 53340
rect 45032 53284 45080 53340
rect 45136 53284 45184 53340
rect 45240 53284 45288 53340
rect 45344 53284 45392 53340
rect 45448 53284 45458 53340
rect 53758 53284 53768 53340
rect 53824 53284 53872 53340
rect 53928 53284 53976 53340
rect 54032 53284 54080 53340
rect 54136 53284 54184 53340
rect 54240 53284 54288 53340
rect 54344 53284 54392 53340
rect 54448 53284 54458 53340
rect 62758 53284 62768 53340
rect 62824 53284 62872 53340
rect 62928 53284 62976 53340
rect 63032 53284 63080 53340
rect 63136 53284 63184 53340
rect 63240 53284 63288 53340
rect 63344 53284 63392 53340
rect 63448 53284 63458 53340
rect 71758 53284 71768 53340
rect 71824 53284 71872 53340
rect 71928 53284 71976 53340
rect 72032 53284 72080 53340
rect 72136 53284 72184 53340
rect 72240 53284 72288 53340
rect 72344 53284 72392 53340
rect 72448 53284 72458 53340
rect 80758 53284 80768 53340
rect 80824 53284 80872 53340
rect 80928 53284 80976 53340
rect 81032 53284 81080 53340
rect 81136 53284 81184 53340
rect 81240 53284 81288 53340
rect 81344 53284 81392 53340
rect 81448 53284 81458 53340
rect 89758 53284 89768 53340
rect 89824 53284 89872 53340
rect 89928 53284 89976 53340
rect 90032 53284 90080 53340
rect 90136 53284 90184 53340
rect 90240 53284 90288 53340
rect 90344 53284 90392 53340
rect 90448 53284 90458 53340
rect 39554 53228 39564 53284
rect 39620 53228 40908 53284
rect 40964 53228 40974 53284
rect 55412 53228 56476 53284
rect 56532 53228 58044 53284
rect 58100 53228 58110 53284
rect 29586 53116 29596 53172
rect 29652 53116 35532 53172
rect 35588 53116 35598 53172
rect 35858 53116 35868 53172
rect 35924 53116 36988 53172
rect 37044 53116 37054 53172
rect 38322 53116 38332 53172
rect 38388 53116 47292 53172
rect 47348 53116 47358 53172
rect 50194 53116 50204 53172
rect 50260 53116 50876 53172
rect 50932 53116 50942 53172
rect 25778 53004 25788 53060
rect 25844 53004 29372 53060
rect 29428 53004 29820 53060
rect 29876 53004 29886 53060
rect 31154 53004 31164 53060
rect 31220 53004 33740 53060
rect 33796 53004 41916 53060
rect 41972 53004 41982 53060
rect 43810 53004 43820 53060
rect 43876 53004 45500 53060
rect 45556 53004 46060 53060
rect 46116 53004 46126 53060
rect 55412 52948 55468 53228
rect 99200 53172 100000 53200
rect 57698 53116 57708 53172
rect 57764 53116 67228 53172
rect 67284 53116 67294 53172
rect 98018 53116 98028 53172
rect 98084 53116 100000 53172
rect 99200 53088 100000 53116
rect 57138 53004 57148 53060
rect 57204 53004 64540 53060
rect 64596 53004 65436 53060
rect 65492 53004 65502 53060
rect 27682 52892 27692 52948
rect 27748 52892 28812 52948
rect 28868 52892 28878 52948
rect 31266 52892 31276 52948
rect 31332 52892 31948 52948
rect 32004 52892 34300 52948
rect 34356 52892 34366 52948
rect 35410 52892 35420 52948
rect 35476 52892 37212 52948
rect 37268 52892 37278 52948
rect 41122 52892 41132 52948
rect 41188 52892 42700 52948
rect 42756 52892 42766 52948
rect 48178 52892 48188 52948
rect 48244 52892 49420 52948
rect 49476 52892 49486 52948
rect 54460 52892 55468 52948
rect 55570 52892 55580 52948
rect 55636 52892 56588 52948
rect 56644 52892 56654 52948
rect 58930 52892 58940 52948
rect 58996 52892 59006 52948
rect 65202 52892 65212 52948
rect 65268 52892 68796 52948
rect 68852 52892 69580 52948
rect 69636 52892 69646 52948
rect 54460 52836 54516 52892
rect 58940 52836 58996 52892
rect 1698 52780 1708 52836
rect 1764 52780 2492 52836
rect 2548 52780 2558 52836
rect 25106 52780 25116 52836
rect 25172 52780 28028 52836
rect 28084 52780 28094 52836
rect 28578 52780 28588 52836
rect 28644 52780 35644 52836
rect 35700 52780 35710 52836
rect 36530 52780 36540 52836
rect 36596 52780 38444 52836
rect 38500 52780 38510 52836
rect 49074 52780 49084 52836
rect 49140 52780 54460 52836
rect 54516 52780 54526 52836
rect 55122 52780 55132 52836
rect 55188 52780 58996 52836
rect 62066 52780 62076 52836
rect 62132 52780 81452 52836
rect 81508 52780 81518 52836
rect 30146 52668 30156 52724
rect 30212 52668 32172 52724
rect 32228 52668 32238 52724
rect 34290 52668 34300 52724
rect 34356 52668 35756 52724
rect 35812 52668 41692 52724
rect 41748 52668 42028 52724
rect 42084 52668 42094 52724
rect 49084 52668 49980 52724
rect 50036 52668 56028 52724
rect 56084 52668 56924 52724
rect 56980 52668 56990 52724
rect 57362 52668 57372 52724
rect 57428 52668 62636 52724
rect 62692 52668 62702 52724
rect 66546 52668 66556 52724
rect 66612 52668 68124 52724
rect 68180 52668 71260 52724
rect 71316 52668 71326 52724
rect 49084 52612 49140 52668
rect 35634 52556 35644 52612
rect 35700 52556 37324 52612
rect 37380 52556 37390 52612
rect 38612 52556 39228 52612
rect 39284 52556 40124 52612
rect 40180 52556 40190 52612
rect 44706 52556 44716 52612
rect 44772 52556 45612 52612
rect 45668 52556 47740 52612
rect 47796 52556 47806 52612
rect 49074 52556 49084 52612
rect 49140 52556 49150 52612
rect 4258 52500 4268 52556
rect 4324 52500 4372 52556
rect 4428 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4788 52556
rect 4844 52500 4892 52556
rect 4948 52500 4958 52556
rect 13258 52500 13268 52556
rect 13324 52500 13372 52556
rect 13428 52500 13476 52556
rect 13532 52500 13580 52556
rect 13636 52500 13684 52556
rect 13740 52500 13788 52556
rect 13844 52500 13892 52556
rect 13948 52500 13958 52556
rect 22258 52500 22268 52556
rect 22324 52500 22372 52556
rect 22428 52500 22476 52556
rect 22532 52500 22580 52556
rect 22636 52500 22684 52556
rect 22740 52500 22788 52556
rect 22844 52500 22892 52556
rect 22948 52500 22958 52556
rect 31258 52500 31268 52556
rect 31324 52500 31372 52556
rect 31428 52500 31476 52556
rect 31532 52500 31580 52556
rect 31636 52500 31684 52556
rect 31740 52500 31788 52556
rect 31844 52500 31892 52556
rect 31948 52500 31958 52556
rect 38612 52500 38668 52556
rect 40258 52500 40268 52556
rect 40324 52500 40372 52556
rect 40428 52500 40476 52556
rect 40532 52500 40580 52556
rect 40636 52500 40684 52556
rect 40740 52500 40788 52556
rect 40844 52500 40892 52556
rect 40948 52500 40958 52556
rect 26852 52444 28588 52500
rect 28644 52444 28654 52500
rect 34402 52444 34412 52500
rect 34468 52444 34972 52500
rect 35028 52444 38668 52500
rect 41458 52444 41468 52500
rect 41524 52444 41692 52500
rect 41748 52444 43932 52500
rect 43988 52444 46172 52500
rect 46228 52444 48748 52500
rect 48804 52444 48814 52500
rect 0 52276 800 52304
rect 26852 52276 26908 52444
rect 49084 52388 49140 52556
rect 49258 52500 49268 52556
rect 49324 52500 49372 52556
rect 49428 52500 49476 52556
rect 49532 52500 49580 52556
rect 49636 52500 49684 52556
rect 49740 52500 49788 52556
rect 49844 52500 49892 52556
rect 49948 52500 49958 52556
rect 58258 52500 58268 52556
rect 58324 52500 58372 52556
rect 58428 52500 58476 52556
rect 58532 52500 58580 52556
rect 58636 52500 58684 52556
rect 58740 52500 58788 52556
rect 58844 52500 58892 52556
rect 58948 52500 58958 52556
rect 67258 52500 67268 52556
rect 67324 52500 67372 52556
rect 67428 52500 67476 52556
rect 67532 52500 67580 52556
rect 67636 52500 67684 52556
rect 67740 52500 67788 52556
rect 67844 52500 67892 52556
rect 67948 52500 67958 52556
rect 76258 52500 76268 52556
rect 76324 52500 76372 52556
rect 76428 52500 76476 52556
rect 76532 52500 76580 52556
rect 76636 52500 76684 52556
rect 76740 52500 76788 52556
rect 76844 52500 76892 52556
rect 76948 52500 76958 52556
rect 85258 52500 85268 52556
rect 85324 52500 85372 52556
rect 85428 52500 85476 52556
rect 85532 52500 85580 52556
rect 85636 52500 85684 52556
rect 85740 52500 85788 52556
rect 85844 52500 85892 52556
rect 85948 52500 85958 52556
rect 94258 52500 94268 52556
rect 94324 52500 94372 52556
rect 94428 52500 94476 52556
rect 94532 52500 94580 52556
rect 94636 52500 94684 52556
rect 94740 52500 94788 52556
rect 94844 52500 94892 52556
rect 94948 52500 94958 52556
rect 50194 52444 50204 52500
rect 50260 52444 50764 52500
rect 50820 52444 57932 52500
rect 57988 52444 57998 52500
rect 28466 52332 28476 52388
rect 28532 52332 31052 52388
rect 31108 52332 31118 52388
rect 32162 52332 32172 52388
rect 32228 52332 35308 52388
rect 35364 52332 35374 52388
rect 41570 52332 41580 52388
rect 41636 52332 49140 52388
rect 49746 52332 49756 52388
rect 49812 52332 50428 52388
rect 50484 52332 52444 52388
rect 52500 52332 53340 52388
rect 53396 52332 55132 52388
rect 55188 52332 55198 52388
rect 56802 52332 56812 52388
rect 56868 52332 57260 52388
rect 57316 52332 58492 52388
rect 58548 52332 58558 52388
rect 0 52220 1708 52276
rect 1764 52220 1774 52276
rect 22978 52220 22988 52276
rect 23044 52220 26908 52276
rect 28354 52220 28364 52276
rect 28420 52220 29260 52276
rect 29316 52220 31276 52276
rect 31332 52220 31342 52276
rect 45948 52220 47180 52276
rect 47236 52220 48300 52276
rect 48356 52220 52108 52276
rect 52164 52220 53788 52276
rect 53844 52220 54348 52276
rect 54404 52220 55020 52276
rect 55076 52220 55086 52276
rect 58146 52220 58156 52276
rect 58212 52220 58604 52276
rect 58660 52220 59052 52276
rect 59108 52220 60508 52276
rect 60564 52220 60574 52276
rect 0 52192 800 52220
rect 45948 52164 46004 52220
rect 28130 52108 28140 52164
rect 28196 52108 28812 52164
rect 28868 52108 30156 52164
rect 30212 52108 30222 52164
rect 30818 52108 30828 52164
rect 30884 52108 32956 52164
rect 33012 52108 34244 52164
rect 35298 52108 35308 52164
rect 35364 52108 36204 52164
rect 36260 52108 36270 52164
rect 42018 52108 42028 52164
rect 42084 52108 43260 52164
rect 43316 52108 43708 52164
rect 43764 52108 45948 52164
rect 46004 52108 46014 52164
rect 46610 52108 46620 52164
rect 46676 52108 49644 52164
rect 49700 52108 49710 52164
rect 55682 52108 55692 52164
rect 55748 52108 56812 52164
rect 56868 52108 56878 52164
rect 58034 52108 58044 52164
rect 58100 52108 61852 52164
rect 61908 52108 63420 52164
rect 63476 52108 63868 52164
rect 63924 52108 65100 52164
rect 65156 52108 65166 52164
rect 34188 52052 34244 52108
rect 26898 51996 26908 52052
rect 26964 51996 27804 52052
rect 27860 51996 27870 52052
rect 34178 51996 34188 52052
rect 34244 51996 37996 52052
rect 38052 51996 38892 52052
rect 38948 51996 39564 52052
rect 39620 51996 39630 52052
rect 46386 51996 46396 52052
rect 46452 51996 46956 52052
rect 47012 51996 47022 52052
rect 55794 51996 55804 52052
rect 55860 51996 56476 52052
rect 56532 51996 56542 52052
rect 26226 51884 26236 51940
rect 26292 51884 27020 51940
rect 27076 51884 27086 51940
rect 46162 51884 46172 51940
rect 46228 51884 46732 51940
rect 46788 51884 47852 51940
rect 47908 51884 47918 51940
rect 8758 51716 8768 51772
rect 8824 51716 8872 51772
rect 8928 51716 8976 51772
rect 9032 51716 9080 51772
rect 9136 51716 9184 51772
rect 9240 51716 9288 51772
rect 9344 51716 9392 51772
rect 9448 51716 9458 51772
rect 17758 51716 17768 51772
rect 17824 51716 17872 51772
rect 17928 51716 17976 51772
rect 18032 51716 18080 51772
rect 18136 51716 18184 51772
rect 18240 51716 18288 51772
rect 18344 51716 18392 51772
rect 18448 51716 18458 51772
rect 26758 51716 26768 51772
rect 26824 51716 26872 51772
rect 26928 51716 26976 51772
rect 27032 51716 27080 51772
rect 27136 51716 27184 51772
rect 27240 51716 27288 51772
rect 27344 51716 27392 51772
rect 27448 51716 27458 51772
rect 35758 51716 35768 51772
rect 35824 51716 35872 51772
rect 35928 51716 35976 51772
rect 36032 51716 36080 51772
rect 36136 51716 36184 51772
rect 36240 51716 36288 51772
rect 36344 51716 36392 51772
rect 36448 51716 36458 51772
rect 44758 51716 44768 51772
rect 44824 51716 44872 51772
rect 44928 51716 44976 51772
rect 45032 51716 45080 51772
rect 45136 51716 45184 51772
rect 45240 51716 45288 51772
rect 45344 51716 45392 51772
rect 45448 51716 45458 51772
rect 53758 51716 53768 51772
rect 53824 51716 53872 51772
rect 53928 51716 53976 51772
rect 54032 51716 54080 51772
rect 54136 51716 54184 51772
rect 54240 51716 54288 51772
rect 54344 51716 54392 51772
rect 54448 51716 54458 51772
rect 62758 51716 62768 51772
rect 62824 51716 62872 51772
rect 62928 51716 62976 51772
rect 63032 51716 63080 51772
rect 63136 51716 63184 51772
rect 63240 51716 63288 51772
rect 63344 51716 63392 51772
rect 63448 51716 63458 51772
rect 71758 51716 71768 51772
rect 71824 51716 71872 51772
rect 71928 51716 71976 51772
rect 72032 51716 72080 51772
rect 72136 51716 72184 51772
rect 72240 51716 72288 51772
rect 72344 51716 72392 51772
rect 72448 51716 72458 51772
rect 80758 51716 80768 51772
rect 80824 51716 80872 51772
rect 80928 51716 80976 51772
rect 81032 51716 81080 51772
rect 81136 51716 81184 51772
rect 81240 51716 81288 51772
rect 81344 51716 81392 51772
rect 81448 51716 81458 51772
rect 89758 51716 89768 51772
rect 89824 51716 89872 51772
rect 89928 51716 89976 51772
rect 90032 51716 90080 51772
rect 90136 51716 90184 51772
rect 90240 51716 90288 51772
rect 90344 51716 90392 51772
rect 90448 51716 90458 51772
rect 2034 51660 2044 51716
rect 2100 51660 5852 51716
rect 5908 51660 5918 51716
rect 38658 51548 38668 51604
rect 38724 51548 39676 51604
rect 39732 51548 40124 51604
rect 40180 51548 44604 51604
rect 44660 51548 44670 51604
rect 90962 51548 90972 51604
rect 91028 51548 97020 51604
rect 97076 51548 97086 51604
rect 39554 51436 39564 51492
rect 39620 51436 40908 51492
rect 40964 51436 41580 51492
rect 41636 51436 41646 51492
rect 71362 51436 71372 51492
rect 71428 51436 72492 51492
rect 72548 51436 72558 51492
rect 99200 51380 100000 51408
rect 36530 51324 36540 51380
rect 36596 51324 38444 51380
rect 38500 51324 39116 51380
rect 39172 51324 41692 51380
rect 41748 51324 41758 51380
rect 42242 51324 42252 51380
rect 42308 51324 46396 51380
rect 46452 51324 46462 51380
rect 46722 51324 46732 51380
rect 46788 51324 47404 51380
rect 47460 51324 47470 51380
rect 97682 51324 97692 51380
rect 97748 51324 100000 51380
rect 99200 51296 100000 51324
rect 54786 51212 54796 51268
rect 54852 51212 61740 51268
rect 61796 51212 62188 51268
rect 62244 51212 62254 51268
rect 74274 51212 74284 51268
rect 74340 51212 76636 51268
rect 76692 51212 79660 51268
rect 79716 51212 79726 51268
rect 0 51156 800 51184
rect 0 51100 1708 51156
rect 1764 51100 2492 51156
rect 2548 51100 2558 51156
rect 0 51072 800 51100
rect 4258 50932 4268 50988
rect 4324 50932 4372 50988
rect 4428 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4788 50988
rect 4844 50932 4892 50988
rect 4948 50932 4958 50988
rect 13258 50932 13268 50988
rect 13324 50932 13372 50988
rect 13428 50932 13476 50988
rect 13532 50932 13580 50988
rect 13636 50932 13684 50988
rect 13740 50932 13788 50988
rect 13844 50932 13892 50988
rect 13948 50932 13958 50988
rect 22258 50932 22268 50988
rect 22324 50932 22372 50988
rect 22428 50932 22476 50988
rect 22532 50932 22580 50988
rect 22636 50932 22684 50988
rect 22740 50932 22788 50988
rect 22844 50932 22892 50988
rect 22948 50932 22958 50988
rect 31258 50932 31268 50988
rect 31324 50932 31372 50988
rect 31428 50932 31476 50988
rect 31532 50932 31580 50988
rect 31636 50932 31684 50988
rect 31740 50932 31788 50988
rect 31844 50932 31892 50988
rect 31948 50932 31958 50988
rect 40258 50932 40268 50988
rect 40324 50932 40372 50988
rect 40428 50932 40476 50988
rect 40532 50932 40580 50988
rect 40636 50932 40684 50988
rect 40740 50932 40788 50988
rect 40844 50932 40892 50988
rect 40948 50932 40958 50988
rect 49258 50932 49268 50988
rect 49324 50932 49372 50988
rect 49428 50932 49476 50988
rect 49532 50932 49580 50988
rect 49636 50932 49684 50988
rect 49740 50932 49788 50988
rect 49844 50932 49892 50988
rect 49948 50932 49958 50988
rect 58258 50932 58268 50988
rect 58324 50932 58372 50988
rect 58428 50932 58476 50988
rect 58532 50932 58580 50988
rect 58636 50932 58684 50988
rect 58740 50932 58788 50988
rect 58844 50932 58892 50988
rect 58948 50932 58958 50988
rect 67258 50932 67268 50988
rect 67324 50932 67372 50988
rect 67428 50932 67476 50988
rect 67532 50932 67580 50988
rect 67636 50932 67684 50988
rect 67740 50932 67788 50988
rect 67844 50932 67892 50988
rect 67948 50932 67958 50988
rect 76258 50932 76268 50988
rect 76324 50932 76372 50988
rect 76428 50932 76476 50988
rect 76532 50932 76580 50988
rect 76636 50932 76684 50988
rect 76740 50932 76788 50988
rect 76844 50932 76892 50988
rect 76948 50932 76958 50988
rect 85258 50932 85268 50988
rect 85324 50932 85372 50988
rect 85428 50932 85476 50988
rect 85532 50932 85580 50988
rect 85636 50932 85684 50988
rect 85740 50932 85788 50988
rect 85844 50932 85892 50988
rect 85948 50932 85958 50988
rect 94258 50932 94268 50988
rect 94324 50932 94372 50988
rect 94428 50932 94476 50988
rect 94532 50932 94580 50988
rect 94636 50932 94684 50988
rect 94740 50932 94788 50988
rect 94844 50932 94892 50988
rect 94948 50932 94958 50988
rect 43586 50764 43596 50820
rect 43652 50596 43708 50820
rect 39890 50540 39900 50596
rect 39956 50540 40796 50596
rect 40852 50540 45500 50596
rect 45556 50540 46172 50596
rect 46228 50540 50428 50596
rect 50484 50540 50494 50596
rect 76514 50540 76524 50596
rect 76580 50540 77308 50596
rect 77364 50540 77374 50596
rect 1922 50428 1932 50484
rect 1988 50428 16156 50484
rect 16212 50428 17276 50484
rect 17332 50428 17342 50484
rect 19618 50428 19628 50484
rect 19684 50428 20524 50484
rect 20580 50428 20860 50484
rect 20916 50428 20926 50484
rect 33730 50428 33740 50484
rect 33796 50428 40460 50484
rect 40516 50428 43596 50484
rect 43652 50428 46060 50484
rect 46116 50428 49084 50484
rect 49140 50428 49150 50484
rect 63298 50428 63308 50484
rect 63364 50428 64540 50484
rect 64596 50428 67228 50484
rect 73154 50428 73164 50484
rect 73220 50428 74284 50484
rect 74340 50428 74956 50484
rect 75012 50428 75022 50484
rect 77970 50428 77980 50484
rect 78036 50428 80444 50484
rect 80500 50428 80510 50484
rect 67172 50372 67228 50428
rect 2034 50316 2044 50372
rect 2100 50316 2828 50372
rect 2884 50316 2894 50372
rect 29474 50316 29484 50372
rect 29540 50316 29932 50372
rect 29988 50316 29998 50372
rect 67172 50316 68124 50372
rect 68180 50316 69244 50372
rect 69300 50316 69310 50372
rect 8758 50148 8768 50204
rect 8824 50148 8872 50204
rect 8928 50148 8976 50204
rect 9032 50148 9080 50204
rect 9136 50148 9184 50204
rect 9240 50148 9288 50204
rect 9344 50148 9392 50204
rect 9448 50148 9458 50204
rect 17758 50148 17768 50204
rect 17824 50148 17872 50204
rect 17928 50148 17976 50204
rect 18032 50148 18080 50204
rect 18136 50148 18184 50204
rect 18240 50148 18288 50204
rect 18344 50148 18392 50204
rect 18448 50148 18458 50204
rect 26758 50148 26768 50204
rect 26824 50148 26872 50204
rect 26928 50148 26976 50204
rect 27032 50148 27080 50204
rect 27136 50148 27184 50204
rect 27240 50148 27288 50204
rect 27344 50148 27392 50204
rect 27448 50148 27458 50204
rect 35758 50148 35768 50204
rect 35824 50148 35872 50204
rect 35928 50148 35976 50204
rect 36032 50148 36080 50204
rect 36136 50148 36184 50204
rect 36240 50148 36288 50204
rect 36344 50148 36392 50204
rect 36448 50148 36458 50204
rect 44758 50148 44768 50204
rect 44824 50148 44872 50204
rect 44928 50148 44976 50204
rect 45032 50148 45080 50204
rect 45136 50148 45184 50204
rect 45240 50148 45288 50204
rect 45344 50148 45392 50204
rect 45448 50148 45458 50204
rect 53758 50148 53768 50204
rect 53824 50148 53872 50204
rect 53928 50148 53976 50204
rect 54032 50148 54080 50204
rect 54136 50148 54184 50204
rect 54240 50148 54288 50204
rect 54344 50148 54392 50204
rect 54448 50148 54458 50204
rect 62758 50148 62768 50204
rect 62824 50148 62872 50204
rect 62928 50148 62976 50204
rect 63032 50148 63080 50204
rect 63136 50148 63184 50204
rect 63240 50148 63288 50204
rect 63344 50148 63392 50204
rect 63448 50148 63458 50204
rect 71758 50148 71768 50204
rect 71824 50148 71872 50204
rect 71928 50148 71976 50204
rect 72032 50148 72080 50204
rect 72136 50148 72184 50204
rect 72240 50148 72288 50204
rect 72344 50148 72392 50204
rect 72448 50148 72458 50204
rect 80758 50148 80768 50204
rect 80824 50148 80872 50204
rect 80928 50148 80976 50204
rect 81032 50148 81080 50204
rect 81136 50148 81184 50204
rect 81240 50148 81288 50204
rect 81344 50148 81392 50204
rect 81448 50148 81458 50204
rect 89758 50148 89768 50204
rect 89824 50148 89872 50204
rect 89928 50148 89976 50204
rect 90032 50148 90080 50204
rect 90136 50148 90184 50204
rect 90240 50148 90288 50204
rect 90344 50148 90392 50204
rect 90448 50148 90458 50204
rect 0 50036 800 50064
rect 0 49980 1708 50036
rect 1764 49980 2492 50036
rect 2548 49980 2558 50036
rect 0 49952 800 49980
rect 10098 49868 10108 49924
rect 10164 49868 11340 49924
rect 11396 49868 14476 49924
rect 14532 49868 14542 49924
rect 37650 49868 37660 49924
rect 37716 49868 41132 49924
rect 41188 49868 41198 49924
rect 50306 49868 50316 49924
rect 50372 49868 51548 49924
rect 51604 49868 51614 49924
rect 10108 49700 10164 49868
rect 25554 49756 25564 49812
rect 25620 49756 26348 49812
rect 26404 49756 29036 49812
rect 29092 49756 29102 49812
rect 38434 49756 38444 49812
rect 38500 49756 38668 49812
rect 64978 49756 64988 49812
rect 65044 49756 65772 49812
rect 65828 49756 65838 49812
rect 75730 49756 75740 49812
rect 75796 49756 77196 49812
rect 77252 49756 77644 49812
rect 77700 49756 77710 49812
rect 38612 49700 38668 49756
rect 8306 49644 8316 49700
rect 8372 49644 10164 49700
rect 29922 49644 29932 49700
rect 29988 49644 31948 49700
rect 32004 49644 32014 49700
rect 38612 49644 39004 49700
rect 39060 49644 42252 49700
rect 42308 49644 42318 49700
rect 60610 49644 60620 49700
rect 60676 49644 61964 49700
rect 62020 49644 62300 49700
rect 62356 49644 71708 49700
rect 71764 49644 72940 49700
rect 72996 49644 76188 49700
rect 76244 49644 77420 49700
rect 77476 49644 77486 49700
rect 90514 49644 90524 49700
rect 90580 49644 92428 49700
rect 92484 49644 95452 49700
rect 95508 49644 95518 49700
rect 8372 49588 8428 49644
rect 99200 49588 100000 49616
rect 5842 49532 5852 49588
rect 5908 49532 8428 49588
rect 35522 49532 35532 49588
rect 35588 49532 42812 49588
rect 42868 49532 61292 49588
rect 61348 49532 62076 49588
rect 62132 49476 62188 49588
rect 62850 49532 62860 49588
rect 62916 49532 64092 49588
rect 64148 49532 64876 49588
rect 64932 49532 64942 49588
rect 65874 49532 65884 49588
rect 65940 49532 68908 49588
rect 68964 49532 68974 49588
rect 98018 49532 98028 49588
rect 98084 49532 100000 49588
rect 99200 49504 100000 49532
rect 62132 49420 63644 49476
rect 63700 49420 63710 49476
rect 4258 49364 4268 49420
rect 4324 49364 4372 49420
rect 4428 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4788 49420
rect 4844 49364 4892 49420
rect 4948 49364 4958 49420
rect 13258 49364 13268 49420
rect 13324 49364 13372 49420
rect 13428 49364 13476 49420
rect 13532 49364 13580 49420
rect 13636 49364 13684 49420
rect 13740 49364 13788 49420
rect 13844 49364 13892 49420
rect 13948 49364 13958 49420
rect 22258 49364 22268 49420
rect 22324 49364 22372 49420
rect 22428 49364 22476 49420
rect 22532 49364 22580 49420
rect 22636 49364 22684 49420
rect 22740 49364 22788 49420
rect 22844 49364 22892 49420
rect 22948 49364 22958 49420
rect 31258 49364 31268 49420
rect 31324 49364 31372 49420
rect 31428 49364 31476 49420
rect 31532 49364 31580 49420
rect 31636 49364 31684 49420
rect 31740 49364 31788 49420
rect 31844 49364 31892 49420
rect 31948 49364 31958 49420
rect 40258 49364 40268 49420
rect 40324 49364 40372 49420
rect 40428 49364 40476 49420
rect 40532 49364 40580 49420
rect 40636 49364 40684 49420
rect 40740 49364 40788 49420
rect 40844 49364 40892 49420
rect 40948 49364 40958 49420
rect 49258 49364 49268 49420
rect 49324 49364 49372 49420
rect 49428 49364 49476 49420
rect 49532 49364 49580 49420
rect 49636 49364 49684 49420
rect 49740 49364 49788 49420
rect 49844 49364 49892 49420
rect 49948 49364 49958 49420
rect 58258 49364 58268 49420
rect 58324 49364 58372 49420
rect 58428 49364 58476 49420
rect 58532 49364 58580 49420
rect 58636 49364 58684 49420
rect 58740 49364 58788 49420
rect 58844 49364 58892 49420
rect 58948 49364 58958 49420
rect 67258 49364 67268 49420
rect 67324 49364 67372 49420
rect 67428 49364 67476 49420
rect 67532 49364 67580 49420
rect 67636 49364 67684 49420
rect 67740 49364 67788 49420
rect 67844 49364 67892 49420
rect 67948 49364 67958 49420
rect 76258 49364 76268 49420
rect 76324 49364 76372 49420
rect 76428 49364 76476 49420
rect 76532 49364 76580 49420
rect 76636 49364 76684 49420
rect 76740 49364 76788 49420
rect 76844 49364 76892 49420
rect 76948 49364 76958 49420
rect 85258 49364 85268 49420
rect 85324 49364 85372 49420
rect 85428 49364 85476 49420
rect 85532 49364 85580 49420
rect 85636 49364 85684 49420
rect 85740 49364 85788 49420
rect 85844 49364 85892 49420
rect 85948 49364 85958 49420
rect 94258 49364 94268 49420
rect 94324 49364 94372 49420
rect 94428 49364 94476 49420
rect 94532 49364 94580 49420
rect 94636 49364 94684 49420
rect 94740 49364 94788 49420
rect 94844 49364 94892 49420
rect 94948 49364 94958 49420
rect 32834 49196 32844 49252
rect 32900 49196 35084 49252
rect 35140 49196 35150 49252
rect 29250 49084 29260 49140
rect 29316 49084 32284 49140
rect 32340 49084 35756 49140
rect 35812 49084 38668 49140
rect 38724 49084 39900 49140
rect 39956 49084 39966 49140
rect 77634 49084 77644 49140
rect 77700 49084 77980 49140
rect 78036 49084 78876 49140
rect 78932 49084 78942 49140
rect 90692 49028 90748 49252
rect 90804 49196 90814 49252
rect 2258 48972 2268 49028
rect 2324 48972 9324 49028
rect 9380 48972 9390 49028
rect 63634 48972 63644 49028
rect 63700 48972 65100 49028
rect 65156 48972 65166 49028
rect 71250 48972 71260 49028
rect 71316 48972 72156 49028
rect 72212 48972 72716 49028
rect 72772 48972 72782 49028
rect 85810 48972 85820 49028
rect 85876 48972 90188 49028
rect 90244 48972 90748 49028
rect 0 48916 800 48944
rect 0 48860 2380 48916
rect 2436 48860 3164 48916
rect 3220 48860 3230 48916
rect 64194 48860 64204 48916
rect 64260 48860 65324 48916
rect 65380 48860 71820 48916
rect 71876 48860 71886 48916
rect 78418 48860 78428 48916
rect 78484 48860 85036 48916
rect 85092 48860 85102 48916
rect 89618 48860 89628 48916
rect 89684 48860 90524 48916
rect 90580 48860 90590 48916
rect 0 48832 800 48860
rect 71820 48804 71876 48860
rect 12450 48748 12460 48804
rect 12516 48748 14924 48804
rect 14980 48748 14990 48804
rect 56354 48748 56364 48804
rect 56420 48748 57372 48804
rect 57428 48748 57438 48804
rect 71820 48748 72660 48804
rect 72604 48692 72660 48748
rect 1698 48636 1708 48692
rect 1764 48636 2492 48692
rect 2548 48636 2558 48692
rect 72604 48636 72940 48692
rect 72996 48636 73006 48692
rect 93090 48636 93100 48692
rect 93156 48636 96236 48692
rect 96292 48636 96302 48692
rect 8758 48580 8768 48636
rect 8824 48580 8872 48636
rect 8928 48580 8976 48636
rect 9032 48580 9080 48636
rect 9136 48580 9184 48636
rect 9240 48580 9288 48636
rect 9344 48580 9392 48636
rect 9448 48580 9458 48636
rect 17758 48580 17768 48636
rect 17824 48580 17872 48636
rect 17928 48580 17976 48636
rect 18032 48580 18080 48636
rect 18136 48580 18184 48636
rect 18240 48580 18288 48636
rect 18344 48580 18392 48636
rect 18448 48580 18458 48636
rect 26758 48580 26768 48636
rect 26824 48580 26872 48636
rect 26928 48580 26976 48636
rect 27032 48580 27080 48636
rect 27136 48580 27184 48636
rect 27240 48580 27288 48636
rect 27344 48580 27392 48636
rect 27448 48580 27458 48636
rect 35758 48580 35768 48636
rect 35824 48580 35872 48636
rect 35928 48580 35976 48636
rect 36032 48580 36080 48636
rect 36136 48580 36184 48636
rect 36240 48580 36288 48636
rect 36344 48580 36392 48636
rect 36448 48580 36458 48636
rect 44758 48580 44768 48636
rect 44824 48580 44872 48636
rect 44928 48580 44976 48636
rect 45032 48580 45080 48636
rect 45136 48580 45184 48636
rect 45240 48580 45288 48636
rect 45344 48580 45392 48636
rect 45448 48580 45458 48636
rect 53758 48580 53768 48636
rect 53824 48580 53872 48636
rect 53928 48580 53976 48636
rect 54032 48580 54080 48636
rect 54136 48580 54184 48636
rect 54240 48580 54288 48636
rect 54344 48580 54392 48636
rect 54448 48580 54458 48636
rect 62758 48580 62768 48636
rect 62824 48580 62872 48636
rect 62928 48580 62976 48636
rect 63032 48580 63080 48636
rect 63136 48580 63184 48636
rect 63240 48580 63288 48636
rect 63344 48580 63392 48636
rect 63448 48580 63458 48636
rect 71758 48580 71768 48636
rect 71824 48580 71872 48636
rect 71928 48580 71976 48636
rect 72032 48580 72080 48636
rect 72136 48580 72184 48636
rect 72240 48580 72288 48636
rect 72344 48580 72392 48636
rect 72448 48580 72458 48636
rect 80758 48580 80768 48636
rect 80824 48580 80872 48636
rect 80928 48580 80976 48636
rect 81032 48580 81080 48636
rect 81136 48580 81184 48636
rect 81240 48580 81288 48636
rect 81344 48580 81392 48636
rect 81448 48580 81458 48636
rect 89758 48580 89768 48636
rect 89824 48580 89872 48636
rect 89928 48580 89976 48636
rect 90032 48580 90080 48636
rect 90136 48580 90184 48636
rect 90240 48580 90288 48636
rect 90344 48580 90392 48636
rect 90448 48580 90458 48636
rect 39890 48412 39900 48468
rect 39956 48412 41020 48468
rect 41076 48412 41086 48468
rect 52322 48412 52332 48468
rect 52388 48412 52668 48468
rect 52724 48412 53228 48468
rect 53284 48412 54460 48468
rect 54516 48412 54526 48468
rect 63858 48412 63868 48468
rect 63924 48412 65548 48468
rect 65604 48412 74060 48468
rect 74116 48412 74620 48468
rect 74676 48412 74686 48468
rect 13570 48300 13580 48356
rect 13636 48300 15036 48356
rect 15092 48300 19852 48356
rect 19908 48300 20300 48356
rect 20356 48300 20366 48356
rect 64530 48300 64540 48356
rect 64596 48300 65100 48356
rect 65156 48300 73612 48356
rect 73668 48300 74172 48356
rect 74228 48300 76468 48356
rect 77186 48300 77196 48356
rect 77252 48300 78316 48356
rect 78372 48300 83692 48356
rect 83748 48300 83758 48356
rect 76412 48244 76468 48300
rect 14018 48188 14028 48244
rect 14084 48188 15820 48244
rect 15876 48188 15886 48244
rect 71698 48188 71708 48244
rect 71764 48188 72380 48244
rect 72436 48188 72446 48244
rect 73490 48188 73500 48244
rect 73556 48188 74396 48244
rect 74452 48188 74462 48244
rect 76402 48188 76412 48244
rect 76468 48188 77420 48244
rect 77476 48188 77486 48244
rect 79538 48188 79548 48244
rect 79604 48188 80556 48244
rect 80612 48188 80622 48244
rect 85138 48188 85148 48244
rect 85204 48188 91196 48244
rect 91252 48188 92316 48244
rect 92372 48188 92382 48244
rect 4722 48076 4732 48132
rect 4788 48076 5628 48132
rect 5684 48076 5694 48132
rect 21074 48076 21084 48132
rect 21140 48076 22092 48132
rect 22148 48076 22158 48132
rect 74610 48076 74620 48132
rect 74676 48076 75964 48132
rect 76020 48076 76972 48132
rect 77028 48076 77038 48132
rect 5282 47964 5292 48020
rect 5348 47964 9660 48020
rect 9716 47964 9726 48020
rect 15474 47964 15484 48020
rect 15540 47964 16492 48020
rect 16548 47964 16558 48020
rect 20738 47964 20748 48020
rect 20804 47964 21420 48020
rect 21476 47964 21486 48020
rect 40002 47964 40012 48020
rect 40068 47964 40460 48020
rect 40516 47964 47740 48020
rect 47796 47964 47806 48020
rect 72930 47964 72940 48020
rect 72996 47964 77420 48020
rect 77476 47964 78092 48020
rect 78148 47964 78158 48020
rect 0 47796 800 47824
rect 4258 47796 4268 47852
rect 4324 47796 4372 47852
rect 4428 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4788 47852
rect 4844 47796 4892 47852
rect 4948 47796 4958 47852
rect 13258 47796 13268 47852
rect 13324 47796 13372 47852
rect 13428 47796 13476 47852
rect 13532 47796 13580 47852
rect 13636 47796 13684 47852
rect 13740 47796 13788 47852
rect 13844 47796 13892 47852
rect 13948 47796 13958 47852
rect 22258 47796 22268 47852
rect 22324 47796 22372 47852
rect 22428 47796 22476 47852
rect 22532 47796 22580 47852
rect 22636 47796 22684 47852
rect 22740 47796 22788 47852
rect 22844 47796 22892 47852
rect 22948 47796 22958 47852
rect 31258 47796 31268 47852
rect 31324 47796 31372 47852
rect 31428 47796 31476 47852
rect 31532 47796 31580 47852
rect 31636 47796 31684 47852
rect 31740 47796 31788 47852
rect 31844 47796 31892 47852
rect 31948 47796 31958 47852
rect 40258 47796 40268 47852
rect 40324 47796 40372 47852
rect 40428 47796 40476 47852
rect 40532 47796 40580 47852
rect 40636 47796 40684 47852
rect 40740 47796 40788 47852
rect 40844 47796 40892 47852
rect 40948 47796 40958 47852
rect 49258 47796 49268 47852
rect 49324 47796 49372 47852
rect 49428 47796 49476 47852
rect 49532 47796 49580 47852
rect 49636 47796 49684 47852
rect 49740 47796 49788 47852
rect 49844 47796 49892 47852
rect 49948 47796 49958 47852
rect 58258 47796 58268 47852
rect 58324 47796 58372 47852
rect 58428 47796 58476 47852
rect 58532 47796 58580 47852
rect 58636 47796 58684 47852
rect 58740 47796 58788 47852
rect 58844 47796 58892 47852
rect 58948 47796 58958 47852
rect 67258 47796 67268 47852
rect 67324 47796 67372 47852
rect 67428 47796 67476 47852
rect 67532 47796 67580 47852
rect 67636 47796 67684 47852
rect 67740 47796 67788 47852
rect 67844 47796 67892 47852
rect 67948 47796 67958 47852
rect 76258 47796 76268 47852
rect 76324 47796 76372 47852
rect 76428 47796 76476 47852
rect 76532 47796 76580 47852
rect 76636 47796 76684 47852
rect 76740 47796 76788 47852
rect 76844 47796 76892 47852
rect 76948 47796 76958 47852
rect 85258 47796 85268 47852
rect 85324 47796 85372 47852
rect 85428 47796 85476 47852
rect 85532 47796 85580 47852
rect 85636 47796 85684 47852
rect 85740 47796 85788 47852
rect 85844 47796 85892 47852
rect 85948 47796 85958 47852
rect 94258 47796 94268 47852
rect 94324 47796 94372 47852
rect 94428 47796 94476 47852
rect 94532 47796 94580 47852
rect 94636 47796 94684 47852
rect 94740 47796 94788 47852
rect 94844 47796 94892 47852
rect 94948 47796 94958 47852
rect 99200 47796 100000 47824
rect 0 47740 1708 47796
rect 1764 47740 1774 47796
rect 98018 47740 98028 47796
rect 98084 47740 100000 47796
rect 0 47712 800 47740
rect 99200 47712 100000 47740
rect 75282 47628 75292 47684
rect 75348 47628 91644 47684
rect 91700 47628 92540 47684
rect 92596 47628 92606 47684
rect 30370 47516 30380 47572
rect 30436 47516 31612 47572
rect 31668 47516 34748 47572
rect 34804 47516 35644 47572
rect 35700 47516 35710 47572
rect 48178 47516 48188 47572
rect 48244 47516 48748 47572
rect 48804 47516 50092 47572
rect 50148 47516 64540 47572
rect 64596 47516 64606 47572
rect 8372 47404 10108 47460
rect 10164 47404 10174 47460
rect 10434 47404 10444 47460
rect 10500 47404 11844 47460
rect 20738 47404 20748 47460
rect 20804 47404 21756 47460
rect 21812 47404 21822 47460
rect 43250 47404 43260 47460
rect 43316 47404 43708 47460
rect 43764 47404 43774 47460
rect 47394 47404 47404 47460
rect 47460 47404 48860 47460
rect 48916 47404 49196 47460
rect 49252 47404 62188 47460
rect 92642 47404 92652 47460
rect 92708 47404 93436 47460
rect 93492 47404 93502 47460
rect 8372 47348 8428 47404
rect 2034 47292 2044 47348
rect 2100 47292 8428 47348
rect 10210 47292 10220 47348
rect 10276 47292 11340 47348
rect 11396 47292 11406 47348
rect 11788 47236 11844 47404
rect 17266 47292 17276 47348
rect 17332 47292 18228 47348
rect 34626 47292 34636 47348
rect 34692 47292 35308 47348
rect 35364 47292 35374 47348
rect 37650 47292 37660 47348
rect 37716 47292 39116 47348
rect 39172 47292 39182 47348
rect 46050 47292 46060 47348
rect 46116 47292 46956 47348
rect 47012 47292 47022 47348
rect 54450 47292 54460 47348
rect 54516 47292 57596 47348
rect 57652 47292 57662 47348
rect 18172 47236 18228 47292
rect 62132 47236 62188 47404
rect 77298 47292 77308 47348
rect 77364 47292 78092 47348
rect 78148 47292 78158 47348
rect 8754 47180 8764 47236
rect 8820 47180 10780 47236
rect 10836 47180 10846 47236
rect 11778 47180 11788 47236
rect 11844 47180 13132 47236
rect 13188 47180 13198 47236
rect 16482 47180 16492 47236
rect 16548 47180 17612 47236
rect 17668 47180 17678 47236
rect 18162 47180 18172 47236
rect 18228 47180 20524 47236
rect 20580 47180 21028 47236
rect 22082 47180 22092 47236
rect 22148 47180 24892 47236
rect 24948 47180 24958 47236
rect 32498 47180 32508 47236
rect 32564 47180 33628 47236
rect 33684 47180 33694 47236
rect 57026 47180 57036 47236
rect 57092 47180 58380 47236
rect 58436 47180 58446 47236
rect 62132 47180 63868 47236
rect 63924 47180 63934 47236
rect 74050 47180 74060 47236
rect 74116 47180 74956 47236
rect 75012 47180 75022 47236
rect 20972 47124 21028 47180
rect 20962 47068 20972 47124
rect 21028 47068 21532 47124
rect 21588 47068 24108 47124
rect 24164 47068 24174 47124
rect 41010 47068 41020 47124
rect 41076 47068 41804 47124
rect 41860 47068 41972 47124
rect 8758 47012 8768 47068
rect 8824 47012 8872 47068
rect 8928 47012 8976 47068
rect 9032 47012 9080 47068
rect 9136 47012 9184 47068
rect 9240 47012 9288 47068
rect 9344 47012 9392 47068
rect 9448 47012 9458 47068
rect 17758 47012 17768 47068
rect 17824 47012 17872 47068
rect 17928 47012 17976 47068
rect 18032 47012 18080 47068
rect 18136 47012 18184 47068
rect 18240 47012 18288 47068
rect 18344 47012 18392 47068
rect 18448 47012 18458 47068
rect 26758 47012 26768 47068
rect 26824 47012 26872 47068
rect 26928 47012 26976 47068
rect 27032 47012 27080 47068
rect 27136 47012 27184 47068
rect 27240 47012 27288 47068
rect 27344 47012 27392 47068
rect 27448 47012 27458 47068
rect 35758 47012 35768 47068
rect 35824 47012 35872 47068
rect 35928 47012 35976 47068
rect 36032 47012 36080 47068
rect 36136 47012 36184 47068
rect 36240 47012 36288 47068
rect 36344 47012 36392 47068
rect 36448 47012 36458 47068
rect 41916 47012 41972 47068
rect 44758 47012 44768 47068
rect 44824 47012 44872 47068
rect 44928 47012 44976 47068
rect 45032 47012 45080 47068
rect 45136 47012 45184 47068
rect 45240 47012 45288 47068
rect 45344 47012 45392 47068
rect 45448 47012 45458 47068
rect 53758 47012 53768 47068
rect 53824 47012 53872 47068
rect 53928 47012 53976 47068
rect 54032 47012 54080 47068
rect 54136 47012 54184 47068
rect 54240 47012 54288 47068
rect 54344 47012 54392 47068
rect 54448 47012 54458 47068
rect 62758 47012 62768 47068
rect 62824 47012 62872 47068
rect 62928 47012 62976 47068
rect 63032 47012 63080 47068
rect 63136 47012 63184 47068
rect 63240 47012 63288 47068
rect 63344 47012 63392 47068
rect 63448 47012 63458 47068
rect 71758 47012 71768 47068
rect 71824 47012 71872 47068
rect 71928 47012 71976 47068
rect 72032 47012 72080 47068
rect 72136 47012 72184 47068
rect 72240 47012 72288 47068
rect 72344 47012 72392 47068
rect 72448 47012 72458 47068
rect 80758 47012 80768 47068
rect 80824 47012 80872 47068
rect 80928 47012 80976 47068
rect 81032 47012 81080 47068
rect 81136 47012 81184 47068
rect 81240 47012 81288 47068
rect 81344 47012 81392 47068
rect 81448 47012 81458 47068
rect 89758 47012 89768 47068
rect 89824 47012 89872 47068
rect 89928 47012 89976 47068
rect 90032 47012 90080 47068
rect 90136 47012 90184 47068
rect 90240 47012 90288 47068
rect 90344 47012 90392 47068
rect 90448 47012 90458 47068
rect 38546 46956 38556 47012
rect 38612 46900 38668 47012
rect 41916 46956 42812 47012
rect 42868 46956 42878 47012
rect 8530 46844 8540 46900
rect 8596 46844 10332 46900
rect 10388 46844 10398 46900
rect 24882 46844 24892 46900
rect 24948 46844 38500 46900
rect 38612 46844 50428 46900
rect 51426 46844 51436 46900
rect 51492 46844 52444 46900
rect 52500 46844 52510 46900
rect 53554 46844 53564 46900
rect 53620 46844 57820 46900
rect 57876 46844 57886 46900
rect 33292 46732 38220 46788
rect 38276 46732 38286 46788
rect 0 46676 800 46704
rect 33292 46676 33348 46732
rect 38444 46676 38500 46844
rect 50372 46788 50428 46844
rect 50372 46732 64988 46788
rect 65044 46732 65436 46788
rect 65492 46732 65502 46788
rect 91970 46732 91980 46788
rect 92036 46732 92540 46788
rect 92596 46732 92606 46788
rect 0 46620 1820 46676
rect 1876 46620 1886 46676
rect 8978 46620 8988 46676
rect 9044 46620 9996 46676
rect 10052 46620 10062 46676
rect 26114 46620 26124 46676
rect 26180 46620 26908 46676
rect 26964 46620 26974 46676
rect 28924 46620 33292 46676
rect 33348 46620 33358 46676
rect 33954 46620 33964 46676
rect 34020 46620 34524 46676
rect 34580 46620 35644 46676
rect 35700 46620 35710 46676
rect 38444 46620 54124 46676
rect 54180 46620 54190 46676
rect 54562 46620 54572 46676
rect 54628 46620 55244 46676
rect 55300 46620 60172 46676
rect 60228 46620 60238 46676
rect 64866 46620 64876 46676
rect 64932 46620 65772 46676
rect 65828 46620 65838 46676
rect 73042 46620 73052 46676
rect 73108 46620 74508 46676
rect 74564 46620 74574 46676
rect 91858 46620 91868 46676
rect 91924 46620 92876 46676
rect 92932 46620 92942 46676
rect 96002 46620 96012 46676
rect 96068 46620 96908 46676
rect 96964 46620 96974 46676
rect 0 46592 800 46620
rect 28924 46564 28980 46620
rect 17602 46508 17612 46564
rect 17668 46508 28980 46564
rect 29138 46508 29148 46564
rect 29204 46508 29820 46564
rect 29876 46508 34972 46564
rect 35028 46508 35038 46564
rect 40226 46508 40236 46564
rect 40292 46508 41020 46564
rect 41076 46508 41580 46564
rect 41636 46508 41646 46564
rect 50372 46508 54236 46564
rect 54292 46508 54302 46564
rect 55346 46508 55356 46564
rect 55412 46508 57260 46564
rect 57316 46508 57326 46564
rect 58258 46508 58268 46564
rect 58324 46508 76636 46564
rect 76692 46508 76702 46564
rect 50372 46452 50428 46508
rect 27234 46396 27244 46452
rect 27300 46396 29484 46452
rect 29540 46396 29550 46452
rect 40002 46396 40012 46452
rect 40068 46396 50428 46452
rect 52210 46396 52220 46452
rect 52276 46396 52892 46452
rect 52948 46396 60060 46452
rect 60116 46396 60126 46452
rect 66770 46396 66780 46452
rect 66836 46396 85484 46452
rect 85540 46396 86380 46452
rect 86436 46396 86446 46452
rect 86930 46396 86940 46452
rect 86996 46396 89628 46452
rect 89684 46396 89694 46452
rect 4258 46228 4268 46284
rect 4324 46228 4372 46284
rect 4428 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4788 46284
rect 4844 46228 4892 46284
rect 4948 46228 4958 46284
rect 13258 46228 13268 46284
rect 13324 46228 13372 46284
rect 13428 46228 13476 46284
rect 13532 46228 13580 46284
rect 13636 46228 13684 46284
rect 13740 46228 13788 46284
rect 13844 46228 13892 46284
rect 13948 46228 13958 46284
rect 22258 46228 22268 46284
rect 22324 46228 22372 46284
rect 22428 46228 22476 46284
rect 22532 46228 22580 46284
rect 22636 46228 22684 46284
rect 22740 46228 22788 46284
rect 22844 46228 22892 46284
rect 22948 46228 22958 46284
rect 31258 46228 31268 46284
rect 31324 46228 31372 46284
rect 31428 46228 31476 46284
rect 31532 46228 31580 46284
rect 31636 46228 31684 46284
rect 31740 46228 31788 46284
rect 31844 46228 31892 46284
rect 31948 46228 31958 46284
rect 40258 46228 40268 46284
rect 40324 46228 40372 46284
rect 40428 46228 40476 46284
rect 40532 46228 40580 46284
rect 40636 46228 40684 46284
rect 40740 46228 40788 46284
rect 40844 46228 40892 46284
rect 40948 46228 40958 46284
rect 49258 46228 49268 46284
rect 49324 46228 49372 46284
rect 49428 46228 49476 46284
rect 49532 46228 49580 46284
rect 49636 46228 49684 46284
rect 49740 46228 49788 46284
rect 49844 46228 49892 46284
rect 49948 46228 49958 46284
rect 58258 46228 58268 46284
rect 58324 46228 58372 46284
rect 58428 46228 58476 46284
rect 58532 46228 58580 46284
rect 58636 46228 58684 46284
rect 58740 46228 58788 46284
rect 58844 46228 58892 46284
rect 58948 46228 58958 46284
rect 67258 46228 67268 46284
rect 67324 46228 67372 46284
rect 67428 46228 67476 46284
rect 67532 46228 67580 46284
rect 67636 46228 67684 46284
rect 67740 46228 67788 46284
rect 67844 46228 67892 46284
rect 67948 46228 67958 46284
rect 76258 46228 76268 46284
rect 76324 46228 76372 46284
rect 76428 46228 76476 46284
rect 76532 46228 76580 46284
rect 76636 46228 76684 46284
rect 76740 46228 76788 46284
rect 76844 46228 76892 46284
rect 76948 46228 76958 46284
rect 85258 46228 85268 46284
rect 85324 46228 85372 46284
rect 85428 46228 85476 46284
rect 85532 46228 85580 46284
rect 85636 46228 85684 46284
rect 85740 46228 85788 46284
rect 85844 46228 85892 46284
rect 85948 46228 85958 46284
rect 94258 46228 94268 46284
rect 94324 46228 94372 46284
rect 94428 46228 94476 46284
rect 94532 46228 94580 46284
rect 94636 46228 94684 46284
rect 94740 46228 94788 46284
rect 94844 46228 94892 46284
rect 94948 46228 94958 46284
rect 54898 46172 54908 46228
rect 54964 46172 55244 46228
rect 55300 46172 55310 46228
rect 31490 46060 31500 46116
rect 31556 46060 32172 46116
rect 32228 46060 32238 46116
rect 36754 46060 36764 46116
rect 36820 46060 39004 46116
rect 39060 46060 39070 46116
rect 50372 46060 55580 46116
rect 55636 46060 56588 46116
rect 56644 46060 56654 46116
rect 50372 46004 50428 46060
rect 99200 46004 100000 46032
rect 13234 45948 13244 46004
rect 13300 45948 50428 46004
rect 79090 45948 79100 46004
rect 79156 45948 79548 46004
rect 79604 45948 82796 46004
rect 82852 45948 82862 46004
rect 98018 45948 98028 46004
rect 98084 45948 100000 46004
rect 99200 45920 100000 45948
rect 39340 45836 40684 45892
rect 40740 45836 41916 45892
rect 41972 45836 41982 45892
rect 47394 45836 47404 45892
rect 47460 45836 49196 45892
rect 49252 45836 49262 45892
rect 54114 45836 54124 45892
rect 54180 45836 55020 45892
rect 55076 45836 55086 45892
rect 64642 45836 64652 45892
rect 64708 45836 65324 45892
rect 65380 45836 65390 45892
rect 72930 45836 72940 45892
rect 72996 45836 75852 45892
rect 75908 45836 77084 45892
rect 77140 45836 77308 45892
rect 77364 45836 77374 45892
rect 79874 45836 79884 45892
rect 79940 45836 80556 45892
rect 80612 45836 80622 45892
rect 39340 45780 39396 45836
rect 28578 45724 28588 45780
rect 28644 45724 29260 45780
rect 29316 45724 30604 45780
rect 30660 45724 33740 45780
rect 33796 45724 33806 45780
rect 35074 45724 35084 45780
rect 35140 45724 38556 45780
rect 38612 45724 39340 45780
rect 39396 45724 39406 45780
rect 40226 45724 40236 45780
rect 40292 45724 41020 45780
rect 41076 45724 41086 45780
rect 56802 45724 56812 45780
rect 56868 45724 58044 45780
rect 58100 45724 58110 45780
rect 62132 45724 73388 45780
rect 73444 45724 73454 45780
rect 78642 45724 78652 45780
rect 78708 45724 79324 45780
rect 79380 45724 79390 45780
rect 89618 45724 89628 45780
rect 89684 45724 96124 45780
rect 96180 45724 96190 45780
rect 62132 45668 62188 45724
rect 38434 45612 38444 45668
rect 38500 45612 39900 45668
rect 39956 45612 39966 45668
rect 43036 45612 47516 45668
rect 47572 45612 47582 45668
rect 54450 45612 54460 45668
rect 54516 45612 55020 45668
rect 55076 45612 56028 45668
rect 56084 45612 56700 45668
rect 56756 45612 56766 45668
rect 56914 45612 56924 45668
rect 56980 45612 62188 45668
rect 62626 45612 62636 45668
rect 62692 45612 64092 45668
rect 64148 45612 64652 45668
rect 64708 45612 64718 45668
rect 70466 45612 70476 45668
rect 70532 45612 71932 45668
rect 71988 45612 73052 45668
rect 73108 45612 73118 45668
rect 77410 45612 77420 45668
rect 77476 45612 78316 45668
rect 78372 45612 83580 45668
rect 83636 45612 83646 45668
rect 89058 45612 89068 45668
rect 89124 45612 89964 45668
rect 90020 45612 91364 45668
rect 92530 45612 92540 45668
rect 92596 45612 95676 45668
rect 95732 45612 96236 45668
rect 96292 45612 96302 45668
rect 0 45556 800 45584
rect 0 45500 1708 45556
rect 1764 45500 2492 45556
rect 2548 45500 2558 45556
rect 0 45472 800 45500
rect 8758 45444 8768 45500
rect 8824 45444 8872 45500
rect 8928 45444 8976 45500
rect 9032 45444 9080 45500
rect 9136 45444 9184 45500
rect 9240 45444 9288 45500
rect 9344 45444 9392 45500
rect 9448 45444 9458 45500
rect 17758 45444 17768 45500
rect 17824 45444 17872 45500
rect 17928 45444 17976 45500
rect 18032 45444 18080 45500
rect 18136 45444 18184 45500
rect 18240 45444 18288 45500
rect 18344 45444 18392 45500
rect 18448 45444 18458 45500
rect 26758 45444 26768 45500
rect 26824 45444 26872 45500
rect 26928 45444 26976 45500
rect 27032 45444 27080 45500
rect 27136 45444 27184 45500
rect 27240 45444 27288 45500
rect 27344 45444 27392 45500
rect 27448 45444 27458 45500
rect 35758 45444 35768 45500
rect 35824 45444 35872 45500
rect 35928 45444 35976 45500
rect 36032 45444 36080 45500
rect 36136 45444 36184 45500
rect 36240 45444 36288 45500
rect 36344 45444 36392 45500
rect 36448 45444 36458 45500
rect 43036 45444 43092 45612
rect 91308 45556 91364 45612
rect 91298 45500 91308 45556
rect 91364 45500 95004 45556
rect 95060 45500 95070 45556
rect 44758 45444 44768 45500
rect 44824 45444 44872 45500
rect 44928 45444 44976 45500
rect 45032 45444 45080 45500
rect 45136 45444 45184 45500
rect 45240 45444 45288 45500
rect 45344 45444 45392 45500
rect 45448 45444 45458 45500
rect 53758 45444 53768 45500
rect 53824 45444 53872 45500
rect 53928 45444 53976 45500
rect 54032 45444 54080 45500
rect 54136 45444 54184 45500
rect 54240 45444 54288 45500
rect 54344 45444 54392 45500
rect 54448 45444 54458 45500
rect 62758 45444 62768 45500
rect 62824 45444 62872 45500
rect 62928 45444 62976 45500
rect 63032 45444 63080 45500
rect 63136 45444 63184 45500
rect 63240 45444 63288 45500
rect 63344 45444 63392 45500
rect 63448 45444 63458 45500
rect 71758 45444 71768 45500
rect 71824 45444 71872 45500
rect 71928 45444 71976 45500
rect 72032 45444 72080 45500
rect 72136 45444 72184 45500
rect 72240 45444 72288 45500
rect 72344 45444 72392 45500
rect 72448 45444 72458 45500
rect 80758 45444 80768 45500
rect 80824 45444 80872 45500
rect 80928 45444 80976 45500
rect 81032 45444 81080 45500
rect 81136 45444 81184 45500
rect 81240 45444 81288 45500
rect 81344 45444 81392 45500
rect 81448 45444 81458 45500
rect 89758 45444 89768 45500
rect 89824 45444 89872 45500
rect 89928 45444 89976 45500
rect 90032 45444 90080 45500
rect 90136 45444 90184 45500
rect 90240 45444 90288 45500
rect 90344 45444 90392 45500
rect 90448 45444 90458 45500
rect 38546 45388 38556 45444
rect 38612 45388 43092 45444
rect 52434 45388 52444 45444
rect 52500 45388 53452 45444
rect 53508 45388 53518 45444
rect 63522 45388 63532 45444
rect 63588 45388 64540 45444
rect 64596 45388 67788 45444
rect 67844 45388 71372 45444
rect 71428 45388 71438 45444
rect 41906 45276 41916 45332
rect 41972 45276 44492 45332
rect 44548 45276 45276 45332
rect 45332 45276 45342 45332
rect 50306 45276 50316 45332
rect 50372 45276 91196 45332
rect 91252 45276 91980 45332
rect 92036 45276 92046 45332
rect 5954 45164 5964 45220
rect 6020 45164 15484 45220
rect 15540 45164 15550 45220
rect 17378 45164 17388 45220
rect 17444 45164 19628 45220
rect 19684 45164 23436 45220
rect 23492 45164 23502 45220
rect 43586 45164 43596 45220
rect 43652 45164 43820 45220
rect 43876 45164 43886 45220
rect 61282 45164 61292 45220
rect 61348 45164 62076 45220
rect 62132 45164 63308 45220
rect 63364 45164 63374 45220
rect 76738 45164 76748 45220
rect 76804 45164 77756 45220
rect 77812 45164 77822 45220
rect 86706 45164 86716 45220
rect 86772 45164 90636 45220
rect 90692 45164 91084 45220
rect 91140 45164 91756 45220
rect 91812 45164 91822 45220
rect 2706 45052 2716 45108
rect 2772 45052 3388 45108
rect 3444 45052 3454 45108
rect 14914 45052 14924 45108
rect 14980 45052 16492 45108
rect 16548 45052 16558 45108
rect 41346 45052 41356 45108
rect 41412 45052 47516 45108
rect 47572 45052 47582 45108
rect 68898 45052 68908 45108
rect 68964 45052 70140 45108
rect 70196 45052 70206 45108
rect 71250 45052 71260 45108
rect 71316 45052 76356 45108
rect 71260 44996 71316 45052
rect 76300 44996 76356 45052
rect 1698 44940 1708 44996
rect 1764 44940 2492 44996
rect 2548 44940 2558 44996
rect 42130 44940 42140 44996
rect 42196 44940 42700 44996
rect 42756 44940 42766 44996
rect 61730 44940 61740 44996
rect 61796 44940 62076 44996
rect 62132 44940 63532 44996
rect 63588 44940 69468 44996
rect 69524 44940 71316 44996
rect 73602 44940 73612 44996
rect 73668 44940 74508 44996
rect 74564 44940 74574 44996
rect 76290 44940 76300 44996
rect 76356 44940 77532 44996
rect 77588 44940 77598 44996
rect 16146 44828 16156 44884
rect 16212 44828 17612 44884
rect 17668 44828 17678 44884
rect 53554 44828 53564 44884
rect 53620 44828 54908 44884
rect 54964 44828 58492 44884
rect 58548 44828 58558 44884
rect 4258 44660 4268 44716
rect 4324 44660 4372 44716
rect 4428 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4788 44716
rect 4844 44660 4892 44716
rect 4948 44660 4958 44716
rect 13258 44660 13268 44716
rect 13324 44660 13372 44716
rect 13428 44660 13476 44716
rect 13532 44660 13580 44716
rect 13636 44660 13684 44716
rect 13740 44660 13788 44716
rect 13844 44660 13892 44716
rect 13948 44660 13958 44716
rect 22258 44660 22268 44716
rect 22324 44660 22372 44716
rect 22428 44660 22476 44716
rect 22532 44660 22580 44716
rect 22636 44660 22684 44716
rect 22740 44660 22788 44716
rect 22844 44660 22892 44716
rect 22948 44660 22958 44716
rect 31258 44660 31268 44716
rect 31324 44660 31372 44716
rect 31428 44660 31476 44716
rect 31532 44660 31580 44716
rect 31636 44660 31684 44716
rect 31740 44660 31788 44716
rect 31844 44660 31892 44716
rect 31948 44660 31958 44716
rect 40258 44660 40268 44716
rect 40324 44660 40372 44716
rect 40428 44660 40476 44716
rect 40532 44660 40580 44716
rect 40636 44660 40684 44716
rect 40740 44660 40788 44716
rect 40844 44660 40892 44716
rect 40948 44660 40958 44716
rect 49258 44660 49268 44716
rect 49324 44660 49372 44716
rect 49428 44660 49476 44716
rect 49532 44660 49580 44716
rect 49636 44660 49684 44716
rect 49740 44660 49788 44716
rect 49844 44660 49892 44716
rect 49948 44660 49958 44716
rect 58258 44660 58268 44716
rect 58324 44660 58372 44716
rect 58428 44660 58476 44716
rect 58532 44660 58580 44716
rect 58636 44660 58684 44716
rect 58740 44660 58788 44716
rect 58844 44660 58892 44716
rect 58948 44660 58958 44716
rect 67258 44660 67268 44716
rect 67324 44660 67372 44716
rect 67428 44660 67476 44716
rect 67532 44660 67580 44716
rect 67636 44660 67684 44716
rect 67740 44660 67788 44716
rect 67844 44660 67892 44716
rect 67948 44660 67958 44716
rect 76258 44660 76268 44716
rect 76324 44660 76372 44716
rect 76428 44660 76476 44716
rect 76532 44660 76580 44716
rect 76636 44660 76684 44716
rect 76740 44660 76788 44716
rect 76844 44660 76892 44716
rect 76948 44660 76958 44716
rect 85258 44660 85268 44716
rect 85324 44660 85372 44716
rect 85428 44660 85476 44716
rect 85532 44660 85580 44716
rect 85636 44660 85684 44716
rect 85740 44660 85788 44716
rect 85844 44660 85892 44716
rect 85948 44660 85958 44716
rect 94258 44660 94268 44716
rect 94324 44660 94372 44716
rect 94428 44660 94476 44716
rect 94532 44660 94580 44716
rect 94636 44660 94684 44716
rect 94740 44660 94788 44716
rect 94844 44660 94892 44716
rect 94948 44660 94958 44716
rect 6514 44492 6524 44548
rect 6580 44492 21420 44548
rect 21476 44492 21486 44548
rect 63074 44492 63084 44548
rect 63140 44492 64428 44548
rect 64484 44492 64494 44548
rect 0 44436 800 44464
rect 0 44380 1708 44436
rect 1764 44380 1774 44436
rect 20066 44380 20076 44436
rect 20132 44380 22540 44436
rect 22596 44380 22606 44436
rect 30594 44380 30604 44436
rect 30660 44380 31052 44436
rect 31108 44380 35084 44436
rect 35140 44380 35980 44436
rect 36036 44380 36046 44436
rect 0 44352 800 44380
rect 9762 44268 9772 44324
rect 9828 44268 11564 44324
rect 11620 44268 13132 44324
rect 13188 44268 13198 44324
rect 46050 44268 46060 44324
rect 46116 44268 47180 44324
rect 47236 44268 48076 44324
rect 48132 44268 48142 44324
rect 54114 44268 54124 44324
rect 54180 44268 54796 44324
rect 54852 44268 55468 44324
rect 55524 44268 55534 44324
rect 55682 44268 55692 44324
rect 55748 44268 57484 44324
rect 57540 44268 58492 44324
rect 58548 44268 69692 44324
rect 69748 44268 71260 44324
rect 71316 44268 71326 44324
rect 73602 44268 73612 44324
rect 73668 44268 74620 44324
rect 74676 44268 75068 44324
rect 75124 44268 75404 44324
rect 75460 44268 75470 44324
rect 99200 44212 100000 44240
rect 7186 44156 7196 44212
rect 7252 44156 14028 44212
rect 14084 44156 17388 44212
rect 17444 44156 17454 44212
rect 34850 44156 34860 44212
rect 34916 44156 35532 44212
rect 35588 44156 35598 44212
rect 40898 44156 40908 44212
rect 40964 44156 41804 44212
rect 41860 44156 42364 44212
rect 42420 44156 43260 44212
rect 43316 44156 43326 44212
rect 47730 44156 47740 44212
rect 47796 44156 48636 44212
rect 48692 44156 48972 44212
rect 49028 44156 49038 44212
rect 51986 44156 51996 44212
rect 52052 44156 54572 44212
rect 54628 44156 54638 44212
rect 55906 44156 55916 44212
rect 55972 44156 56924 44212
rect 56980 44156 57260 44212
rect 57316 44156 57326 44212
rect 65202 44156 65212 44212
rect 65268 44156 65884 44212
rect 65940 44156 65950 44212
rect 78306 44156 78316 44212
rect 78372 44156 79772 44212
rect 79828 44156 79838 44212
rect 98018 44156 98028 44212
rect 98084 44156 100000 44212
rect 99200 44128 100000 44156
rect 8978 44044 8988 44100
rect 9044 44044 9772 44100
rect 9828 44044 9838 44100
rect 17938 44044 17948 44100
rect 18004 44044 19796 44100
rect 22194 44044 22204 44100
rect 22260 44044 23100 44100
rect 23156 44044 24220 44100
rect 24276 44044 33796 44100
rect 49858 44044 49868 44100
rect 49924 44044 52892 44100
rect 52948 44044 52958 44100
rect 56690 44044 56700 44100
rect 56756 44044 57932 44100
rect 57988 44044 57998 44100
rect 63522 44044 63532 44100
rect 63588 44044 64652 44100
rect 64708 44044 64718 44100
rect 73042 44044 73052 44100
rect 73108 44044 73118 44100
rect 73266 44044 73276 44100
rect 73332 44044 76636 44100
rect 76692 44044 77308 44100
rect 77364 44044 77374 44100
rect 8758 43876 8768 43932
rect 8824 43876 8872 43932
rect 8928 43876 8976 43932
rect 9032 43876 9080 43932
rect 9136 43876 9184 43932
rect 9240 43876 9288 43932
rect 9344 43876 9392 43932
rect 9448 43876 9458 43932
rect 17758 43876 17768 43932
rect 17824 43876 17872 43932
rect 17928 43876 17976 43932
rect 18032 43876 18080 43932
rect 18136 43876 18184 43932
rect 18240 43876 18288 43932
rect 18344 43876 18392 43932
rect 18448 43876 18458 43932
rect 19740 43764 19796 44044
rect 26758 43876 26768 43932
rect 26824 43876 26872 43932
rect 26928 43876 26976 43932
rect 27032 43876 27080 43932
rect 27136 43876 27184 43932
rect 27240 43876 27288 43932
rect 27344 43876 27392 43932
rect 27448 43876 27458 43932
rect 33740 43876 33796 44044
rect 73052 43988 73108 44044
rect 73052 43932 73948 43988
rect 74004 43932 74956 43988
rect 75012 43932 75022 43988
rect 35758 43876 35768 43932
rect 35824 43876 35872 43932
rect 35928 43876 35976 43932
rect 36032 43876 36080 43932
rect 36136 43876 36184 43932
rect 36240 43876 36288 43932
rect 36344 43876 36392 43932
rect 36448 43876 36458 43932
rect 44758 43876 44768 43932
rect 44824 43876 44872 43932
rect 44928 43876 44976 43932
rect 45032 43876 45080 43932
rect 45136 43876 45184 43932
rect 45240 43876 45288 43932
rect 45344 43876 45392 43932
rect 45448 43876 45458 43932
rect 53758 43876 53768 43932
rect 53824 43876 53872 43932
rect 53928 43876 53976 43932
rect 54032 43876 54080 43932
rect 54136 43876 54184 43932
rect 54240 43876 54288 43932
rect 54344 43876 54392 43932
rect 54448 43876 54458 43932
rect 62758 43876 62768 43932
rect 62824 43876 62872 43932
rect 62928 43876 62976 43932
rect 63032 43876 63080 43932
rect 63136 43876 63184 43932
rect 63240 43876 63288 43932
rect 63344 43876 63392 43932
rect 63448 43876 63458 43932
rect 71758 43876 71768 43932
rect 71824 43876 71872 43932
rect 71928 43876 71976 43932
rect 72032 43876 72080 43932
rect 72136 43876 72184 43932
rect 72240 43876 72288 43932
rect 72344 43876 72392 43932
rect 72448 43876 72458 43932
rect 80758 43876 80768 43932
rect 80824 43876 80872 43932
rect 80928 43876 80976 43932
rect 81032 43876 81080 43932
rect 81136 43876 81184 43932
rect 81240 43876 81288 43932
rect 81344 43876 81392 43932
rect 81448 43876 81458 43932
rect 89758 43876 89768 43932
rect 89824 43876 89872 43932
rect 89928 43876 89976 43932
rect 90032 43876 90080 43932
rect 90136 43876 90184 43932
rect 90240 43876 90288 43932
rect 90344 43876 90392 43932
rect 90448 43876 90458 43932
rect 33730 43820 33740 43876
rect 33796 43820 33806 43876
rect 8306 43708 8316 43764
rect 8372 43708 9436 43764
rect 9492 43708 9502 43764
rect 19740 43708 31948 43764
rect 32004 43708 32014 43764
rect 56802 43708 56812 43764
rect 56868 43708 57708 43764
rect 57764 43708 60172 43764
rect 60228 43708 60238 43764
rect 63410 43708 63420 43764
rect 63476 43708 64092 43764
rect 64148 43708 64158 43764
rect 80098 43708 80108 43764
rect 80164 43708 81340 43764
rect 81396 43708 81406 43764
rect 88386 43708 88396 43764
rect 88452 43708 90860 43764
rect 90916 43708 92316 43764
rect 92372 43708 92382 43764
rect 5730 43596 5740 43652
rect 5796 43596 6300 43652
rect 6356 43596 12348 43652
rect 12404 43596 12414 43652
rect 20738 43596 20748 43652
rect 20804 43596 21756 43652
rect 21812 43596 21822 43652
rect 32050 43596 32060 43652
rect 32116 43596 33068 43652
rect 33124 43596 33134 43652
rect 43250 43596 43260 43652
rect 43316 43596 45836 43652
rect 45892 43596 46396 43652
rect 46452 43596 47628 43652
rect 47684 43596 47694 43652
rect 52770 43596 52780 43652
rect 52836 43596 53228 43652
rect 53284 43596 53900 43652
rect 53956 43596 56028 43652
rect 56084 43596 57820 43652
rect 57876 43596 59388 43652
rect 59444 43596 60956 43652
rect 61012 43596 61022 43652
rect 71698 43596 71708 43652
rect 71764 43596 72492 43652
rect 72548 43596 73164 43652
rect 73220 43596 73230 43652
rect 76962 43596 76972 43652
rect 77028 43596 77420 43652
rect 77476 43596 84476 43652
rect 84532 43596 84542 43652
rect 29250 43484 29260 43540
rect 29316 43484 29932 43540
rect 29988 43484 35196 43540
rect 35252 43484 35262 43540
rect 65426 43484 65436 43540
rect 65492 43484 67004 43540
rect 67060 43484 67070 43540
rect 70690 43484 70700 43540
rect 70756 43484 72380 43540
rect 72436 43484 72446 43540
rect 31938 43372 31948 43428
rect 32004 43372 32508 43428
rect 32564 43372 38444 43428
rect 38500 43372 38510 43428
rect 64530 43372 64540 43428
rect 64596 43372 65548 43428
rect 65604 43372 66332 43428
rect 66388 43372 66398 43428
rect 71250 43372 71260 43428
rect 71316 43372 72716 43428
rect 72772 43372 72782 43428
rect 90962 43372 90972 43428
rect 91028 43372 94556 43428
rect 94612 43372 94622 43428
rect 0 43316 800 43344
rect 0 43260 1820 43316
rect 1876 43260 1886 43316
rect 5954 43260 5964 43316
rect 6020 43260 8428 43316
rect 27234 43260 27244 43316
rect 27300 43260 29596 43316
rect 29652 43260 29662 43316
rect 31714 43260 31724 43316
rect 31780 43260 32116 43316
rect 75282 43260 75292 43316
rect 75348 43260 77196 43316
rect 77252 43260 77262 43316
rect 0 43232 800 43260
rect 4258 43092 4268 43148
rect 4324 43092 4372 43148
rect 4428 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4788 43148
rect 4844 43092 4892 43148
rect 4948 43092 4958 43148
rect 8372 42980 8428 43260
rect 13258 43092 13268 43148
rect 13324 43092 13372 43148
rect 13428 43092 13476 43148
rect 13532 43092 13580 43148
rect 13636 43092 13684 43148
rect 13740 43092 13788 43148
rect 13844 43092 13892 43148
rect 13948 43092 13958 43148
rect 22258 43092 22268 43148
rect 22324 43092 22372 43148
rect 22428 43092 22476 43148
rect 22532 43092 22580 43148
rect 22636 43092 22684 43148
rect 22740 43092 22788 43148
rect 22844 43092 22892 43148
rect 22948 43092 22958 43148
rect 31258 43092 31268 43148
rect 31324 43092 31372 43148
rect 31428 43092 31476 43148
rect 31532 43092 31580 43148
rect 31636 43092 31684 43148
rect 31740 43092 31788 43148
rect 31844 43092 31892 43148
rect 31948 43092 31958 43148
rect 32060 42980 32116 43260
rect 40258 43092 40268 43148
rect 40324 43092 40372 43148
rect 40428 43092 40476 43148
rect 40532 43092 40580 43148
rect 40636 43092 40684 43148
rect 40740 43092 40788 43148
rect 40844 43092 40892 43148
rect 40948 43092 40958 43148
rect 49258 43092 49268 43148
rect 49324 43092 49372 43148
rect 49428 43092 49476 43148
rect 49532 43092 49580 43148
rect 49636 43092 49684 43148
rect 49740 43092 49788 43148
rect 49844 43092 49892 43148
rect 49948 43092 49958 43148
rect 58258 43092 58268 43148
rect 58324 43092 58372 43148
rect 58428 43092 58476 43148
rect 58532 43092 58580 43148
rect 58636 43092 58684 43148
rect 58740 43092 58788 43148
rect 58844 43092 58892 43148
rect 58948 43092 58958 43148
rect 67258 43092 67268 43148
rect 67324 43092 67372 43148
rect 67428 43092 67476 43148
rect 67532 43092 67580 43148
rect 67636 43092 67684 43148
rect 67740 43092 67788 43148
rect 67844 43092 67892 43148
rect 67948 43092 67958 43148
rect 76258 43092 76268 43148
rect 76324 43092 76372 43148
rect 76428 43092 76476 43148
rect 76532 43092 76580 43148
rect 76636 43092 76684 43148
rect 76740 43092 76788 43148
rect 76844 43092 76892 43148
rect 76948 43092 76958 43148
rect 85258 43092 85268 43148
rect 85324 43092 85372 43148
rect 85428 43092 85476 43148
rect 85532 43092 85580 43148
rect 85636 43092 85684 43148
rect 85740 43092 85788 43148
rect 85844 43092 85892 43148
rect 85948 43092 85958 43148
rect 94258 43092 94268 43148
rect 94324 43092 94372 43148
rect 94428 43092 94476 43148
rect 94532 43092 94580 43148
rect 94636 43092 94684 43148
rect 94740 43092 94788 43148
rect 94844 43092 94892 43148
rect 94948 43092 94958 43148
rect 8372 42924 13580 42980
rect 13636 42924 13646 42980
rect 31602 42924 31612 42980
rect 31668 42924 32116 42980
rect 34178 42924 34188 42980
rect 34244 42924 35084 42980
rect 35140 42924 35868 42980
rect 35924 42924 35934 42980
rect 92754 42924 92764 42980
rect 92820 42924 95340 42980
rect 95396 42924 95406 42980
rect 13234 42812 13244 42868
rect 13300 42812 14028 42868
rect 14084 42812 14094 42868
rect 19516 42812 20748 42868
rect 20804 42812 20814 42868
rect 28242 42812 28252 42868
rect 28308 42812 28588 42868
rect 28644 42812 29372 42868
rect 29428 42812 30828 42868
rect 30884 42812 31164 42868
rect 31220 42812 31230 42868
rect 60946 42812 60956 42868
rect 61012 42812 61852 42868
rect 61908 42812 62188 42868
rect 64978 42812 64988 42868
rect 65044 42812 65660 42868
rect 65716 42812 66668 42868
rect 66724 42812 66734 42868
rect 90692 42812 96236 42868
rect 96292 42812 96302 42868
rect 19516 42756 19572 42812
rect 12236 42700 13804 42756
rect 13860 42700 15148 42756
rect 15204 42700 18956 42756
rect 19012 42700 19516 42756
rect 19572 42700 19582 42756
rect 20178 42700 20188 42756
rect 20244 42700 21868 42756
rect 21924 42700 21934 42756
rect 12236 42532 12292 42700
rect 12674 42588 12684 42644
rect 12740 42588 14700 42644
rect 14756 42588 14766 42644
rect 15586 42588 15596 42644
rect 15652 42588 19404 42644
rect 19460 42588 19470 42644
rect 26226 42588 26236 42644
rect 26292 42588 26908 42644
rect 26964 42588 26974 42644
rect 62132 42532 62188 42812
rect 66434 42700 66444 42756
rect 66500 42700 67900 42756
rect 67956 42700 73948 42756
rect 73892 42532 73948 42700
rect 90692 42532 90748 42812
rect 10322 42476 10332 42532
rect 10388 42476 12236 42532
rect 12292 42476 12302 42532
rect 12898 42476 12908 42532
rect 12964 42476 13804 42532
rect 13860 42476 13870 42532
rect 14354 42476 14364 42532
rect 14420 42476 15260 42532
rect 15316 42476 16940 42532
rect 16996 42476 17006 42532
rect 62132 42476 64988 42532
rect 65044 42476 69356 42532
rect 69412 42476 72492 42532
rect 72548 42476 72558 42532
rect 73892 42476 74508 42532
rect 74564 42476 75404 42532
rect 75460 42476 77084 42532
rect 77140 42476 77150 42532
rect 88834 42476 88844 42532
rect 88900 42476 90076 42532
rect 90132 42476 90748 42532
rect 92306 42476 92316 42532
rect 92372 42476 93100 42532
rect 93156 42476 93166 42532
rect 99200 42420 100000 42448
rect 98018 42364 98028 42420
rect 98084 42364 100000 42420
rect 8758 42308 8768 42364
rect 8824 42308 8872 42364
rect 8928 42308 8976 42364
rect 9032 42308 9080 42364
rect 9136 42308 9184 42364
rect 9240 42308 9288 42364
rect 9344 42308 9392 42364
rect 9448 42308 9458 42364
rect 17758 42308 17768 42364
rect 17824 42308 17872 42364
rect 17928 42308 17976 42364
rect 18032 42308 18080 42364
rect 18136 42308 18184 42364
rect 18240 42308 18288 42364
rect 18344 42308 18392 42364
rect 18448 42308 18458 42364
rect 26758 42308 26768 42364
rect 26824 42308 26872 42364
rect 26928 42308 26976 42364
rect 27032 42308 27080 42364
rect 27136 42308 27184 42364
rect 27240 42308 27288 42364
rect 27344 42308 27392 42364
rect 27448 42308 27458 42364
rect 35758 42308 35768 42364
rect 35824 42308 35872 42364
rect 35928 42308 35976 42364
rect 36032 42308 36080 42364
rect 36136 42308 36184 42364
rect 36240 42308 36288 42364
rect 36344 42308 36392 42364
rect 36448 42308 36458 42364
rect 44758 42308 44768 42364
rect 44824 42308 44872 42364
rect 44928 42308 44976 42364
rect 45032 42308 45080 42364
rect 45136 42308 45184 42364
rect 45240 42308 45288 42364
rect 45344 42308 45392 42364
rect 45448 42308 45458 42364
rect 53758 42308 53768 42364
rect 53824 42308 53872 42364
rect 53928 42308 53976 42364
rect 54032 42308 54080 42364
rect 54136 42308 54184 42364
rect 54240 42308 54288 42364
rect 54344 42308 54392 42364
rect 54448 42308 54458 42364
rect 62758 42308 62768 42364
rect 62824 42308 62872 42364
rect 62928 42308 62976 42364
rect 63032 42308 63080 42364
rect 63136 42308 63184 42364
rect 63240 42308 63288 42364
rect 63344 42308 63392 42364
rect 63448 42308 63458 42364
rect 71758 42308 71768 42364
rect 71824 42308 71872 42364
rect 71928 42308 71976 42364
rect 72032 42308 72080 42364
rect 72136 42308 72184 42364
rect 72240 42308 72288 42364
rect 72344 42308 72392 42364
rect 72448 42308 72458 42364
rect 80758 42308 80768 42364
rect 80824 42308 80872 42364
rect 80928 42308 80976 42364
rect 81032 42308 81080 42364
rect 81136 42308 81184 42364
rect 81240 42308 81288 42364
rect 81344 42308 81392 42364
rect 81448 42308 81458 42364
rect 89758 42308 89768 42364
rect 89824 42308 89872 42364
rect 89928 42308 89976 42364
rect 90032 42308 90080 42364
rect 90136 42308 90184 42364
rect 90240 42308 90288 42364
rect 90344 42308 90392 42364
rect 90448 42308 90458 42364
rect 99200 42336 100000 42364
rect 0 42196 800 42224
rect 0 42140 1708 42196
rect 1764 42140 2492 42196
rect 2548 42140 2558 42196
rect 6178 42140 6188 42196
rect 6244 42140 6748 42196
rect 6804 42140 6814 42196
rect 66994 42140 67004 42196
rect 67060 42140 74620 42196
rect 74676 42140 74686 42196
rect 0 42112 800 42140
rect 21858 42028 21868 42084
rect 21924 42028 24444 42084
rect 24500 42028 38780 42084
rect 38836 42028 38846 42084
rect 49074 42028 49084 42084
rect 49140 42028 49644 42084
rect 49700 42028 49710 42084
rect 77970 42028 77980 42084
rect 78036 42028 79100 42084
rect 79156 42028 79166 42084
rect 16370 41916 16380 41972
rect 16436 41916 17500 41972
rect 17556 41916 19740 41972
rect 19796 41916 21532 41972
rect 21588 41916 21980 41972
rect 22036 41916 23548 41972
rect 23604 41916 23614 41972
rect 39554 41916 39564 41972
rect 39620 41916 41020 41972
rect 41076 41916 41086 41972
rect 42354 41916 42364 41972
rect 42420 41916 44492 41972
rect 44548 41916 44558 41972
rect 55122 41916 55132 41972
rect 55188 41916 55580 41972
rect 55636 41916 55646 41972
rect 56914 41916 56924 41972
rect 56980 41916 56990 41972
rect 66994 41916 67004 41972
rect 67060 41916 67788 41972
rect 67844 41916 67854 41972
rect 75730 41916 75740 41972
rect 75796 41916 76860 41972
rect 76916 41916 78204 41972
rect 78260 41916 78270 41972
rect 80546 41916 80556 41972
rect 80612 41916 80892 41972
rect 80948 41916 81676 41972
rect 81732 41916 83468 41972
rect 83524 41916 83534 41972
rect 87154 41916 87164 41972
rect 87220 41916 89180 41972
rect 89236 41916 89246 41972
rect 56924 41860 56980 41916
rect 51090 41804 51100 41860
rect 51156 41804 53788 41860
rect 53844 41804 53854 41860
rect 54898 41804 54908 41860
rect 54964 41804 56028 41860
rect 56084 41804 57484 41860
rect 57540 41804 57550 41860
rect 72258 41804 72268 41860
rect 72324 41804 73500 41860
rect 73556 41804 76412 41860
rect 76468 41804 77868 41860
rect 77924 41804 77934 41860
rect 53788 41748 53844 41804
rect 6290 41692 6300 41748
rect 6356 41692 17612 41748
rect 17668 41692 17678 41748
rect 53788 41692 55020 41748
rect 55076 41692 56140 41748
rect 56196 41692 56206 41748
rect 55458 41580 55468 41636
rect 55524 41580 57596 41636
rect 57652 41580 57662 41636
rect 4258 41524 4268 41580
rect 4324 41524 4372 41580
rect 4428 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4788 41580
rect 4844 41524 4892 41580
rect 4948 41524 4958 41580
rect 13258 41524 13268 41580
rect 13324 41524 13372 41580
rect 13428 41524 13476 41580
rect 13532 41524 13580 41580
rect 13636 41524 13684 41580
rect 13740 41524 13788 41580
rect 13844 41524 13892 41580
rect 13948 41524 13958 41580
rect 22258 41524 22268 41580
rect 22324 41524 22372 41580
rect 22428 41524 22476 41580
rect 22532 41524 22580 41580
rect 22636 41524 22684 41580
rect 22740 41524 22788 41580
rect 22844 41524 22892 41580
rect 22948 41524 22958 41580
rect 31258 41524 31268 41580
rect 31324 41524 31372 41580
rect 31428 41524 31476 41580
rect 31532 41524 31580 41580
rect 31636 41524 31684 41580
rect 31740 41524 31788 41580
rect 31844 41524 31892 41580
rect 31948 41524 31958 41580
rect 40258 41524 40268 41580
rect 40324 41524 40372 41580
rect 40428 41524 40476 41580
rect 40532 41524 40580 41580
rect 40636 41524 40684 41580
rect 40740 41524 40788 41580
rect 40844 41524 40892 41580
rect 40948 41524 40958 41580
rect 49258 41524 49268 41580
rect 49324 41524 49372 41580
rect 49428 41524 49476 41580
rect 49532 41524 49580 41580
rect 49636 41524 49684 41580
rect 49740 41524 49788 41580
rect 49844 41524 49892 41580
rect 49948 41524 49958 41580
rect 58258 41524 58268 41580
rect 58324 41524 58372 41580
rect 58428 41524 58476 41580
rect 58532 41524 58580 41580
rect 58636 41524 58684 41580
rect 58740 41524 58788 41580
rect 58844 41524 58892 41580
rect 58948 41524 58958 41580
rect 67258 41524 67268 41580
rect 67324 41524 67372 41580
rect 67428 41524 67476 41580
rect 67532 41524 67580 41580
rect 67636 41524 67684 41580
rect 67740 41524 67788 41580
rect 67844 41524 67892 41580
rect 67948 41524 67958 41580
rect 76258 41524 76268 41580
rect 76324 41524 76372 41580
rect 76428 41524 76476 41580
rect 76532 41524 76580 41580
rect 76636 41524 76684 41580
rect 76740 41524 76788 41580
rect 76844 41524 76892 41580
rect 76948 41524 76958 41580
rect 85258 41524 85268 41580
rect 85324 41524 85372 41580
rect 85428 41524 85476 41580
rect 85532 41524 85580 41580
rect 85636 41524 85684 41580
rect 85740 41524 85788 41580
rect 85844 41524 85892 41580
rect 85948 41524 85958 41580
rect 94258 41524 94268 41580
rect 94324 41524 94372 41580
rect 94428 41524 94476 41580
rect 94532 41524 94580 41580
rect 94636 41524 94684 41580
rect 94740 41524 94788 41580
rect 94844 41524 94892 41580
rect 94948 41524 94958 41580
rect 2034 41356 2044 41412
rect 2100 41356 5964 41412
rect 6020 41356 6030 41412
rect 13122 41356 13132 41412
rect 13188 41356 53340 41412
rect 53396 41356 58716 41412
rect 58772 41356 58782 41412
rect 59266 41356 59276 41412
rect 59332 41356 73948 41412
rect 76738 41356 76748 41412
rect 76804 41356 78652 41412
rect 78708 41356 81564 41412
rect 81620 41356 81630 41412
rect 41458 41244 41468 41300
rect 41524 41244 42140 41300
rect 42196 41244 42364 41300
rect 42420 41244 42430 41300
rect 57586 41244 57596 41300
rect 57652 41244 72268 41300
rect 72324 41244 72334 41300
rect 35298 41132 35308 41188
rect 35364 41132 35868 41188
rect 35924 41132 35934 41188
rect 44258 41132 44268 41188
rect 44324 41132 45276 41188
rect 45332 41132 45342 41188
rect 57026 41132 57036 41188
rect 57092 41132 61740 41188
rect 61796 41132 61806 41188
rect 64642 41132 64652 41188
rect 64708 41132 65212 41188
rect 65268 41132 65278 41188
rect 0 41076 800 41104
rect 0 41020 2380 41076
rect 2436 41020 2446 41076
rect 18498 41020 18508 41076
rect 18564 41020 19068 41076
rect 19124 41020 22652 41076
rect 22708 41020 37100 41076
rect 37156 41020 37166 41076
rect 42018 41020 42028 41076
rect 42084 41020 49532 41076
rect 49588 41020 49598 41076
rect 50978 41020 50988 41076
rect 51044 41020 53564 41076
rect 53620 41020 53630 41076
rect 54674 41020 54684 41076
rect 54740 41020 55356 41076
rect 55412 41020 57820 41076
rect 57876 41020 57886 41076
rect 60498 41020 60508 41076
rect 60564 41020 61964 41076
rect 62020 41020 71372 41076
rect 71428 41020 71438 41076
rect 0 40992 800 41020
rect 8372 40908 9324 40964
rect 9380 40908 9660 40964
rect 9716 40908 12348 40964
rect 12404 40908 12414 40964
rect 33394 40908 33404 40964
rect 33460 40908 34188 40964
rect 34244 40908 34254 40964
rect 34962 40908 34972 40964
rect 35028 40908 39900 40964
rect 39956 40908 39966 40964
rect 62066 40908 62076 40964
rect 62132 40908 65996 40964
rect 66052 40908 67116 40964
rect 67172 40908 67182 40964
rect 4722 40572 4732 40628
rect 4788 40572 5852 40628
rect 5908 40572 6636 40628
rect 6692 40572 8316 40628
rect 8372 40572 8428 40908
rect 73892 40852 73948 41356
rect 76178 41132 76188 41188
rect 76244 41132 76580 41188
rect 76524 41076 76580 41132
rect 74162 41020 74172 41076
rect 74228 41020 74732 41076
rect 74788 41020 76300 41076
rect 76356 41020 76366 41076
rect 76524 41020 76860 41076
rect 76916 41020 76926 41076
rect 75618 40908 75628 40964
rect 75684 40908 76412 40964
rect 76468 40908 76478 40964
rect 77634 40908 77644 40964
rect 77700 40908 78540 40964
rect 78596 40908 80892 40964
rect 80948 40908 80958 40964
rect 30370 40796 30380 40852
rect 30436 40796 31612 40852
rect 31668 40796 32172 40852
rect 32228 40796 33292 40852
rect 33348 40796 35196 40852
rect 35252 40796 35262 40852
rect 73892 40796 76300 40852
rect 76356 40796 76366 40852
rect 8758 40740 8768 40796
rect 8824 40740 8872 40796
rect 8928 40740 8976 40796
rect 9032 40740 9080 40796
rect 9136 40740 9184 40796
rect 9240 40740 9288 40796
rect 9344 40740 9392 40796
rect 9448 40740 9458 40796
rect 17758 40740 17768 40796
rect 17824 40740 17872 40796
rect 17928 40740 17976 40796
rect 18032 40740 18080 40796
rect 18136 40740 18184 40796
rect 18240 40740 18288 40796
rect 18344 40740 18392 40796
rect 18448 40740 18458 40796
rect 26758 40740 26768 40796
rect 26824 40740 26872 40796
rect 26928 40740 26976 40796
rect 27032 40740 27080 40796
rect 27136 40740 27184 40796
rect 27240 40740 27288 40796
rect 27344 40740 27392 40796
rect 27448 40740 27458 40796
rect 35758 40740 35768 40796
rect 35824 40740 35872 40796
rect 35928 40740 35976 40796
rect 36032 40740 36080 40796
rect 36136 40740 36184 40796
rect 36240 40740 36288 40796
rect 36344 40740 36392 40796
rect 36448 40740 36458 40796
rect 44758 40740 44768 40796
rect 44824 40740 44872 40796
rect 44928 40740 44976 40796
rect 45032 40740 45080 40796
rect 45136 40740 45184 40796
rect 45240 40740 45288 40796
rect 45344 40740 45392 40796
rect 45448 40740 45458 40796
rect 53758 40740 53768 40796
rect 53824 40740 53872 40796
rect 53928 40740 53976 40796
rect 54032 40740 54080 40796
rect 54136 40740 54184 40796
rect 54240 40740 54288 40796
rect 54344 40740 54392 40796
rect 54448 40740 54458 40796
rect 62758 40740 62768 40796
rect 62824 40740 62872 40796
rect 62928 40740 62976 40796
rect 63032 40740 63080 40796
rect 63136 40740 63184 40796
rect 63240 40740 63288 40796
rect 63344 40740 63392 40796
rect 63448 40740 63458 40796
rect 71758 40740 71768 40796
rect 71824 40740 71872 40796
rect 71928 40740 71976 40796
rect 72032 40740 72080 40796
rect 72136 40740 72184 40796
rect 72240 40740 72288 40796
rect 72344 40740 72392 40796
rect 72448 40740 72458 40796
rect 80758 40740 80768 40796
rect 80824 40740 80872 40796
rect 80928 40740 80976 40796
rect 81032 40740 81080 40796
rect 81136 40740 81184 40796
rect 81240 40740 81288 40796
rect 81344 40740 81392 40796
rect 81448 40740 81458 40796
rect 89758 40740 89768 40796
rect 89824 40740 89872 40796
rect 89928 40740 89976 40796
rect 90032 40740 90080 40796
rect 90136 40740 90184 40796
rect 90240 40740 90288 40796
rect 90344 40740 90392 40796
rect 90448 40740 90458 40796
rect 84130 40684 84140 40740
rect 84196 40684 85708 40740
rect 85652 40628 85708 40684
rect 99200 40628 100000 40656
rect 21074 40572 21084 40628
rect 21140 40572 21980 40628
rect 22036 40572 22988 40628
rect 23044 40572 23054 40628
rect 33730 40572 33740 40628
rect 33796 40572 38556 40628
rect 38612 40572 38622 40628
rect 38994 40572 39004 40628
rect 39060 40572 68124 40628
rect 68180 40572 68190 40628
rect 71586 40572 71596 40628
rect 71652 40572 72268 40628
rect 72324 40572 72334 40628
rect 85362 40572 85372 40628
rect 85428 40572 85438 40628
rect 85652 40572 85932 40628
rect 85988 40572 96236 40628
rect 96292 40572 96302 40628
rect 98018 40572 98028 40628
rect 98084 40572 100000 40628
rect 85372 40516 85428 40572
rect 99200 40544 100000 40572
rect 30146 40460 30156 40516
rect 30212 40460 30604 40516
rect 30660 40460 30940 40516
rect 30996 40460 31006 40516
rect 34850 40460 34860 40516
rect 34916 40460 36092 40516
rect 36148 40460 36158 40516
rect 41570 40460 41580 40516
rect 41636 40460 42700 40516
rect 42756 40460 42766 40516
rect 45938 40460 45948 40516
rect 46004 40460 48412 40516
rect 48468 40460 48478 40516
rect 53218 40460 53228 40516
rect 53284 40460 54796 40516
rect 54852 40460 54862 40516
rect 66098 40460 66108 40516
rect 66164 40460 67452 40516
rect 67508 40460 67518 40516
rect 85372 40460 86268 40516
rect 86324 40460 86828 40516
rect 86884 40460 86894 40516
rect 89506 40460 89516 40516
rect 89572 40460 90748 40516
rect 90804 40460 94780 40516
rect 94836 40460 94846 40516
rect 16930 40348 16940 40404
rect 16996 40348 17500 40404
rect 17556 40348 17566 40404
rect 28914 40348 28924 40404
rect 28980 40348 29596 40404
rect 29652 40348 35420 40404
rect 35476 40348 35486 40404
rect 49074 40348 49084 40404
rect 49140 40348 49420 40404
rect 49476 40348 49486 40404
rect 50082 40348 50092 40404
rect 50148 40348 50652 40404
rect 50708 40348 50718 40404
rect 53106 40348 53116 40404
rect 53172 40348 54012 40404
rect 54068 40348 55692 40404
rect 55748 40348 55758 40404
rect 57698 40348 57708 40404
rect 57764 40348 58604 40404
rect 58660 40348 58670 40404
rect 65538 40348 65548 40404
rect 65604 40348 66556 40404
rect 66612 40348 66622 40404
rect 71698 40348 71708 40404
rect 71764 40348 73948 40404
rect 74004 40348 74014 40404
rect 76962 40348 76972 40404
rect 77028 40348 77756 40404
rect 77812 40348 77822 40404
rect 91644 40348 95340 40404
rect 95396 40348 96124 40404
rect 96180 40348 96190 40404
rect 28242 40236 28252 40292
rect 28308 40236 29036 40292
rect 29092 40236 29102 40292
rect 40338 40236 40348 40292
rect 40404 40236 41244 40292
rect 41300 40236 41310 40292
rect 54562 40236 54572 40292
rect 54628 40236 55356 40292
rect 55412 40236 55422 40292
rect 74162 40236 74172 40292
rect 74228 40236 75068 40292
rect 75124 40236 75134 40292
rect 78082 40236 78092 40292
rect 78148 40236 87500 40292
rect 87556 40236 87566 40292
rect 91644 40180 91700 40348
rect 12460 40124 13580 40180
rect 13636 40124 16828 40180
rect 16884 40124 16894 40180
rect 26786 40124 26796 40180
rect 26852 40124 29260 40180
rect 29316 40124 29326 40180
rect 66882 40124 66892 40180
rect 66948 40124 67676 40180
rect 67732 40124 67742 40180
rect 69682 40124 69692 40180
rect 69748 40124 91084 40180
rect 91140 40124 91150 40180
rect 91634 40124 91644 40180
rect 91700 40124 91710 40180
rect 0 39956 800 39984
rect 4258 39956 4268 40012
rect 4324 39956 4372 40012
rect 4428 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4788 40012
rect 4844 39956 4892 40012
rect 4948 39956 4958 40012
rect 12460 39956 12516 40124
rect 13258 39956 13268 40012
rect 13324 39956 13372 40012
rect 13428 39956 13476 40012
rect 13532 39956 13580 40012
rect 13636 39956 13684 40012
rect 13740 39956 13788 40012
rect 13844 39956 13892 40012
rect 13948 39956 13958 40012
rect 22258 39956 22268 40012
rect 22324 39956 22372 40012
rect 22428 39956 22476 40012
rect 22532 39956 22580 40012
rect 22636 39956 22684 40012
rect 22740 39956 22788 40012
rect 22844 39956 22892 40012
rect 22948 39956 22958 40012
rect 31258 39956 31268 40012
rect 31324 39956 31372 40012
rect 31428 39956 31476 40012
rect 31532 39956 31580 40012
rect 31636 39956 31684 40012
rect 31740 39956 31788 40012
rect 31844 39956 31892 40012
rect 31948 39956 31958 40012
rect 40258 39956 40268 40012
rect 40324 39956 40372 40012
rect 40428 39956 40476 40012
rect 40532 39956 40580 40012
rect 40636 39956 40684 40012
rect 40740 39956 40788 40012
rect 40844 39956 40892 40012
rect 40948 39956 40958 40012
rect 49258 39956 49268 40012
rect 49324 39956 49372 40012
rect 49428 39956 49476 40012
rect 49532 39956 49580 40012
rect 49636 39956 49684 40012
rect 49740 39956 49788 40012
rect 49844 39956 49892 40012
rect 49948 39956 49958 40012
rect 58258 39956 58268 40012
rect 58324 39956 58372 40012
rect 58428 39956 58476 40012
rect 58532 39956 58580 40012
rect 58636 39956 58684 40012
rect 58740 39956 58788 40012
rect 58844 39956 58892 40012
rect 58948 39956 58958 40012
rect 67258 39956 67268 40012
rect 67324 39956 67372 40012
rect 67428 39956 67476 40012
rect 67532 39956 67580 40012
rect 67636 39956 67684 40012
rect 67740 39956 67788 40012
rect 67844 39956 67892 40012
rect 67948 39956 67958 40012
rect 76258 39956 76268 40012
rect 76324 39956 76372 40012
rect 76428 39956 76476 40012
rect 76532 39956 76580 40012
rect 76636 39956 76684 40012
rect 76740 39956 76788 40012
rect 76844 39956 76892 40012
rect 76948 39956 76958 40012
rect 85258 39956 85268 40012
rect 85324 39956 85372 40012
rect 85428 39956 85476 40012
rect 85532 39956 85580 40012
rect 85636 39956 85684 40012
rect 85740 39956 85788 40012
rect 85844 39956 85892 40012
rect 85948 39956 85958 40012
rect 94258 39956 94268 40012
rect 94324 39956 94372 40012
rect 94428 39956 94476 40012
rect 94532 39956 94580 40012
rect 94636 39956 94684 40012
rect 94740 39956 94788 40012
rect 94844 39956 94892 40012
rect 94948 39956 94958 40012
rect 0 39900 1708 39956
rect 1764 39900 3164 39956
rect 3220 39900 3230 39956
rect 12450 39900 12460 39956
rect 12516 39900 12526 39956
rect 0 39872 800 39900
rect 31826 39788 31836 39844
rect 31892 39788 33068 39844
rect 33124 39788 33134 39844
rect 64642 39788 64652 39844
rect 64708 39788 65324 39844
rect 65380 39788 68348 39844
rect 68404 39788 69020 39844
rect 69076 39788 75964 39844
rect 76020 39788 77756 39844
rect 77812 39788 77822 39844
rect 36540 39676 82124 39732
rect 82180 39676 82190 39732
rect 36540 39620 36596 39676
rect 9090 39564 9100 39620
rect 9156 39564 15484 39620
rect 15540 39564 15550 39620
rect 36530 39564 36540 39620
rect 36596 39564 36606 39620
rect 37314 39564 37324 39620
rect 37380 39564 73948 39620
rect 83010 39564 83020 39620
rect 83076 39564 83916 39620
rect 83972 39564 83982 39620
rect 84914 39564 84924 39620
rect 84980 39564 87164 39620
rect 87220 39564 87230 39620
rect 73892 39508 73948 39564
rect 12786 39452 12796 39508
rect 12852 39452 13468 39508
rect 13524 39452 13534 39508
rect 36194 39452 36204 39508
rect 36260 39452 36988 39508
rect 37044 39452 37054 39508
rect 66882 39452 66892 39508
rect 66948 39452 68460 39508
rect 68516 39452 68526 39508
rect 73892 39452 84364 39508
rect 84420 39452 84812 39508
rect 84868 39452 84878 39508
rect 2034 39340 2044 39396
rect 2100 39340 11788 39396
rect 11844 39340 11854 39396
rect 13346 39340 13356 39396
rect 13412 39340 14140 39396
rect 14196 39340 14206 39396
rect 35858 39340 35868 39396
rect 35924 39340 36316 39396
rect 36372 39340 36382 39396
rect 42578 39340 42588 39396
rect 42644 39340 52220 39396
rect 52276 39340 52556 39396
rect 52612 39340 52622 39396
rect 85810 39340 85820 39396
rect 85876 39340 90300 39396
rect 90356 39340 96236 39396
rect 96292 39340 96302 39396
rect 8758 39172 8768 39228
rect 8824 39172 8872 39228
rect 8928 39172 8976 39228
rect 9032 39172 9080 39228
rect 9136 39172 9184 39228
rect 9240 39172 9288 39228
rect 9344 39172 9392 39228
rect 9448 39172 9458 39228
rect 17758 39172 17768 39228
rect 17824 39172 17872 39228
rect 17928 39172 17976 39228
rect 18032 39172 18080 39228
rect 18136 39172 18184 39228
rect 18240 39172 18288 39228
rect 18344 39172 18392 39228
rect 18448 39172 18458 39228
rect 26758 39172 26768 39228
rect 26824 39172 26872 39228
rect 26928 39172 26976 39228
rect 27032 39172 27080 39228
rect 27136 39172 27184 39228
rect 27240 39172 27288 39228
rect 27344 39172 27392 39228
rect 27448 39172 27458 39228
rect 35758 39172 35768 39228
rect 35824 39172 35872 39228
rect 35928 39172 35976 39228
rect 36032 39172 36080 39228
rect 36136 39172 36184 39228
rect 36240 39172 36288 39228
rect 36344 39172 36392 39228
rect 36448 39172 36458 39228
rect 44758 39172 44768 39228
rect 44824 39172 44872 39228
rect 44928 39172 44976 39228
rect 45032 39172 45080 39228
rect 45136 39172 45184 39228
rect 45240 39172 45288 39228
rect 45344 39172 45392 39228
rect 45448 39172 45458 39228
rect 53758 39172 53768 39228
rect 53824 39172 53872 39228
rect 53928 39172 53976 39228
rect 54032 39172 54080 39228
rect 54136 39172 54184 39228
rect 54240 39172 54288 39228
rect 54344 39172 54392 39228
rect 54448 39172 54458 39228
rect 62758 39172 62768 39228
rect 62824 39172 62872 39228
rect 62928 39172 62976 39228
rect 63032 39172 63080 39228
rect 63136 39172 63184 39228
rect 63240 39172 63288 39228
rect 63344 39172 63392 39228
rect 63448 39172 63458 39228
rect 71758 39172 71768 39228
rect 71824 39172 71872 39228
rect 71928 39172 71976 39228
rect 72032 39172 72080 39228
rect 72136 39172 72184 39228
rect 72240 39172 72288 39228
rect 72344 39172 72392 39228
rect 72448 39172 72458 39228
rect 80758 39172 80768 39228
rect 80824 39172 80872 39228
rect 80928 39172 80976 39228
rect 81032 39172 81080 39228
rect 81136 39172 81184 39228
rect 81240 39172 81288 39228
rect 81344 39172 81392 39228
rect 81448 39172 81458 39228
rect 89758 39172 89768 39228
rect 89824 39172 89872 39228
rect 89928 39172 89976 39228
rect 90032 39172 90080 39228
rect 90136 39172 90184 39228
rect 90240 39172 90288 39228
rect 90344 39172 90392 39228
rect 90448 39172 90458 39228
rect 16258 39004 16268 39060
rect 16324 39004 17500 39060
rect 17556 39004 17566 39060
rect 35186 39004 35196 39060
rect 35252 39004 50428 39060
rect 50530 39004 50540 39060
rect 50596 39004 52892 39060
rect 52948 39004 52958 39060
rect 60946 39004 60956 39060
rect 61012 39004 65548 39060
rect 65604 39004 65614 39060
rect 66658 39004 66668 39060
rect 66724 39004 67788 39060
rect 67844 39004 75404 39060
rect 75460 39004 75470 39060
rect 77186 39004 77196 39060
rect 77252 39004 77262 39060
rect 77746 39004 77756 39060
rect 77812 39004 78540 39060
rect 78596 39004 78606 39060
rect 82674 39004 82684 39060
rect 82740 39004 83468 39060
rect 83524 39004 84476 39060
rect 84532 39004 85260 39060
rect 85316 39004 85326 39060
rect 89730 39004 89740 39060
rect 89796 39004 90860 39060
rect 90916 39004 91364 39060
rect 43586 38892 43596 38948
rect 43652 38892 43820 38948
rect 43876 38892 43886 38948
rect 47730 38892 47740 38948
rect 47796 38892 49084 38948
rect 49140 38892 49150 38948
rect 0 38836 800 38864
rect 50372 38836 50428 39004
rect 66668 38948 66724 39004
rect 77196 38948 77252 39004
rect 91308 38948 91364 39004
rect 52658 38892 52668 38948
rect 52724 38892 53900 38948
rect 53956 38892 53966 38948
rect 58034 38892 58044 38948
rect 58100 38892 66724 38948
rect 66994 38892 67004 38948
rect 67060 38892 68012 38948
rect 68068 38892 68078 38948
rect 77196 38892 77420 38948
rect 77476 38892 77486 38948
rect 83906 38892 83916 38948
rect 83972 38892 84700 38948
rect 84756 38892 84766 38948
rect 89058 38892 89068 38948
rect 89124 38892 90188 38948
rect 90244 38892 90972 38948
rect 91028 38892 91038 38948
rect 91298 38892 91308 38948
rect 91364 38892 91374 38948
rect 99200 38836 100000 38864
rect 0 38780 1820 38836
rect 1876 38780 1886 38836
rect 50372 38780 60172 38836
rect 60228 38780 60956 38836
rect 61012 38780 61022 38836
rect 64530 38780 64540 38836
rect 64596 38780 67228 38836
rect 67284 38780 69020 38836
rect 69076 38780 69086 38836
rect 74834 38780 74844 38836
rect 74900 38780 79604 38836
rect 98018 38780 98028 38836
rect 98084 38780 100000 38836
rect 0 38752 800 38780
rect 76860 38724 76916 38780
rect 79548 38724 79604 38780
rect 99200 38752 100000 38780
rect 16818 38668 16828 38724
rect 16884 38668 35644 38724
rect 35700 38668 35710 38724
rect 76850 38668 76860 38724
rect 76916 38668 76926 38724
rect 77186 38668 77196 38724
rect 77252 38668 77868 38724
rect 77924 38668 77934 38724
rect 79538 38668 79548 38724
rect 79604 38668 80500 38724
rect 80444 38612 80500 38668
rect 41234 38556 41244 38612
rect 41300 38556 44492 38612
rect 44548 38556 45276 38612
rect 45332 38556 45342 38612
rect 55794 38556 55804 38612
rect 55860 38556 56700 38612
rect 56756 38556 57820 38612
rect 57876 38556 57886 38612
rect 80444 38556 87164 38612
rect 87220 38556 87230 38612
rect 4258 38388 4268 38444
rect 4324 38388 4372 38444
rect 4428 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4788 38444
rect 4844 38388 4892 38444
rect 4948 38388 4958 38444
rect 13258 38388 13268 38444
rect 13324 38388 13372 38444
rect 13428 38388 13476 38444
rect 13532 38388 13580 38444
rect 13636 38388 13684 38444
rect 13740 38388 13788 38444
rect 13844 38388 13892 38444
rect 13948 38388 13958 38444
rect 22258 38388 22268 38444
rect 22324 38388 22372 38444
rect 22428 38388 22476 38444
rect 22532 38388 22580 38444
rect 22636 38388 22684 38444
rect 22740 38388 22788 38444
rect 22844 38388 22892 38444
rect 22948 38388 22958 38444
rect 31258 38388 31268 38444
rect 31324 38388 31372 38444
rect 31428 38388 31476 38444
rect 31532 38388 31580 38444
rect 31636 38388 31684 38444
rect 31740 38388 31788 38444
rect 31844 38388 31892 38444
rect 31948 38388 31958 38444
rect 40258 38388 40268 38444
rect 40324 38388 40372 38444
rect 40428 38388 40476 38444
rect 40532 38388 40580 38444
rect 40636 38388 40684 38444
rect 40740 38388 40788 38444
rect 40844 38388 40892 38444
rect 40948 38388 40958 38444
rect 49258 38388 49268 38444
rect 49324 38388 49372 38444
rect 49428 38388 49476 38444
rect 49532 38388 49580 38444
rect 49636 38388 49684 38444
rect 49740 38388 49788 38444
rect 49844 38388 49892 38444
rect 49948 38388 49958 38444
rect 58258 38388 58268 38444
rect 58324 38388 58372 38444
rect 58428 38388 58476 38444
rect 58532 38388 58580 38444
rect 58636 38388 58684 38444
rect 58740 38388 58788 38444
rect 58844 38388 58892 38444
rect 58948 38388 58958 38444
rect 67258 38388 67268 38444
rect 67324 38388 67372 38444
rect 67428 38388 67476 38444
rect 67532 38388 67580 38444
rect 67636 38388 67684 38444
rect 67740 38388 67788 38444
rect 67844 38388 67892 38444
rect 67948 38388 67958 38444
rect 76258 38388 76268 38444
rect 76324 38388 76372 38444
rect 76428 38388 76476 38444
rect 76532 38388 76580 38444
rect 76636 38388 76684 38444
rect 76740 38388 76788 38444
rect 76844 38388 76892 38444
rect 76948 38388 76958 38444
rect 85258 38388 85268 38444
rect 85324 38388 85372 38444
rect 85428 38388 85476 38444
rect 85532 38388 85580 38444
rect 85636 38388 85684 38444
rect 85740 38388 85788 38444
rect 85844 38388 85892 38444
rect 85948 38388 85958 38444
rect 94258 38388 94268 38444
rect 94324 38388 94372 38444
rect 94428 38388 94476 38444
rect 94532 38388 94580 38444
rect 94636 38388 94684 38444
rect 94740 38388 94788 38444
rect 94844 38388 94892 38444
rect 94948 38388 94958 38444
rect 63858 38332 63868 38388
rect 63924 38332 64428 38388
rect 64484 38332 66108 38388
rect 66164 38332 66174 38388
rect 17266 38220 17276 38276
rect 17332 38220 33404 38276
rect 33460 38220 38332 38276
rect 38388 38220 38398 38276
rect 41346 38220 41356 38276
rect 41412 38220 42028 38276
rect 42084 38220 48076 38276
rect 48132 38220 48142 38276
rect 50194 38220 50204 38276
rect 50260 38220 67788 38276
rect 67844 38220 68572 38276
rect 68628 38220 68638 38276
rect 75394 38220 75404 38276
rect 75460 38220 77196 38276
rect 77252 38220 77262 38276
rect 29922 38108 29932 38164
rect 29988 38108 42364 38164
rect 42420 38108 42430 38164
rect 51538 38108 51548 38164
rect 51604 38108 89068 38164
rect 89124 38108 89134 38164
rect 20738 37996 20748 38052
rect 20804 37996 21868 38052
rect 21924 37996 21934 38052
rect 28354 37996 28364 38052
rect 28420 37996 30156 38052
rect 30212 37996 30222 38052
rect 38434 37996 38444 38052
rect 38500 37996 48188 38052
rect 48244 37996 48254 38052
rect 48402 37996 48412 38052
rect 48468 37996 49756 38052
rect 49812 37996 49822 38052
rect 52546 37996 52556 38052
rect 52612 37996 67228 38052
rect 67284 37996 67294 38052
rect 68562 37996 68572 38052
rect 68628 37996 75628 38052
rect 75684 37996 75694 38052
rect 78530 37996 78540 38052
rect 78596 37996 79324 38052
rect 79380 37996 79390 38052
rect 87490 37996 87500 38052
rect 87556 37996 90972 38052
rect 91028 37996 91038 38052
rect 28466 37884 28476 37940
rect 28532 37884 32956 37940
rect 33012 37884 34860 37940
rect 34916 37884 34926 37940
rect 59266 37884 59276 37940
rect 59332 37884 60620 37940
rect 60676 37884 60686 37940
rect 61730 37884 61740 37940
rect 61796 37884 68348 37940
rect 68404 37884 68414 37940
rect 68572 37884 72380 37940
rect 72436 37884 73948 37940
rect 74004 37884 74014 37940
rect 74274 37884 74284 37940
rect 74340 37884 76300 37940
rect 76356 37884 76366 37940
rect 84130 37884 84140 37940
rect 84196 37884 84980 37940
rect 5282 37772 5292 37828
rect 5348 37772 20188 37828
rect 20244 37772 20254 37828
rect 24994 37772 25004 37828
rect 25060 37772 37100 37828
rect 37156 37772 37166 37828
rect 41458 37772 41468 37828
rect 41524 37772 41916 37828
rect 41972 37772 43372 37828
rect 43428 37772 43438 37828
rect 46050 37772 46060 37828
rect 46116 37772 47180 37828
rect 47236 37772 48748 37828
rect 48804 37772 48814 37828
rect 54562 37772 54572 37828
rect 54628 37772 56364 37828
rect 56420 37772 56430 37828
rect 59938 37772 59948 37828
rect 60004 37772 60508 37828
rect 60564 37772 61180 37828
rect 61236 37772 61246 37828
rect 66434 37772 66444 37828
rect 66500 37772 67116 37828
rect 67172 37772 67676 37828
rect 67732 37772 67742 37828
rect 0 37716 800 37744
rect 68572 37716 68628 37884
rect 84924 37828 84980 37884
rect 71922 37772 71932 37828
rect 71988 37772 72604 37828
rect 72660 37772 72670 37828
rect 74946 37772 74956 37828
rect 75012 37772 76188 37828
rect 76244 37772 76254 37828
rect 77522 37772 77532 37828
rect 77588 37772 78316 37828
rect 78372 37772 82460 37828
rect 82516 37772 82526 37828
rect 83458 37772 83468 37828
rect 83524 37772 84252 37828
rect 84308 37772 84318 37828
rect 84914 37772 84924 37828
rect 84980 37772 85484 37828
rect 85540 37772 85932 37828
rect 85988 37772 85998 37828
rect 0 37660 1708 37716
rect 1764 37660 2492 37716
rect 2548 37660 2558 37716
rect 20514 37660 20524 37716
rect 20580 37660 21644 37716
rect 21700 37660 21710 37716
rect 66098 37660 66108 37716
rect 66164 37660 68628 37716
rect 0 37632 800 37660
rect 8758 37604 8768 37660
rect 8824 37604 8872 37660
rect 8928 37604 8976 37660
rect 9032 37604 9080 37660
rect 9136 37604 9184 37660
rect 9240 37604 9288 37660
rect 9344 37604 9392 37660
rect 9448 37604 9458 37660
rect 17758 37604 17768 37660
rect 17824 37604 17872 37660
rect 17928 37604 17976 37660
rect 18032 37604 18080 37660
rect 18136 37604 18184 37660
rect 18240 37604 18288 37660
rect 18344 37604 18392 37660
rect 18448 37604 18458 37660
rect 26758 37604 26768 37660
rect 26824 37604 26872 37660
rect 26928 37604 26976 37660
rect 27032 37604 27080 37660
rect 27136 37604 27184 37660
rect 27240 37604 27288 37660
rect 27344 37604 27392 37660
rect 27448 37604 27458 37660
rect 35758 37604 35768 37660
rect 35824 37604 35872 37660
rect 35928 37604 35976 37660
rect 36032 37604 36080 37660
rect 36136 37604 36184 37660
rect 36240 37604 36288 37660
rect 36344 37604 36392 37660
rect 36448 37604 36458 37660
rect 44758 37604 44768 37660
rect 44824 37604 44872 37660
rect 44928 37604 44976 37660
rect 45032 37604 45080 37660
rect 45136 37604 45184 37660
rect 45240 37604 45288 37660
rect 45344 37604 45392 37660
rect 45448 37604 45458 37660
rect 53758 37604 53768 37660
rect 53824 37604 53872 37660
rect 53928 37604 53976 37660
rect 54032 37604 54080 37660
rect 54136 37604 54184 37660
rect 54240 37604 54288 37660
rect 54344 37604 54392 37660
rect 54448 37604 54458 37660
rect 62758 37604 62768 37660
rect 62824 37604 62872 37660
rect 62928 37604 62976 37660
rect 63032 37604 63080 37660
rect 63136 37604 63184 37660
rect 63240 37604 63288 37660
rect 63344 37604 63392 37660
rect 63448 37604 63458 37660
rect 71758 37604 71768 37660
rect 71824 37604 71872 37660
rect 71928 37604 71976 37660
rect 72032 37604 72080 37660
rect 72136 37604 72184 37660
rect 72240 37604 72288 37660
rect 72344 37604 72392 37660
rect 72448 37604 72458 37660
rect 80758 37604 80768 37660
rect 80824 37604 80872 37660
rect 80928 37604 80976 37660
rect 81032 37604 81080 37660
rect 81136 37604 81184 37660
rect 81240 37604 81288 37660
rect 81344 37604 81392 37660
rect 81448 37604 81458 37660
rect 89758 37604 89768 37660
rect 89824 37604 89872 37660
rect 89928 37604 89976 37660
rect 90032 37604 90080 37660
rect 90136 37604 90184 37660
rect 90240 37604 90288 37660
rect 90344 37604 90392 37660
rect 90448 37604 90458 37660
rect 36540 37548 40460 37604
rect 40516 37548 41244 37604
rect 41300 37548 41916 37604
rect 41972 37548 41982 37604
rect 57922 37548 57932 37604
rect 57988 37548 60956 37604
rect 61012 37548 61022 37604
rect 68198 37548 68236 37604
rect 68292 37548 68908 37604
rect 68964 37548 68974 37604
rect 36540 37492 36596 37548
rect 7298 37436 7308 37492
rect 7364 37436 18396 37492
rect 18452 37436 19740 37492
rect 19796 37436 19806 37492
rect 34850 37436 34860 37492
rect 34916 37436 36596 37492
rect 37314 37436 37324 37492
rect 37380 37436 73948 37492
rect 76850 37436 76860 37492
rect 76916 37436 77532 37492
rect 77588 37436 77598 37492
rect 86818 37436 86828 37492
rect 86884 37436 88060 37492
rect 88116 37436 89516 37492
rect 89572 37436 89582 37492
rect 73892 37380 73948 37436
rect 5842 37324 5852 37380
rect 5908 37324 8428 37380
rect 8642 37324 8652 37380
rect 8708 37324 9660 37380
rect 9716 37324 9726 37380
rect 10546 37324 10556 37380
rect 10612 37324 10622 37380
rect 29138 37324 29148 37380
rect 29204 37324 29820 37380
rect 29876 37324 29886 37380
rect 37986 37324 37996 37380
rect 38052 37324 39228 37380
rect 39284 37324 39294 37380
rect 41682 37324 41692 37380
rect 41748 37324 43204 37380
rect 43362 37324 43372 37380
rect 43428 37324 46396 37380
rect 46452 37324 46462 37380
rect 53218 37324 53228 37380
rect 53284 37324 54572 37380
rect 54628 37324 54638 37380
rect 73892 37324 83468 37380
rect 83524 37324 83534 37380
rect 8372 37268 8428 37324
rect 10556 37268 10612 37324
rect 43148 37268 43204 37324
rect 8372 37212 10612 37268
rect 21298 37212 21308 37268
rect 21364 37212 25004 37268
rect 25060 37212 25070 37268
rect 27682 37212 27692 37268
rect 27748 37212 29708 37268
rect 29764 37212 35084 37268
rect 35140 37212 35150 37268
rect 39778 37212 39788 37268
rect 39844 37212 41020 37268
rect 41076 37212 41086 37268
rect 42018 37212 42028 37268
rect 42084 37212 42094 37268
rect 43148 37212 45612 37268
rect 45668 37212 45678 37268
rect 42028 37156 42084 37212
rect 35634 37100 35644 37156
rect 35700 37100 36036 37156
rect 36866 37100 36876 37156
rect 36932 37100 39116 37156
rect 39172 37100 39564 37156
rect 39620 37100 41972 37156
rect 42028 37100 42700 37156
rect 42756 37100 43036 37156
rect 43092 37100 44156 37156
rect 44212 37100 44222 37156
rect 48962 37100 48972 37156
rect 49028 37100 50316 37156
rect 50372 37100 50428 37156
rect 50484 37100 51212 37156
rect 51268 37100 51278 37156
rect 54002 37100 54012 37156
rect 54068 37100 55244 37156
rect 55300 37100 55310 37156
rect 57474 37100 57484 37156
rect 57540 37100 63868 37156
rect 63924 37100 63934 37156
rect 75282 37100 75292 37156
rect 75348 37100 76188 37156
rect 76244 37100 77756 37156
rect 77812 37100 77822 37156
rect 35980 37044 36036 37100
rect 41916 37044 41972 37100
rect 99200 37044 100000 37072
rect 6066 36988 6076 37044
rect 6132 36988 6804 37044
rect 9986 36988 9996 37044
rect 10052 36988 11900 37044
rect 11956 36988 11966 37044
rect 20738 36988 20748 37044
rect 20804 36988 21084 37044
rect 21140 36988 24220 37044
rect 24276 36988 24286 37044
rect 29138 36988 29148 37044
rect 29204 36988 29932 37044
rect 29988 36988 29998 37044
rect 31714 36988 31724 37044
rect 31780 36988 32116 37044
rect 34290 36988 34300 37044
rect 34356 36988 35084 37044
rect 35140 36988 35756 37044
rect 35812 36988 35822 37044
rect 35980 36988 41692 37044
rect 41748 36988 41758 37044
rect 41916 36988 51100 37044
rect 51156 36988 51166 37044
rect 53890 36988 53900 37044
rect 53956 36988 59948 37044
rect 60004 36988 60014 37044
rect 66882 36988 66892 37044
rect 66948 36988 67228 37044
rect 67284 36988 68684 37044
rect 68740 36988 68750 37044
rect 85362 36988 85372 37044
rect 85428 36988 87500 37044
rect 87556 36988 96236 37044
rect 96292 36988 96302 37044
rect 98018 36988 98028 37044
rect 98084 36988 100000 37044
rect 6748 36932 6804 36988
rect 6738 36876 6748 36932
rect 6804 36876 6814 36932
rect 10098 36876 10108 36932
rect 10164 36876 11340 36932
rect 11396 36876 11406 36932
rect 19618 36876 19628 36932
rect 19684 36876 20524 36932
rect 20580 36876 20590 36932
rect 4258 36820 4268 36876
rect 4324 36820 4372 36876
rect 4428 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4788 36876
rect 4844 36820 4892 36876
rect 4948 36820 4958 36876
rect 13258 36820 13268 36876
rect 13324 36820 13372 36876
rect 13428 36820 13476 36876
rect 13532 36820 13580 36876
rect 13636 36820 13684 36876
rect 13740 36820 13788 36876
rect 13844 36820 13892 36876
rect 13948 36820 13958 36876
rect 22258 36820 22268 36876
rect 22324 36820 22372 36876
rect 22428 36820 22476 36876
rect 22532 36820 22580 36876
rect 22636 36820 22684 36876
rect 22740 36820 22788 36876
rect 22844 36820 22892 36876
rect 22948 36820 22958 36876
rect 31258 36820 31268 36876
rect 31324 36820 31372 36876
rect 31428 36820 31476 36876
rect 31532 36820 31580 36876
rect 31636 36820 31684 36876
rect 31740 36820 31788 36876
rect 31844 36820 31892 36876
rect 31948 36820 31958 36876
rect 32060 36708 32116 36988
rect 99200 36960 100000 36988
rect 50194 36876 50204 36932
rect 50260 36876 51436 36932
rect 51492 36876 51502 36932
rect 52098 36876 52108 36932
rect 52164 36876 56812 36932
rect 56868 36876 56878 36932
rect 69458 36876 69468 36932
rect 69524 36876 75740 36932
rect 75796 36876 75806 36932
rect 40258 36820 40268 36876
rect 40324 36820 40372 36876
rect 40428 36820 40476 36876
rect 40532 36820 40580 36876
rect 40636 36820 40684 36876
rect 40740 36820 40788 36876
rect 40844 36820 40892 36876
rect 40948 36820 40958 36876
rect 49258 36820 49268 36876
rect 49324 36820 49372 36876
rect 49428 36820 49476 36876
rect 49532 36820 49580 36876
rect 49636 36820 49684 36876
rect 49740 36820 49788 36876
rect 49844 36820 49892 36876
rect 49948 36820 49958 36876
rect 58258 36820 58268 36876
rect 58324 36820 58372 36876
rect 58428 36820 58476 36876
rect 58532 36820 58580 36876
rect 58636 36820 58684 36876
rect 58740 36820 58788 36876
rect 58844 36820 58892 36876
rect 58948 36820 58958 36876
rect 67258 36820 67268 36876
rect 67324 36820 67372 36876
rect 67428 36820 67476 36876
rect 67532 36820 67580 36876
rect 67636 36820 67684 36876
rect 67740 36820 67788 36876
rect 67844 36820 67892 36876
rect 67948 36820 67958 36876
rect 76258 36820 76268 36876
rect 76324 36820 76372 36876
rect 76428 36820 76476 36876
rect 76532 36820 76580 36876
rect 76636 36820 76684 36876
rect 76740 36820 76788 36876
rect 76844 36820 76892 36876
rect 76948 36820 76958 36876
rect 85258 36820 85268 36876
rect 85324 36820 85372 36876
rect 85428 36820 85476 36876
rect 85532 36820 85580 36876
rect 85636 36820 85684 36876
rect 85740 36820 85788 36876
rect 85844 36820 85892 36876
rect 85948 36820 85958 36876
rect 94258 36820 94268 36876
rect 94324 36820 94372 36876
rect 94428 36820 94476 36876
rect 94532 36820 94580 36876
rect 94636 36820 94684 36876
rect 94740 36820 94788 36876
rect 94844 36820 94892 36876
rect 94948 36820 94958 36876
rect 51986 36764 51996 36820
rect 52052 36764 53004 36820
rect 53060 36764 53070 36820
rect 68786 36764 68796 36820
rect 68852 36764 69580 36820
rect 69636 36764 69646 36820
rect 17602 36652 17612 36708
rect 17668 36652 18620 36708
rect 18676 36652 18956 36708
rect 19012 36652 20748 36708
rect 20804 36652 20814 36708
rect 31602 36652 31612 36708
rect 31668 36652 32116 36708
rect 36866 36652 36876 36708
rect 36932 36652 84252 36708
rect 84308 36652 84318 36708
rect 0 36596 800 36624
rect 0 36540 1708 36596
rect 1764 36540 3276 36596
rect 3332 36540 3342 36596
rect 49746 36540 49756 36596
rect 49812 36540 50876 36596
rect 50932 36540 52444 36596
rect 52500 36540 52780 36596
rect 52836 36540 52846 36596
rect 64866 36540 64876 36596
rect 64932 36540 65548 36596
rect 65604 36540 67452 36596
rect 67508 36540 68796 36596
rect 68852 36540 68862 36596
rect 73490 36540 73500 36596
rect 73556 36540 77196 36596
rect 77252 36540 77262 36596
rect 0 36512 800 36540
rect 12338 36428 12348 36484
rect 12404 36428 37100 36484
rect 37156 36428 37166 36484
rect 37314 36428 37324 36484
rect 37380 36428 77980 36484
rect 78036 36428 78046 36484
rect 37100 36372 37156 36428
rect 16146 36316 16156 36372
rect 16212 36316 17500 36372
rect 17556 36316 18508 36372
rect 18564 36316 36764 36372
rect 36820 36316 36830 36372
rect 37100 36316 37660 36372
rect 37716 36316 37726 36372
rect 52770 36316 52780 36372
rect 52836 36316 56028 36372
rect 56084 36316 56094 36372
rect 57362 36316 57372 36372
rect 57428 36316 65436 36372
rect 65492 36316 65502 36372
rect 67778 36316 67788 36372
rect 67844 36316 69468 36372
rect 69524 36316 69534 36372
rect 81554 36316 81564 36372
rect 81620 36316 96236 36372
rect 96292 36316 96302 36372
rect 5058 36204 5068 36260
rect 5124 36204 5628 36260
rect 5684 36204 5964 36260
rect 6020 36204 6300 36260
rect 6356 36204 6636 36260
rect 6692 36204 8428 36260
rect 8484 36204 11564 36260
rect 11620 36204 11630 36260
rect 30034 36204 30044 36260
rect 30100 36204 31164 36260
rect 31220 36204 34300 36260
rect 34356 36204 34366 36260
rect 42914 36204 42924 36260
rect 42980 36204 44044 36260
rect 44100 36204 53900 36260
rect 53956 36204 53966 36260
rect 78418 36204 78428 36260
rect 78484 36204 78988 36260
rect 79044 36204 84812 36260
rect 84868 36204 84878 36260
rect 89282 36204 89292 36260
rect 89348 36204 91868 36260
rect 91924 36204 91934 36260
rect 45938 36092 45948 36148
rect 46004 36092 46396 36148
rect 46452 36092 46462 36148
rect 51538 36092 51548 36148
rect 51604 36092 53452 36148
rect 53508 36092 53518 36148
rect 8758 36036 8768 36092
rect 8824 36036 8872 36092
rect 8928 36036 8976 36092
rect 9032 36036 9080 36092
rect 9136 36036 9184 36092
rect 9240 36036 9288 36092
rect 9344 36036 9392 36092
rect 9448 36036 9458 36092
rect 17758 36036 17768 36092
rect 17824 36036 17872 36092
rect 17928 36036 17976 36092
rect 18032 36036 18080 36092
rect 18136 36036 18184 36092
rect 18240 36036 18288 36092
rect 18344 36036 18392 36092
rect 18448 36036 18458 36092
rect 26758 36036 26768 36092
rect 26824 36036 26872 36092
rect 26928 36036 26976 36092
rect 27032 36036 27080 36092
rect 27136 36036 27184 36092
rect 27240 36036 27288 36092
rect 27344 36036 27392 36092
rect 27448 36036 27458 36092
rect 35758 36036 35768 36092
rect 35824 36036 35872 36092
rect 35928 36036 35976 36092
rect 36032 36036 36080 36092
rect 36136 36036 36184 36092
rect 36240 36036 36288 36092
rect 36344 36036 36392 36092
rect 36448 36036 36458 36092
rect 44758 36036 44768 36092
rect 44824 36036 44872 36092
rect 44928 36036 44976 36092
rect 45032 36036 45080 36092
rect 45136 36036 45184 36092
rect 45240 36036 45288 36092
rect 45344 36036 45392 36092
rect 45448 36036 45458 36092
rect 53758 36036 53768 36092
rect 53824 36036 53872 36092
rect 53928 36036 53976 36092
rect 54032 36036 54080 36092
rect 54136 36036 54184 36092
rect 54240 36036 54288 36092
rect 54344 36036 54392 36092
rect 54448 36036 54458 36092
rect 62758 36036 62768 36092
rect 62824 36036 62872 36092
rect 62928 36036 62976 36092
rect 63032 36036 63080 36092
rect 63136 36036 63184 36092
rect 63240 36036 63288 36092
rect 63344 36036 63392 36092
rect 63448 36036 63458 36092
rect 71758 36036 71768 36092
rect 71824 36036 71872 36092
rect 71928 36036 71976 36092
rect 72032 36036 72080 36092
rect 72136 36036 72184 36092
rect 72240 36036 72288 36092
rect 72344 36036 72392 36092
rect 72448 36036 72458 36092
rect 80758 36036 80768 36092
rect 80824 36036 80872 36092
rect 80928 36036 80976 36092
rect 81032 36036 81080 36092
rect 81136 36036 81184 36092
rect 81240 36036 81288 36092
rect 81344 36036 81392 36092
rect 81448 36036 81458 36092
rect 89758 36036 89768 36092
rect 89824 36036 89872 36092
rect 89928 36036 89976 36092
rect 90032 36036 90080 36092
rect 90136 36036 90184 36092
rect 90240 36036 90288 36092
rect 90344 36036 90392 36092
rect 90448 36036 90458 36092
rect 68114 35980 68124 36036
rect 68180 35980 68460 36036
rect 68516 35980 68526 36036
rect 92418 35980 92428 36036
rect 92484 35980 93828 36036
rect 93772 35924 93828 35980
rect 36754 35868 36764 35924
rect 36820 35868 37324 35924
rect 37380 35868 37390 35924
rect 53554 35868 53564 35924
rect 53620 35868 57148 35924
rect 57204 35868 57214 35924
rect 69570 35868 69580 35924
rect 69636 35868 71932 35924
rect 71988 35868 71998 35924
rect 73714 35868 73724 35924
rect 73780 35868 78428 35924
rect 78484 35868 78494 35924
rect 89506 35868 89516 35924
rect 89572 35868 92988 35924
rect 93044 35868 93054 35924
rect 93762 35868 93772 35924
rect 93828 35868 96124 35924
rect 96180 35868 96190 35924
rect 2034 35756 2044 35812
rect 2100 35756 2380 35812
rect 2436 35756 2446 35812
rect 8372 35756 20300 35812
rect 20356 35756 20366 35812
rect 47730 35756 47740 35812
rect 47796 35756 49084 35812
rect 49140 35756 49150 35812
rect 80210 35756 80220 35812
rect 80276 35756 81564 35812
rect 81620 35756 81630 35812
rect 84924 35756 85484 35812
rect 85540 35756 85550 35812
rect 8372 35700 8428 35756
rect 84924 35700 84980 35756
rect 89964 35700 90020 35868
rect 6178 35644 6188 35700
rect 6244 35644 8428 35700
rect 15362 35644 15372 35700
rect 15428 35644 16716 35700
rect 16772 35644 16782 35700
rect 35858 35644 35868 35700
rect 35924 35644 36652 35700
rect 36708 35644 36988 35700
rect 37044 35644 37054 35700
rect 39330 35644 39340 35700
rect 39396 35644 53788 35700
rect 53844 35644 53854 35700
rect 56018 35644 56028 35700
rect 56084 35644 57148 35700
rect 57204 35644 64540 35700
rect 64596 35644 64606 35700
rect 68198 35644 68236 35700
rect 68292 35644 68302 35700
rect 78866 35644 78876 35700
rect 78932 35644 79996 35700
rect 80052 35644 80062 35700
rect 84578 35644 84588 35700
rect 84644 35644 84980 35700
rect 85250 35644 85260 35700
rect 85316 35644 86156 35700
rect 86212 35644 86222 35700
rect 89954 35644 89964 35700
rect 90020 35644 90030 35700
rect 45042 35532 45052 35588
rect 45108 35532 46508 35588
rect 46564 35532 47068 35588
rect 47124 35532 47134 35588
rect 53442 35532 53452 35588
rect 53508 35532 56700 35588
rect 56756 35532 57820 35588
rect 57876 35532 57886 35588
rect 84914 35532 84924 35588
rect 84980 35532 84990 35588
rect 0 35476 800 35504
rect 0 35420 1708 35476
rect 1764 35420 1774 35476
rect 46610 35420 46620 35476
rect 46676 35420 47180 35476
rect 47236 35420 47246 35476
rect 74722 35420 74732 35476
rect 74788 35420 80332 35476
rect 80388 35420 80398 35476
rect 0 35392 800 35420
rect 84924 35364 84980 35532
rect 85138 35420 85148 35476
rect 85204 35420 86044 35476
rect 86100 35420 86110 35476
rect 46274 35308 46284 35364
rect 46340 35308 46350 35364
rect 68338 35308 68348 35364
rect 68404 35308 68908 35364
rect 68964 35308 68974 35364
rect 78082 35308 78092 35364
rect 78148 35308 79100 35364
rect 79156 35308 79166 35364
rect 80770 35308 80780 35364
rect 80836 35308 85092 35364
rect 4258 35252 4268 35308
rect 4324 35252 4372 35308
rect 4428 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4788 35308
rect 4844 35252 4892 35308
rect 4948 35252 4958 35308
rect 13258 35252 13268 35308
rect 13324 35252 13372 35308
rect 13428 35252 13476 35308
rect 13532 35252 13580 35308
rect 13636 35252 13684 35308
rect 13740 35252 13788 35308
rect 13844 35252 13892 35308
rect 13948 35252 13958 35308
rect 22258 35252 22268 35308
rect 22324 35252 22372 35308
rect 22428 35252 22476 35308
rect 22532 35252 22580 35308
rect 22636 35252 22684 35308
rect 22740 35252 22788 35308
rect 22844 35252 22892 35308
rect 22948 35252 22958 35308
rect 31258 35252 31268 35308
rect 31324 35252 31372 35308
rect 31428 35252 31476 35308
rect 31532 35252 31580 35308
rect 31636 35252 31684 35308
rect 31740 35252 31788 35308
rect 31844 35252 31892 35308
rect 31948 35252 31958 35308
rect 40258 35252 40268 35308
rect 40324 35252 40372 35308
rect 40428 35252 40476 35308
rect 40532 35252 40580 35308
rect 40636 35252 40684 35308
rect 40740 35252 40788 35308
rect 40844 35252 40892 35308
rect 40948 35252 40958 35308
rect 46284 35252 46340 35308
rect 49258 35252 49268 35308
rect 49324 35252 49372 35308
rect 49428 35252 49476 35308
rect 49532 35252 49580 35308
rect 49636 35252 49684 35308
rect 49740 35252 49788 35308
rect 49844 35252 49892 35308
rect 49948 35252 49958 35308
rect 58258 35252 58268 35308
rect 58324 35252 58372 35308
rect 58428 35252 58476 35308
rect 58532 35252 58580 35308
rect 58636 35252 58684 35308
rect 58740 35252 58788 35308
rect 58844 35252 58892 35308
rect 58948 35252 58958 35308
rect 67258 35252 67268 35308
rect 67324 35252 67372 35308
rect 67428 35252 67476 35308
rect 67532 35252 67580 35308
rect 67636 35252 67684 35308
rect 67740 35252 67788 35308
rect 67844 35252 67892 35308
rect 67948 35252 67958 35308
rect 76258 35252 76268 35308
rect 76324 35252 76372 35308
rect 76428 35252 76476 35308
rect 76532 35252 76580 35308
rect 76636 35252 76684 35308
rect 76740 35252 76788 35308
rect 76844 35252 76892 35308
rect 76948 35252 76958 35308
rect 46284 35196 46620 35252
rect 46676 35196 46686 35252
rect 85036 35140 85092 35308
rect 85258 35252 85268 35308
rect 85324 35252 85372 35308
rect 85428 35252 85476 35308
rect 85532 35252 85580 35308
rect 85636 35252 85684 35308
rect 85740 35252 85788 35308
rect 85844 35252 85892 35308
rect 85948 35252 85958 35308
rect 94258 35252 94268 35308
rect 94324 35252 94372 35308
rect 94428 35252 94476 35308
rect 94532 35252 94580 35308
rect 94636 35252 94684 35308
rect 94740 35252 94788 35308
rect 94844 35252 94892 35308
rect 94948 35252 94958 35308
rect 99200 35252 100000 35280
rect 97682 35196 97692 35252
rect 97748 35196 100000 35252
rect 99200 35168 100000 35196
rect 38882 35084 38892 35140
rect 38948 35084 39900 35140
rect 39956 35084 50316 35140
rect 50372 35084 50382 35140
rect 85036 35084 85372 35140
rect 85428 35084 85438 35140
rect 35298 34972 35308 35028
rect 35364 34972 40796 35028
rect 40852 34972 46620 35028
rect 46676 34972 50988 35028
rect 51044 34972 52108 35028
rect 52164 34972 52668 35028
rect 52724 34972 52734 35028
rect 54114 34972 54124 35028
rect 54180 34972 64316 35028
rect 64372 34972 64382 35028
rect 2146 34860 2156 34916
rect 2212 34860 6076 34916
rect 6132 34860 6142 34916
rect 37202 34860 37212 34916
rect 37268 34860 38668 34916
rect 38724 34860 41244 34916
rect 41300 34860 41310 34916
rect 46050 34860 46060 34916
rect 46116 34860 57540 34916
rect 57698 34860 57708 34916
rect 57764 34860 58940 34916
rect 58996 34860 59006 34916
rect 73892 34860 89068 34916
rect 89124 34860 89134 34916
rect 57484 34804 57540 34860
rect 73892 34804 73948 34860
rect 20962 34748 20972 34804
rect 21028 34748 24892 34804
rect 24948 34748 35756 34804
rect 35812 34748 35822 34804
rect 39106 34748 39116 34804
rect 39172 34748 44604 34804
rect 44660 34748 44940 34804
rect 44996 34748 45006 34804
rect 47058 34748 47068 34804
rect 47124 34748 48412 34804
rect 48468 34748 49084 34804
rect 49140 34748 49150 34804
rect 50306 34748 50316 34804
rect 50372 34748 54796 34804
rect 54852 34748 57204 34804
rect 57484 34748 61516 34804
rect 61572 34748 61582 34804
rect 64642 34748 64652 34804
rect 64708 34748 73948 34804
rect 77634 34748 77644 34804
rect 77700 34748 80780 34804
rect 80836 34748 80846 34804
rect 85810 34748 85820 34804
rect 85876 34748 88172 34804
rect 88228 34748 96236 34804
rect 96292 34748 96302 34804
rect 39116 34692 39172 34748
rect 2034 34636 2044 34692
rect 2100 34636 2716 34692
rect 2772 34636 2782 34692
rect 30930 34636 30940 34692
rect 30996 34636 36204 34692
rect 36260 34636 39172 34692
rect 44604 34636 45388 34692
rect 45444 34636 46844 34692
rect 46900 34636 48972 34692
rect 49028 34636 49308 34692
rect 49364 34636 49868 34692
rect 49924 34636 50428 34692
rect 50484 34636 50494 34692
rect 51090 34636 51100 34692
rect 51156 34636 51660 34692
rect 51716 34636 51726 34692
rect 53218 34636 53228 34692
rect 53284 34636 54684 34692
rect 54740 34636 55524 34692
rect 44604 34580 44660 34636
rect 36978 34524 36988 34580
rect 37044 34524 44660 34580
rect 55468 34580 55524 34636
rect 57148 34580 57204 34748
rect 66994 34636 67004 34692
rect 67060 34636 67900 34692
rect 67956 34636 71148 34692
rect 71204 34636 71214 34692
rect 75170 34636 75180 34692
rect 75236 34636 75852 34692
rect 75908 34636 76412 34692
rect 76468 34636 76478 34692
rect 55468 34524 56868 34580
rect 57148 34524 60732 34580
rect 60788 34524 60798 34580
rect 8758 34468 8768 34524
rect 8824 34468 8872 34524
rect 8928 34468 8976 34524
rect 9032 34468 9080 34524
rect 9136 34468 9184 34524
rect 9240 34468 9288 34524
rect 9344 34468 9392 34524
rect 9448 34468 9458 34524
rect 17758 34468 17768 34524
rect 17824 34468 17872 34524
rect 17928 34468 17976 34524
rect 18032 34468 18080 34524
rect 18136 34468 18184 34524
rect 18240 34468 18288 34524
rect 18344 34468 18392 34524
rect 18448 34468 18458 34524
rect 26758 34468 26768 34524
rect 26824 34468 26872 34524
rect 26928 34468 26976 34524
rect 27032 34468 27080 34524
rect 27136 34468 27184 34524
rect 27240 34468 27288 34524
rect 27344 34468 27392 34524
rect 27448 34468 27458 34524
rect 35758 34468 35768 34524
rect 35824 34468 35872 34524
rect 35928 34468 35976 34524
rect 36032 34468 36080 34524
rect 36136 34468 36184 34524
rect 36240 34468 36288 34524
rect 36344 34468 36392 34524
rect 36448 34468 36458 34524
rect 44758 34468 44768 34524
rect 44824 34468 44872 34524
rect 44928 34468 44976 34524
rect 45032 34468 45080 34524
rect 45136 34468 45184 34524
rect 45240 34468 45288 34524
rect 45344 34468 45392 34524
rect 45448 34468 45458 34524
rect 53758 34468 53768 34524
rect 53824 34468 53872 34524
rect 53928 34468 53976 34524
rect 54032 34468 54080 34524
rect 54136 34468 54184 34524
rect 54240 34468 54288 34524
rect 54344 34468 54392 34524
rect 54448 34468 54458 34524
rect 56812 34468 56868 34524
rect 62758 34468 62768 34524
rect 62824 34468 62872 34524
rect 62928 34468 62976 34524
rect 63032 34468 63080 34524
rect 63136 34468 63184 34524
rect 63240 34468 63288 34524
rect 63344 34468 63392 34524
rect 63448 34468 63458 34524
rect 71758 34468 71768 34524
rect 71824 34468 71872 34524
rect 71928 34468 71976 34524
rect 72032 34468 72080 34524
rect 72136 34468 72184 34524
rect 72240 34468 72288 34524
rect 72344 34468 72392 34524
rect 72448 34468 72458 34524
rect 80758 34468 80768 34524
rect 80824 34468 80872 34524
rect 80928 34468 80976 34524
rect 81032 34468 81080 34524
rect 81136 34468 81184 34524
rect 81240 34468 81288 34524
rect 81344 34468 81392 34524
rect 81448 34468 81458 34524
rect 89758 34468 89768 34524
rect 89824 34468 89872 34524
rect 89928 34468 89976 34524
rect 90032 34468 90080 34524
rect 90136 34468 90184 34524
rect 90240 34468 90288 34524
rect 90344 34468 90392 34524
rect 90448 34468 90458 34524
rect 1810 34412 1820 34468
rect 1876 34412 2380 34468
rect 2436 34412 2446 34468
rect 39554 34412 39564 34468
rect 39620 34412 40124 34468
rect 40180 34412 41468 34468
rect 41524 34412 41534 34468
rect 56812 34412 58156 34468
rect 58212 34412 58222 34468
rect 0 34356 800 34384
rect 0 34300 1708 34356
rect 1764 34300 2940 34356
rect 2996 34300 3006 34356
rect 35522 34300 35532 34356
rect 35588 34300 72492 34356
rect 72548 34300 72558 34356
rect 74498 34300 74508 34356
rect 74564 34300 75740 34356
rect 75796 34300 76188 34356
rect 76244 34300 76254 34356
rect 76402 34300 76412 34356
rect 76468 34300 84364 34356
rect 84420 34300 87388 34356
rect 87444 34300 87454 34356
rect 0 34272 800 34300
rect 4722 34188 4732 34244
rect 4788 34188 5628 34244
rect 5684 34188 5694 34244
rect 12002 34188 12012 34244
rect 12068 34188 14028 34244
rect 14084 34188 14094 34244
rect 46274 34188 46284 34244
rect 46340 34188 46620 34244
rect 46676 34188 55356 34244
rect 55412 34188 57372 34244
rect 57428 34188 57438 34244
rect 61618 34188 61628 34244
rect 61684 34188 62972 34244
rect 63028 34188 68012 34244
rect 68068 34188 68078 34244
rect 76514 34188 76524 34244
rect 76580 34188 76590 34244
rect 85362 34188 85372 34244
rect 85428 34188 85932 34244
rect 85988 34188 85998 34244
rect 76524 34132 76580 34188
rect 13234 34076 13244 34132
rect 13300 34076 36428 34132
rect 36484 34076 36494 34132
rect 47394 34076 47404 34132
rect 47460 34076 48524 34132
rect 48580 34076 49756 34132
rect 49812 34076 49822 34132
rect 50082 34076 50092 34132
rect 50148 34076 52332 34132
rect 52388 34076 52398 34132
rect 73378 34076 73388 34132
rect 73444 34076 74284 34132
rect 74340 34076 74350 34132
rect 76524 34076 96572 34132
rect 96628 34076 97020 34132
rect 97076 34076 97086 34132
rect 5282 33964 5292 34020
rect 5348 33964 19516 34020
rect 19572 33964 19582 34020
rect 30146 33964 30156 34020
rect 30212 33964 31388 34020
rect 31444 33964 31454 34020
rect 32162 33964 32172 34020
rect 32228 33964 33404 34020
rect 33460 33964 33470 34020
rect 29698 33852 29708 33908
rect 29764 33852 35308 33908
rect 35364 33852 35374 33908
rect 41234 33852 41244 33908
rect 41300 33852 44940 33908
rect 44996 33852 45006 33908
rect 4258 33684 4268 33740
rect 4324 33684 4372 33740
rect 4428 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4788 33740
rect 4844 33684 4892 33740
rect 4948 33684 4958 33740
rect 13258 33684 13268 33740
rect 13324 33684 13372 33740
rect 13428 33684 13476 33740
rect 13532 33684 13580 33740
rect 13636 33684 13684 33740
rect 13740 33684 13788 33740
rect 13844 33684 13892 33740
rect 13948 33684 13958 33740
rect 22258 33684 22268 33740
rect 22324 33684 22372 33740
rect 22428 33684 22476 33740
rect 22532 33684 22580 33740
rect 22636 33684 22684 33740
rect 22740 33684 22788 33740
rect 22844 33684 22892 33740
rect 22948 33684 22958 33740
rect 31258 33684 31268 33740
rect 31324 33684 31372 33740
rect 31428 33684 31476 33740
rect 31532 33684 31580 33740
rect 31636 33684 31684 33740
rect 31740 33684 31788 33740
rect 31844 33684 31892 33740
rect 31948 33684 31958 33740
rect 40258 33684 40268 33740
rect 40324 33684 40372 33740
rect 40428 33684 40476 33740
rect 40532 33684 40580 33740
rect 40636 33684 40684 33740
rect 40740 33684 40788 33740
rect 40844 33684 40892 33740
rect 40948 33684 40958 33740
rect 49258 33684 49268 33740
rect 49324 33684 49372 33740
rect 49428 33684 49476 33740
rect 49532 33684 49580 33740
rect 49636 33684 49684 33740
rect 49740 33684 49788 33740
rect 49844 33684 49892 33740
rect 49948 33684 49958 33740
rect 58258 33684 58268 33740
rect 58324 33684 58372 33740
rect 58428 33684 58476 33740
rect 58532 33684 58580 33740
rect 58636 33684 58684 33740
rect 58740 33684 58788 33740
rect 58844 33684 58892 33740
rect 58948 33684 58958 33740
rect 67258 33684 67268 33740
rect 67324 33684 67372 33740
rect 67428 33684 67476 33740
rect 67532 33684 67580 33740
rect 67636 33684 67684 33740
rect 67740 33684 67788 33740
rect 67844 33684 67892 33740
rect 67948 33684 67958 33740
rect 76258 33684 76268 33740
rect 76324 33684 76372 33740
rect 76428 33684 76476 33740
rect 76532 33684 76580 33740
rect 76636 33684 76684 33740
rect 76740 33684 76788 33740
rect 76844 33684 76892 33740
rect 76948 33684 76958 33740
rect 85258 33684 85268 33740
rect 85324 33684 85372 33740
rect 85428 33684 85476 33740
rect 85532 33684 85580 33740
rect 85636 33684 85684 33740
rect 85740 33684 85788 33740
rect 85844 33684 85892 33740
rect 85948 33684 85958 33740
rect 94258 33684 94268 33740
rect 94324 33684 94372 33740
rect 94428 33684 94476 33740
rect 94532 33684 94580 33740
rect 94636 33684 94684 33740
rect 94740 33684 94788 33740
rect 94844 33684 94892 33740
rect 94948 33684 94958 33740
rect 8642 33628 8652 33684
rect 8708 33628 12012 33684
rect 12068 33628 12078 33684
rect 63634 33628 63644 33684
rect 63700 33628 64652 33684
rect 64708 33628 64718 33684
rect 66098 33628 66108 33684
rect 66164 33628 67004 33684
rect 67060 33628 67070 33684
rect 38434 33516 38444 33572
rect 38500 33516 39228 33572
rect 39284 33516 39294 33572
rect 44146 33516 44156 33572
rect 44212 33516 44604 33572
rect 44660 33516 50428 33572
rect 61058 33516 61068 33572
rect 61124 33516 62524 33572
rect 62580 33516 62590 33572
rect 50372 33460 50428 33516
rect 99200 33460 100000 33488
rect 10098 33404 10108 33460
rect 10164 33404 14588 33460
rect 14644 33404 19068 33460
rect 19124 33404 19628 33460
rect 19684 33404 19694 33460
rect 44706 33404 44716 33460
rect 44772 33404 45948 33460
rect 46004 33404 47852 33460
rect 47908 33404 48860 33460
rect 48916 33404 48926 33460
rect 50372 33404 60844 33460
rect 60900 33404 62076 33460
rect 62132 33404 62142 33460
rect 97682 33404 97692 33460
rect 97748 33404 100000 33460
rect 99200 33376 100000 33404
rect 9538 33292 9548 33348
rect 9604 33292 15372 33348
rect 15428 33292 15438 33348
rect 45154 33292 45164 33348
rect 45220 33292 46172 33348
rect 46228 33292 46238 33348
rect 61842 33292 61852 33348
rect 61908 33292 62412 33348
rect 62468 33292 62478 33348
rect 73042 33292 73052 33348
rect 73108 33292 74508 33348
rect 74564 33292 75068 33348
rect 75124 33292 75134 33348
rect 0 33236 800 33264
rect 0 33180 1708 33236
rect 1764 33180 2492 33236
rect 2548 33180 2558 33236
rect 48738 33180 48748 33236
rect 48804 33180 59836 33236
rect 59892 33180 59902 33236
rect 0 33152 800 33180
rect 32498 33068 32508 33124
rect 32564 33068 35868 33124
rect 35924 33068 35934 33124
rect 44930 33068 44940 33124
rect 44996 33068 46396 33124
rect 46452 33068 48300 33124
rect 48356 33068 48366 33124
rect 50418 33068 50428 33124
rect 50484 33068 60284 33124
rect 60340 33068 60350 33124
rect 63186 33068 63196 33124
rect 63252 33068 63756 33124
rect 63812 33068 66668 33124
rect 66724 33068 66734 33124
rect 50428 33012 50484 33068
rect 48178 32956 48188 33012
rect 48244 32956 50484 33012
rect 8758 32900 8768 32956
rect 8824 32900 8872 32956
rect 8928 32900 8976 32956
rect 9032 32900 9080 32956
rect 9136 32900 9184 32956
rect 9240 32900 9288 32956
rect 9344 32900 9392 32956
rect 9448 32900 9458 32956
rect 17758 32900 17768 32956
rect 17824 32900 17872 32956
rect 17928 32900 17976 32956
rect 18032 32900 18080 32956
rect 18136 32900 18184 32956
rect 18240 32900 18288 32956
rect 18344 32900 18392 32956
rect 18448 32900 18458 32956
rect 26758 32900 26768 32956
rect 26824 32900 26872 32956
rect 26928 32900 26976 32956
rect 27032 32900 27080 32956
rect 27136 32900 27184 32956
rect 27240 32900 27288 32956
rect 27344 32900 27392 32956
rect 27448 32900 27458 32956
rect 35758 32900 35768 32956
rect 35824 32900 35872 32956
rect 35928 32900 35976 32956
rect 36032 32900 36080 32956
rect 36136 32900 36184 32956
rect 36240 32900 36288 32956
rect 36344 32900 36392 32956
rect 36448 32900 36458 32956
rect 44758 32900 44768 32956
rect 44824 32900 44872 32956
rect 44928 32900 44976 32956
rect 45032 32900 45080 32956
rect 45136 32900 45184 32956
rect 45240 32900 45288 32956
rect 45344 32900 45392 32956
rect 45448 32900 45458 32956
rect 53758 32900 53768 32956
rect 53824 32900 53872 32956
rect 53928 32900 53976 32956
rect 54032 32900 54080 32956
rect 54136 32900 54184 32956
rect 54240 32900 54288 32956
rect 54344 32900 54392 32956
rect 54448 32900 54458 32956
rect 62758 32900 62768 32956
rect 62824 32900 62872 32956
rect 62928 32900 62976 32956
rect 63032 32900 63080 32956
rect 63136 32900 63184 32956
rect 63240 32900 63288 32956
rect 63344 32900 63392 32956
rect 63448 32900 63458 32956
rect 71758 32900 71768 32956
rect 71824 32900 71872 32956
rect 71928 32900 71976 32956
rect 72032 32900 72080 32956
rect 72136 32900 72184 32956
rect 72240 32900 72288 32956
rect 72344 32900 72392 32956
rect 72448 32900 72458 32956
rect 80758 32900 80768 32956
rect 80824 32900 80872 32956
rect 80928 32900 80976 32956
rect 81032 32900 81080 32956
rect 81136 32900 81184 32956
rect 81240 32900 81288 32956
rect 81344 32900 81392 32956
rect 81448 32900 81458 32956
rect 89758 32900 89768 32956
rect 89824 32900 89872 32956
rect 89928 32900 89976 32956
rect 90032 32900 90080 32956
rect 90136 32900 90184 32956
rect 90240 32900 90288 32956
rect 90344 32900 90392 32956
rect 90448 32900 90458 32956
rect 39890 32732 39900 32788
rect 39956 32732 41020 32788
rect 41076 32732 41580 32788
rect 41636 32732 42364 32788
rect 42420 32732 42924 32788
rect 42980 32732 42990 32788
rect 54562 32732 54572 32788
rect 54628 32732 55244 32788
rect 55300 32732 55692 32788
rect 55748 32732 56364 32788
rect 56420 32732 57148 32788
rect 57204 32732 57820 32788
rect 57876 32732 61068 32788
rect 61124 32732 61134 32788
rect 8372 32620 8540 32676
rect 8596 32620 12348 32676
rect 12404 32620 12414 32676
rect 15138 32620 15148 32676
rect 15204 32620 16156 32676
rect 16212 32620 16222 32676
rect 20290 32620 20300 32676
rect 20356 32620 23436 32676
rect 23492 32620 23502 32676
rect 26852 32620 35980 32676
rect 36036 32620 36046 32676
rect 39778 32620 39788 32676
rect 39844 32620 41468 32676
rect 41524 32620 41534 32676
rect 55412 32620 56028 32676
rect 56084 32620 57260 32676
rect 57316 32620 57326 32676
rect 59826 32620 59836 32676
rect 59892 32620 63308 32676
rect 63364 32620 68236 32676
rect 68292 32620 68302 32676
rect 8372 32564 8428 32620
rect 5618 32508 5628 32564
rect 5684 32508 8428 32564
rect 9090 32508 9100 32564
rect 9156 32508 9996 32564
rect 10052 32508 10062 32564
rect 26852 32340 26908 32620
rect 30034 32508 30044 32564
rect 30100 32508 38668 32564
rect 40226 32508 40236 32564
rect 40292 32508 43820 32564
rect 43876 32508 43886 32564
rect 50082 32508 50092 32564
rect 50148 32508 50876 32564
rect 50932 32508 50942 32564
rect 53106 32508 53116 32564
rect 53172 32508 53788 32564
rect 53844 32508 53854 32564
rect 38612 32452 38668 32508
rect 55412 32452 55468 32620
rect 57026 32508 57036 32564
rect 57092 32508 59164 32564
rect 59220 32508 61740 32564
rect 61796 32508 61806 32564
rect 62132 32508 62972 32564
rect 63028 32508 64540 32564
rect 64596 32508 64606 32564
rect 62132 32452 62188 32508
rect 29026 32396 29036 32452
rect 29092 32396 30156 32452
rect 30212 32396 32508 32452
rect 32564 32396 32574 32452
rect 38612 32396 44492 32452
rect 44548 32396 53340 32452
rect 53396 32396 55468 32452
rect 60274 32396 60284 32452
rect 60340 32396 62188 32452
rect 14578 32284 14588 32340
rect 14644 32284 15484 32340
rect 15540 32284 15550 32340
rect 20402 32284 20412 32340
rect 20468 32284 24220 32340
rect 24276 32284 26908 32340
rect 38546 32284 38556 32340
rect 38612 32284 39900 32340
rect 39956 32284 41804 32340
rect 41860 32284 41870 32340
rect 51202 32284 51212 32340
rect 51268 32284 53452 32340
rect 53508 32284 53518 32340
rect 0 32116 800 32144
rect 4258 32116 4268 32172
rect 4324 32116 4372 32172
rect 4428 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4788 32172
rect 4844 32116 4892 32172
rect 4948 32116 4958 32172
rect 13258 32116 13268 32172
rect 13324 32116 13372 32172
rect 13428 32116 13476 32172
rect 13532 32116 13580 32172
rect 13636 32116 13684 32172
rect 13740 32116 13788 32172
rect 13844 32116 13892 32172
rect 13948 32116 13958 32172
rect 22258 32116 22268 32172
rect 22324 32116 22372 32172
rect 22428 32116 22476 32172
rect 22532 32116 22580 32172
rect 22636 32116 22684 32172
rect 22740 32116 22788 32172
rect 22844 32116 22892 32172
rect 22948 32116 22958 32172
rect 31258 32116 31268 32172
rect 31324 32116 31372 32172
rect 31428 32116 31476 32172
rect 31532 32116 31580 32172
rect 31636 32116 31684 32172
rect 31740 32116 31788 32172
rect 31844 32116 31892 32172
rect 31948 32116 31958 32172
rect 40258 32116 40268 32172
rect 40324 32116 40372 32172
rect 40428 32116 40476 32172
rect 40532 32116 40580 32172
rect 40636 32116 40684 32172
rect 40740 32116 40788 32172
rect 40844 32116 40892 32172
rect 40948 32116 40958 32172
rect 49258 32116 49268 32172
rect 49324 32116 49372 32172
rect 49428 32116 49476 32172
rect 49532 32116 49580 32172
rect 49636 32116 49684 32172
rect 49740 32116 49788 32172
rect 49844 32116 49892 32172
rect 49948 32116 49958 32172
rect 58258 32116 58268 32172
rect 58324 32116 58372 32172
rect 58428 32116 58476 32172
rect 58532 32116 58580 32172
rect 58636 32116 58684 32172
rect 58740 32116 58788 32172
rect 58844 32116 58892 32172
rect 58948 32116 58958 32172
rect 67258 32116 67268 32172
rect 67324 32116 67372 32172
rect 67428 32116 67476 32172
rect 67532 32116 67580 32172
rect 67636 32116 67684 32172
rect 67740 32116 67788 32172
rect 67844 32116 67892 32172
rect 67948 32116 67958 32172
rect 76258 32116 76268 32172
rect 76324 32116 76372 32172
rect 76428 32116 76476 32172
rect 76532 32116 76580 32172
rect 76636 32116 76684 32172
rect 76740 32116 76788 32172
rect 76844 32116 76892 32172
rect 76948 32116 76958 32172
rect 85258 32116 85268 32172
rect 85324 32116 85372 32172
rect 85428 32116 85476 32172
rect 85532 32116 85580 32172
rect 85636 32116 85684 32172
rect 85740 32116 85788 32172
rect 85844 32116 85892 32172
rect 85948 32116 85958 32172
rect 94258 32116 94268 32172
rect 94324 32116 94372 32172
rect 94428 32116 94476 32172
rect 94532 32116 94580 32172
rect 94636 32116 94684 32172
rect 94740 32116 94788 32172
rect 94844 32116 94892 32172
rect 94948 32116 94958 32172
rect 0 32060 1708 32116
rect 1764 32060 2492 32116
rect 2548 32060 2558 32116
rect 45836 32060 47124 32116
rect 53106 32060 53116 32116
rect 53172 32060 54460 32116
rect 54516 32060 54526 32116
rect 0 32032 800 32060
rect 45836 32004 45892 32060
rect 47068 32004 47124 32060
rect 53116 32004 53172 32060
rect 1810 31948 1820 32004
rect 1876 31948 2212 32004
rect 41682 31948 41692 32004
rect 41748 31948 42364 32004
rect 42420 31948 45612 32004
rect 45668 31948 45678 32004
rect 45826 31948 45836 32004
rect 45892 31948 45902 32004
rect 46162 31948 46172 32004
rect 46228 31948 46844 32004
rect 46900 31948 46910 32004
rect 47068 31948 53172 32004
rect 62514 31948 62524 32004
rect 62580 31948 64092 32004
rect 64148 31948 64158 32004
rect 2156 31892 2212 31948
rect 2156 31836 3276 31892
rect 3332 31836 3342 31892
rect 9202 31836 9212 31892
rect 9268 31836 30604 31892
rect 30660 31836 30670 31892
rect 44034 31836 44044 31892
rect 44100 31836 46396 31892
rect 46452 31836 46462 31892
rect 63522 31836 63532 31892
rect 63588 31836 64428 31892
rect 64484 31836 67004 31892
rect 67060 31836 67900 31892
rect 67956 31836 68572 31892
rect 68628 31836 68638 31892
rect 70690 31836 70700 31892
rect 70756 31836 72940 31892
rect 72996 31836 73006 31892
rect 2594 31724 2604 31780
rect 2660 31724 6076 31780
rect 6132 31724 6142 31780
rect 27122 31724 27132 31780
rect 27188 31724 28140 31780
rect 28196 31724 28206 31780
rect 41458 31724 41468 31780
rect 41524 31724 42700 31780
rect 42756 31724 42766 31780
rect 43362 31724 43372 31780
rect 43428 31724 44828 31780
rect 44884 31724 44894 31780
rect 99200 31668 100000 31696
rect 16706 31612 16716 31668
rect 16772 31612 18060 31668
rect 18116 31612 35868 31668
rect 35924 31612 36316 31668
rect 36372 31612 36382 31668
rect 36530 31612 36540 31668
rect 36596 31612 65100 31668
rect 65156 31612 65166 31668
rect 72930 31612 72940 31668
rect 72996 31612 74060 31668
rect 74116 31612 74126 31668
rect 98018 31612 98028 31668
rect 98084 31612 100000 31668
rect 99200 31584 100000 31612
rect 1698 31500 1708 31556
rect 1764 31500 2940 31556
rect 2996 31500 3006 31556
rect 17490 31500 17500 31556
rect 17556 31500 18396 31556
rect 18452 31500 19964 31556
rect 20020 31500 20030 31556
rect 26450 31500 26460 31556
rect 26516 31500 27468 31556
rect 27524 31500 27534 31556
rect 38882 31500 38892 31556
rect 38948 31500 39788 31556
rect 39844 31500 40684 31556
rect 40740 31500 40750 31556
rect 43810 31500 43820 31556
rect 43876 31500 45388 31556
rect 45444 31500 45454 31556
rect 55346 31500 55356 31556
rect 55412 31500 56476 31556
rect 56532 31500 56542 31556
rect 64642 31500 64652 31556
rect 64708 31500 65324 31556
rect 65380 31500 66556 31556
rect 66612 31500 66622 31556
rect 68898 31500 68908 31556
rect 68964 31500 71148 31556
rect 71204 31500 72156 31556
rect 72212 31500 72222 31556
rect 74386 31500 74396 31556
rect 74452 31500 96684 31556
rect 96740 31500 96750 31556
rect 66556 31444 66612 31500
rect 66556 31388 69020 31444
rect 69076 31388 69916 31444
rect 69972 31388 70700 31444
rect 70756 31388 70766 31444
rect 8758 31332 8768 31388
rect 8824 31332 8872 31388
rect 8928 31332 8976 31388
rect 9032 31332 9080 31388
rect 9136 31332 9184 31388
rect 9240 31332 9288 31388
rect 9344 31332 9392 31388
rect 9448 31332 9458 31388
rect 17758 31332 17768 31388
rect 17824 31332 17872 31388
rect 17928 31332 17976 31388
rect 18032 31332 18080 31388
rect 18136 31332 18184 31388
rect 18240 31332 18288 31388
rect 18344 31332 18392 31388
rect 18448 31332 18458 31388
rect 26758 31332 26768 31388
rect 26824 31332 26872 31388
rect 26928 31332 26976 31388
rect 27032 31332 27080 31388
rect 27136 31332 27184 31388
rect 27240 31332 27288 31388
rect 27344 31332 27392 31388
rect 27448 31332 27458 31388
rect 35758 31332 35768 31388
rect 35824 31332 35872 31388
rect 35928 31332 35976 31388
rect 36032 31332 36080 31388
rect 36136 31332 36184 31388
rect 36240 31332 36288 31388
rect 36344 31332 36392 31388
rect 36448 31332 36458 31388
rect 44758 31332 44768 31388
rect 44824 31332 44872 31388
rect 44928 31332 44976 31388
rect 45032 31332 45080 31388
rect 45136 31332 45184 31388
rect 45240 31332 45288 31388
rect 45344 31332 45392 31388
rect 45448 31332 45458 31388
rect 53758 31332 53768 31388
rect 53824 31332 53872 31388
rect 53928 31332 53976 31388
rect 54032 31332 54080 31388
rect 54136 31332 54184 31388
rect 54240 31332 54288 31388
rect 54344 31332 54392 31388
rect 54448 31332 54458 31388
rect 62758 31332 62768 31388
rect 62824 31332 62872 31388
rect 62928 31332 62976 31388
rect 63032 31332 63080 31388
rect 63136 31332 63184 31388
rect 63240 31332 63288 31388
rect 63344 31332 63392 31388
rect 63448 31332 63458 31388
rect 71758 31332 71768 31388
rect 71824 31332 71872 31388
rect 71928 31332 71976 31388
rect 72032 31332 72080 31388
rect 72136 31332 72184 31388
rect 72240 31332 72288 31388
rect 72344 31332 72392 31388
rect 72448 31332 72458 31388
rect 80758 31332 80768 31388
rect 80824 31332 80872 31388
rect 80928 31332 80976 31388
rect 81032 31332 81080 31388
rect 81136 31332 81184 31388
rect 81240 31332 81288 31388
rect 81344 31332 81392 31388
rect 81448 31332 81458 31388
rect 89758 31332 89768 31388
rect 89824 31332 89872 31388
rect 89928 31332 89976 31388
rect 90032 31332 90080 31388
rect 90136 31332 90184 31388
rect 90240 31332 90288 31388
rect 90344 31332 90392 31388
rect 90448 31332 90458 31388
rect 1810 31164 1820 31220
rect 1876 31164 2380 31220
rect 2436 31164 2446 31220
rect 36866 31164 36876 31220
rect 36932 31164 55468 31220
rect 65090 31164 65100 31220
rect 65156 31164 65996 31220
rect 66052 31164 66062 31220
rect 55412 31108 55468 31164
rect 55412 31052 69468 31108
rect 69524 31052 69534 31108
rect 0 30996 800 31024
rect 0 30940 1708 30996
rect 1764 30940 1774 30996
rect 8372 30940 20412 30996
rect 20468 30940 21644 30996
rect 21700 30940 21710 30996
rect 32162 30940 32172 30996
rect 32228 30940 33516 30996
rect 33572 30940 33582 30996
rect 45042 30940 45052 30996
rect 45108 30940 45724 30996
rect 45780 30940 47180 30996
rect 47236 30940 47246 30996
rect 65202 30940 65212 30996
rect 65268 30940 65436 30996
rect 65492 30940 65502 30996
rect 70354 30940 70364 30996
rect 70420 30940 72268 30996
rect 72324 30940 72334 30996
rect 0 30912 800 30940
rect 8372 30884 8428 30940
rect 3266 30828 3276 30884
rect 3332 30828 8428 30884
rect 31714 30828 31724 30884
rect 31780 30828 33180 30884
rect 33236 30828 33246 30884
rect 46274 30828 46284 30884
rect 46340 30828 46956 30884
rect 47012 30828 47022 30884
rect 27906 30716 27916 30772
rect 27972 30716 29932 30772
rect 29988 30716 37100 30772
rect 37156 30716 37166 30772
rect 4258 30548 4268 30604
rect 4324 30548 4372 30604
rect 4428 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4788 30604
rect 4844 30548 4892 30604
rect 4948 30548 4958 30604
rect 13258 30548 13268 30604
rect 13324 30548 13372 30604
rect 13428 30548 13476 30604
rect 13532 30548 13580 30604
rect 13636 30548 13684 30604
rect 13740 30548 13788 30604
rect 13844 30548 13892 30604
rect 13948 30548 13958 30604
rect 22258 30548 22268 30604
rect 22324 30548 22372 30604
rect 22428 30548 22476 30604
rect 22532 30548 22580 30604
rect 22636 30548 22684 30604
rect 22740 30548 22788 30604
rect 22844 30548 22892 30604
rect 22948 30548 22958 30604
rect 31258 30548 31268 30604
rect 31324 30548 31372 30604
rect 31428 30548 31476 30604
rect 31532 30548 31580 30604
rect 31636 30548 31684 30604
rect 31740 30548 31788 30604
rect 31844 30548 31892 30604
rect 31948 30548 31958 30604
rect 40258 30548 40268 30604
rect 40324 30548 40372 30604
rect 40428 30548 40476 30604
rect 40532 30548 40580 30604
rect 40636 30548 40684 30604
rect 40740 30548 40788 30604
rect 40844 30548 40892 30604
rect 40948 30548 40958 30604
rect 49258 30548 49268 30604
rect 49324 30548 49372 30604
rect 49428 30548 49476 30604
rect 49532 30548 49580 30604
rect 49636 30548 49684 30604
rect 49740 30548 49788 30604
rect 49844 30548 49892 30604
rect 49948 30548 49958 30604
rect 58258 30548 58268 30604
rect 58324 30548 58372 30604
rect 58428 30548 58476 30604
rect 58532 30548 58580 30604
rect 58636 30548 58684 30604
rect 58740 30548 58788 30604
rect 58844 30548 58892 30604
rect 58948 30548 58958 30604
rect 67258 30548 67268 30604
rect 67324 30548 67372 30604
rect 67428 30548 67476 30604
rect 67532 30548 67580 30604
rect 67636 30548 67684 30604
rect 67740 30548 67788 30604
rect 67844 30548 67892 30604
rect 67948 30548 67958 30604
rect 76258 30548 76268 30604
rect 76324 30548 76372 30604
rect 76428 30548 76476 30604
rect 76532 30548 76580 30604
rect 76636 30548 76684 30604
rect 76740 30548 76788 30604
rect 76844 30548 76892 30604
rect 76948 30548 76958 30604
rect 85258 30548 85268 30604
rect 85324 30548 85372 30604
rect 85428 30548 85476 30604
rect 85532 30548 85580 30604
rect 85636 30548 85684 30604
rect 85740 30548 85788 30604
rect 85844 30548 85892 30604
rect 85948 30548 85958 30604
rect 94258 30548 94268 30604
rect 94324 30548 94372 30604
rect 94428 30548 94476 30604
rect 94532 30548 94580 30604
rect 94636 30548 94684 30604
rect 94740 30548 94788 30604
rect 94844 30548 94892 30604
rect 94948 30548 94958 30604
rect 15922 30268 15932 30324
rect 15988 30268 16828 30324
rect 16884 30268 16894 30324
rect 19954 30268 19964 30324
rect 20020 30268 20188 30324
rect 44146 30268 44156 30324
rect 44212 30268 44492 30324
rect 44548 30268 44558 30324
rect 2594 30156 2604 30212
rect 2660 30156 9436 30212
rect 9492 30156 9502 30212
rect 20132 30100 20188 30268
rect 25442 30156 25452 30212
rect 25508 30156 26236 30212
rect 26292 30156 27244 30212
rect 27300 30156 30268 30212
rect 30324 30156 30940 30212
rect 30996 30156 31006 30212
rect 32722 30156 32732 30212
rect 32788 30156 33068 30212
rect 33124 30156 35868 30212
rect 35924 30156 35934 30212
rect 36978 30156 36988 30212
rect 37044 30156 38780 30212
rect 38836 30156 38846 30212
rect 42130 30156 42140 30212
rect 42196 30156 44044 30212
rect 44100 30156 45052 30212
rect 45108 30156 45724 30212
rect 45780 30156 46508 30212
rect 46564 30156 46844 30212
rect 46900 30156 46910 30212
rect 47058 30156 47068 30212
rect 47124 30156 49756 30212
rect 49812 30156 49822 30212
rect 66658 30156 66668 30212
rect 66724 30156 68572 30212
rect 68628 30156 72492 30212
rect 72548 30156 72558 30212
rect 77410 30156 77420 30212
rect 77476 30156 83468 30212
rect 83524 30156 84476 30212
rect 84532 30156 91308 30212
rect 91364 30156 91374 30212
rect 14690 30044 14700 30100
rect 14756 30044 16268 30100
rect 16324 30044 16334 30100
rect 20132 30044 21532 30100
rect 21588 30044 22428 30100
rect 22484 30044 23996 30100
rect 24052 30044 24062 30100
rect 42466 30044 42476 30100
rect 42532 30044 43596 30100
rect 43652 30044 44604 30100
rect 44660 30044 44940 30100
rect 44996 30044 45006 30100
rect 46162 30044 46172 30100
rect 46228 30044 49196 30100
rect 49252 30044 49262 30100
rect 72818 30044 72828 30100
rect 72884 30044 96684 30100
rect 96740 30044 96750 30100
rect 9986 29932 9996 29988
rect 10052 29932 12012 29988
rect 12068 29932 12078 29988
rect 43698 29932 43708 29988
rect 43764 29932 59052 29988
rect 59108 29932 61628 29988
rect 61684 29932 61694 29988
rect 0 29876 800 29904
rect 99200 29876 100000 29904
rect 0 29820 1708 29876
rect 1764 29820 2492 29876
rect 2548 29820 2558 29876
rect 98018 29820 98028 29876
rect 98084 29820 100000 29876
rect 0 29792 800 29820
rect 8758 29764 8768 29820
rect 8824 29764 8872 29820
rect 8928 29764 8976 29820
rect 9032 29764 9080 29820
rect 9136 29764 9184 29820
rect 9240 29764 9288 29820
rect 9344 29764 9392 29820
rect 9448 29764 9458 29820
rect 17758 29764 17768 29820
rect 17824 29764 17872 29820
rect 17928 29764 17976 29820
rect 18032 29764 18080 29820
rect 18136 29764 18184 29820
rect 18240 29764 18288 29820
rect 18344 29764 18392 29820
rect 18448 29764 18458 29820
rect 26758 29764 26768 29820
rect 26824 29764 26872 29820
rect 26928 29764 26976 29820
rect 27032 29764 27080 29820
rect 27136 29764 27184 29820
rect 27240 29764 27288 29820
rect 27344 29764 27392 29820
rect 27448 29764 27458 29820
rect 35758 29764 35768 29820
rect 35824 29764 35872 29820
rect 35928 29764 35976 29820
rect 36032 29764 36080 29820
rect 36136 29764 36184 29820
rect 36240 29764 36288 29820
rect 36344 29764 36392 29820
rect 36448 29764 36458 29820
rect 44758 29764 44768 29820
rect 44824 29764 44872 29820
rect 44928 29764 44976 29820
rect 45032 29764 45080 29820
rect 45136 29764 45184 29820
rect 45240 29764 45288 29820
rect 45344 29764 45392 29820
rect 45448 29764 45458 29820
rect 53758 29764 53768 29820
rect 53824 29764 53872 29820
rect 53928 29764 53976 29820
rect 54032 29764 54080 29820
rect 54136 29764 54184 29820
rect 54240 29764 54288 29820
rect 54344 29764 54392 29820
rect 54448 29764 54458 29820
rect 62758 29764 62768 29820
rect 62824 29764 62872 29820
rect 62928 29764 62976 29820
rect 63032 29764 63080 29820
rect 63136 29764 63184 29820
rect 63240 29764 63288 29820
rect 63344 29764 63392 29820
rect 63448 29764 63458 29820
rect 71758 29764 71768 29820
rect 71824 29764 71872 29820
rect 71928 29764 71976 29820
rect 72032 29764 72080 29820
rect 72136 29764 72184 29820
rect 72240 29764 72288 29820
rect 72344 29764 72392 29820
rect 72448 29764 72458 29820
rect 80758 29764 80768 29820
rect 80824 29764 80872 29820
rect 80928 29764 80976 29820
rect 81032 29764 81080 29820
rect 81136 29764 81184 29820
rect 81240 29764 81288 29820
rect 81344 29764 81392 29820
rect 81448 29764 81458 29820
rect 89758 29764 89768 29820
rect 89824 29764 89872 29820
rect 89928 29764 89976 29820
rect 90032 29764 90080 29820
rect 90136 29764 90184 29820
rect 90240 29764 90288 29820
rect 90344 29764 90392 29820
rect 90448 29764 90458 29820
rect 99200 29792 100000 29820
rect 40002 29708 40012 29764
rect 40068 29708 44156 29764
rect 44212 29708 44222 29764
rect 49298 29708 49308 29764
rect 49364 29708 50540 29764
rect 50596 29708 50606 29764
rect 5282 29596 5292 29652
rect 5348 29596 26572 29652
rect 26628 29596 26638 29652
rect 33170 29596 33180 29652
rect 33236 29596 36652 29652
rect 36708 29596 61628 29652
rect 61684 29596 61694 29652
rect 69010 29596 69020 29652
rect 69076 29596 69692 29652
rect 69748 29596 69758 29652
rect 44146 29484 44156 29540
rect 44212 29484 46396 29540
rect 46452 29484 46462 29540
rect 53218 29484 53228 29540
rect 53284 29484 54236 29540
rect 54292 29484 55244 29540
rect 55300 29484 55310 29540
rect 56914 29484 56924 29540
rect 56980 29484 57596 29540
rect 57652 29484 64652 29540
rect 64708 29484 64718 29540
rect 2370 29372 2380 29428
rect 2436 29372 17724 29428
rect 17780 29372 18956 29428
rect 19012 29372 19022 29428
rect 44706 29372 44716 29428
rect 44772 29372 45500 29428
rect 45556 29372 46060 29428
rect 46116 29372 46956 29428
rect 47012 29372 47022 29428
rect 54898 29372 54908 29428
rect 54964 29372 56812 29428
rect 56868 29372 56878 29428
rect 69234 29372 69244 29428
rect 69300 29372 70476 29428
rect 70532 29372 70542 29428
rect 75394 29372 75404 29428
rect 75460 29372 75852 29428
rect 75908 29372 77420 29428
rect 77476 29372 77486 29428
rect 6066 29260 6076 29316
rect 6132 29260 13020 29316
rect 13076 29260 16156 29316
rect 16212 29260 16222 29316
rect 43250 29260 43260 29316
rect 43316 29260 44044 29316
rect 44100 29260 45836 29316
rect 45892 29260 45902 29316
rect 68338 29260 68348 29316
rect 68404 29260 68572 29316
rect 68628 29260 68638 29316
rect 41682 29148 41692 29204
rect 41748 29148 42140 29204
rect 42196 29148 42206 29204
rect 49746 29148 49756 29204
rect 49812 29148 53676 29204
rect 53732 29148 53742 29204
rect 4258 28980 4268 29036
rect 4324 28980 4372 29036
rect 4428 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4788 29036
rect 4844 28980 4892 29036
rect 4948 28980 4958 29036
rect 13258 28980 13268 29036
rect 13324 28980 13372 29036
rect 13428 28980 13476 29036
rect 13532 28980 13580 29036
rect 13636 28980 13684 29036
rect 13740 28980 13788 29036
rect 13844 28980 13892 29036
rect 13948 28980 13958 29036
rect 22258 28980 22268 29036
rect 22324 28980 22372 29036
rect 22428 28980 22476 29036
rect 22532 28980 22580 29036
rect 22636 28980 22684 29036
rect 22740 28980 22788 29036
rect 22844 28980 22892 29036
rect 22948 28980 22958 29036
rect 31258 28980 31268 29036
rect 31324 28980 31372 29036
rect 31428 28980 31476 29036
rect 31532 28980 31580 29036
rect 31636 28980 31684 29036
rect 31740 28980 31788 29036
rect 31844 28980 31892 29036
rect 31948 28980 31958 29036
rect 40258 28980 40268 29036
rect 40324 28980 40372 29036
rect 40428 28980 40476 29036
rect 40532 28980 40580 29036
rect 40636 28980 40684 29036
rect 40740 28980 40788 29036
rect 40844 28980 40892 29036
rect 40948 28980 40958 29036
rect 49258 28980 49268 29036
rect 49324 28980 49372 29036
rect 49428 28980 49476 29036
rect 49532 28980 49580 29036
rect 49636 28980 49684 29036
rect 49740 28980 49788 29036
rect 49844 28980 49892 29036
rect 49948 28980 49958 29036
rect 58258 28980 58268 29036
rect 58324 28980 58372 29036
rect 58428 28980 58476 29036
rect 58532 28980 58580 29036
rect 58636 28980 58684 29036
rect 58740 28980 58788 29036
rect 58844 28980 58892 29036
rect 58948 28980 58958 29036
rect 67258 28980 67268 29036
rect 67324 28980 67372 29036
rect 67428 28980 67476 29036
rect 67532 28980 67580 29036
rect 67636 28980 67684 29036
rect 67740 28980 67788 29036
rect 67844 28980 67892 29036
rect 67948 28980 67958 29036
rect 76258 28980 76268 29036
rect 76324 28980 76372 29036
rect 76428 28980 76476 29036
rect 76532 28980 76580 29036
rect 76636 28980 76684 29036
rect 76740 28980 76788 29036
rect 76844 28980 76892 29036
rect 76948 28980 76958 29036
rect 85258 28980 85268 29036
rect 85324 28980 85372 29036
rect 85428 28980 85476 29036
rect 85532 28980 85580 29036
rect 85636 28980 85684 29036
rect 85740 28980 85788 29036
rect 85844 28980 85892 29036
rect 85948 28980 85958 29036
rect 94258 28980 94268 29036
rect 94324 28980 94372 29036
rect 94428 28980 94476 29036
rect 94532 28980 94580 29036
rect 94636 28980 94684 29036
rect 94740 28980 94788 29036
rect 94844 28980 94892 29036
rect 94948 28980 94958 29036
rect 16930 28812 16940 28868
rect 16996 28812 60732 28868
rect 60788 28812 60798 28868
rect 61730 28812 61740 28868
rect 61796 28812 76076 28868
rect 76132 28812 76142 28868
rect 0 28756 800 28784
rect 0 28700 1708 28756
rect 1764 28700 2492 28756
rect 2548 28700 2558 28756
rect 21970 28700 21980 28756
rect 22036 28700 24220 28756
rect 24276 28700 25452 28756
rect 25508 28700 25518 28756
rect 25890 28700 25900 28756
rect 25956 28700 26852 28756
rect 29586 28700 29596 28756
rect 29652 28700 30268 28756
rect 30324 28700 30334 28756
rect 37314 28700 37324 28756
rect 37380 28700 68348 28756
rect 68404 28700 68414 28756
rect 0 28672 800 28700
rect 26796 28644 26852 28700
rect 2034 28588 2044 28644
rect 2100 28588 7644 28644
rect 7700 28588 7710 28644
rect 24434 28588 24444 28644
rect 24500 28588 26236 28644
rect 26292 28588 26302 28644
rect 26786 28588 26796 28644
rect 26852 28588 28812 28644
rect 28868 28588 28878 28644
rect 30034 28588 30044 28644
rect 30100 28588 30110 28644
rect 44370 28588 44380 28644
rect 44436 28588 45836 28644
rect 45892 28588 45902 28644
rect 60722 28588 60732 28644
rect 60788 28588 61124 28644
rect 61282 28588 61292 28644
rect 61348 28588 62972 28644
rect 63028 28588 63038 28644
rect 63186 28588 63196 28644
rect 63252 28588 63532 28644
rect 63588 28588 64428 28644
rect 64484 28588 64494 28644
rect 64754 28588 64764 28644
rect 64820 28588 68124 28644
rect 68180 28588 68190 28644
rect 70690 28588 70700 28644
rect 70756 28588 71932 28644
rect 71988 28588 72380 28644
rect 72436 28588 72446 28644
rect 72706 28588 72716 28644
rect 72772 28588 96572 28644
rect 96628 28588 97020 28644
rect 97076 28588 97086 28644
rect 30044 28532 30100 28588
rect 61068 28532 61124 28588
rect 28242 28476 28252 28532
rect 28308 28476 29260 28532
rect 29316 28476 32060 28532
rect 32116 28476 32126 28532
rect 55010 28476 55020 28532
rect 55076 28476 56924 28532
rect 56980 28476 56990 28532
rect 61068 28476 61180 28532
rect 61236 28476 61246 28532
rect 29138 28364 29148 28420
rect 29204 28364 30940 28420
rect 30996 28364 31006 28420
rect 61058 28364 61068 28420
rect 61124 28364 61628 28420
rect 61684 28364 61694 28420
rect 62626 28364 62636 28420
rect 62692 28364 63084 28420
rect 63140 28364 63150 28420
rect 76178 28364 76188 28420
rect 76244 28364 77756 28420
rect 77812 28364 77822 28420
rect 8758 28196 8768 28252
rect 8824 28196 8872 28252
rect 8928 28196 8976 28252
rect 9032 28196 9080 28252
rect 9136 28196 9184 28252
rect 9240 28196 9288 28252
rect 9344 28196 9392 28252
rect 9448 28196 9458 28252
rect 17758 28196 17768 28252
rect 17824 28196 17872 28252
rect 17928 28196 17976 28252
rect 18032 28196 18080 28252
rect 18136 28196 18184 28252
rect 18240 28196 18288 28252
rect 18344 28196 18392 28252
rect 18448 28196 18458 28252
rect 26758 28196 26768 28252
rect 26824 28196 26872 28252
rect 26928 28196 26976 28252
rect 27032 28196 27080 28252
rect 27136 28196 27184 28252
rect 27240 28196 27288 28252
rect 27344 28196 27392 28252
rect 27448 28196 27458 28252
rect 35758 28196 35768 28252
rect 35824 28196 35872 28252
rect 35928 28196 35976 28252
rect 36032 28196 36080 28252
rect 36136 28196 36184 28252
rect 36240 28196 36288 28252
rect 36344 28196 36392 28252
rect 36448 28196 36458 28252
rect 44758 28196 44768 28252
rect 44824 28196 44872 28252
rect 44928 28196 44976 28252
rect 45032 28196 45080 28252
rect 45136 28196 45184 28252
rect 45240 28196 45288 28252
rect 45344 28196 45392 28252
rect 45448 28196 45458 28252
rect 53758 28196 53768 28252
rect 53824 28196 53872 28252
rect 53928 28196 53976 28252
rect 54032 28196 54080 28252
rect 54136 28196 54184 28252
rect 54240 28196 54288 28252
rect 54344 28196 54392 28252
rect 54448 28196 54458 28252
rect 62758 28196 62768 28252
rect 62824 28196 62872 28252
rect 62928 28196 62976 28252
rect 63032 28196 63080 28252
rect 63136 28196 63184 28252
rect 63240 28196 63288 28252
rect 63344 28196 63392 28252
rect 63448 28196 63458 28252
rect 71758 28196 71768 28252
rect 71824 28196 71872 28252
rect 71928 28196 71976 28252
rect 72032 28196 72080 28252
rect 72136 28196 72184 28252
rect 72240 28196 72288 28252
rect 72344 28196 72392 28252
rect 72448 28196 72458 28252
rect 80758 28196 80768 28252
rect 80824 28196 80872 28252
rect 80928 28196 80976 28252
rect 81032 28196 81080 28252
rect 81136 28196 81184 28252
rect 81240 28196 81288 28252
rect 81344 28196 81392 28252
rect 81448 28196 81458 28252
rect 89758 28196 89768 28252
rect 89824 28196 89872 28252
rect 89928 28196 89976 28252
rect 90032 28196 90080 28252
rect 90136 28196 90184 28252
rect 90240 28196 90288 28252
rect 90344 28196 90392 28252
rect 90448 28196 90458 28252
rect 32050 28140 32060 28196
rect 32116 28140 33068 28196
rect 33124 28140 33134 28196
rect 99200 28084 100000 28112
rect 5058 28028 5068 28084
rect 5124 28028 6748 28084
rect 6804 28028 6814 28084
rect 13010 28028 13020 28084
rect 13076 28028 13804 28084
rect 13860 28028 17388 28084
rect 17444 28028 61180 28084
rect 61236 28028 61246 28084
rect 62132 28028 96348 28084
rect 96404 28028 96414 28084
rect 97682 28028 97692 28084
rect 97748 28028 100000 28084
rect 6748 27972 6804 28028
rect 62132 27972 62188 28028
rect 99200 28000 100000 28028
rect 6748 27916 9996 27972
rect 10052 27916 10062 27972
rect 34850 27916 34860 27972
rect 34916 27916 35196 27972
rect 35252 27916 37996 27972
rect 38052 27916 38062 27972
rect 51762 27916 51772 27972
rect 51828 27916 52892 27972
rect 52948 27916 53676 27972
rect 53732 27916 53742 27972
rect 57250 27916 57260 27972
rect 57316 27916 60172 27972
rect 60228 27916 62188 27972
rect 65650 27916 65660 27972
rect 65716 27916 66332 27972
rect 66388 27916 66398 27972
rect 70802 27916 70812 27972
rect 70868 27916 71260 27972
rect 71316 27916 73052 27972
rect 73108 27916 73118 27972
rect 12226 27804 12236 27860
rect 12292 27804 15148 27860
rect 15204 27804 15214 27860
rect 24658 27804 24668 27860
rect 24724 27804 25676 27860
rect 25732 27804 25742 27860
rect 48066 27804 48076 27860
rect 48132 27804 49196 27860
rect 49252 27804 49262 27860
rect 75954 27804 75964 27860
rect 76020 27804 76524 27860
rect 76580 27804 76590 27860
rect 46386 27692 46396 27748
rect 46452 27692 46844 27748
rect 46900 27692 52444 27748
rect 52500 27692 52510 27748
rect 57922 27692 57932 27748
rect 57988 27692 73164 27748
rect 73220 27692 73612 27748
rect 73668 27692 73678 27748
rect 0 27636 800 27664
rect 0 27580 1708 27636
rect 1764 27580 1774 27636
rect 28802 27580 28812 27636
rect 28868 27580 61740 27636
rect 61796 27580 61806 27636
rect 63634 27580 63644 27636
rect 63700 27580 65660 27636
rect 65716 27580 65726 27636
rect 77522 27580 77532 27636
rect 77588 27580 79660 27636
rect 79716 27580 84028 27636
rect 84084 27580 84094 27636
rect 0 27552 800 27580
rect 4258 27412 4268 27468
rect 4324 27412 4372 27468
rect 4428 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4788 27468
rect 4844 27412 4892 27468
rect 4948 27412 4958 27468
rect 13258 27412 13268 27468
rect 13324 27412 13372 27468
rect 13428 27412 13476 27468
rect 13532 27412 13580 27468
rect 13636 27412 13684 27468
rect 13740 27412 13788 27468
rect 13844 27412 13892 27468
rect 13948 27412 13958 27468
rect 22258 27412 22268 27468
rect 22324 27412 22372 27468
rect 22428 27412 22476 27468
rect 22532 27412 22580 27468
rect 22636 27412 22684 27468
rect 22740 27412 22788 27468
rect 22844 27412 22892 27468
rect 22948 27412 22958 27468
rect 31258 27412 31268 27468
rect 31324 27412 31372 27468
rect 31428 27412 31476 27468
rect 31532 27412 31580 27468
rect 31636 27412 31684 27468
rect 31740 27412 31788 27468
rect 31844 27412 31892 27468
rect 31948 27412 31958 27468
rect 40258 27412 40268 27468
rect 40324 27412 40372 27468
rect 40428 27412 40476 27468
rect 40532 27412 40580 27468
rect 40636 27412 40684 27468
rect 40740 27412 40788 27468
rect 40844 27412 40892 27468
rect 40948 27412 40958 27468
rect 49258 27412 49268 27468
rect 49324 27412 49372 27468
rect 49428 27412 49476 27468
rect 49532 27412 49580 27468
rect 49636 27412 49684 27468
rect 49740 27412 49788 27468
rect 49844 27412 49892 27468
rect 49948 27412 49958 27468
rect 58258 27412 58268 27468
rect 58324 27412 58372 27468
rect 58428 27412 58476 27468
rect 58532 27412 58580 27468
rect 58636 27412 58684 27468
rect 58740 27412 58788 27468
rect 58844 27412 58892 27468
rect 58948 27412 58958 27468
rect 67258 27412 67268 27468
rect 67324 27412 67372 27468
rect 67428 27412 67476 27468
rect 67532 27412 67580 27468
rect 67636 27412 67684 27468
rect 67740 27412 67788 27468
rect 67844 27412 67892 27468
rect 67948 27412 67958 27468
rect 76258 27412 76268 27468
rect 76324 27412 76372 27468
rect 76428 27412 76476 27468
rect 76532 27412 76580 27468
rect 76636 27412 76684 27468
rect 76740 27412 76788 27468
rect 76844 27412 76892 27468
rect 76948 27412 76958 27468
rect 85258 27412 85268 27468
rect 85324 27412 85372 27468
rect 85428 27412 85476 27468
rect 85532 27412 85580 27468
rect 85636 27412 85684 27468
rect 85740 27412 85788 27468
rect 85844 27412 85892 27468
rect 85948 27412 85958 27468
rect 94258 27412 94268 27468
rect 94324 27412 94372 27468
rect 94428 27412 94476 27468
rect 94532 27412 94580 27468
rect 94636 27412 94684 27468
rect 94740 27412 94788 27468
rect 94844 27412 94892 27468
rect 94948 27412 94958 27468
rect 5618 27244 5628 27300
rect 5684 27244 29932 27300
rect 29988 27244 30492 27300
rect 30548 27244 30558 27300
rect 32050 27244 32060 27300
rect 32116 27244 32620 27300
rect 32676 27244 59948 27300
rect 60004 27244 60620 27300
rect 60676 27244 60686 27300
rect 66322 27244 66332 27300
rect 66388 27244 67228 27300
rect 67284 27244 67294 27300
rect 67554 27244 67564 27300
rect 67620 27244 96572 27300
rect 96628 27244 96638 27300
rect 15138 27132 15148 27188
rect 15204 27132 20748 27188
rect 20804 27132 21980 27188
rect 22036 27132 22046 27188
rect 29474 27132 29484 27188
rect 29540 27132 30380 27188
rect 30436 27132 30446 27188
rect 37538 27132 37548 27188
rect 37604 27132 38108 27188
rect 38164 27132 38780 27188
rect 38836 27132 54572 27188
rect 54628 27132 54638 27188
rect 60844 27132 72604 27188
rect 72660 27132 72670 27188
rect 75954 27132 75964 27188
rect 76020 27132 76412 27188
rect 76468 27132 76478 27188
rect 60844 27076 60900 27132
rect 1698 27020 1708 27076
rect 1764 27020 2492 27076
rect 2548 27020 2558 27076
rect 21746 27020 21756 27076
rect 21812 27020 23100 27076
rect 23156 27020 23166 27076
rect 31154 27020 31164 27076
rect 31220 27020 32060 27076
rect 32116 27020 32126 27076
rect 56914 27020 56924 27076
rect 56980 27020 57820 27076
rect 57876 27020 57886 27076
rect 60834 27020 60844 27076
rect 60900 27020 60910 27076
rect 62738 27020 62748 27076
rect 62804 27020 63868 27076
rect 63924 27020 63934 27076
rect 16594 26908 16604 26964
rect 16660 26908 17612 26964
rect 17668 26908 17678 26964
rect 29698 26908 29708 26964
rect 29764 26908 30156 26964
rect 30212 26908 35196 26964
rect 35252 26908 35262 26964
rect 60498 26908 60508 26964
rect 60564 26908 60574 26964
rect 61730 26908 61740 26964
rect 61796 26908 62300 26964
rect 62356 26908 62366 26964
rect 73042 26908 73052 26964
rect 73108 26908 73892 26964
rect 60508 26852 60564 26908
rect 73836 26852 73892 26908
rect 12002 26796 12012 26852
rect 12068 26796 36988 26852
rect 37044 26796 37054 26852
rect 53554 26796 53564 26852
rect 53620 26796 57036 26852
rect 57092 26796 57102 26852
rect 59938 26796 59948 26852
rect 60004 26796 61068 26852
rect 61124 26796 61134 26852
rect 61394 26796 61404 26852
rect 61460 26796 67116 26852
rect 67172 26796 67182 26852
rect 73836 26796 74508 26852
rect 74564 26796 74574 26852
rect 56018 26684 56028 26740
rect 56084 26684 58044 26740
rect 58100 26684 59612 26740
rect 59668 26684 62300 26740
rect 62356 26684 62366 26740
rect 66770 26684 66780 26740
rect 66836 26684 68908 26740
rect 68964 26684 70476 26740
rect 70532 26684 70542 26740
rect 8758 26628 8768 26684
rect 8824 26628 8872 26684
rect 8928 26628 8976 26684
rect 9032 26628 9080 26684
rect 9136 26628 9184 26684
rect 9240 26628 9288 26684
rect 9344 26628 9392 26684
rect 9448 26628 9458 26684
rect 17758 26628 17768 26684
rect 17824 26628 17872 26684
rect 17928 26628 17976 26684
rect 18032 26628 18080 26684
rect 18136 26628 18184 26684
rect 18240 26628 18288 26684
rect 18344 26628 18392 26684
rect 18448 26628 18458 26684
rect 26758 26628 26768 26684
rect 26824 26628 26872 26684
rect 26928 26628 26976 26684
rect 27032 26628 27080 26684
rect 27136 26628 27184 26684
rect 27240 26628 27288 26684
rect 27344 26628 27392 26684
rect 27448 26628 27458 26684
rect 35758 26628 35768 26684
rect 35824 26628 35872 26684
rect 35928 26628 35976 26684
rect 36032 26628 36080 26684
rect 36136 26628 36184 26684
rect 36240 26628 36288 26684
rect 36344 26628 36392 26684
rect 36448 26628 36458 26684
rect 44758 26628 44768 26684
rect 44824 26628 44872 26684
rect 44928 26628 44976 26684
rect 45032 26628 45080 26684
rect 45136 26628 45184 26684
rect 45240 26628 45288 26684
rect 45344 26628 45392 26684
rect 45448 26628 45458 26684
rect 53758 26628 53768 26684
rect 53824 26628 53872 26684
rect 53928 26628 53976 26684
rect 54032 26628 54080 26684
rect 54136 26628 54184 26684
rect 54240 26628 54288 26684
rect 54344 26628 54392 26684
rect 54448 26628 54458 26684
rect 62758 26628 62768 26684
rect 62824 26628 62872 26684
rect 62928 26628 62976 26684
rect 63032 26628 63080 26684
rect 63136 26628 63184 26684
rect 63240 26628 63288 26684
rect 63344 26628 63392 26684
rect 63448 26628 63458 26684
rect 71758 26628 71768 26684
rect 71824 26628 71872 26684
rect 71928 26628 71976 26684
rect 72032 26628 72080 26684
rect 72136 26628 72184 26684
rect 72240 26628 72288 26684
rect 72344 26628 72392 26684
rect 72448 26628 72458 26684
rect 80758 26628 80768 26684
rect 80824 26628 80872 26684
rect 80928 26628 80976 26684
rect 81032 26628 81080 26684
rect 81136 26628 81184 26684
rect 81240 26628 81288 26684
rect 81344 26628 81392 26684
rect 81448 26628 81458 26684
rect 89758 26628 89768 26684
rect 89824 26628 89872 26684
rect 89928 26628 89976 26684
rect 90032 26628 90080 26684
rect 90136 26628 90184 26684
rect 90240 26628 90288 26684
rect 90344 26628 90392 26684
rect 90448 26628 90458 26684
rect 0 26516 800 26544
rect 0 26460 2604 26516
rect 2660 26460 2670 26516
rect 17602 26460 17612 26516
rect 17668 26460 19180 26516
rect 19236 26460 19628 26516
rect 19684 26460 22316 26516
rect 22372 26460 22382 26516
rect 23090 26460 23100 26516
rect 23156 26460 59612 26516
rect 59668 26460 60060 26516
rect 60116 26460 60126 26516
rect 0 26432 800 26460
rect 52882 26348 52892 26404
rect 52948 26348 53452 26404
rect 53508 26348 53788 26404
rect 53844 26348 53854 26404
rect 58482 26348 58492 26404
rect 58548 26348 59948 26404
rect 60004 26348 60014 26404
rect 67172 26348 67340 26404
rect 67396 26348 68124 26404
rect 68180 26348 72716 26404
rect 72772 26348 73500 26404
rect 73556 26348 76524 26404
rect 76580 26348 77084 26404
rect 77140 26348 77150 26404
rect 84242 26348 84252 26404
rect 84308 26348 96908 26404
rect 96964 26348 96974 26404
rect 26450 26236 26460 26292
rect 26516 26236 27244 26292
rect 27300 26236 27310 26292
rect 48402 26236 48412 26292
rect 48468 26236 50428 26292
rect 50484 26236 50494 26292
rect 57026 26236 57036 26292
rect 57092 26236 57932 26292
rect 57988 26236 57998 26292
rect 62290 26236 62300 26292
rect 62356 26236 64540 26292
rect 64596 26236 65436 26292
rect 65492 26236 65502 26292
rect 67106 26124 67116 26180
rect 67172 26124 67228 26348
rect 99200 26292 100000 26320
rect 73154 26236 73164 26292
rect 73220 26236 74172 26292
rect 74228 26236 74238 26292
rect 75740 26236 77644 26292
rect 77700 26236 77710 26292
rect 97682 26236 97692 26292
rect 97748 26236 100000 26292
rect 75740 26180 75796 26236
rect 99200 26208 100000 26236
rect 74498 26124 74508 26180
rect 74564 26124 75740 26180
rect 75796 26124 75806 26180
rect 75954 26124 75964 26180
rect 76020 26124 77980 26180
rect 78036 26124 78876 26180
rect 78932 26124 78942 26180
rect 60050 26012 60060 26068
rect 60116 26012 76076 26068
rect 76132 26012 76142 26068
rect 4258 25844 4268 25900
rect 4324 25844 4372 25900
rect 4428 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4788 25900
rect 4844 25844 4892 25900
rect 4948 25844 4958 25900
rect 13258 25844 13268 25900
rect 13324 25844 13372 25900
rect 13428 25844 13476 25900
rect 13532 25844 13580 25900
rect 13636 25844 13684 25900
rect 13740 25844 13788 25900
rect 13844 25844 13892 25900
rect 13948 25844 13958 25900
rect 22258 25844 22268 25900
rect 22324 25844 22372 25900
rect 22428 25844 22476 25900
rect 22532 25844 22580 25900
rect 22636 25844 22684 25900
rect 22740 25844 22788 25900
rect 22844 25844 22892 25900
rect 22948 25844 22958 25900
rect 31258 25844 31268 25900
rect 31324 25844 31372 25900
rect 31428 25844 31476 25900
rect 31532 25844 31580 25900
rect 31636 25844 31684 25900
rect 31740 25844 31788 25900
rect 31844 25844 31892 25900
rect 31948 25844 31958 25900
rect 40258 25844 40268 25900
rect 40324 25844 40372 25900
rect 40428 25844 40476 25900
rect 40532 25844 40580 25900
rect 40636 25844 40684 25900
rect 40740 25844 40788 25900
rect 40844 25844 40892 25900
rect 40948 25844 40958 25900
rect 49258 25844 49268 25900
rect 49324 25844 49372 25900
rect 49428 25844 49476 25900
rect 49532 25844 49580 25900
rect 49636 25844 49684 25900
rect 49740 25844 49788 25900
rect 49844 25844 49892 25900
rect 49948 25844 49958 25900
rect 58258 25844 58268 25900
rect 58324 25844 58372 25900
rect 58428 25844 58476 25900
rect 58532 25844 58580 25900
rect 58636 25844 58684 25900
rect 58740 25844 58788 25900
rect 58844 25844 58892 25900
rect 58948 25844 58958 25900
rect 67258 25844 67268 25900
rect 67324 25844 67372 25900
rect 67428 25844 67476 25900
rect 67532 25844 67580 25900
rect 67636 25844 67684 25900
rect 67740 25844 67788 25900
rect 67844 25844 67892 25900
rect 67948 25844 67958 25900
rect 76258 25844 76268 25900
rect 76324 25844 76372 25900
rect 76428 25844 76476 25900
rect 76532 25844 76580 25900
rect 76636 25844 76684 25900
rect 76740 25844 76788 25900
rect 76844 25844 76892 25900
rect 76948 25844 76958 25900
rect 85258 25844 85268 25900
rect 85324 25844 85372 25900
rect 85428 25844 85476 25900
rect 85532 25844 85580 25900
rect 85636 25844 85684 25900
rect 85740 25844 85788 25900
rect 85844 25844 85892 25900
rect 85948 25844 85958 25900
rect 94258 25844 94268 25900
rect 94324 25844 94372 25900
rect 94428 25844 94476 25900
rect 94532 25844 94580 25900
rect 94636 25844 94684 25900
rect 94740 25844 94788 25900
rect 94844 25844 94892 25900
rect 94948 25844 94958 25900
rect 2034 25676 2044 25732
rect 2100 25676 16156 25732
rect 16212 25676 16222 25732
rect 5842 25564 5852 25620
rect 5908 25564 25676 25620
rect 25732 25564 26124 25620
rect 26180 25564 26190 25620
rect 57138 25564 57148 25620
rect 57204 25564 58044 25620
rect 58100 25564 58110 25620
rect 65314 25564 65324 25620
rect 65380 25564 65772 25620
rect 65828 25564 65838 25620
rect 78866 25564 78876 25620
rect 2146 25452 2156 25508
rect 2212 25452 6076 25508
rect 6132 25452 6142 25508
rect 25330 25452 25340 25508
rect 25396 25452 26236 25508
rect 26292 25452 26302 25508
rect 26898 25452 26908 25508
rect 26964 25452 28252 25508
rect 28308 25452 28318 25508
rect 43138 25452 43148 25508
rect 43204 25452 54572 25508
rect 54628 25452 54638 25508
rect 62962 25452 62972 25508
rect 63028 25452 64988 25508
rect 65044 25452 65054 25508
rect 77410 25452 77420 25508
rect 77476 25452 78764 25508
rect 78820 25452 78830 25508
rect 0 25396 800 25424
rect 78932 25396 78988 25620
rect 0 25340 1708 25396
rect 1764 25340 2492 25396
rect 2548 25340 2558 25396
rect 11106 25340 11116 25396
rect 11172 25340 11564 25396
rect 11620 25340 12348 25396
rect 12404 25340 12414 25396
rect 33058 25340 33068 25396
rect 33124 25340 34188 25396
rect 34244 25340 34254 25396
rect 34850 25340 34860 25396
rect 34916 25340 43260 25396
rect 43316 25340 43326 25396
rect 43810 25340 43820 25396
rect 43876 25340 45276 25396
rect 45332 25340 45342 25396
rect 75058 25340 75068 25396
rect 75124 25340 75964 25396
rect 76020 25340 76030 25396
rect 78932 25340 81116 25396
rect 81172 25340 81182 25396
rect 0 25312 800 25340
rect 11330 25228 11340 25284
rect 11396 25228 12684 25284
rect 12740 25228 15148 25284
rect 15204 25228 15214 25284
rect 26450 25228 26460 25284
rect 26516 25228 27692 25284
rect 27748 25228 27758 25284
rect 34066 25228 34076 25284
rect 34132 25228 34972 25284
rect 35028 25228 42700 25284
rect 42756 25228 42766 25284
rect 44268 25228 47628 25284
rect 47684 25228 47694 25284
rect 62514 25228 62524 25284
rect 62580 25228 63308 25284
rect 63364 25228 67116 25284
rect 67172 25228 67182 25284
rect 74498 25228 74508 25284
rect 74564 25228 74956 25284
rect 75012 25228 75022 25284
rect 44268 25172 44324 25228
rect 43922 25116 43932 25172
rect 43988 25116 44268 25172
rect 44324 25116 44334 25172
rect 8758 25060 8768 25116
rect 8824 25060 8872 25116
rect 8928 25060 8976 25116
rect 9032 25060 9080 25116
rect 9136 25060 9184 25116
rect 9240 25060 9288 25116
rect 9344 25060 9392 25116
rect 9448 25060 9458 25116
rect 17758 25060 17768 25116
rect 17824 25060 17872 25116
rect 17928 25060 17976 25116
rect 18032 25060 18080 25116
rect 18136 25060 18184 25116
rect 18240 25060 18288 25116
rect 18344 25060 18392 25116
rect 18448 25060 18458 25116
rect 26758 25060 26768 25116
rect 26824 25060 26872 25116
rect 26928 25060 26976 25116
rect 27032 25060 27080 25116
rect 27136 25060 27184 25116
rect 27240 25060 27288 25116
rect 27344 25060 27392 25116
rect 27448 25060 27458 25116
rect 35758 25060 35768 25116
rect 35824 25060 35872 25116
rect 35928 25060 35976 25116
rect 36032 25060 36080 25116
rect 36136 25060 36184 25116
rect 36240 25060 36288 25116
rect 36344 25060 36392 25116
rect 36448 25060 36458 25116
rect 44758 25060 44768 25116
rect 44824 25060 44872 25116
rect 44928 25060 44976 25116
rect 45032 25060 45080 25116
rect 45136 25060 45184 25116
rect 45240 25060 45288 25116
rect 45344 25060 45392 25116
rect 45448 25060 45458 25116
rect 53758 25060 53768 25116
rect 53824 25060 53872 25116
rect 53928 25060 53976 25116
rect 54032 25060 54080 25116
rect 54136 25060 54184 25116
rect 54240 25060 54288 25116
rect 54344 25060 54392 25116
rect 54448 25060 54458 25116
rect 62758 25060 62768 25116
rect 62824 25060 62872 25116
rect 62928 25060 62976 25116
rect 63032 25060 63080 25116
rect 63136 25060 63184 25116
rect 63240 25060 63288 25116
rect 63344 25060 63392 25116
rect 63448 25060 63458 25116
rect 71758 25060 71768 25116
rect 71824 25060 71872 25116
rect 71928 25060 71976 25116
rect 72032 25060 72080 25116
rect 72136 25060 72184 25116
rect 72240 25060 72288 25116
rect 72344 25060 72392 25116
rect 72448 25060 72458 25116
rect 80758 25060 80768 25116
rect 80824 25060 80872 25116
rect 80928 25060 80976 25116
rect 81032 25060 81080 25116
rect 81136 25060 81184 25116
rect 81240 25060 81288 25116
rect 81344 25060 81392 25116
rect 81448 25060 81458 25116
rect 89758 25060 89768 25116
rect 89824 25060 89872 25116
rect 89928 25060 89976 25116
rect 90032 25060 90080 25116
rect 90136 25060 90184 25116
rect 90240 25060 90288 25116
rect 90344 25060 90392 25116
rect 90448 25060 90458 25116
rect 30482 25004 30492 25060
rect 30548 25004 32060 25060
rect 32116 25004 32126 25060
rect 5282 24892 5292 24948
rect 5348 24892 10556 24948
rect 10612 24892 10622 24948
rect 11890 24892 11900 24948
rect 11956 24892 13244 24948
rect 13300 24892 13310 24948
rect 28578 24892 28588 24948
rect 28644 24892 30156 24948
rect 30212 24892 60172 24948
rect 60228 24892 60620 24948
rect 60676 24892 60686 24948
rect 66322 24892 66332 24948
rect 66388 24892 67004 24948
rect 67060 24892 67070 24948
rect 68786 24892 68796 24948
rect 68852 24892 70252 24948
rect 70308 24892 71148 24948
rect 71204 24892 71214 24948
rect 78082 24892 78092 24948
rect 78148 24892 81900 24948
rect 81956 24892 83132 24948
rect 83188 24892 83198 24948
rect 4722 24780 4732 24836
rect 4788 24780 5068 24836
rect 5124 24780 5740 24836
rect 5796 24780 6076 24836
rect 6132 24780 8428 24836
rect 8484 24780 8494 24836
rect 29362 24780 29372 24836
rect 29428 24780 30492 24836
rect 30548 24780 30558 24836
rect 35186 24780 35196 24836
rect 35252 24780 35868 24836
rect 35924 24780 35934 24836
rect 41570 24780 41580 24836
rect 41636 24780 43932 24836
rect 43988 24780 43998 24836
rect 74386 24780 74396 24836
rect 74452 24780 75740 24836
rect 75796 24780 75806 24836
rect 33842 24668 33852 24724
rect 33908 24668 34748 24724
rect 34804 24668 36652 24724
rect 36708 24668 59388 24724
rect 59444 24668 59454 24724
rect 99200 24500 100000 24528
rect 39218 24444 39228 24500
rect 39284 24444 40124 24500
rect 40180 24444 40190 24500
rect 60610 24444 60620 24500
rect 60676 24444 62076 24500
rect 62132 24444 62142 24500
rect 98018 24444 98028 24500
rect 98084 24444 100000 24500
rect 99200 24416 100000 24444
rect 0 24276 800 24304
rect 4258 24276 4268 24332
rect 4324 24276 4372 24332
rect 4428 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4788 24332
rect 4844 24276 4892 24332
rect 4948 24276 4958 24332
rect 13258 24276 13268 24332
rect 13324 24276 13372 24332
rect 13428 24276 13476 24332
rect 13532 24276 13580 24332
rect 13636 24276 13684 24332
rect 13740 24276 13788 24332
rect 13844 24276 13892 24332
rect 13948 24276 13958 24332
rect 22258 24276 22268 24332
rect 22324 24276 22372 24332
rect 22428 24276 22476 24332
rect 22532 24276 22580 24332
rect 22636 24276 22684 24332
rect 22740 24276 22788 24332
rect 22844 24276 22892 24332
rect 22948 24276 22958 24332
rect 31258 24276 31268 24332
rect 31324 24276 31372 24332
rect 31428 24276 31476 24332
rect 31532 24276 31580 24332
rect 31636 24276 31684 24332
rect 31740 24276 31788 24332
rect 31844 24276 31892 24332
rect 31948 24276 31958 24332
rect 40258 24276 40268 24332
rect 40324 24276 40372 24332
rect 40428 24276 40476 24332
rect 40532 24276 40580 24332
rect 40636 24276 40684 24332
rect 40740 24276 40788 24332
rect 40844 24276 40892 24332
rect 40948 24276 40958 24332
rect 49258 24276 49268 24332
rect 49324 24276 49372 24332
rect 49428 24276 49476 24332
rect 49532 24276 49580 24332
rect 49636 24276 49684 24332
rect 49740 24276 49788 24332
rect 49844 24276 49892 24332
rect 49948 24276 49958 24332
rect 58258 24276 58268 24332
rect 58324 24276 58372 24332
rect 58428 24276 58476 24332
rect 58532 24276 58580 24332
rect 58636 24276 58684 24332
rect 58740 24276 58788 24332
rect 58844 24276 58892 24332
rect 58948 24276 58958 24332
rect 67258 24276 67268 24332
rect 67324 24276 67372 24332
rect 67428 24276 67476 24332
rect 67532 24276 67580 24332
rect 67636 24276 67684 24332
rect 67740 24276 67788 24332
rect 67844 24276 67892 24332
rect 67948 24276 67958 24332
rect 76258 24276 76268 24332
rect 76324 24276 76372 24332
rect 76428 24276 76476 24332
rect 76532 24276 76580 24332
rect 76636 24276 76684 24332
rect 76740 24276 76788 24332
rect 76844 24276 76892 24332
rect 76948 24276 76958 24332
rect 85258 24276 85268 24332
rect 85324 24276 85372 24332
rect 85428 24276 85476 24332
rect 85532 24276 85580 24332
rect 85636 24276 85684 24332
rect 85740 24276 85788 24332
rect 85844 24276 85892 24332
rect 85948 24276 85958 24332
rect 94258 24276 94268 24332
rect 94324 24276 94372 24332
rect 94428 24276 94476 24332
rect 94532 24276 94580 24332
rect 94636 24276 94684 24332
rect 94740 24276 94788 24332
rect 94844 24276 94892 24332
rect 94948 24276 94958 24332
rect 0 24220 1708 24276
rect 1764 24220 3612 24276
rect 3668 24220 3678 24276
rect 0 24192 800 24220
rect 10770 24108 10780 24164
rect 10836 24108 38108 24164
rect 38164 24108 38174 24164
rect 15138 23996 15148 24052
rect 15204 23996 16380 24052
rect 16436 23996 61180 24052
rect 61236 23996 61246 24052
rect 75730 23884 75740 23940
rect 75796 23884 76300 23940
rect 76356 23884 76366 23940
rect 9650 23772 9660 23828
rect 9716 23772 32620 23828
rect 32676 23772 33068 23828
rect 33124 23772 33134 23828
rect 59714 23772 59724 23828
rect 59780 23772 60508 23828
rect 60564 23772 61068 23828
rect 61124 23772 61134 23828
rect 64642 23772 64652 23828
rect 64708 23772 65548 23828
rect 65604 23772 65614 23828
rect 12450 23660 12460 23716
rect 12516 23660 15596 23716
rect 15652 23660 15662 23716
rect 19282 23660 19292 23716
rect 19348 23660 21420 23716
rect 21476 23660 21486 23716
rect 21634 23660 21644 23716
rect 21700 23660 22540 23716
rect 22596 23660 22606 23716
rect 40226 23660 40236 23716
rect 40292 23660 42364 23716
rect 42420 23660 60284 23716
rect 60340 23660 60350 23716
rect 61394 23660 61404 23716
rect 61460 23660 73500 23716
rect 73556 23660 73566 23716
rect 38770 23548 38780 23604
rect 38836 23548 40012 23604
rect 40068 23548 41580 23604
rect 41636 23548 41646 23604
rect 65202 23548 65212 23604
rect 65268 23548 66332 23604
rect 66388 23548 66398 23604
rect 8758 23492 8768 23548
rect 8824 23492 8872 23548
rect 8928 23492 8976 23548
rect 9032 23492 9080 23548
rect 9136 23492 9184 23548
rect 9240 23492 9288 23548
rect 9344 23492 9392 23548
rect 9448 23492 9458 23548
rect 17758 23492 17768 23548
rect 17824 23492 17872 23548
rect 17928 23492 17976 23548
rect 18032 23492 18080 23548
rect 18136 23492 18184 23548
rect 18240 23492 18288 23548
rect 18344 23492 18392 23548
rect 18448 23492 18458 23548
rect 26758 23492 26768 23548
rect 26824 23492 26872 23548
rect 26928 23492 26976 23548
rect 27032 23492 27080 23548
rect 27136 23492 27184 23548
rect 27240 23492 27288 23548
rect 27344 23492 27392 23548
rect 27448 23492 27458 23548
rect 35758 23492 35768 23548
rect 35824 23492 35872 23548
rect 35928 23492 35976 23548
rect 36032 23492 36080 23548
rect 36136 23492 36184 23548
rect 36240 23492 36288 23548
rect 36344 23492 36392 23548
rect 36448 23492 36458 23548
rect 44758 23492 44768 23548
rect 44824 23492 44872 23548
rect 44928 23492 44976 23548
rect 45032 23492 45080 23548
rect 45136 23492 45184 23548
rect 45240 23492 45288 23548
rect 45344 23492 45392 23548
rect 45448 23492 45458 23548
rect 53758 23492 53768 23548
rect 53824 23492 53872 23548
rect 53928 23492 53976 23548
rect 54032 23492 54080 23548
rect 54136 23492 54184 23548
rect 54240 23492 54288 23548
rect 54344 23492 54392 23548
rect 54448 23492 54458 23548
rect 62758 23492 62768 23548
rect 62824 23492 62872 23548
rect 62928 23492 62976 23548
rect 63032 23492 63080 23548
rect 63136 23492 63184 23548
rect 63240 23492 63288 23548
rect 63344 23492 63392 23548
rect 63448 23492 63458 23548
rect 71758 23492 71768 23548
rect 71824 23492 71872 23548
rect 71928 23492 71976 23548
rect 72032 23492 72080 23548
rect 72136 23492 72184 23548
rect 72240 23492 72288 23548
rect 72344 23492 72392 23548
rect 72448 23492 72458 23548
rect 80758 23492 80768 23548
rect 80824 23492 80872 23548
rect 80928 23492 80976 23548
rect 81032 23492 81080 23548
rect 81136 23492 81184 23548
rect 81240 23492 81288 23548
rect 81344 23492 81392 23548
rect 81448 23492 81458 23548
rect 89758 23492 89768 23548
rect 89824 23492 89872 23548
rect 89928 23492 89976 23548
rect 90032 23492 90080 23548
rect 90136 23492 90184 23548
rect 90240 23492 90288 23548
rect 90344 23492 90392 23548
rect 90448 23492 90458 23548
rect 2370 23436 2380 23492
rect 2436 23436 3164 23492
rect 3220 23436 3230 23492
rect 2034 23324 2044 23380
rect 2100 23324 26348 23380
rect 26404 23324 27132 23380
rect 27188 23324 27198 23380
rect 32274 23324 32284 23380
rect 32340 23324 32620 23380
rect 32676 23324 33628 23380
rect 33684 23324 37996 23380
rect 38052 23324 38062 23380
rect 60722 23324 60732 23380
rect 60788 23324 60798 23380
rect 65986 23324 65996 23380
rect 66052 23324 67004 23380
rect 67060 23324 69468 23380
rect 69524 23324 69804 23380
rect 69860 23324 69870 23380
rect 76626 23324 76636 23380
rect 76692 23324 96572 23380
rect 96628 23324 96638 23380
rect 60732 23268 60788 23324
rect 5282 23212 5292 23268
rect 5348 23212 10220 23268
rect 10276 23212 10286 23268
rect 19618 23212 19628 23268
rect 19684 23212 20300 23268
rect 20356 23212 21756 23268
rect 21812 23212 23436 23268
rect 23492 23212 23502 23268
rect 60732 23212 67228 23268
rect 72146 23212 72156 23268
rect 72212 23212 72940 23268
rect 72996 23212 73006 23268
rect 73714 23212 73724 23268
rect 73780 23212 74508 23268
rect 74564 23212 74574 23268
rect 77746 23212 77756 23268
rect 77812 23212 77822 23268
rect 82562 23212 82572 23268
rect 82628 23212 85036 23268
rect 85092 23212 85708 23268
rect 85764 23212 85774 23268
rect 0 23156 800 23184
rect 67172 23156 67228 23212
rect 77756 23156 77812 23212
rect 0 23100 2156 23156
rect 2212 23100 2222 23156
rect 22194 23100 22204 23156
rect 22260 23100 23100 23156
rect 23156 23100 24220 23156
rect 24276 23100 45164 23156
rect 45220 23100 46060 23156
rect 46116 23100 46126 23156
rect 62962 23100 62972 23156
rect 63028 23100 64204 23156
rect 64260 23100 64270 23156
rect 67172 23100 77812 23156
rect 78418 23100 78428 23156
rect 78484 23100 80220 23156
rect 80276 23100 80286 23156
rect 82114 23100 82124 23156
rect 82180 23100 83356 23156
rect 83412 23100 83422 23156
rect 0 23072 800 23100
rect 30258 22876 30268 22932
rect 30324 22876 38668 22932
rect 38724 22876 38734 22932
rect 69346 22876 69356 22932
rect 69412 22876 70588 22932
rect 70644 22876 70654 22932
rect 4258 22708 4268 22764
rect 4324 22708 4372 22764
rect 4428 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4788 22764
rect 4844 22708 4892 22764
rect 4948 22708 4958 22764
rect 13258 22708 13268 22764
rect 13324 22708 13372 22764
rect 13428 22708 13476 22764
rect 13532 22708 13580 22764
rect 13636 22708 13684 22764
rect 13740 22708 13788 22764
rect 13844 22708 13892 22764
rect 13948 22708 13958 22764
rect 22258 22708 22268 22764
rect 22324 22708 22372 22764
rect 22428 22708 22476 22764
rect 22532 22708 22580 22764
rect 22636 22708 22684 22764
rect 22740 22708 22788 22764
rect 22844 22708 22892 22764
rect 22948 22708 22958 22764
rect 31258 22708 31268 22764
rect 31324 22708 31372 22764
rect 31428 22708 31476 22764
rect 31532 22708 31580 22764
rect 31636 22708 31684 22764
rect 31740 22708 31788 22764
rect 31844 22708 31892 22764
rect 31948 22708 31958 22764
rect 40258 22708 40268 22764
rect 40324 22708 40372 22764
rect 40428 22708 40476 22764
rect 40532 22708 40580 22764
rect 40636 22708 40684 22764
rect 40740 22708 40788 22764
rect 40844 22708 40892 22764
rect 40948 22708 40958 22764
rect 49258 22708 49268 22764
rect 49324 22708 49372 22764
rect 49428 22708 49476 22764
rect 49532 22708 49580 22764
rect 49636 22708 49684 22764
rect 49740 22708 49788 22764
rect 49844 22708 49892 22764
rect 49948 22708 49958 22764
rect 58258 22708 58268 22764
rect 58324 22708 58372 22764
rect 58428 22708 58476 22764
rect 58532 22708 58580 22764
rect 58636 22708 58684 22764
rect 58740 22708 58788 22764
rect 58844 22708 58892 22764
rect 58948 22708 58958 22764
rect 67258 22708 67268 22764
rect 67324 22708 67372 22764
rect 67428 22708 67476 22764
rect 67532 22708 67580 22764
rect 67636 22708 67684 22764
rect 67740 22708 67788 22764
rect 67844 22708 67892 22764
rect 67948 22708 67958 22764
rect 76258 22708 76268 22764
rect 76324 22708 76372 22764
rect 76428 22708 76476 22764
rect 76532 22708 76580 22764
rect 76636 22708 76684 22764
rect 76740 22708 76788 22764
rect 76844 22708 76892 22764
rect 76948 22708 76958 22764
rect 85258 22708 85268 22764
rect 85324 22708 85372 22764
rect 85428 22708 85476 22764
rect 85532 22708 85580 22764
rect 85636 22708 85684 22764
rect 85740 22708 85788 22764
rect 85844 22708 85892 22764
rect 85948 22708 85958 22764
rect 94258 22708 94268 22764
rect 94324 22708 94372 22764
rect 94428 22708 94476 22764
rect 94532 22708 94580 22764
rect 94636 22708 94684 22764
rect 94740 22708 94788 22764
rect 94844 22708 94892 22764
rect 94948 22708 94958 22764
rect 99200 22708 100000 22736
rect 98018 22652 98028 22708
rect 98084 22652 100000 22708
rect 99200 22624 100000 22652
rect 46274 22540 46284 22596
rect 46340 22540 81452 22596
rect 81508 22540 81518 22596
rect 8418 22428 8428 22484
rect 8484 22428 9548 22484
rect 9604 22428 9614 22484
rect 38098 22428 38108 22484
rect 38164 22428 38556 22484
rect 38612 22428 38622 22484
rect 68562 22428 68572 22484
rect 68628 22428 69916 22484
rect 69972 22428 73724 22484
rect 73780 22428 73790 22484
rect 75058 22428 75068 22484
rect 75124 22428 75628 22484
rect 75684 22428 76300 22484
rect 76356 22428 77756 22484
rect 77812 22428 77822 22484
rect 2818 22316 2828 22372
rect 2884 22316 6076 22372
rect 6132 22316 6142 22372
rect 33618 22316 33628 22372
rect 33684 22316 34636 22372
rect 34692 22316 34702 22372
rect 60050 22316 60060 22372
rect 60116 22316 68348 22372
rect 68404 22316 68414 22372
rect 68572 22260 68628 22428
rect 75394 22316 75404 22372
rect 75460 22316 82572 22372
rect 82628 22316 82638 22372
rect 9874 22204 9884 22260
rect 9940 22204 10780 22260
rect 10836 22204 10846 22260
rect 28578 22204 28588 22260
rect 28644 22204 29708 22260
rect 29764 22204 29774 22260
rect 67106 22204 67116 22260
rect 67172 22204 68628 22260
rect 82674 22204 82684 22260
rect 82740 22204 84588 22260
rect 84644 22204 84654 22260
rect 84802 22204 84812 22260
rect 84868 22204 86492 22260
rect 86548 22204 86558 22260
rect 11666 22092 11676 22148
rect 11732 22092 14588 22148
rect 14644 22092 14654 22148
rect 33394 22092 33404 22148
rect 33460 22092 34188 22148
rect 34244 22092 34254 22148
rect 77746 22092 77756 22148
rect 77812 22092 80892 22148
rect 80948 22092 80958 22148
rect 0 22036 800 22064
rect 0 21980 1708 22036
rect 1764 21980 2940 22036
rect 2996 21980 3006 22036
rect 74834 21980 74844 22036
rect 74900 21980 75404 22036
rect 75460 21980 75470 22036
rect 0 21952 800 21980
rect 8758 21924 8768 21980
rect 8824 21924 8872 21980
rect 8928 21924 8976 21980
rect 9032 21924 9080 21980
rect 9136 21924 9184 21980
rect 9240 21924 9288 21980
rect 9344 21924 9392 21980
rect 9448 21924 9458 21980
rect 17758 21924 17768 21980
rect 17824 21924 17872 21980
rect 17928 21924 17976 21980
rect 18032 21924 18080 21980
rect 18136 21924 18184 21980
rect 18240 21924 18288 21980
rect 18344 21924 18392 21980
rect 18448 21924 18458 21980
rect 26758 21924 26768 21980
rect 26824 21924 26872 21980
rect 26928 21924 26976 21980
rect 27032 21924 27080 21980
rect 27136 21924 27184 21980
rect 27240 21924 27288 21980
rect 27344 21924 27392 21980
rect 27448 21924 27458 21980
rect 35758 21924 35768 21980
rect 35824 21924 35872 21980
rect 35928 21924 35976 21980
rect 36032 21924 36080 21980
rect 36136 21924 36184 21980
rect 36240 21924 36288 21980
rect 36344 21924 36392 21980
rect 36448 21924 36458 21980
rect 44758 21924 44768 21980
rect 44824 21924 44872 21980
rect 44928 21924 44976 21980
rect 45032 21924 45080 21980
rect 45136 21924 45184 21980
rect 45240 21924 45288 21980
rect 45344 21924 45392 21980
rect 45448 21924 45458 21980
rect 53758 21924 53768 21980
rect 53824 21924 53872 21980
rect 53928 21924 53976 21980
rect 54032 21924 54080 21980
rect 54136 21924 54184 21980
rect 54240 21924 54288 21980
rect 54344 21924 54392 21980
rect 54448 21924 54458 21980
rect 62758 21924 62768 21980
rect 62824 21924 62872 21980
rect 62928 21924 62976 21980
rect 63032 21924 63080 21980
rect 63136 21924 63184 21980
rect 63240 21924 63288 21980
rect 63344 21924 63392 21980
rect 63448 21924 63458 21980
rect 71758 21924 71768 21980
rect 71824 21924 71872 21980
rect 71928 21924 71976 21980
rect 72032 21924 72080 21980
rect 72136 21924 72184 21980
rect 72240 21924 72288 21980
rect 72344 21924 72392 21980
rect 72448 21924 72458 21980
rect 80758 21924 80768 21980
rect 80824 21924 80872 21980
rect 80928 21924 80976 21980
rect 81032 21924 81080 21980
rect 81136 21924 81184 21980
rect 81240 21924 81288 21980
rect 81344 21924 81392 21980
rect 81448 21924 81458 21980
rect 89758 21924 89768 21980
rect 89824 21924 89872 21980
rect 89928 21924 89976 21980
rect 90032 21924 90080 21980
rect 90136 21924 90184 21980
rect 90240 21924 90288 21980
rect 90344 21924 90392 21980
rect 90448 21924 90458 21980
rect 9090 21756 9100 21812
rect 9156 21756 12460 21812
rect 12516 21756 13020 21812
rect 13076 21756 13086 21812
rect 14802 21756 14812 21812
rect 14868 21756 15596 21812
rect 15652 21756 20076 21812
rect 20132 21756 23100 21812
rect 23156 21756 23166 21812
rect 28354 21756 28364 21812
rect 28420 21756 29036 21812
rect 29092 21756 29102 21812
rect 30594 21756 30604 21812
rect 30660 21756 31948 21812
rect 32004 21756 33124 21812
rect 39890 21756 39900 21812
rect 39956 21756 43372 21812
rect 43428 21756 43438 21812
rect 43652 21756 43820 21812
rect 43876 21756 43886 21812
rect 66658 21756 66668 21812
rect 66724 21756 96572 21812
rect 96628 21756 96638 21812
rect 33068 21700 33124 21756
rect 13794 21644 13804 21700
rect 13860 21644 15148 21700
rect 15204 21644 15214 21700
rect 33058 21644 33068 21700
rect 33124 21644 36204 21700
rect 36260 21644 36270 21700
rect 43652 21588 43708 21756
rect 64642 21644 64652 21700
rect 64708 21644 65100 21700
rect 65156 21644 68124 21700
rect 68180 21644 69468 21700
rect 69524 21644 70364 21700
rect 70420 21644 70430 21700
rect 75170 21644 75180 21700
rect 75236 21644 75740 21700
rect 75796 21644 77756 21700
rect 77812 21644 77822 21700
rect 1922 21532 1932 21588
rect 1988 21532 10668 21588
rect 10724 21532 10734 21588
rect 14354 21532 14364 21588
rect 14420 21532 16156 21588
rect 16212 21532 16222 21588
rect 38994 21532 39004 21588
rect 39060 21532 42924 21588
rect 42980 21532 43708 21588
rect 70364 21588 70420 21644
rect 70364 21532 73500 21588
rect 73556 21532 75292 21588
rect 75348 21532 75852 21588
rect 75908 21532 78764 21588
rect 78820 21532 80556 21588
rect 80612 21532 81004 21588
rect 81060 21532 81564 21588
rect 81620 21532 81630 21588
rect 1698 21420 1708 21476
rect 1764 21420 2492 21476
rect 2548 21420 2558 21476
rect 2706 21420 2716 21476
rect 2772 21420 27020 21476
rect 27076 21420 29372 21476
rect 29428 21420 29438 21476
rect 43586 21420 43596 21476
rect 43652 21420 45612 21476
rect 45668 21420 46956 21476
rect 47012 21420 47022 21476
rect 32498 21308 32508 21364
rect 32564 21308 33628 21364
rect 33684 21308 33694 21364
rect 43810 21308 43820 21364
rect 43876 21308 84364 21364
rect 84420 21308 84430 21364
rect 80434 21196 80444 21252
rect 80500 21196 81676 21252
rect 81732 21196 82684 21252
rect 82740 21196 82750 21252
rect 4258 21140 4268 21196
rect 4324 21140 4372 21196
rect 4428 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4788 21196
rect 4844 21140 4892 21196
rect 4948 21140 4958 21196
rect 13258 21140 13268 21196
rect 13324 21140 13372 21196
rect 13428 21140 13476 21196
rect 13532 21140 13580 21196
rect 13636 21140 13684 21196
rect 13740 21140 13788 21196
rect 13844 21140 13892 21196
rect 13948 21140 13958 21196
rect 22258 21140 22268 21196
rect 22324 21140 22372 21196
rect 22428 21140 22476 21196
rect 22532 21140 22580 21196
rect 22636 21140 22684 21196
rect 22740 21140 22788 21196
rect 22844 21140 22892 21196
rect 22948 21140 22958 21196
rect 31258 21140 31268 21196
rect 31324 21140 31372 21196
rect 31428 21140 31476 21196
rect 31532 21140 31580 21196
rect 31636 21140 31684 21196
rect 31740 21140 31788 21196
rect 31844 21140 31892 21196
rect 31948 21140 31958 21196
rect 40258 21140 40268 21196
rect 40324 21140 40372 21196
rect 40428 21140 40476 21196
rect 40532 21140 40580 21196
rect 40636 21140 40684 21196
rect 40740 21140 40788 21196
rect 40844 21140 40892 21196
rect 40948 21140 40958 21196
rect 49258 21140 49268 21196
rect 49324 21140 49372 21196
rect 49428 21140 49476 21196
rect 49532 21140 49580 21196
rect 49636 21140 49684 21196
rect 49740 21140 49788 21196
rect 49844 21140 49892 21196
rect 49948 21140 49958 21196
rect 58258 21140 58268 21196
rect 58324 21140 58372 21196
rect 58428 21140 58476 21196
rect 58532 21140 58580 21196
rect 58636 21140 58684 21196
rect 58740 21140 58788 21196
rect 58844 21140 58892 21196
rect 58948 21140 58958 21196
rect 67258 21140 67268 21196
rect 67324 21140 67372 21196
rect 67428 21140 67476 21196
rect 67532 21140 67580 21196
rect 67636 21140 67684 21196
rect 67740 21140 67788 21196
rect 67844 21140 67892 21196
rect 67948 21140 67958 21196
rect 76258 21140 76268 21196
rect 76324 21140 76372 21196
rect 76428 21140 76476 21196
rect 76532 21140 76580 21196
rect 76636 21140 76684 21196
rect 76740 21140 76788 21196
rect 76844 21140 76892 21196
rect 76948 21140 76958 21196
rect 85258 21140 85268 21196
rect 85324 21140 85372 21196
rect 85428 21140 85476 21196
rect 85532 21140 85580 21196
rect 85636 21140 85684 21196
rect 85740 21140 85788 21196
rect 85844 21140 85892 21196
rect 85948 21140 85958 21196
rect 94258 21140 94268 21196
rect 94324 21140 94372 21196
rect 94428 21140 94476 21196
rect 94532 21140 94580 21196
rect 94636 21140 94684 21196
rect 94740 21140 94788 21196
rect 94844 21140 94892 21196
rect 94948 21140 94958 21196
rect 4610 20972 4620 21028
rect 4676 20972 5852 21028
rect 5908 20972 26572 21028
rect 26628 20972 27356 21028
rect 27412 20972 29148 21028
rect 29204 20972 29214 21028
rect 30146 20972 30156 21028
rect 30212 20972 39004 21028
rect 39060 20972 42140 21028
rect 42196 20972 42206 21028
rect 56018 20972 56028 21028
rect 56084 20972 56700 21028
rect 56756 20972 56766 21028
rect 64530 20972 64540 21028
rect 64596 20972 65212 21028
rect 65268 20972 65884 21028
rect 65940 20972 65950 21028
rect 0 20916 800 20944
rect 99200 20916 100000 20944
rect 0 20860 1708 20916
rect 1764 20860 1774 20916
rect 15810 20860 15820 20916
rect 15876 20860 16828 20916
rect 16884 20860 18396 20916
rect 18452 20860 55468 20916
rect 55524 20860 56140 20916
rect 56196 20860 56206 20916
rect 64642 20860 64652 20916
rect 64708 20860 65548 20916
rect 65604 20860 65614 20916
rect 68674 20860 68684 20916
rect 68740 20860 73724 20916
rect 73780 20860 74172 20916
rect 74228 20860 74238 20916
rect 98018 20860 98028 20916
rect 98084 20860 100000 20916
rect 0 20832 800 20860
rect 99200 20832 100000 20860
rect 2034 20748 2044 20804
rect 2100 20748 6748 20804
rect 6804 20748 6814 20804
rect 14578 20748 14588 20804
rect 14644 20748 15260 20804
rect 15316 20748 15326 20804
rect 22978 20748 22988 20804
rect 23044 20748 24052 20804
rect 24210 20748 24220 20804
rect 24276 20748 28588 20804
rect 28644 20748 28654 20804
rect 31892 20748 32620 20804
rect 32676 20748 33740 20804
rect 33796 20748 33806 20804
rect 39218 20748 39228 20804
rect 39284 20748 40124 20804
rect 40180 20748 40190 20804
rect 55412 20748 56028 20804
rect 56084 20748 56094 20804
rect 56354 20748 56364 20804
rect 56420 20748 72044 20804
rect 72100 20748 72110 20804
rect 23996 20692 24052 20748
rect 31892 20692 31948 20748
rect 55412 20692 55468 20748
rect 17826 20636 17836 20692
rect 17892 20636 18732 20692
rect 18788 20636 18798 20692
rect 22418 20636 22428 20692
rect 22484 20636 23436 20692
rect 23492 20636 23502 20692
rect 23986 20636 23996 20692
rect 24052 20636 31948 20692
rect 34402 20636 34412 20692
rect 34468 20636 36988 20692
rect 37044 20636 43932 20692
rect 43988 20636 43998 20692
rect 46946 20636 46956 20692
rect 47012 20636 55468 20692
rect 24546 20524 24556 20580
rect 24612 20524 25340 20580
rect 25396 20524 25406 20580
rect 44146 20524 44156 20580
rect 44212 20524 55468 20580
rect 71362 20524 71372 20580
rect 71428 20524 72156 20580
rect 72212 20524 72222 20580
rect 72482 20524 72492 20580
rect 72548 20524 73052 20580
rect 73108 20524 74956 20580
rect 75012 20524 75022 20580
rect 85026 20524 85036 20580
rect 85092 20524 86156 20580
rect 86212 20524 86222 20580
rect 8758 20356 8768 20412
rect 8824 20356 8872 20412
rect 8928 20356 8976 20412
rect 9032 20356 9080 20412
rect 9136 20356 9184 20412
rect 9240 20356 9288 20412
rect 9344 20356 9392 20412
rect 9448 20356 9458 20412
rect 17758 20356 17768 20412
rect 17824 20356 17872 20412
rect 17928 20356 17976 20412
rect 18032 20356 18080 20412
rect 18136 20356 18184 20412
rect 18240 20356 18288 20412
rect 18344 20356 18392 20412
rect 18448 20356 18458 20412
rect 26758 20356 26768 20412
rect 26824 20356 26872 20412
rect 26928 20356 26976 20412
rect 27032 20356 27080 20412
rect 27136 20356 27184 20412
rect 27240 20356 27288 20412
rect 27344 20356 27392 20412
rect 27448 20356 27458 20412
rect 35758 20356 35768 20412
rect 35824 20356 35872 20412
rect 35928 20356 35976 20412
rect 36032 20356 36080 20412
rect 36136 20356 36184 20412
rect 36240 20356 36288 20412
rect 36344 20356 36392 20412
rect 36448 20356 36458 20412
rect 44758 20356 44768 20412
rect 44824 20356 44872 20412
rect 44928 20356 44976 20412
rect 45032 20356 45080 20412
rect 45136 20356 45184 20412
rect 45240 20356 45288 20412
rect 45344 20356 45392 20412
rect 45448 20356 45458 20412
rect 53758 20356 53768 20412
rect 53824 20356 53872 20412
rect 53928 20356 53976 20412
rect 54032 20356 54080 20412
rect 54136 20356 54184 20412
rect 54240 20356 54288 20412
rect 54344 20356 54392 20412
rect 54448 20356 54458 20412
rect 55412 20244 55468 20524
rect 62758 20356 62768 20412
rect 62824 20356 62872 20412
rect 62928 20356 62976 20412
rect 63032 20356 63080 20412
rect 63136 20356 63184 20412
rect 63240 20356 63288 20412
rect 63344 20356 63392 20412
rect 63448 20356 63458 20412
rect 71758 20356 71768 20412
rect 71824 20356 71872 20412
rect 71928 20356 71976 20412
rect 72032 20356 72080 20412
rect 72136 20356 72184 20412
rect 72240 20356 72288 20412
rect 72344 20356 72392 20412
rect 72448 20356 72458 20412
rect 80758 20356 80768 20412
rect 80824 20356 80872 20412
rect 80928 20356 80976 20412
rect 81032 20356 81080 20412
rect 81136 20356 81184 20412
rect 81240 20356 81288 20412
rect 81344 20356 81392 20412
rect 81448 20356 81458 20412
rect 89758 20356 89768 20412
rect 89824 20356 89872 20412
rect 89928 20356 89976 20412
rect 90032 20356 90080 20412
rect 90136 20356 90184 20412
rect 90240 20356 90288 20412
rect 90344 20356 90392 20412
rect 90448 20356 90458 20412
rect 28578 20188 28588 20244
rect 28644 20188 40236 20244
rect 40292 20188 40302 20244
rect 55412 20188 76300 20244
rect 76356 20188 76366 20244
rect 80098 20188 80108 20244
rect 80164 20188 81900 20244
rect 81956 20188 81966 20244
rect 5282 20076 5292 20132
rect 5348 20076 10444 20132
rect 10500 20076 10510 20132
rect 27794 20076 27804 20132
rect 27860 20076 28476 20132
rect 28532 20076 29372 20132
rect 29428 20076 30604 20132
rect 30660 20076 30670 20132
rect 73378 20076 73388 20132
rect 73444 20076 74396 20132
rect 74452 20076 74462 20132
rect 78082 20076 78092 20132
rect 78148 20076 79772 20132
rect 79828 20076 79838 20132
rect 81554 20076 81564 20132
rect 81620 20076 82908 20132
rect 82964 20076 83356 20132
rect 83412 20076 84252 20132
rect 84308 20076 85372 20132
rect 85428 20076 85438 20132
rect 85586 20076 85596 20132
rect 85652 20076 89068 20132
rect 89124 20076 89134 20132
rect 4498 19964 4508 20020
rect 4564 19964 6076 20020
rect 6132 19964 6142 20020
rect 40450 19964 40460 20020
rect 40516 19964 43708 20020
rect 76962 19964 76972 20020
rect 77028 19964 77980 20020
rect 78036 19964 78046 20020
rect 81666 19964 81676 20020
rect 81732 19964 83020 20020
rect 83076 19964 83086 20020
rect 5058 19852 5068 19908
rect 5124 19852 5740 19908
rect 5796 19852 7308 19908
rect 7364 19852 17500 19908
rect 17556 19852 17566 19908
rect 0 19796 800 19824
rect 43652 19796 43708 19964
rect 74946 19852 74956 19908
rect 75012 19852 76524 19908
rect 76580 19852 77420 19908
rect 77476 19852 80668 19908
rect 80724 19852 84700 19908
rect 84756 19852 85036 19908
rect 85092 19852 85102 19908
rect 0 19740 1708 19796
rect 1764 19740 1774 19796
rect 43652 19740 80444 19796
rect 80500 19740 81004 19796
rect 81060 19740 81070 19796
rect 0 19712 800 19740
rect 4258 19572 4268 19628
rect 4324 19572 4372 19628
rect 4428 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4788 19628
rect 4844 19572 4892 19628
rect 4948 19572 4958 19628
rect 13258 19572 13268 19628
rect 13324 19572 13372 19628
rect 13428 19572 13476 19628
rect 13532 19572 13580 19628
rect 13636 19572 13684 19628
rect 13740 19572 13788 19628
rect 13844 19572 13892 19628
rect 13948 19572 13958 19628
rect 22258 19572 22268 19628
rect 22324 19572 22372 19628
rect 22428 19572 22476 19628
rect 22532 19572 22580 19628
rect 22636 19572 22684 19628
rect 22740 19572 22788 19628
rect 22844 19572 22892 19628
rect 22948 19572 22958 19628
rect 31258 19572 31268 19628
rect 31324 19572 31372 19628
rect 31428 19572 31476 19628
rect 31532 19572 31580 19628
rect 31636 19572 31684 19628
rect 31740 19572 31788 19628
rect 31844 19572 31892 19628
rect 31948 19572 31958 19628
rect 40258 19572 40268 19628
rect 40324 19572 40372 19628
rect 40428 19572 40476 19628
rect 40532 19572 40580 19628
rect 40636 19572 40684 19628
rect 40740 19572 40788 19628
rect 40844 19572 40892 19628
rect 40948 19572 40958 19628
rect 49258 19572 49268 19628
rect 49324 19572 49372 19628
rect 49428 19572 49476 19628
rect 49532 19572 49580 19628
rect 49636 19572 49684 19628
rect 49740 19572 49788 19628
rect 49844 19572 49892 19628
rect 49948 19572 49958 19628
rect 58258 19572 58268 19628
rect 58324 19572 58372 19628
rect 58428 19572 58476 19628
rect 58532 19572 58580 19628
rect 58636 19572 58684 19628
rect 58740 19572 58788 19628
rect 58844 19572 58892 19628
rect 58948 19572 58958 19628
rect 67258 19572 67268 19628
rect 67324 19572 67372 19628
rect 67428 19572 67476 19628
rect 67532 19572 67580 19628
rect 67636 19572 67684 19628
rect 67740 19572 67788 19628
rect 67844 19572 67892 19628
rect 67948 19572 67958 19628
rect 76258 19572 76268 19628
rect 76324 19572 76372 19628
rect 76428 19572 76476 19628
rect 76532 19572 76580 19628
rect 76636 19572 76684 19628
rect 76740 19572 76788 19628
rect 76844 19572 76892 19628
rect 76948 19572 76958 19628
rect 85258 19572 85268 19628
rect 85324 19572 85372 19628
rect 85428 19572 85476 19628
rect 85532 19572 85580 19628
rect 85636 19572 85684 19628
rect 85740 19572 85788 19628
rect 85844 19572 85892 19628
rect 85948 19572 85958 19628
rect 94258 19572 94268 19628
rect 94324 19572 94372 19628
rect 94428 19572 94476 19628
rect 94532 19572 94580 19628
rect 94636 19572 94684 19628
rect 94740 19572 94788 19628
rect 94844 19572 94892 19628
rect 94948 19572 94958 19628
rect 2370 19404 2380 19460
rect 2436 19404 18508 19460
rect 18564 19404 19292 19460
rect 19348 19404 19358 19460
rect 74386 19404 74396 19460
rect 74452 19404 75180 19460
rect 75236 19404 75246 19460
rect 1698 19292 1708 19348
rect 1764 19292 3164 19348
rect 3220 19292 3230 19348
rect 73826 19292 73836 19348
rect 73892 19292 74732 19348
rect 74788 19292 75628 19348
rect 75684 19292 79212 19348
rect 79268 19292 79278 19348
rect 40002 19180 40012 19236
rect 40068 19180 44268 19236
rect 44324 19180 44334 19236
rect 99200 19124 100000 19152
rect 71474 19068 71484 19124
rect 71540 19068 96684 19124
rect 96740 19068 96750 19124
rect 98018 19068 98028 19124
rect 98084 19068 100000 19124
rect 99200 19040 100000 19068
rect 2034 18956 2044 19012
rect 2100 18956 2828 19012
rect 2884 18956 2894 19012
rect 79202 18956 79212 19012
rect 79268 18956 79660 19012
rect 79716 18956 82796 19012
rect 82852 18956 82862 19012
rect 85138 18956 85148 19012
rect 85204 18956 88284 19012
rect 88340 18956 88350 19012
rect 8758 18788 8768 18844
rect 8824 18788 8872 18844
rect 8928 18788 8976 18844
rect 9032 18788 9080 18844
rect 9136 18788 9184 18844
rect 9240 18788 9288 18844
rect 9344 18788 9392 18844
rect 9448 18788 9458 18844
rect 17758 18788 17768 18844
rect 17824 18788 17872 18844
rect 17928 18788 17976 18844
rect 18032 18788 18080 18844
rect 18136 18788 18184 18844
rect 18240 18788 18288 18844
rect 18344 18788 18392 18844
rect 18448 18788 18458 18844
rect 26758 18788 26768 18844
rect 26824 18788 26872 18844
rect 26928 18788 26976 18844
rect 27032 18788 27080 18844
rect 27136 18788 27184 18844
rect 27240 18788 27288 18844
rect 27344 18788 27392 18844
rect 27448 18788 27458 18844
rect 35758 18788 35768 18844
rect 35824 18788 35872 18844
rect 35928 18788 35976 18844
rect 36032 18788 36080 18844
rect 36136 18788 36184 18844
rect 36240 18788 36288 18844
rect 36344 18788 36392 18844
rect 36448 18788 36458 18844
rect 44758 18788 44768 18844
rect 44824 18788 44872 18844
rect 44928 18788 44976 18844
rect 45032 18788 45080 18844
rect 45136 18788 45184 18844
rect 45240 18788 45288 18844
rect 45344 18788 45392 18844
rect 45448 18788 45458 18844
rect 53758 18788 53768 18844
rect 53824 18788 53872 18844
rect 53928 18788 53976 18844
rect 54032 18788 54080 18844
rect 54136 18788 54184 18844
rect 54240 18788 54288 18844
rect 54344 18788 54392 18844
rect 54448 18788 54458 18844
rect 62758 18788 62768 18844
rect 62824 18788 62872 18844
rect 62928 18788 62976 18844
rect 63032 18788 63080 18844
rect 63136 18788 63184 18844
rect 63240 18788 63288 18844
rect 63344 18788 63392 18844
rect 63448 18788 63458 18844
rect 71758 18788 71768 18844
rect 71824 18788 71872 18844
rect 71928 18788 71976 18844
rect 72032 18788 72080 18844
rect 72136 18788 72184 18844
rect 72240 18788 72288 18844
rect 72344 18788 72392 18844
rect 72448 18788 72458 18844
rect 80758 18788 80768 18844
rect 80824 18788 80872 18844
rect 80928 18788 80976 18844
rect 81032 18788 81080 18844
rect 81136 18788 81184 18844
rect 81240 18788 81288 18844
rect 81344 18788 81392 18844
rect 81448 18788 81458 18844
rect 89758 18788 89768 18844
rect 89824 18788 89872 18844
rect 89928 18788 89976 18844
rect 90032 18788 90080 18844
rect 90136 18788 90184 18844
rect 90240 18788 90288 18844
rect 90344 18788 90392 18844
rect 90448 18788 90458 18844
rect 0 18676 800 18704
rect 0 18620 2268 18676
rect 2324 18620 2716 18676
rect 2772 18620 2782 18676
rect 0 18592 800 18620
rect 89058 18508 89068 18564
rect 89124 18508 89964 18564
rect 90020 18508 90030 18564
rect 4258 18004 4268 18060
rect 4324 18004 4372 18060
rect 4428 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4788 18060
rect 4844 18004 4892 18060
rect 4948 18004 4958 18060
rect 13258 18004 13268 18060
rect 13324 18004 13372 18060
rect 13428 18004 13476 18060
rect 13532 18004 13580 18060
rect 13636 18004 13684 18060
rect 13740 18004 13788 18060
rect 13844 18004 13892 18060
rect 13948 18004 13958 18060
rect 22258 18004 22268 18060
rect 22324 18004 22372 18060
rect 22428 18004 22476 18060
rect 22532 18004 22580 18060
rect 22636 18004 22684 18060
rect 22740 18004 22788 18060
rect 22844 18004 22892 18060
rect 22948 18004 22958 18060
rect 31258 18004 31268 18060
rect 31324 18004 31372 18060
rect 31428 18004 31476 18060
rect 31532 18004 31580 18060
rect 31636 18004 31684 18060
rect 31740 18004 31788 18060
rect 31844 18004 31892 18060
rect 31948 18004 31958 18060
rect 40258 18004 40268 18060
rect 40324 18004 40372 18060
rect 40428 18004 40476 18060
rect 40532 18004 40580 18060
rect 40636 18004 40684 18060
rect 40740 18004 40788 18060
rect 40844 18004 40892 18060
rect 40948 18004 40958 18060
rect 49258 18004 49268 18060
rect 49324 18004 49372 18060
rect 49428 18004 49476 18060
rect 49532 18004 49580 18060
rect 49636 18004 49684 18060
rect 49740 18004 49788 18060
rect 49844 18004 49892 18060
rect 49948 18004 49958 18060
rect 58258 18004 58268 18060
rect 58324 18004 58372 18060
rect 58428 18004 58476 18060
rect 58532 18004 58580 18060
rect 58636 18004 58684 18060
rect 58740 18004 58788 18060
rect 58844 18004 58892 18060
rect 58948 18004 58958 18060
rect 67258 18004 67268 18060
rect 67324 18004 67372 18060
rect 67428 18004 67476 18060
rect 67532 18004 67580 18060
rect 67636 18004 67684 18060
rect 67740 18004 67788 18060
rect 67844 18004 67892 18060
rect 67948 18004 67958 18060
rect 76258 18004 76268 18060
rect 76324 18004 76372 18060
rect 76428 18004 76476 18060
rect 76532 18004 76580 18060
rect 76636 18004 76684 18060
rect 76740 18004 76788 18060
rect 76844 18004 76892 18060
rect 76948 18004 76958 18060
rect 85258 18004 85268 18060
rect 85324 18004 85372 18060
rect 85428 18004 85476 18060
rect 85532 18004 85580 18060
rect 85636 18004 85684 18060
rect 85740 18004 85788 18060
rect 85844 18004 85892 18060
rect 85948 18004 85958 18060
rect 94258 18004 94268 18060
rect 94324 18004 94372 18060
rect 94428 18004 94476 18060
rect 94532 18004 94580 18060
rect 94636 18004 94684 18060
rect 94740 18004 94788 18060
rect 94844 18004 94892 18060
rect 94948 18004 94958 18060
rect 83570 17612 83580 17668
rect 83636 17612 85708 17668
rect 85764 17612 85774 17668
rect 0 17556 800 17584
rect 0 17500 1708 17556
rect 1764 17500 2492 17556
rect 2548 17500 2558 17556
rect 0 17472 800 17500
rect 83682 17388 83692 17444
rect 83748 17388 96684 17444
rect 96740 17388 96750 17444
rect 99200 17332 100000 17360
rect 98018 17276 98028 17332
rect 98084 17276 100000 17332
rect 8758 17220 8768 17276
rect 8824 17220 8872 17276
rect 8928 17220 8976 17276
rect 9032 17220 9080 17276
rect 9136 17220 9184 17276
rect 9240 17220 9288 17276
rect 9344 17220 9392 17276
rect 9448 17220 9458 17276
rect 17758 17220 17768 17276
rect 17824 17220 17872 17276
rect 17928 17220 17976 17276
rect 18032 17220 18080 17276
rect 18136 17220 18184 17276
rect 18240 17220 18288 17276
rect 18344 17220 18392 17276
rect 18448 17220 18458 17276
rect 26758 17220 26768 17276
rect 26824 17220 26872 17276
rect 26928 17220 26976 17276
rect 27032 17220 27080 17276
rect 27136 17220 27184 17276
rect 27240 17220 27288 17276
rect 27344 17220 27392 17276
rect 27448 17220 27458 17276
rect 35758 17220 35768 17276
rect 35824 17220 35872 17276
rect 35928 17220 35976 17276
rect 36032 17220 36080 17276
rect 36136 17220 36184 17276
rect 36240 17220 36288 17276
rect 36344 17220 36392 17276
rect 36448 17220 36458 17276
rect 44758 17220 44768 17276
rect 44824 17220 44872 17276
rect 44928 17220 44976 17276
rect 45032 17220 45080 17276
rect 45136 17220 45184 17276
rect 45240 17220 45288 17276
rect 45344 17220 45392 17276
rect 45448 17220 45458 17276
rect 53758 17220 53768 17276
rect 53824 17220 53872 17276
rect 53928 17220 53976 17276
rect 54032 17220 54080 17276
rect 54136 17220 54184 17276
rect 54240 17220 54288 17276
rect 54344 17220 54392 17276
rect 54448 17220 54458 17276
rect 62758 17220 62768 17276
rect 62824 17220 62872 17276
rect 62928 17220 62976 17276
rect 63032 17220 63080 17276
rect 63136 17220 63184 17276
rect 63240 17220 63288 17276
rect 63344 17220 63392 17276
rect 63448 17220 63458 17276
rect 71758 17220 71768 17276
rect 71824 17220 71872 17276
rect 71928 17220 71976 17276
rect 72032 17220 72080 17276
rect 72136 17220 72184 17276
rect 72240 17220 72288 17276
rect 72344 17220 72392 17276
rect 72448 17220 72458 17276
rect 80758 17220 80768 17276
rect 80824 17220 80872 17276
rect 80928 17220 80976 17276
rect 81032 17220 81080 17276
rect 81136 17220 81184 17276
rect 81240 17220 81288 17276
rect 81344 17220 81392 17276
rect 81448 17220 81458 17276
rect 89758 17220 89768 17276
rect 89824 17220 89872 17276
rect 89928 17220 89976 17276
rect 90032 17220 90080 17276
rect 90136 17220 90184 17276
rect 90240 17220 90288 17276
rect 90344 17220 90392 17276
rect 90448 17220 90458 17276
rect 99200 17248 100000 17276
rect 0 16436 800 16464
rect 4258 16436 4268 16492
rect 4324 16436 4372 16492
rect 4428 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4788 16492
rect 4844 16436 4892 16492
rect 4948 16436 4958 16492
rect 13258 16436 13268 16492
rect 13324 16436 13372 16492
rect 13428 16436 13476 16492
rect 13532 16436 13580 16492
rect 13636 16436 13684 16492
rect 13740 16436 13788 16492
rect 13844 16436 13892 16492
rect 13948 16436 13958 16492
rect 22258 16436 22268 16492
rect 22324 16436 22372 16492
rect 22428 16436 22476 16492
rect 22532 16436 22580 16492
rect 22636 16436 22684 16492
rect 22740 16436 22788 16492
rect 22844 16436 22892 16492
rect 22948 16436 22958 16492
rect 31258 16436 31268 16492
rect 31324 16436 31372 16492
rect 31428 16436 31476 16492
rect 31532 16436 31580 16492
rect 31636 16436 31684 16492
rect 31740 16436 31788 16492
rect 31844 16436 31892 16492
rect 31948 16436 31958 16492
rect 40258 16436 40268 16492
rect 40324 16436 40372 16492
rect 40428 16436 40476 16492
rect 40532 16436 40580 16492
rect 40636 16436 40684 16492
rect 40740 16436 40788 16492
rect 40844 16436 40892 16492
rect 40948 16436 40958 16492
rect 49258 16436 49268 16492
rect 49324 16436 49372 16492
rect 49428 16436 49476 16492
rect 49532 16436 49580 16492
rect 49636 16436 49684 16492
rect 49740 16436 49788 16492
rect 49844 16436 49892 16492
rect 49948 16436 49958 16492
rect 58258 16436 58268 16492
rect 58324 16436 58372 16492
rect 58428 16436 58476 16492
rect 58532 16436 58580 16492
rect 58636 16436 58684 16492
rect 58740 16436 58788 16492
rect 58844 16436 58892 16492
rect 58948 16436 58958 16492
rect 67258 16436 67268 16492
rect 67324 16436 67372 16492
rect 67428 16436 67476 16492
rect 67532 16436 67580 16492
rect 67636 16436 67684 16492
rect 67740 16436 67788 16492
rect 67844 16436 67892 16492
rect 67948 16436 67958 16492
rect 76258 16436 76268 16492
rect 76324 16436 76372 16492
rect 76428 16436 76476 16492
rect 76532 16436 76580 16492
rect 76636 16436 76684 16492
rect 76740 16436 76788 16492
rect 76844 16436 76892 16492
rect 76948 16436 76958 16492
rect 85258 16436 85268 16492
rect 85324 16436 85372 16492
rect 85428 16436 85476 16492
rect 85532 16436 85580 16492
rect 85636 16436 85684 16492
rect 85740 16436 85788 16492
rect 85844 16436 85892 16492
rect 85948 16436 85958 16492
rect 94258 16436 94268 16492
rect 94324 16436 94372 16492
rect 94428 16436 94476 16492
rect 94532 16436 94580 16492
rect 94636 16436 94684 16492
rect 94740 16436 94788 16492
rect 94844 16436 94892 16492
rect 94948 16436 94958 16492
rect 0 16380 1708 16436
rect 1764 16380 2492 16436
rect 2548 16380 2558 16436
rect 0 16352 800 16380
rect 66210 16044 66220 16100
rect 66276 16044 96684 16100
rect 96740 16044 96750 16100
rect 8758 15652 8768 15708
rect 8824 15652 8872 15708
rect 8928 15652 8976 15708
rect 9032 15652 9080 15708
rect 9136 15652 9184 15708
rect 9240 15652 9288 15708
rect 9344 15652 9392 15708
rect 9448 15652 9458 15708
rect 17758 15652 17768 15708
rect 17824 15652 17872 15708
rect 17928 15652 17976 15708
rect 18032 15652 18080 15708
rect 18136 15652 18184 15708
rect 18240 15652 18288 15708
rect 18344 15652 18392 15708
rect 18448 15652 18458 15708
rect 26758 15652 26768 15708
rect 26824 15652 26872 15708
rect 26928 15652 26976 15708
rect 27032 15652 27080 15708
rect 27136 15652 27184 15708
rect 27240 15652 27288 15708
rect 27344 15652 27392 15708
rect 27448 15652 27458 15708
rect 35758 15652 35768 15708
rect 35824 15652 35872 15708
rect 35928 15652 35976 15708
rect 36032 15652 36080 15708
rect 36136 15652 36184 15708
rect 36240 15652 36288 15708
rect 36344 15652 36392 15708
rect 36448 15652 36458 15708
rect 44758 15652 44768 15708
rect 44824 15652 44872 15708
rect 44928 15652 44976 15708
rect 45032 15652 45080 15708
rect 45136 15652 45184 15708
rect 45240 15652 45288 15708
rect 45344 15652 45392 15708
rect 45448 15652 45458 15708
rect 53758 15652 53768 15708
rect 53824 15652 53872 15708
rect 53928 15652 53976 15708
rect 54032 15652 54080 15708
rect 54136 15652 54184 15708
rect 54240 15652 54288 15708
rect 54344 15652 54392 15708
rect 54448 15652 54458 15708
rect 62758 15652 62768 15708
rect 62824 15652 62872 15708
rect 62928 15652 62976 15708
rect 63032 15652 63080 15708
rect 63136 15652 63184 15708
rect 63240 15652 63288 15708
rect 63344 15652 63392 15708
rect 63448 15652 63458 15708
rect 71758 15652 71768 15708
rect 71824 15652 71872 15708
rect 71928 15652 71976 15708
rect 72032 15652 72080 15708
rect 72136 15652 72184 15708
rect 72240 15652 72288 15708
rect 72344 15652 72392 15708
rect 72448 15652 72458 15708
rect 80758 15652 80768 15708
rect 80824 15652 80872 15708
rect 80928 15652 80976 15708
rect 81032 15652 81080 15708
rect 81136 15652 81184 15708
rect 81240 15652 81288 15708
rect 81344 15652 81392 15708
rect 81448 15652 81458 15708
rect 89758 15652 89768 15708
rect 89824 15652 89872 15708
rect 89928 15652 89976 15708
rect 90032 15652 90080 15708
rect 90136 15652 90184 15708
rect 90240 15652 90288 15708
rect 90344 15652 90392 15708
rect 90448 15652 90458 15708
rect 99200 15540 100000 15568
rect 98018 15484 98028 15540
rect 98084 15484 100000 15540
rect 99200 15456 100000 15484
rect 0 15232 800 15344
rect 41234 15148 41244 15204
rect 41300 15148 43036 15204
rect 43092 15148 43102 15204
rect 4258 14868 4268 14924
rect 4324 14868 4372 14924
rect 4428 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4788 14924
rect 4844 14868 4892 14924
rect 4948 14868 4958 14924
rect 13258 14868 13268 14924
rect 13324 14868 13372 14924
rect 13428 14868 13476 14924
rect 13532 14868 13580 14924
rect 13636 14868 13684 14924
rect 13740 14868 13788 14924
rect 13844 14868 13892 14924
rect 13948 14868 13958 14924
rect 22258 14868 22268 14924
rect 22324 14868 22372 14924
rect 22428 14868 22476 14924
rect 22532 14868 22580 14924
rect 22636 14868 22684 14924
rect 22740 14868 22788 14924
rect 22844 14868 22892 14924
rect 22948 14868 22958 14924
rect 31258 14868 31268 14924
rect 31324 14868 31372 14924
rect 31428 14868 31476 14924
rect 31532 14868 31580 14924
rect 31636 14868 31684 14924
rect 31740 14868 31788 14924
rect 31844 14868 31892 14924
rect 31948 14868 31958 14924
rect 40258 14868 40268 14924
rect 40324 14868 40372 14924
rect 40428 14868 40476 14924
rect 40532 14868 40580 14924
rect 40636 14868 40684 14924
rect 40740 14868 40788 14924
rect 40844 14868 40892 14924
rect 40948 14868 40958 14924
rect 49258 14868 49268 14924
rect 49324 14868 49372 14924
rect 49428 14868 49476 14924
rect 49532 14868 49580 14924
rect 49636 14868 49684 14924
rect 49740 14868 49788 14924
rect 49844 14868 49892 14924
rect 49948 14868 49958 14924
rect 58258 14868 58268 14924
rect 58324 14868 58372 14924
rect 58428 14868 58476 14924
rect 58532 14868 58580 14924
rect 58636 14868 58684 14924
rect 58740 14868 58788 14924
rect 58844 14868 58892 14924
rect 58948 14868 58958 14924
rect 67258 14868 67268 14924
rect 67324 14868 67372 14924
rect 67428 14868 67476 14924
rect 67532 14868 67580 14924
rect 67636 14868 67684 14924
rect 67740 14868 67788 14924
rect 67844 14868 67892 14924
rect 67948 14868 67958 14924
rect 76258 14868 76268 14924
rect 76324 14868 76372 14924
rect 76428 14868 76476 14924
rect 76532 14868 76580 14924
rect 76636 14868 76684 14924
rect 76740 14868 76788 14924
rect 76844 14868 76892 14924
rect 76948 14868 76958 14924
rect 85258 14868 85268 14924
rect 85324 14868 85372 14924
rect 85428 14868 85476 14924
rect 85532 14868 85580 14924
rect 85636 14868 85684 14924
rect 85740 14868 85788 14924
rect 85844 14868 85892 14924
rect 85948 14868 85958 14924
rect 94258 14868 94268 14924
rect 94324 14868 94372 14924
rect 94428 14868 94476 14924
rect 94532 14868 94580 14924
rect 94636 14868 94684 14924
rect 94740 14868 94788 14924
rect 94844 14868 94892 14924
rect 94948 14868 94958 14924
rect 20738 14476 20748 14532
rect 20804 14476 21420 14532
rect 21476 14476 21486 14532
rect 45938 14476 45948 14532
rect 46004 14476 46732 14532
rect 46788 14476 46798 14532
rect 68338 14476 68348 14532
rect 68404 14476 70028 14532
rect 70084 14476 70094 14532
rect 80546 14476 80556 14532
rect 80612 14476 83020 14532
rect 83076 14476 90860 14532
rect 90916 14476 90926 14532
rect 96898 14476 96908 14532
rect 96964 14476 96974 14532
rect 96908 14420 96964 14476
rect 44258 14364 44268 14420
rect 44324 14364 47068 14420
rect 47124 14364 47134 14420
rect 83122 14364 83132 14420
rect 83188 14364 96964 14420
rect 27682 14252 27692 14308
rect 27748 14252 52108 14308
rect 52164 14252 52174 14308
rect 82226 14252 82236 14308
rect 82292 14252 88172 14308
rect 88228 14252 88238 14308
rect 0 14112 800 14224
rect 8758 14084 8768 14140
rect 8824 14084 8872 14140
rect 8928 14084 8976 14140
rect 9032 14084 9080 14140
rect 9136 14084 9184 14140
rect 9240 14084 9288 14140
rect 9344 14084 9392 14140
rect 9448 14084 9458 14140
rect 17758 14084 17768 14140
rect 17824 14084 17872 14140
rect 17928 14084 17976 14140
rect 18032 14084 18080 14140
rect 18136 14084 18184 14140
rect 18240 14084 18288 14140
rect 18344 14084 18392 14140
rect 18448 14084 18458 14140
rect 26758 14084 26768 14140
rect 26824 14084 26872 14140
rect 26928 14084 26976 14140
rect 27032 14084 27080 14140
rect 27136 14084 27184 14140
rect 27240 14084 27288 14140
rect 27344 14084 27392 14140
rect 27448 14084 27458 14140
rect 35758 14084 35768 14140
rect 35824 14084 35872 14140
rect 35928 14084 35976 14140
rect 36032 14084 36080 14140
rect 36136 14084 36184 14140
rect 36240 14084 36288 14140
rect 36344 14084 36392 14140
rect 36448 14084 36458 14140
rect 44758 14084 44768 14140
rect 44824 14084 44872 14140
rect 44928 14084 44976 14140
rect 45032 14084 45080 14140
rect 45136 14084 45184 14140
rect 45240 14084 45288 14140
rect 45344 14084 45392 14140
rect 45448 14084 45458 14140
rect 53758 14084 53768 14140
rect 53824 14084 53872 14140
rect 53928 14084 53976 14140
rect 54032 14084 54080 14140
rect 54136 14084 54184 14140
rect 54240 14084 54288 14140
rect 54344 14084 54392 14140
rect 54448 14084 54458 14140
rect 62758 14084 62768 14140
rect 62824 14084 62872 14140
rect 62928 14084 62976 14140
rect 63032 14084 63080 14140
rect 63136 14084 63184 14140
rect 63240 14084 63288 14140
rect 63344 14084 63392 14140
rect 63448 14084 63458 14140
rect 71758 14084 71768 14140
rect 71824 14084 71872 14140
rect 71928 14084 71976 14140
rect 72032 14084 72080 14140
rect 72136 14084 72184 14140
rect 72240 14084 72288 14140
rect 72344 14084 72392 14140
rect 72448 14084 72458 14140
rect 80758 14084 80768 14140
rect 80824 14084 80872 14140
rect 80928 14084 80976 14140
rect 81032 14084 81080 14140
rect 81136 14084 81184 14140
rect 81240 14084 81288 14140
rect 81344 14084 81392 14140
rect 81448 14084 81458 14140
rect 89758 14084 89768 14140
rect 89824 14084 89872 14140
rect 89928 14084 89976 14140
rect 90032 14084 90080 14140
rect 90136 14084 90184 14140
rect 90240 14084 90288 14140
rect 90344 14084 90392 14140
rect 90448 14084 90458 14140
rect 77746 14028 77756 14084
rect 77812 14028 78428 14084
rect 78484 14028 78494 14084
rect 2034 13916 2044 13972
rect 2100 13916 9660 13972
rect 9716 13916 9726 13972
rect 48962 13916 48972 13972
rect 49028 13916 53004 13972
rect 53060 13916 55580 13972
rect 55636 13916 55646 13972
rect 50372 13804 51660 13860
rect 51716 13804 52444 13860
rect 52500 13804 55132 13860
rect 55188 13804 55198 13860
rect 70802 13804 70812 13860
rect 70868 13804 72268 13860
rect 72324 13804 72334 13860
rect 77746 13804 77756 13860
rect 77812 13804 80220 13860
rect 80276 13804 80286 13860
rect 50372 13748 50428 13804
rect 99200 13748 100000 13776
rect 45378 13692 45388 13748
rect 45444 13692 46172 13748
rect 46228 13692 50428 13748
rect 54562 13692 54572 13748
rect 54628 13692 65548 13748
rect 65604 13692 65614 13748
rect 68338 13692 68348 13748
rect 68404 13692 74060 13748
rect 74116 13692 77308 13748
rect 77364 13692 77374 13748
rect 78642 13692 78652 13748
rect 78708 13692 80108 13748
rect 80164 13692 80174 13748
rect 80434 13692 80444 13748
rect 80500 13692 81788 13748
rect 81844 13692 81854 13748
rect 98018 13692 98028 13748
rect 98084 13692 100000 13748
rect 99200 13664 100000 13692
rect 46050 13580 46060 13636
rect 46116 13580 52332 13636
rect 52388 13580 52398 13636
rect 74834 13580 74844 13636
rect 74900 13580 75516 13636
rect 75572 13580 79324 13636
rect 79380 13580 82796 13636
rect 82852 13580 83580 13636
rect 83636 13580 83646 13636
rect 58930 13468 58940 13524
rect 58996 13468 60284 13524
rect 60340 13468 60350 13524
rect 4258 13300 4268 13356
rect 4324 13300 4372 13356
rect 4428 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4788 13356
rect 4844 13300 4892 13356
rect 4948 13300 4958 13356
rect 13258 13300 13268 13356
rect 13324 13300 13372 13356
rect 13428 13300 13476 13356
rect 13532 13300 13580 13356
rect 13636 13300 13684 13356
rect 13740 13300 13788 13356
rect 13844 13300 13892 13356
rect 13948 13300 13958 13356
rect 22258 13300 22268 13356
rect 22324 13300 22372 13356
rect 22428 13300 22476 13356
rect 22532 13300 22580 13356
rect 22636 13300 22684 13356
rect 22740 13300 22788 13356
rect 22844 13300 22892 13356
rect 22948 13300 22958 13356
rect 31258 13300 31268 13356
rect 31324 13300 31372 13356
rect 31428 13300 31476 13356
rect 31532 13300 31580 13356
rect 31636 13300 31684 13356
rect 31740 13300 31788 13356
rect 31844 13300 31892 13356
rect 31948 13300 31958 13356
rect 40258 13300 40268 13356
rect 40324 13300 40372 13356
rect 40428 13300 40476 13356
rect 40532 13300 40580 13356
rect 40636 13300 40684 13356
rect 40740 13300 40788 13356
rect 40844 13300 40892 13356
rect 40948 13300 40958 13356
rect 49258 13300 49268 13356
rect 49324 13300 49372 13356
rect 49428 13300 49476 13356
rect 49532 13300 49580 13356
rect 49636 13300 49684 13356
rect 49740 13300 49788 13356
rect 49844 13300 49892 13356
rect 49948 13300 49958 13356
rect 58258 13300 58268 13356
rect 58324 13300 58372 13356
rect 58428 13300 58476 13356
rect 58532 13300 58580 13356
rect 58636 13300 58684 13356
rect 58740 13300 58788 13356
rect 58844 13300 58892 13356
rect 58948 13300 58958 13356
rect 67258 13300 67268 13356
rect 67324 13300 67372 13356
rect 67428 13300 67476 13356
rect 67532 13300 67580 13356
rect 67636 13300 67684 13356
rect 67740 13300 67788 13356
rect 67844 13300 67892 13356
rect 67948 13300 67958 13356
rect 76258 13300 76268 13356
rect 76324 13300 76372 13356
rect 76428 13300 76476 13356
rect 76532 13300 76580 13356
rect 76636 13300 76684 13356
rect 76740 13300 76788 13356
rect 76844 13300 76892 13356
rect 76948 13300 76958 13356
rect 85258 13300 85268 13356
rect 85324 13300 85372 13356
rect 85428 13300 85476 13356
rect 85532 13300 85580 13356
rect 85636 13300 85684 13356
rect 85740 13300 85788 13356
rect 85844 13300 85892 13356
rect 85948 13300 85958 13356
rect 94258 13300 94268 13356
rect 94324 13300 94372 13356
rect 94428 13300 94476 13356
rect 94532 13300 94580 13356
rect 94636 13300 94684 13356
rect 94740 13300 94788 13356
rect 94844 13300 94892 13356
rect 94948 13300 94958 13356
rect 0 13076 800 13104
rect 0 13020 1708 13076
rect 1764 13020 2492 13076
rect 2548 13020 2558 13076
rect 0 12992 800 13020
rect 47170 12908 47180 12964
rect 47236 12908 50428 12964
rect 47730 12796 47740 12852
rect 47796 12796 49532 12852
rect 49588 12796 49598 12852
rect 50372 12684 50428 12908
rect 50484 12684 50876 12740
rect 50932 12684 51324 12740
rect 51380 12684 51390 12740
rect 73826 12684 73836 12740
rect 73892 12684 74284 12740
rect 74340 12684 81788 12740
rect 81844 12684 81854 12740
rect 78866 12572 78876 12628
rect 8758 12516 8768 12572
rect 8824 12516 8872 12572
rect 8928 12516 8976 12572
rect 9032 12516 9080 12572
rect 9136 12516 9184 12572
rect 9240 12516 9288 12572
rect 9344 12516 9392 12572
rect 9448 12516 9458 12572
rect 17758 12516 17768 12572
rect 17824 12516 17872 12572
rect 17928 12516 17976 12572
rect 18032 12516 18080 12572
rect 18136 12516 18184 12572
rect 18240 12516 18288 12572
rect 18344 12516 18392 12572
rect 18448 12516 18458 12572
rect 26758 12516 26768 12572
rect 26824 12516 26872 12572
rect 26928 12516 26976 12572
rect 27032 12516 27080 12572
rect 27136 12516 27184 12572
rect 27240 12516 27288 12572
rect 27344 12516 27392 12572
rect 27448 12516 27458 12572
rect 35758 12516 35768 12572
rect 35824 12516 35872 12572
rect 35928 12516 35976 12572
rect 36032 12516 36080 12572
rect 36136 12516 36184 12572
rect 36240 12516 36288 12572
rect 36344 12516 36392 12572
rect 36448 12516 36458 12572
rect 44758 12516 44768 12572
rect 44824 12516 44872 12572
rect 44928 12516 44976 12572
rect 45032 12516 45080 12572
rect 45136 12516 45184 12572
rect 45240 12516 45288 12572
rect 45344 12516 45392 12572
rect 45448 12516 45458 12572
rect 53758 12516 53768 12572
rect 53824 12516 53872 12572
rect 53928 12516 53976 12572
rect 54032 12516 54080 12572
rect 54136 12516 54184 12572
rect 54240 12516 54288 12572
rect 54344 12516 54392 12572
rect 54448 12516 54458 12572
rect 62758 12516 62768 12572
rect 62824 12516 62872 12572
rect 62928 12516 62976 12572
rect 63032 12516 63080 12572
rect 63136 12516 63184 12572
rect 63240 12516 63288 12572
rect 63344 12516 63392 12572
rect 63448 12516 63458 12572
rect 71758 12516 71768 12572
rect 71824 12516 71872 12572
rect 71928 12516 71976 12572
rect 72032 12516 72080 12572
rect 72136 12516 72184 12572
rect 72240 12516 72288 12572
rect 72344 12516 72392 12572
rect 72448 12516 72458 12572
rect 78932 12404 78988 12628
rect 80758 12516 80768 12572
rect 80824 12516 80872 12572
rect 80928 12516 80976 12572
rect 81032 12516 81080 12572
rect 81136 12516 81184 12572
rect 81240 12516 81288 12572
rect 81344 12516 81392 12572
rect 81448 12516 81458 12572
rect 89758 12516 89768 12572
rect 89824 12516 89872 12572
rect 89928 12516 89976 12572
rect 90032 12516 90080 12572
rect 90136 12516 90184 12572
rect 90240 12516 90288 12572
rect 90344 12516 90392 12572
rect 90448 12516 90458 12572
rect 57810 12348 57820 12404
rect 57876 12348 59052 12404
rect 59108 12348 59118 12404
rect 78932 12348 81620 12404
rect 81564 12292 81620 12348
rect 2034 12236 2044 12292
rect 2100 12236 33292 12292
rect 33348 12236 33358 12292
rect 46834 12236 46844 12292
rect 46900 12236 48860 12292
rect 48916 12236 48926 12292
rect 72818 12236 72828 12292
rect 72884 12236 81396 12292
rect 81554 12236 81564 12292
rect 81620 12236 81630 12292
rect 82348 12236 96572 12292
rect 96628 12236 96638 12292
rect 81340 12180 81396 12236
rect 82348 12180 82404 12236
rect 46498 12124 46508 12180
rect 46564 12124 48748 12180
rect 48804 12124 48814 12180
rect 78932 12124 80108 12180
rect 80164 12124 80174 12180
rect 81340 12124 82404 12180
rect 82562 12124 82572 12180
rect 82628 12124 91196 12180
rect 91252 12124 91262 12180
rect 30930 12012 30940 12068
rect 30996 12012 44380 12068
rect 44436 12012 47180 12068
rect 47236 12012 48188 12068
rect 48244 12012 48254 12068
rect 71362 12012 71372 12068
rect 71428 12012 72492 12068
rect 72548 12012 72558 12068
rect 78866 12012 78876 12068
rect 78932 12012 78988 12124
rect 81890 12012 81900 12068
rect 81956 12012 83804 12068
rect 83860 12012 86044 12068
rect 86100 12012 86110 12068
rect 0 11956 800 11984
rect 99200 11956 100000 11984
rect 0 11900 1708 11956
rect 1764 11900 2492 11956
rect 2548 11900 2558 11956
rect 98018 11900 98028 11956
rect 98084 11900 100000 11956
rect 0 11872 800 11900
rect 99200 11872 100000 11900
rect 4258 11732 4268 11788
rect 4324 11732 4372 11788
rect 4428 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4788 11788
rect 4844 11732 4892 11788
rect 4948 11732 4958 11788
rect 13258 11732 13268 11788
rect 13324 11732 13372 11788
rect 13428 11732 13476 11788
rect 13532 11732 13580 11788
rect 13636 11732 13684 11788
rect 13740 11732 13788 11788
rect 13844 11732 13892 11788
rect 13948 11732 13958 11788
rect 22258 11732 22268 11788
rect 22324 11732 22372 11788
rect 22428 11732 22476 11788
rect 22532 11732 22580 11788
rect 22636 11732 22684 11788
rect 22740 11732 22788 11788
rect 22844 11732 22892 11788
rect 22948 11732 22958 11788
rect 31258 11732 31268 11788
rect 31324 11732 31372 11788
rect 31428 11732 31476 11788
rect 31532 11732 31580 11788
rect 31636 11732 31684 11788
rect 31740 11732 31788 11788
rect 31844 11732 31892 11788
rect 31948 11732 31958 11788
rect 40258 11732 40268 11788
rect 40324 11732 40372 11788
rect 40428 11732 40476 11788
rect 40532 11732 40580 11788
rect 40636 11732 40684 11788
rect 40740 11732 40788 11788
rect 40844 11732 40892 11788
rect 40948 11732 40958 11788
rect 49258 11732 49268 11788
rect 49324 11732 49372 11788
rect 49428 11732 49476 11788
rect 49532 11732 49580 11788
rect 49636 11732 49684 11788
rect 49740 11732 49788 11788
rect 49844 11732 49892 11788
rect 49948 11732 49958 11788
rect 58258 11732 58268 11788
rect 58324 11732 58372 11788
rect 58428 11732 58476 11788
rect 58532 11732 58580 11788
rect 58636 11732 58684 11788
rect 58740 11732 58788 11788
rect 58844 11732 58892 11788
rect 58948 11732 58958 11788
rect 67258 11732 67268 11788
rect 67324 11732 67372 11788
rect 67428 11732 67476 11788
rect 67532 11732 67580 11788
rect 67636 11732 67684 11788
rect 67740 11732 67788 11788
rect 67844 11732 67892 11788
rect 67948 11732 67958 11788
rect 76258 11732 76268 11788
rect 76324 11732 76372 11788
rect 76428 11732 76476 11788
rect 76532 11732 76580 11788
rect 76636 11732 76684 11788
rect 76740 11732 76788 11788
rect 76844 11732 76892 11788
rect 76948 11732 76958 11788
rect 85258 11732 85268 11788
rect 85324 11732 85372 11788
rect 85428 11732 85476 11788
rect 85532 11732 85580 11788
rect 85636 11732 85684 11788
rect 85740 11732 85788 11788
rect 85844 11732 85892 11788
rect 85948 11732 85958 11788
rect 94258 11732 94268 11788
rect 94324 11732 94372 11788
rect 94428 11732 94476 11788
rect 94532 11732 94580 11788
rect 94636 11732 94684 11788
rect 94740 11732 94788 11788
rect 94844 11732 94892 11788
rect 94948 11732 94958 11788
rect 67554 11564 67564 11620
rect 67620 11564 68348 11620
rect 68404 11564 68414 11620
rect 44594 11452 44604 11508
rect 44660 11452 45612 11508
rect 45668 11452 45678 11508
rect 61282 11452 61292 11508
rect 61348 11452 62188 11508
rect 62244 11452 63644 11508
rect 63700 11452 63710 11508
rect 31154 11340 31164 11396
rect 31220 11340 39004 11396
rect 39060 11340 39070 11396
rect 58146 11340 58156 11396
rect 58212 11340 65772 11396
rect 65828 11340 65838 11396
rect 37650 11228 37660 11284
rect 37716 11228 41020 11284
rect 41076 11228 41086 11284
rect 43026 11228 43036 11284
rect 43092 11228 47068 11284
rect 47124 11228 47134 11284
rect 2034 11116 2044 11172
rect 2100 11116 25788 11172
rect 25844 11116 25854 11172
rect 59378 11116 59388 11172
rect 59444 11116 60620 11172
rect 60676 11116 61068 11172
rect 61124 11116 61134 11172
rect 81442 11116 81452 11172
rect 81508 11116 82124 11172
rect 82180 11116 82190 11172
rect 8758 10948 8768 11004
rect 8824 10948 8872 11004
rect 8928 10948 8976 11004
rect 9032 10948 9080 11004
rect 9136 10948 9184 11004
rect 9240 10948 9288 11004
rect 9344 10948 9392 11004
rect 9448 10948 9458 11004
rect 17758 10948 17768 11004
rect 17824 10948 17872 11004
rect 17928 10948 17976 11004
rect 18032 10948 18080 11004
rect 18136 10948 18184 11004
rect 18240 10948 18288 11004
rect 18344 10948 18392 11004
rect 18448 10948 18458 11004
rect 26758 10948 26768 11004
rect 26824 10948 26872 11004
rect 26928 10948 26976 11004
rect 27032 10948 27080 11004
rect 27136 10948 27184 11004
rect 27240 10948 27288 11004
rect 27344 10948 27392 11004
rect 27448 10948 27458 11004
rect 35758 10948 35768 11004
rect 35824 10948 35872 11004
rect 35928 10948 35976 11004
rect 36032 10948 36080 11004
rect 36136 10948 36184 11004
rect 36240 10948 36288 11004
rect 36344 10948 36392 11004
rect 36448 10948 36458 11004
rect 44758 10948 44768 11004
rect 44824 10948 44872 11004
rect 44928 10948 44976 11004
rect 45032 10948 45080 11004
rect 45136 10948 45184 11004
rect 45240 10948 45288 11004
rect 45344 10948 45392 11004
rect 45448 10948 45458 11004
rect 53758 10948 53768 11004
rect 53824 10948 53872 11004
rect 53928 10948 53976 11004
rect 54032 10948 54080 11004
rect 54136 10948 54184 11004
rect 54240 10948 54288 11004
rect 54344 10948 54392 11004
rect 54448 10948 54458 11004
rect 62758 10948 62768 11004
rect 62824 10948 62872 11004
rect 62928 10948 62976 11004
rect 63032 10948 63080 11004
rect 63136 10948 63184 11004
rect 63240 10948 63288 11004
rect 63344 10948 63392 11004
rect 63448 10948 63458 11004
rect 71758 10948 71768 11004
rect 71824 10948 71872 11004
rect 71928 10948 71976 11004
rect 72032 10948 72080 11004
rect 72136 10948 72184 11004
rect 72240 10948 72288 11004
rect 72344 10948 72392 11004
rect 72448 10948 72458 11004
rect 80758 10948 80768 11004
rect 80824 10948 80872 11004
rect 80928 10948 80976 11004
rect 81032 10948 81080 11004
rect 81136 10948 81184 11004
rect 81240 10948 81288 11004
rect 81344 10948 81392 11004
rect 81448 10948 81458 11004
rect 89758 10948 89768 11004
rect 89824 10948 89872 11004
rect 89928 10948 89976 11004
rect 90032 10948 90080 11004
rect 90136 10948 90184 11004
rect 90240 10948 90288 11004
rect 90344 10948 90392 11004
rect 90448 10948 90458 11004
rect 0 10836 800 10864
rect 0 10780 1708 10836
rect 1764 10780 2492 10836
rect 2548 10780 2558 10836
rect 0 10752 800 10780
rect 75058 10668 75068 10724
rect 75124 10668 76076 10724
rect 76132 10668 76142 10724
rect 78194 10668 78204 10724
rect 78260 10668 96684 10724
rect 96740 10668 96750 10724
rect 82226 10332 82236 10388
rect 82292 10332 88956 10388
rect 89012 10332 89022 10388
rect 4258 10164 4268 10220
rect 4324 10164 4372 10220
rect 4428 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4788 10220
rect 4844 10164 4892 10220
rect 4948 10164 4958 10220
rect 13258 10164 13268 10220
rect 13324 10164 13372 10220
rect 13428 10164 13476 10220
rect 13532 10164 13580 10220
rect 13636 10164 13684 10220
rect 13740 10164 13788 10220
rect 13844 10164 13892 10220
rect 13948 10164 13958 10220
rect 22258 10164 22268 10220
rect 22324 10164 22372 10220
rect 22428 10164 22476 10220
rect 22532 10164 22580 10220
rect 22636 10164 22684 10220
rect 22740 10164 22788 10220
rect 22844 10164 22892 10220
rect 22948 10164 22958 10220
rect 31258 10164 31268 10220
rect 31324 10164 31372 10220
rect 31428 10164 31476 10220
rect 31532 10164 31580 10220
rect 31636 10164 31684 10220
rect 31740 10164 31788 10220
rect 31844 10164 31892 10220
rect 31948 10164 31958 10220
rect 40258 10164 40268 10220
rect 40324 10164 40372 10220
rect 40428 10164 40476 10220
rect 40532 10164 40580 10220
rect 40636 10164 40684 10220
rect 40740 10164 40788 10220
rect 40844 10164 40892 10220
rect 40948 10164 40958 10220
rect 49258 10164 49268 10220
rect 49324 10164 49372 10220
rect 49428 10164 49476 10220
rect 49532 10164 49580 10220
rect 49636 10164 49684 10220
rect 49740 10164 49788 10220
rect 49844 10164 49892 10220
rect 49948 10164 49958 10220
rect 58258 10164 58268 10220
rect 58324 10164 58372 10220
rect 58428 10164 58476 10220
rect 58532 10164 58580 10220
rect 58636 10164 58684 10220
rect 58740 10164 58788 10220
rect 58844 10164 58892 10220
rect 58948 10164 58958 10220
rect 67258 10164 67268 10220
rect 67324 10164 67372 10220
rect 67428 10164 67476 10220
rect 67532 10164 67580 10220
rect 67636 10164 67684 10220
rect 67740 10164 67788 10220
rect 67844 10164 67892 10220
rect 67948 10164 67958 10220
rect 76258 10164 76268 10220
rect 76324 10164 76372 10220
rect 76428 10164 76476 10220
rect 76532 10164 76580 10220
rect 76636 10164 76684 10220
rect 76740 10164 76788 10220
rect 76844 10164 76892 10220
rect 76948 10164 76958 10220
rect 85258 10164 85268 10220
rect 85324 10164 85372 10220
rect 85428 10164 85476 10220
rect 85532 10164 85580 10220
rect 85636 10164 85684 10220
rect 85740 10164 85788 10220
rect 85844 10164 85892 10220
rect 85948 10164 85958 10220
rect 94258 10164 94268 10220
rect 94324 10164 94372 10220
rect 94428 10164 94476 10220
rect 94532 10164 94580 10220
rect 94636 10164 94684 10220
rect 94740 10164 94788 10220
rect 94844 10164 94892 10220
rect 94948 10164 94958 10220
rect 99200 10164 100000 10192
rect 51090 10108 51100 10164
rect 51156 10108 54684 10164
rect 54740 10108 54750 10164
rect 63634 10108 63644 10164
rect 63700 10108 65996 10164
rect 66052 10108 66062 10164
rect 98018 10108 98028 10164
rect 98084 10108 100000 10164
rect 99200 10080 100000 10108
rect 52098 9996 52108 10052
rect 52164 9996 59276 10052
rect 59332 9996 59342 10052
rect 85138 9996 85148 10052
rect 85204 9996 88060 10052
rect 88116 9996 88126 10052
rect 45042 9884 45052 9940
rect 45108 9884 46172 9940
rect 46228 9884 46238 9940
rect 37426 9772 37436 9828
rect 37492 9772 39004 9828
rect 39060 9772 39070 9828
rect 0 9716 800 9744
rect 0 9660 1708 9716
rect 1764 9660 2492 9716
rect 2548 9660 2558 9716
rect 28466 9660 28476 9716
rect 28532 9660 31948 9716
rect 32004 9660 35532 9716
rect 35588 9660 35598 9716
rect 40002 9660 40012 9716
rect 40068 9660 41020 9716
rect 41076 9660 41086 9716
rect 82786 9660 82796 9716
rect 82852 9660 84364 9716
rect 84420 9660 84430 9716
rect 0 9632 800 9660
rect 2034 9548 2044 9604
rect 2100 9548 28028 9604
rect 28084 9548 28094 9604
rect 45154 9548 45164 9604
rect 45220 9548 45668 9604
rect 8758 9380 8768 9436
rect 8824 9380 8872 9436
rect 8928 9380 8976 9436
rect 9032 9380 9080 9436
rect 9136 9380 9184 9436
rect 9240 9380 9288 9436
rect 9344 9380 9392 9436
rect 9448 9380 9458 9436
rect 17758 9380 17768 9436
rect 17824 9380 17872 9436
rect 17928 9380 17976 9436
rect 18032 9380 18080 9436
rect 18136 9380 18184 9436
rect 18240 9380 18288 9436
rect 18344 9380 18392 9436
rect 18448 9380 18458 9436
rect 26758 9380 26768 9436
rect 26824 9380 26872 9436
rect 26928 9380 26976 9436
rect 27032 9380 27080 9436
rect 27136 9380 27184 9436
rect 27240 9380 27288 9436
rect 27344 9380 27392 9436
rect 27448 9380 27458 9436
rect 35758 9380 35768 9436
rect 35824 9380 35872 9436
rect 35928 9380 35976 9436
rect 36032 9380 36080 9436
rect 36136 9380 36184 9436
rect 36240 9380 36288 9436
rect 36344 9380 36392 9436
rect 36448 9380 36458 9436
rect 44758 9380 44768 9436
rect 44824 9380 44872 9436
rect 44928 9380 44976 9436
rect 45032 9380 45080 9436
rect 45136 9380 45184 9436
rect 45240 9380 45288 9436
rect 45344 9380 45392 9436
rect 45448 9380 45458 9436
rect 42466 9324 42476 9380
rect 42532 9324 43708 9380
rect 43764 9324 43774 9380
rect 45612 9268 45668 9548
rect 53758 9380 53768 9436
rect 53824 9380 53872 9436
rect 53928 9380 53976 9436
rect 54032 9380 54080 9436
rect 54136 9380 54184 9436
rect 54240 9380 54288 9436
rect 54344 9380 54392 9436
rect 54448 9380 54458 9436
rect 62758 9380 62768 9436
rect 62824 9380 62872 9436
rect 62928 9380 62976 9436
rect 63032 9380 63080 9436
rect 63136 9380 63184 9436
rect 63240 9380 63288 9436
rect 63344 9380 63392 9436
rect 63448 9380 63458 9436
rect 71758 9380 71768 9436
rect 71824 9380 71872 9436
rect 71928 9380 71976 9436
rect 72032 9380 72080 9436
rect 72136 9380 72184 9436
rect 72240 9380 72288 9436
rect 72344 9380 72392 9436
rect 72448 9380 72458 9436
rect 80758 9380 80768 9436
rect 80824 9380 80872 9436
rect 80928 9380 80976 9436
rect 81032 9380 81080 9436
rect 81136 9380 81184 9436
rect 81240 9380 81288 9436
rect 81344 9380 81392 9436
rect 81448 9380 81458 9436
rect 89758 9380 89768 9436
rect 89824 9380 89872 9436
rect 89928 9380 89976 9436
rect 90032 9380 90080 9436
rect 90136 9380 90184 9436
rect 90240 9380 90288 9436
rect 90344 9380 90392 9436
rect 90448 9380 90458 9436
rect 36418 9212 36428 9268
rect 36484 9212 37212 9268
rect 37268 9212 37278 9268
rect 45378 9212 45388 9268
rect 45444 9212 45668 9268
rect 87378 9212 87388 9268
rect 87444 9212 96684 9268
rect 96740 9212 96750 9268
rect 77186 9100 77196 9156
rect 77252 9100 80668 9156
rect 80724 9100 80734 9156
rect 30034 8988 30044 9044
rect 30100 8988 31836 9044
rect 31892 8988 35308 9044
rect 35364 8988 35374 9044
rect 73602 8988 73612 9044
rect 73668 8988 76076 9044
rect 76132 8988 79100 9044
rect 79156 8988 79166 9044
rect 81890 8988 81900 9044
rect 81956 8988 84028 9044
rect 84084 8988 87500 9044
rect 87556 8988 87566 9044
rect 42690 8876 42700 8932
rect 42756 8876 44156 8932
rect 44212 8876 45836 8932
rect 45892 8876 45902 8932
rect 70914 8876 70924 8932
rect 70980 8876 72492 8932
rect 72548 8876 72558 8932
rect 0 8512 800 8624
rect 4258 8596 4268 8652
rect 4324 8596 4372 8652
rect 4428 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4788 8652
rect 4844 8596 4892 8652
rect 4948 8596 4958 8652
rect 13258 8596 13268 8652
rect 13324 8596 13372 8652
rect 13428 8596 13476 8652
rect 13532 8596 13580 8652
rect 13636 8596 13684 8652
rect 13740 8596 13788 8652
rect 13844 8596 13892 8652
rect 13948 8596 13958 8652
rect 22258 8596 22268 8652
rect 22324 8596 22372 8652
rect 22428 8596 22476 8652
rect 22532 8596 22580 8652
rect 22636 8596 22684 8652
rect 22740 8596 22788 8652
rect 22844 8596 22892 8652
rect 22948 8596 22958 8652
rect 31258 8596 31268 8652
rect 31324 8596 31372 8652
rect 31428 8596 31476 8652
rect 31532 8596 31580 8652
rect 31636 8596 31684 8652
rect 31740 8596 31788 8652
rect 31844 8596 31892 8652
rect 31948 8596 31958 8652
rect 40258 8596 40268 8652
rect 40324 8596 40372 8652
rect 40428 8596 40476 8652
rect 40532 8596 40580 8652
rect 40636 8596 40684 8652
rect 40740 8596 40788 8652
rect 40844 8596 40892 8652
rect 40948 8596 40958 8652
rect 49258 8596 49268 8652
rect 49324 8596 49372 8652
rect 49428 8596 49476 8652
rect 49532 8596 49580 8652
rect 49636 8596 49684 8652
rect 49740 8596 49788 8652
rect 49844 8596 49892 8652
rect 49948 8596 49958 8652
rect 58258 8596 58268 8652
rect 58324 8596 58372 8652
rect 58428 8596 58476 8652
rect 58532 8596 58580 8652
rect 58636 8596 58684 8652
rect 58740 8596 58788 8652
rect 58844 8596 58892 8652
rect 58948 8596 58958 8652
rect 67258 8596 67268 8652
rect 67324 8596 67372 8652
rect 67428 8596 67476 8652
rect 67532 8596 67580 8652
rect 67636 8596 67684 8652
rect 67740 8596 67788 8652
rect 67844 8596 67892 8652
rect 67948 8596 67958 8652
rect 76258 8596 76268 8652
rect 76324 8596 76372 8652
rect 76428 8596 76476 8652
rect 76532 8596 76580 8652
rect 76636 8596 76684 8652
rect 76740 8596 76788 8652
rect 76844 8596 76892 8652
rect 76948 8596 76958 8652
rect 85258 8596 85268 8652
rect 85324 8596 85372 8652
rect 85428 8596 85476 8652
rect 85532 8596 85580 8652
rect 85636 8596 85684 8652
rect 85740 8596 85788 8652
rect 85844 8596 85892 8652
rect 85948 8596 85958 8652
rect 94258 8596 94268 8652
rect 94324 8596 94372 8652
rect 94428 8596 94476 8652
rect 94532 8596 94580 8652
rect 94636 8596 94684 8652
rect 94740 8596 94788 8652
rect 94844 8596 94892 8652
rect 94948 8596 94958 8652
rect 99200 8372 100000 8400
rect 49858 8316 49868 8372
rect 49924 8316 50316 8372
rect 50372 8316 50382 8372
rect 56130 8316 56140 8372
rect 56196 8316 57820 8372
rect 57876 8316 57886 8372
rect 58818 8316 58828 8372
rect 58884 8316 62412 8372
rect 62468 8316 62478 8372
rect 88946 8316 88956 8372
rect 89012 8316 90748 8372
rect 90804 8316 90814 8372
rect 97682 8316 97692 8372
rect 97748 8316 100000 8372
rect 99200 8288 100000 8316
rect 46274 8204 46284 8260
rect 46340 8204 48748 8260
rect 48804 8204 48814 8260
rect 61954 8204 61964 8260
rect 62020 8204 66220 8260
rect 66276 8204 66286 8260
rect 34290 8092 34300 8148
rect 34356 8092 37436 8148
rect 37492 8092 37502 8148
rect 44034 8092 44044 8148
rect 44100 8092 44828 8148
rect 44884 8092 44894 8148
rect 46162 8092 46172 8148
rect 46228 8092 54684 8148
rect 54740 8092 54750 8148
rect 71026 8092 71036 8148
rect 71092 8092 76412 8148
rect 76468 8092 76478 8148
rect 46274 7980 46284 8036
rect 46340 7980 48972 8036
rect 49028 7980 49038 8036
rect 63074 7980 63084 8036
rect 63140 7980 72828 8036
rect 72884 7980 72894 8036
rect 66210 7868 66220 7924
rect 66276 7868 70812 7924
rect 70868 7868 70878 7924
rect 8758 7812 8768 7868
rect 8824 7812 8872 7868
rect 8928 7812 8976 7868
rect 9032 7812 9080 7868
rect 9136 7812 9184 7868
rect 9240 7812 9288 7868
rect 9344 7812 9392 7868
rect 9448 7812 9458 7868
rect 17758 7812 17768 7868
rect 17824 7812 17872 7868
rect 17928 7812 17976 7868
rect 18032 7812 18080 7868
rect 18136 7812 18184 7868
rect 18240 7812 18288 7868
rect 18344 7812 18392 7868
rect 18448 7812 18458 7868
rect 26758 7812 26768 7868
rect 26824 7812 26872 7868
rect 26928 7812 26976 7868
rect 27032 7812 27080 7868
rect 27136 7812 27184 7868
rect 27240 7812 27288 7868
rect 27344 7812 27392 7868
rect 27448 7812 27458 7868
rect 35758 7812 35768 7868
rect 35824 7812 35872 7868
rect 35928 7812 35976 7868
rect 36032 7812 36080 7868
rect 36136 7812 36184 7868
rect 36240 7812 36288 7868
rect 36344 7812 36392 7868
rect 36448 7812 36458 7868
rect 44758 7812 44768 7868
rect 44824 7812 44872 7868
rect 44928 7812 44976 7868
rect 45032 7812 45080 7868
rect 45136 7812 45184 7868
rect 45240 7812 45288 7868
rect 45344 7812 45392 7868
rect 45448 7812 45458 7868
rect 53758 7812 53768 7868
rect 53824 7812 53872 7868
rect 53928 7812 53976 7868
rect 54032 7812 54080 7868
rect 54136 7812 54184 7868
rect 54240 7812 54288 7868
rect 54344 7812 54392 7868
rect 54448 7812 54458 7868
rect 62758 7812 62768 7868
rect 62824 7812 62872 7868
rect 62928 7812 62976 7868
rect 63032 7812 63080 7868
rect 63136 7812 63184 7868
rect 63240 7812 63288 7868
rect 63344 7812 63392 7868
rect 63448 7812 63458 7868
rect 71758 7812 71768 7868
rect 71824 7812 71872 7868
rect 71928 7812 71976 7868
rect 72032 7812 72080 7868
rect 72136 7812 72184 7868
rect 72240 7812 72288 7868
rect 72344 7812 72392 7868
rect 72448 7812 72458 7868
rect 80758 7812 80768 7868
rect 80824 7812 80872 7868
rect 80928 7812 80976 7868
rect 81032 7812 81080 7868
rect 81136 7812 81184 7868
rect 81240 7812 81288 7868
rect 81344 7812 81392 7868
rect 81448 7812 81458 7868
rect 89758 7812 89768 7868
rect 89824 7812 89872 7868
rect 89928 7812 89976 7868
rect 90032 7812 90080 7868
rect 90136 7812 90184 7868
rect 90240 7812 90288 7868
rect 90344 7812 90392 7868
rect 90448 7812 90458 7868
rect 50194 7756 50204 7812
rect 50260 7756 50428 7812
rect 48850 7644 48860 7700
rect 48916 7644 49868 7700
rect 49924 7644 49934 7700
rect 34626 7532 34636 7588
rect 34692 7532 37212 7588
rect 37268 7532 37278 7588
rect 0 7392 800 7504
rect 32498 7420 32508 7476
rect 32564 7420 35084 7476
rect 35140 7420 35150 7476
rect 38612 7420 42140 7476
rect 42196 7420 42206 7476
rect 38612 7364 38668 7420
rect 38322 7308 38332 7364
rect 38388 7308 38668 7364
rect 44146 7308 44156 7364
rect 44212 7308 48076 7364
rect 48132 7308 48142 7364
rect 41010 7196 41020 7252
rect 41076 7196 42364 7252
rect 42420 7196 42430 7252
rect 4258 7028 4268 7084
rect 4324 7028 4372 7084
rect 4428 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4788 7084
rect 4844 7028 4892 7084
rect 4948 7028 4958 7084
rect 13258 7028 13268 7084
rect 13324 7028 13372 7084
rect 13428 7028 13476 7084
rect 13532 7028 13580 7084
rect 13636 7028 13684 7084
rect 13740 7028 13788 7084
rect 13844 7028 13892 7084
rect 13948 7028 13958 7084
rect 22258 7028 22268 7084
rect 22324 7028 22372 7084
rect 22428 7028 22476 7084
rect 22532 7028 22580 7084
rect 22636 7028 22684 7084
rect 22740 7028 22788 7084
rect 22844 7028 22892 7084
rect 22948 7028 22958 7084
rect 31258 7028 31268 7084
rect 31324 7028 31372 7084
rect 31428 7028 31476 7084
rect 31532 7028 31580 7084
rect 31636 7028 31684 7084
rect 31740 7028 31788 7084
rect 31844 7028 31892 7084
rect 31948 7028 31958 7084
rect 40258 7028 40268 7084
rect 40324 7028 40372 7084
rect 40428 7028 40476 7084
rect 40532 7028 40580 7084
rect 40636 7028 40684 7084
rect 40740 7028 40788 7084
rect 40844 7028 40892 7084
rect 40948 7028 40958 7084
rect 49258 7028 49268 7084
rect 49324 7028 49372 7084
rect 49428 7028 49476 7084
rect 49532 7028 49580 7084
rect 49636 7028 49684 7084
rect 49740 7028 49788 7084
rect 49844 7028 49892 7084
rect 49948 7028 49958 7084
rect 34738 6860 34748 6916
rect 34804 6860 37324 6916
rect 37380 6860 37390 6916
rect 48626 6860 48636 6916
rect 48692 6860 49084 6916
rect 49140 6860 49150 6916
rect 50372 6804 50428 7756
rect 51202 7644 51212 7700
rect 51268 7644 54684 7700
rect 54740 7644 54750 7700
rect 51874 7532 51884 7588
rect 51940 7532 55412 7588
rect 59154 7532 59164 7588
rect 59220 7532 66444 7588
rect 66500 7532 66510 7588
rect 55356 7476 55412 7532
rect 51986 7420 51996 7476
rect 52052 7420 52780 7476
rect 52836 7420 52846 7476
rect 55346 7420 55356 7476
rect 55412 7420 56588 7476
rect 56644 7420 56654 7476
rect 77186 7420 77196 7476
rect 77252 7420 83916 7476
rect 83972 7420 83982 7476
rect 61170 7084 61180 7140
rect 61236 7084 64428 7140
rect 64484 7084 64494 7140
rect 68114 7084 68124 7140
rect 68180 7084 73948 7140
rect 58258 7028 58268 7084
rect 58324 7028 58372 7084
rect 58428 7028 58476 7084
rect 58532 7028 58580 7084
rect 58636 7028 58684 7084
rect 58740 7028 58788 7084
rect 58844 7028 58892 7084
rect 58948 7028 58958 7084
rect 67258 7028 67268 7084
rect 67324 7028 67372 7084
rect 67428 7028 67476 7084
rect 67532 7028 67580 7084
rect 67636 7028 67684 7084
rect 67740 7028 67788 7084
rect 67844 7028 67892 7084
rect 67948 7028 67958 7084
rect 70130 6972 70140 7028
rect 70196 6972 70206 7028
rect 70140 6804 70196 6972
rect 73892 6916 73948 7084
rect 76258 7028 76268 7084
rect 76324 7028 76372 7084
rect 76428 7028 76476 7084
rect 76532 7028 76580 7084
rect 76636 7028 76684 7084
rect 76740 7028 76788 7084
rect 76844 7028 76892 7084
rect 76948 7028 76958 7084
rect 85258 7028 85268 7084
rect 85324 7028 85372 7084
rect 85428 7028 85476 7084
rect 85532 7028 85580 7084
rect 85636 7028 85684 7084
rect 85740 7028 85788 7084
rect 85844 7028 85892 7084
rect 85948 7028 85958 7084
rect 94258 7028 94268 7084
rect 94324 7028 94372 7084
rect 94428 7028 94476 7084
rect 94532 7028 94580 7084
rect 94636 7028 94684 7084
rect 94740 7028 94788 7084
rect 94844 7028 94892 7084
rect 94948 7028 94958 7084
rect 73892 6860 74620 6916
rect 74676 6860 74686 6916
rect 33506 6748 33516 6804
rect 33572 6748 33964 6804
rect 34020 6748 34030 6804
rect 40114 6748 40124 6804
rect 40180 6748 41916 6804
rect 41972 6748 47068 6804
rect 47124 6748 47134 6804
rect 50372 6748 58828 6804
rect 58884 6748 58894 6804
rect 70140 6748 77084 6804
rect 77140 6748 77150 6804
rect 81666 6748 81676 6804
rect 81732 6748 87948 6804
rect 88004 6748 88014 6804
rect 25106 6636 25116 6692
rect 25172 6636 25900 6692
rect 25956 6636 25966 6692
rect 28354 6636 28364 6692
rect 28420 6636 30716 6692
rect 30772 6636 30782 6692
rect 40898 6636 40908 6692
rect 40964 6636 45388 6692
rect 45444 6636 45454 6692
rect 45826 6636 45836 6692
rect 45892 6636 50092 6692
rect 50148 6636 50158 6692
rect 58034 6636 58044 6692
rect 58100 6636 60508 6692
rect 60564 6636 60574 6692
rect 62132 6636 62412 6692
rect 62468 6636 62478 6692
rect 62626 6636 62636 6692
rect 62692 6636 65548 6692
rect 65604 6636 65614 6692
rect 71138 6636 71148 6692
rect 71204 6636 73948 6692
rect 74004 6636 74014 6692
rect 78932 6636 82124 6692
rect 82180 6636 82190 6692
rect 82674 6636 82684 6692
rect 82740 6636 84028 6692
rect 84084 6636 84094 6692
rect 90514 6636 90524 6692
rect 90580 6636 96684 6692
rect 96740 6636 96750 6692
rect 62132 6580 62188 6636
rect 34402 6524 34412 6580
rect 34468 6524 41244 6580
rect 41300 6524 41310 6580
rect 49970 6524 49980 6580
rect 50036 6524 54908 6580
rect 54964 6524 54974 6580
rect 59042 6524 59052 6580
rect 59108 6524 62188 6580
rect 65426 6524 65436 6580
rect 65492 6524 69020 6580
rect 69076 6524 69086 6580
rect 75506 6524 75516 6580
rect 75572 6524 78204 6580
rect 78260 6524 78270 6580
rect 26786 6412 26796 6468
rect 26852 6412 29372 6468
rect 29428 6412 41468 6468
rect 41524 6412 41534 6468
rect 45378 6412 45388 6468
rect 45444 6412 46060 6468
rect 46116 6412 46126 6468
rect 49298 6412 49308 6468
rect 49364 6412 53788 6468
rect 53844 6412 53854 6468
rect 70812 6412 71596 6468
rect 71652 6412 73948 6468
rect 74004 6412 74014 6468
rect 74498 6412 74508 6468
rect 74564 6412 75404 6468
rect 75460 6412 75470 6468
rect 0 6356 800 6384
rect 0 6300 1708 6356
rect 1764 6300 1774 6356
rect 27580 6300 34972 6356
rect 35028 6300 35038 6356
rect 59826 6300 59836 6356
rect 59892 6300 62188 6356
rect 62244 6300 62254 6356
rect 0 6272 800 6300
rect 8758 6244 8768 6300
rect 8824 6244 8872 6300
rect 8928 6244 8976 6300
rect 9032 6244 9080 6300
rect 9136 6244 9184 6300
rect 9240 6244 9288 6300
rect 9344 6244 9392 6300
rect 9448 6244 9458 6300
rect 17758 6244 17768 6300
rect 17824 6244 17872 6300
rect 17928 6244 17976 6300
rect 18032 6244 18080 6300
rect 18136 6244 18184 6300
rect 18240 6244 18288 6300
rect 18344 6244 18392 6300
rect 18448 6244 18458 6300
rect 26758 6244 26768 6300
rect 26824 6244 26872 6300
rect 26928 6244 26976 6300
rect 27032 6244 27080 6300
rect 27136 6244 27184 6300
rect 27240 6244 27288 6300
rect 27344 6244 27392 6300
rect 27448 6244 27458 6300
rect 27580 6132 27636 6300
rect 35758 6244 35768 6300
rect 35824 6244 35872 6300
rect 35928 6244 35976 6300
rect 36032 6244 36080 6300
rect 36136 6244 36184 6300
rect 36240 6244 36288 6300
rect 36344 6244 36392 6300
rect 36448 6244 36458 6300
rect 44758 6244 44768 6300
rect 44824 6244 44872 6300
rect 44928 6244 44976 6300
rect 45032 6244 45080 6300
rect 45136 6244 45184 6300
rect 45240 6244 45288 6300
rect 45344 6244 45392 6300
rect 45448 6244 45458 6300
rect 53758 6244 53768 6300
rect 53824 6244 53872 6300
rect 53928 6244 53976 6300
rect 54032 6244 54080 6300
rect 54136 6244 54184 6300
rect 54240 6244 54288 6300
rect 54344 6244 54392 6300
rect 54448 6244 54458 6300
rect 62758 6244 62768 6300
rect 62824 6244 62872 6300
rect 62928 6244 62976 6300
rect 63032 6244 63080 6300
rect 63136 6244 63184 6300
rect 63240 6244 63288 6300
rect 63344 6244 63392 6300
rect 63448 6244 63458 6300
rect 70812 6244 70868 6412
rect 71758 6244 71768 6300
rect 71824 6244 71872 6300
rect 71928 6244 71976 6300
rect 72032 6244 72080 6300
rect 72136 6244 72184 6300
rect 72240 6244 72288 6300
rect 72344 6244 72392 6300
rect 72448 6244 72458 6300
rect 33730 6188 33740 6244
rect 33796 6188 34300 6244
rect 34356 6188 34366 6244
rect 70802 6188 70812 6244
rect 70868 6188 70878 6244
rect 78932 6132 78988 6636
rect 99200 6580 100000 6608
rect 81778 6524 81788 6580
rect 81844 6524 86156 6580
rect 86212 6524 86222 6580
rect 98018 6524 98028 6580
rect 98084 6524 100000 6580
rect 99200 6496 100000 6524
rect 81666 6412 81676 6468
rect 81732 6412 82348 6468
rect 82404 6412 82414 6468
rect 80758 6244 80768 6300
rect 80824 6244 80872 6300
rect 80928 6244 80976 6300
rect 81032 6244 81080 6300
rect 81136 6244 81184 6300
rect 81240 6244 81288 6300
rect 81344 6244 81392 6300
rect 81448 6244 81458 6300
rect 89758 6244 89768 6300
rect 89824 6244 89872 6300
rect 89928 6244 89976 6300
rect 90032 6244 90080 6300
rect 90136 6244 90184 6300
rect 90240 6244 90288 6300
rect 90344 6244 90392 6300
rect 90448 6244 90458 6300
rect 2258 6076 2268 6132
rect 2324 6076 27636 6132
rect 33842 6076 33852 6132
rect 33908 6076 33918 6132
rect 41682 6076 41692 6132
rect 41748 6076 42028 6132
rect 42084 6076 42588 6132
rect 42644 6076 44940 6132
rect 44996 6076 48860 6132
rect 48916 6076 48926 6132
rect 50082 6076 50092 6132
rect 50148 6076 50428 6132
rect 50484 6076 50494 6132
rect 71698 6076 71708 6132
rect 71764 6076 74844 6132
rect 74900 6076 74910 6132
rect 78530 6076 78540 6132
rect 78596 6076 78988 6132
rect 33852 6020 33908 6076
rect 8372 5964 33908 6020
rect 35634 5964 35644 6020
rect 35700 5964 46396 6020
rect 46452 5964 46462 6020
rect 69682 5964 69692 6020
rect 69748 5964 72492 6020
rect 72548 5964 76188 6020
rect 76244 5964 76254 6020
rect 8372 5796 8428 5964
rect 33394 5852 33404 5908
rect 33460 5852 33852 5908
rect 33908 5852 33918 5908
rect 48178 5852 48188 5908
rect 48244 5852 54572 5908
rect 54628 5852 54638 5908
rect 78932 5852 80108 5908
rect 80164 5852 80174 5908
rect 78932 5796 78988 5852
rect 2258 5740 2268 5796
rect 2324 5740 8428 5796
rect 70802 5740 70812 5796
rect 70868 5740 78988 5796
rect 46274 5628 46284 5684
rect 46340 5628 48972 5684
rect 49028 5628 49038 5684
rect 70914 5628 70924 5684
rect 70980 5628 72604 5684
rect 72660 5628 72670 5684
rect 4258 5460 4268 5516
rect 4324 5460 4372 5516
rect 4428 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4788 5516
rect 4844 5460 4892 5516
rect 4948 5460 4958 5516
rect 13258 5460 13268 5516
rect 13324 5460 13372 5516
rect 13428 5460 13476 5516
rect 13532 5460 13580 5516
rect 13636 5460 13684 5516
rect 13740 5460 13788 5516
rect 13844 5460 13892 5516
rect 13948 5460 13958 5516
rect 22258 5460 22268 5516
rect 22324 5460 22372 5516
rect 22428 5460 22476 5516
rect 22532 5460 22580 5516
rect 22636 5460 22684 5516
rect 22740 5460 22788 5516
rect 22844 5460 22892 5516
rect 22948 5460 22958 5516
rect 31258 5460 31268 5516
rect 31324 5460 31372 5516
rect 31428 5460 31476 5516
rect 31532 5460 31580 5516
rect 31636 5460 31684 5516
rect 31740 5460 31788 5516
rect 31844 5460 31892 5516
rect 31948 5460 31958 5516
rect 40258 5460 40268 5516
rect 40324 5460 40372 5516
rect 40428 5460 40476 5516
rect 40532 5460 40580 5516
rect 40636 5460 40684 5516
rect 40740 5460 40788 5516
rect 40844 5460 40892 5516
rect 40948 5460 40958 5516
rect 49258 5460 49268 5516
rect 49324 5460 49372 5516
rect 49428 5460 49476 5516
rect 49532 5460 49580 5516
rect 49636 5460 49684 5516
rect 49740 5460 49788 5516
rect 49844 5460 49892 5516
rect 49948 5460 49958 5516
rect 58258 5460 58268 5516
rect 58324 5460 58372 5516
rect 58428 5460 58476 5516
rect 58532 5460 58580 5516
rect 58636 5460 58684 5516
rect 58740 5460 58788 5516
rect 58844 5460 58892 5516
rect 58948 5460 58958 5516
rect 67258 5460 67268 5516
rect 67324 5460 67372 5516
rect 67428 5460 67476 5516
rect 67532 5460 67580 5516
rect 67636 5460 67684 5516
rect 67740 5460 67788 5516
rect 67844 5460 67892 5516
rect 67948 5460 67958 5516
rect 76258 5460 76268 5516
rect 76324 5460 76372 5516
rect 76428 5460 76476 5516
rect 76532 5460 76580 5516
rect 76636 5460 76684 5516
rect 76740 5460 76788 5516
rect 76844 5460 76892 5516
rect 76948 5460 76958 5516
rect 85258 5460 85268 5516
rect 85324 5460 85372 5516
rect 85428 5460 85476 5516
rect 85532 5460 85580 5516
rect 85636 5460 85684 5516
rect 85740 5460 85788 5516
rect 85844 5460 85892 5516
rect 85948 5460 85958 5516
rect 94258 5460 94268 5516
rect 94324 5460 94372 5516
rect 94428 5460 94476 5516
rect 94532 5460 94580 5516
rect 94636 5460 94684 5516
rect 94740 5460 94788 5516
rect 94844 5460 94892 5516
rect 94948 5460 94958 5516
rect 34962 5404 34972 5460
rect 35028 5404 36540 5460
rect 36596 5404 37996 5460
rect 38052 5404 38780 5460
rect 38836 5404 38846 5460
rect 70700 5404 74508 5460
rect 74564 5404 74574 5460
rect 77298 5404 77308 5460
rect 77364 5404 77980 5460
rect 78036 5404 78046 5460
rect 80434 5404 80444 5460
rect 80500 5404 82628 5460
rect 33282 5292 33292 5348
rect 33348 5292 35420 5348
rect 35476 5292 35486 5348
rect 36418 5292 36428 5348
rect 36484 5292 42308 5348
rect 53442 5292 53452 5348
rect 53508 5292 57428 5348
rect 57922 5292 57932 5348
rect 57988 5292 58716 5348
rect 58772 5292 64652 5348
rect 64708 5292 64718 5348
rect 0 5236 800 5264
rect 42252 5236 42308 5292
rect 57372 5236 57428 5292
rect 0 5180 1820 5236
rect 1876 5180 1886 5236
rect 26562 5180 26572 5236
rect 26628 5180 34076 5236
rect 34132 5180 34142 5236
rect 34402 5180 34412 5236
rect 34468 5180 41692 5236
rect 41748 5180 41758 5236
rect 42242 5180 42252 5236
rect 42308 5180 42924 5236
rect 42980 5180 42990 5236
rect 44370 5180 44380 5236
rect 44436 5180 44940 5236
rect 44996 5180 45006 5236
rect 51762 5180 51772 5236
rect 51828 5180 53228 5236
rect 53284 5180 57148 5236
rect 57204 5180 57214 5236
rect 57372 5180 60732 5236
rect 60788 5180 60798 5236
rect 0 5152 800 5180
rect 27906 5068 27916 5124
rect 27972 5068 34748 5124
rect 34804 5068 34814 5124
rect 41906 5068 41916 5124
rect 41972 5068 42812 5124
rect 42868 5068 42878 5124
rect 48290 5068 48300 5124
rect 48356 5068 49868 5124
rect 49924 5068 49934 5124
rect 59154 5068 59164 5124
rect 59220 5068 68348 5124
rect 68404 5068 68414 5124
rect 30146 4956 30156 5012
rect 30212 4956 33852 5012
rect 33908 4956 33918 5012
rect 39218 4956 39228 5012
rect 39284 4956 42476 5012
rect 42532 4956 42542 5012
rect 45266 4956 45276 5012
rect 45332 4956 49420 5012
rect 49476 4956 49486 5012
rect 59574 4956 59612 5012
rect 59668 4956 59678 5012
rect 62132 4956 67340 5012
rect 67396 4956 68236 5012
rect 68292 4956 70028 5012
rect 70084 4956 70094 5012
rect 62132 4900 62188 4956
rect 70700 4900 70756 5404
rect 82572 5348 82628 5404
rect 71362 5292 71372 5348
rect 71428 5292 81564 5348
rect 81620 5292 81630 5348
rect 82572 5292 96572 5348
rect 96628 5292 96638 5348
rect 74498 5180 74508 5236
rect 74564 5180 80668 5236
rect 80724 5180 82124 5236
rect 82180 5180 84700 5236
rect 84756 5180 84766 5236
rect 73714 5068 73724 5124
rect 73780 5068 81676 5124
rect 81732 5068 81742 5124
rect 81890 5068 81900 5124
rect 81956 5068 82460 5124
rect 82516 5068 82526 5124
rect 41570 4844 41580 4900
rect 41636 4844 43484 4900
rect 43540 4844 43550 4900
rect 46610 4844 46620 4900
rect 46676 4844 50764 4900
rect 50820 4844 50830 4900
rect 59378 4844 59388 4900
rect 59444 4844 62188 4900
rect 62636 4844 70700 4900
rect 70756 4844 70766 4900
rect 41458 4732 41468 4788
rect 41524 4732 42140 4788
rect 42196 4732 42206 4788
rect 44594 4732 44604 4788
rect 44660 4732 44670 4788
rect 8758 4676 8768 4732
rect 8824 4676 8872 4732
rect 8928 4676 8976 4732
rect 9032 4676 9080 4732
rect 9136 4676 9184 4732
rect 9240 4676 9288 4732
rect 9344 4676 9392 4732
rect 9448 4676 9458 4732
rect 17758 4676 17768 4732
rect 17824 4676 17872 4732
rect 17928 4676 17976 4732
rect 18032 4676 18080 4732
rect 18136 4676 18184 4732
rect 18240 4676 18288 4732
rect 18344 4676 18392 4732
rect 18448 4676 18458 4732
rect 26758 4676 26768 4732
rect 26824 4676 26872 4732
rect 26928 4676 26976 4732
rect 27032 4676 27080 4732
rect 27136 4676 27184 4732
rect 27240 4676 27288 4732
rect 27344 4676 27392 4732
rect 27448 4676 27458 4732
rect 35758 4676 35768 4732
rect 35824 4676 35872 4732
rect 35928 4676 35976 4732
rect 36032 4676 36080 4732
rect 36136 4676 36184 4732
rect 36240 4676 36288 4732
rect 36344 4676 36392 4732
rect 36448 4676 36458 4732
rect 44604 4676 44660 4732
rect 44758 4676 44768 4732
rect 44824 4676 44872 4732
rect 44928 4676 44976 4732
rect 45032 4676 45080 4732
rect 45136 4676 45184 4732
rect 45240 4676 45288 4732
rect 45344 4676 45392 4732
rect 45448 4676 45458 4732
rect 53758 4676 53768 4732
rect 53824 4676 53872 4732
rect 53928 4676 53976 4732
rect 54032 4676 54080 4732
rect 54136 4676 54184 4732
rect 54240 4676 54288 4732
rect 54344 4676 54392 4732
rect 54448 4676 54458 4732
rect 62636 4676 62692 4844
rect 99200 4788 100000 4816
rect 97682 4732 97692 4788
rect 97748 4732 100000 4788
rect 62758 4676 62768 4732
rect 62824 4676 62872 4732
rect 62928 4676 62976 4732
rect 63032 4676 63080 4732
rect 63136 4676 63184 4732
rect 63240 4676 63288 4732
rect 63344 4676 63392 4732
rect 63448 4676 63458 4732
rect 71758 4676 71768 4732
rect 71824 4676 71872 4732
rect 71928 4676 71976 4732
rect 72032 4676 72080 4732
rect 72136 4676 72184 4732
rect 72240 4676 72288 4732
rect 72344 4676 72392 4732
rect 72448 4676 72458 4732
rect 80758 4676 80768 4732
rect 80824 4676 80872 4732
rect 80928 4676 80976 4732
rect 81032 4676 81080 4732
rect 81136 4676 81184 4732
rect 81240 4676 81288 4732
rect 81344 4676 81392 4732
rect 81448 4676 81458 4732
rect 89758 4676 89768 4732
rect 89824 4676 89872 4732
rect 89928 4676 89976 4732
rect 90032 4676 90080 4732
rect 90136 4676 90184 4732
rect 90240 4676 90288 4732
rect 90344 4676 90392 4732
rect 90448 4676 90458 4732
rect 99200 4704 100000 4732
rect 38612 4620 41132 4676
rect 41188 4620 41198 4676
rect 41570 4620 41580 4676
rect 41636 4620 44660 4676
rect 62132 4620 62692 4676
rect 38612 4564 38668 4620
rect 62132 4564 62188 4620
rect 30156 4508 38668 4564
rect 40114 4508 40124 4564
rect 40180 4508 42364 4564
rect 42420 4508 42430 4564
rect 50372 4508 52332 4564
rect 52388 4508 62188 4564
rect 63186 4508 63196 4564
rect 63252 4508 65324 4564
rect 65380 4508 65390 4564
rect 73892 4508 79996 4564
rect 80052 4508 80062 4564
rect 86258 4508 86268 4564
rect 86324 4508 96684 4564
rect 96740 4508 96750 4564
rect 30156 4452 30212 4508
rect 50372 4452 50428 4508
rect 73892 4452 73948 4508
rect 30146 4396 30156 4452
rect 30212 4396 30222 4452
rect 38322 4396 38332 4452
rect 38388 4396 43148 4452
rect 43204 4396 43214 4452
rect 49746 4396 49756 4452
rect 49812 4396 49980 4452
rect 50036 4396 50204 4452
rect 50260 4396 50428 4452
rect 52770 4396 52780 4452
rect 52836 4396 52846 4452
rect 62300 4396 62748 4452
rect 62804 4396 73948 4452
rect 75590 4396 75628 4452
rect 75684 4396 75694 4452
rect 75852 4396 78316 4452
rect 78372 4396 78876 4452
rect 78932 4396 78942 4452
rect 52780 4340 52836 4396
rect 62300 4340 62356 4396
rect 75852 4340 75908 4396
rect 32498 4284 32508 4340
rect 32564 4284 33852 4340
rect 33908 4284 34188 4340
rect 34244 4284 34254 4340
rect 34626 4284 34636 4340
rect 34692 4284 35196 4340
rect 35252 4284 35262 4340
rect 40226 4284 40236 4340
rect 40292 4284 43820 4340
rect 43876 4284 43886 4340
rect 48178 4284 48188 4340
rect 48244 4284 52836 4340
rect 59266 4284 59276 4340
rect 59332 4284 62356 4340
rect 73266 4284 73276 4340
rect 73332 4284 75908 4340
rect 77858 4284 77868 4340
rect 77924 4284 79436 4340
rect 79492 4284 79502 4340
rect 34636 4228 34692 4284
rect 33058 4172 33068 4228
rect 33124 4172 34692 4228
rect 41122 4172 41132 4228
rect 41188 4172 41804 4228
rect 41860 4172 41870 4228
rect 60274 4172 60284 4228
rect 60340 4172 62188 4228
rect 62244 4172 62254 4228
rect 71698 4172 71708 4228
rect 71764 4172 75292 4228
rect 75348 4172 75358 4228
rect 77634 4172 77644 4228
rect 77700 4172 79212 4228
rect 79268 4172 79278 4228
rect 85922 4172 85932 4228
rect 85988 4172 86156 4228
rect 86212 4172 86222 4228
rect 0 4116 800 4144
rect 0 4060 20748 4116
rect 20804 4060 20814 4116
rect 38770 4060 38780 4116
rect 38836 4060 42028 4116
rect 42084 4060 42094 4116
rect 48514 4060 48524 4116
rect 48580 4060 49196 4116
rect 49252 4060 51436 4116
rect 51492 4060 57484 4116
rect 57540 4060 59388 4116
rect 59444 4060 59454 4116
rect 70018 4060 70028 4116
rect 70084 4060 71596 4116
rect 71652 4060 73948 4116
rect 74386 4060 74396 4116
rect 74452 4060 78876 4116
rect 78932 4060 78942 4116
rect 0 4032 800 4060
rect 4258 3892 4268 3948
rect 4324 3892 4372 3948
rect 4428 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4788 3948
rect 4844 3892 4892 3948
rect 4948 3892 4958 3948
rect 13258 3892 13268 3948
rect 13324 3892 13372 3948
rect 13428 3892 13476 3948
rect 13532 3892 13580 3948
rect 13636 3892 13684 3948
rect 13740 3892 13788 3948
rect 13844 3892 13892 3948
rect 13948 3892 13958 3948
rect 22258 3892 22268 3948
rect 22324 3892 22372 3948
rect 22428 3892 22476 3948
rect 22532 3892 22580 3948
rect 22636 3892 22684 3948
rect 22740 3892 22788 3948
rect 22844 3892 22892 3948
rect 22948 3892 22958 3948
rect 31258 3892 31268 3948
rect 31324 3892 31372 3948
rect 31428 3892 31476 3948
rect 31532 3892 31580 3948
rect 31636 3892 31684 3948
rect 31740 3892 31788 3948
rect 31844 3892 31892 3948
rect 31948 3892 31958 3948
rect 40258 3892 40268 3948
rect 40324 3892 40372 3948
rect 40428 3892 40476 3948
rect 40532 3892 40580 3948
rect 40636 3892 40684 3948
rect 40740 3892 40788 3948
rect 40844 3892 40892 3948
rect 40948 3892 40958 3948
rect 49258 3892 49268 3948
rect 49324 3892 49372 3948
rect 49428 3892 49476 3948
rect 49532 3892 49580 3948
rect 49636 3892 49684 3948
rect 49740 3892 49788 3948
rect 49844 3892 49892 3948
rect 49948 3892 49958 3948
rect 58258 3892 58268 3948
rect 58324 3892 58372 3948
rect 58428 3892 58476 3948
rect 58532 3892 58580 3948
rect 58636 3892 58684 3948
rect 58740 3892 58788 3948
rect 58844 3892 58892 3948
rect 58948 3892 58958 3948
rect 67258 3892 67268 3948
rect 67324 3892 67372 3948
rect 67428 3892 67476 3948
rect 67532 3892 67580 3948
rect 67636 3892 67684 3948
rect 67740 3892 67788 3948
rect 67844 3892 67892 3948
rect 67948 3892 67958 3948
rect 38210 3836 38220 3892
rect 38276 3836 38286 3892
rect 60162 3836 60172 3892
rect 60228 3836 61740 3892
rect 61796 3836 61806 3892
rect 25890 3724 25900 3780
rect 25956 3724 28812 3780
rect 28868 3724 33292 3780
rect 33348 3724 33358 3780
rect 38220 3668 38276 3836
rect 17826 3612 17836 3668
rect 17892 3612 38276 3668
rect 38332 3724 39116 3780
rect 39172 3724 41020 3780
rect 41076 3724 41468 3780
rect 41524 3724 42252 3780
rect 42308 3724 42318 3780
rect 42578 3724 42588 3780
rect 42644 3724 45276 3780
rect 45332 3724 45342 3780
rect 50194 3724 50204 3780
rect 50260 3724 50428 3780
rect 56690 3724 56700 3780
rect 56756 3724 59052 3780
rect 59108 3724 59118 3780
rect 60834 3724 60844 3780
rect 60900 3724 63532 3780
rect 63588 3724 63598 3780
rect 68450 3724 68460 3780
rect 68516 3724 69580 3780
rect 69636 3724 69646 3780
rect 38332 3556 38388 3724
rect 50372 3668 50428 3724
rect 73892 3668 73948 4060
rect 76258 3892 76268 3948
rect 76324 3892 76372 3948
rect 76428 3892 76476 3948
rect 76532 3892 76580 3948
rect 76636 3892 76684 3948
rect 76740 3892 76788 3948
rect 76844 3892 76892 3948
rect 76948 3892 76958 3948
rect 85258 3892 85268 3948
rect 85324 3892 85372 3948
rect 85428 3892 85476 3948
rect 85532 3892 85580 3948
rect 85636 3892 85684 3948
rect 85740 3892 85788 3948
rect 85844 3892 85892 3948
rect 85948 3892 85958 3948
rect 94258 3892 94268 3948
rect 94324 3892 94372 3948
rect 94428 3892 94476 3948
rect 94532 3892 94580 3948
rect 94636 3892 94684 3948
rect 94740 3892 94788 3948
rect 94844 3892 94892 3948
rect 94948 3892 94958 3948
rect 74946 3724 74956 3780
rect 75012 3724 96348 3780
rect 96404 3724 96908 3780
rect 96964 3724 96974 3780
rect 38658 3612 38668 3668
rect 38724 3612 40908 3668
rect 40964 3612 40974 3668
rect 50372 3612 52444 3668
rect 52500 3612 55468 3668
rect 55524 3612 55534 3668
rect 58156 3612 59836 3668
rect 59892 3612 60732 3668
rect 60788 3612 62748 3668
rect 62804 3612 62814 3668
rect 70354 3612 70364 3668
rect 70420 3612 71036 3668
rect 71092 3612 71102 3668
rect 73892 3612 74284 3668
rect 74340 3612 78092 3668
rect 78148 3612 78158 3668
rect 83234 3612 83244 3668
rect 83300 3612 94164 3668
rect 58156 3556 58212 3612
rect 31714 3500 31724 3556
rect 31780 3500 32508 3556
rect 32564 3500 32574 3556
rect 34738 3500 34748 3556
rect 34804 3500 36092 3556
rect 36148 3500 37436 3556
rect 37492 3500 37884 3556
rect 37940 3500 37950 3556
rect 38322 3500 38332 3556
rect 38388 3500 38398 3556
rect 40338 3500 40348 3556
rect 40404 3500 41580 3556
rect 41636 3500 41646 3556
rect 43026 3500 43036 3556
rect 43092 3500 44940 3556
rect 44996 3500 45006 3556
rect 46386 3500 46396 3556
rect 46452 3500 49308 3556
rect 49364 3500 49374 3556
rect 50418 3500 50428 3556
rect 50484 3500 54572 3556
rect 54628 3500 55020 3556
rect 55076 3500 55086 3556
rect 58146 3500 58156 3556
rect 58212 3500 58222 3556
rect 61282 3500 61292 3556
rect 61348 3500 63196 3556
rect 63252 3500 63262 3556
rect 71586 3500 71596 3556
rect 71652 3500 73948 3556
rect 82898 3500 82908 3556
rect 82964 3500 86156 3556
rect 86212 3500 86222 3556
rect 73892 3444 73948 3500
rect 94108 3444 94164 3612
rect 38546 3388 38556 3444
rect 38612 3388 39004 3444
rect 39060 3388 39788 3444
rect 39844 3388 39854 3444
rect 42578 3388 42588 3444
rect 42644 3388 42980 3444
rect 42924 3332 42980 3388
rect 43372 3388 43820 3444
rect 43876 3388 43886 3444
rect 46722 3388 46732 3444
rect 46788 3388 48860 3444
rect 48916 3388 49420 3444
rect 49476 3388 52668 3444
rect 52724 3388 67452 3444
rect 67508 3388 69692 3444
rect 69748 3388 71932 3444
rect 71988 3388 73276 3444
rect 73332 3388 73342 3444
rect 73892 3388 74396 3444
rect 74452 3388 74462 3444
rect 75842 3388 75852 3444
rect 75908 3388 83244 3444
rect 83300 3388 83310 3444
rect 94098 3388 94108 3444
rect 94164 3388 94174 3444
rect 43372 3332 43428 3388
rect 42924 3276 43428 3332
rect 43652 3276 43932 3332
rect 43988 3276 43998 3332
rect 76178 3276 76188 3332
rect 76244 3276 81900 3332
rect 81956 3276 81966 3332
rect 43652 3220 43708 3276
rect 42690 3164 42700 3220
rect 42756 3164 43708 3220
rect 8758 3108 8768 3164
rect 8824 3108 8872 3164
rect 8928 3108 8976 3164
rect 9032 3108 9080 3164
rect 9136 3108 9184 3164
rect 9240 3108 9288 3164
rect 9344 3108 9392 3164
rect 9448 3108 9458 3164
rect 17758 3108 17768 3164
rect 17824 3108 17872 3164
rect 17928 3108 17976 3164
rect 18032 3108 18080 3164
rect 18136 3108 18184 3164
rect 18240 3108 18288 3164
rect 18344 3108 18392 3164
rect 18448 3108 18458 3164
rect 26758 3108 26768 3164
rect 26824 3108 26872 3164
rect 26928 3108 26976 3164
rect 27032 3108 27080 3164
rect 27136 3108 27184 3164
rect 27240 3108 27288 3164
rect 27344 3108 27392 3164
rect 27448 3108 27458 3164
rect 35758 3108 35768 3164
rect 35824 3108 35872 3164
rect 35928 3108 35976 3164
rect 36032 3108 36080 3164
rect 36136 3108 36184 3164
rect 36240 3108 36288 3164
rect 36344 3108 36392 3164
rect 36448 3108 36458 3164
rect 44758 3108 44768 3164
rect 44824 3108 44872 3164
rect 44928 3108 44976 3164
rect 45032 3108 45080 3164
rect 45136 3108 45184 3164
rect 45240 3108 45288 3164
rect 45344 3108 45392 3164
rect 45448 3108 45458 3164
rect 53758 3108 53768 3164
rect 53824 3108 53872 3164
rect 53928 3108 53976 3164
rect 54032 3108 54080 3164
rect 54136 3108 54184 3164
rect 54240 3108 54288 3164
rect 54344 3108 54392 3164
rect 54448 3108 54458 3164
rect 62758 3108 62768 3164
rect 62824 3108 62872 3164
rect 62928 3108 62976 3164
rect 63032 3108 63080 3164
rect 63136 3108 63184 3164
rect 63240 3108 63288 3164
rect 63344 3108 63392 3164
rect 63448 3108 63458 3164
rect 71758 3108 71768 3164
rect 71824 3108 71872 3164
rect 71928 3108 71976 3164
rect 72032 3108 72080 3164
rect 72136 3108 72184 3164
rect 72240 3108 72288 3164
rect 72344 3108 72392 3164
rect 72448 3108 72458 3164
rect 80758 3108 80768 3164
rect 80824 3108 80872 3164
rect 80928 3108 80976 3164
rect 81032 3108 81080 3164
rect 81136 3108 81184 3164
rect 81240 3108 81288 3164
rect 81344 3108 81392 3164
rect 81448 3108 81458 3164
rect 89758 3108 89768 3164
rect 89824 3108 89872 3164
rect 89928 3108 89976 3164
rect 90032 3108 90080 3164
rect 90136 3108 90184 3164
rect 90240 3108 90288 3164
rect 90344 3108 90392 3164
rect 90448 3108 90458 3164
rect 99200 2996 100000 3024
rect 97682 2940 97692 2996
rect 97748 2940 100000 2996
rect 99200 2912 100000 2940
rect 99200 1204 100000 1232
rect 97794 1148 97804 1204
rect 97860 1148 100000 1204
rect 99200 1120 100000 1148
<< via3 >>
rect 8768 56420 8824 56476
rect 8872 56420 8928 56476
rect 8976 56420 9032 56476
rect 9080 56420 9136 56476
rect 9184 56420 9240 56476
rect 9288 56420 9344 56476
rect 9392 56420 9448 56476
rect 17768 56420 17824 56476
rect 17872 56420 17928 56476
rect 17976 56420 18032 56476
rect 18080 56420 18136 56476
rect 18184 56420 18240 56476
rect 18288 56420 18344 56476
rect 18392 56420 18448 56476
rect 26768 56420 26824 56476
rect 26872 56420 26928 56476
rect 26976 56420 27032 56476
rect 27080 56420 27136 56476
rect 27184 56420 27240 56476
rect 27288 56420 27344 56476
rect 27392 56420 27448 56476
rect 35768 56420 35824 56476
rect 35872 56420 35928 56476
rect 35976 56420 36032 56476
rect 36080 56420 36136 56476
rect 36184 56420 36240 56476
rect 36288 56420 36344 56476
rect 36392 56420 36448 56476
rect 44768 56420 44824 56476
rect 44872 56420 44928 56476
rect 44976 56420 45032 56476
rect 45080 56420 45136 56476
rect 45184 56420 45240 56476
rect 45288 56420 45344 56476
rect 45392 56420 45448 56476
rect 53768 56420 53824 56476
rect 53872 56420 53928 56476
rect 53976 56420 54032 56476
rect 54080 56420 54136 56476
rect 54184 56420 54240 56476
rect 54288 56420 54344 56476
rect 54392 56420 54448 56476
rect 62768 56420 62824 56476
rect 62872 56420 62928 56476
rect 62976 56420 63032 56476
rect 63080 56420 63136 56476
rect 63184 56420 63240 56476
rect 63288 56420 63344 56476
rect 63392 56420 63448 56476
rect 71768 56420 71824 56476
rect 71872 56420 71928 56476
rect 71976 56420 72032 56476
rect 72080 56420 72136 56476
rect 72184 56420 72240 56476
rect 72288 56420 72344 56476
rect 72392 56420 72448 56476
rect 80768 56420 80824 56476
rect 80872 56420 80928 56476
rect 80976 56420 81032 56476
rect 81080 56420 81136 56476
rect 81184 56420 81240 56476
rect 81288 56420 81344 56476
rect 81392 56420 81448 56476
rect 89768 56420 89824 56476
rect 89872 56420 89928 56476
rect 89976 56420 90032 56476
rect 90080 56420 90136 56476
rect 90184 56420 90240 56476
rect 90288 56420 90344 56476
rect 90392 56420 90448 56476
rect 4268 55636 4324 55692
rect 4372 55636 4428 55692
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 4788 55636 4844 55692
rect 4892 55636 4948 55692
rect 13268 55636 13324 55692
rect 13372 55636 13428 55692
rect 13476 55636 13532 55692
rect 13580 55636 13636 55692
rect 13684 55636 13740 55692
rect 13788 55636 13844 55692
rect 13892 55636 13948 55692
rect 22268 55636 22324 55692
rect 22372 55636 22428 55692
rect 22476 55636 22532 55692
rect 22580 55636 22636 55692
rect 22684 55636 22740 55692
rect 22788 55636 22844 55692
rect 22892 55636 22948 55692
rect 31268 55636 31324 55692
rect 31372 55636 31428 55692
rect 31476 55636 31532 55692
rect 31580 55636 31636 55692
rect 31684 55636 31740 55692
rect 31788 55636 31844 55692
rect 31892 55636 31948 55692
rect 40268 55636 40324 55692
rect 40372 55636 40428 55692
rect 40476 55636 40532 55692
rect 40580 55636 40636 55692
rect 40684 55636 40740 55692
rect 40788 55636 40844 55692
rect 40892 55636 40948 55692
rect 49268 55636 49324 55692
rect 49372 55636 49428 55692
rect 49476 55636 49532 55692
rect 49580 55636 49636 55692
rect 49684 55636 49740 55692
rect 49788 55636 49844 55692
rect 49892 55636 49948 55692
rect 58268 55636 58324 55692
rect 58372 55636 58428 55692
rect 58476 55636 58532 55692
rect 58580 55636 58636 55692
rect 58684 55636 58740 55692
rect 58788 55636 58844 55692
rect 58892 55636 58948 55692
rect 67268 55636 67324 55692
rect 67372 55636 67428 55692
rect 67476 55636 67532 55692
rect 67580 55636 67636 55692
rect 67684 55636 67740 55692
rect 67788 55636 67844 55692
rect 67892 55636 67948 55692
rect 76268 55636 76324 55692
rect 76372 55636 76428 55692
rect 76476 55636 76532 55692
rect 76580 55636 76636 55692
rect 76684 55636 76740 55692
rect 76788 55636 76844 55692
rect 76892 55636 76948 55692
rect 85268 55636 85324 55692
rect 85372 55636 85428 55692
rect 85476 55636 85532 55692
rect 85580 55636 85636 55692
rect 85684 55636 85740 55692
rect 85788 55636 85844 55692
rect 85892 55636 85948 55692
rect 94268 55636 94324 55692
rect 94372 55636 94428 55692
rect 94476 55636 94532 55692
rect 94580 55636 94636 55692
rect 94684 55636 94740 55692
rect 94788 55636 94844 55692
rect 94892 55636 94948 55692
rect 8768 54852 8824 54908
rect 8872 54852 8928 54908
rect 8976 54852 9032 54908
rect 9080 54852 9136 54908
rect 9184 54852 9240 54908
rect 9288 54852 9344 54908
rect 9392 54852 9448 54908
rect 17768 54852 17824 54908
rect 17872 54852 17928 54908
rect 17976 54852 18032 54908
rect 18080 54852 18136 54908
rect 18184 54852 18240 54908
rect 18288 54852 18344 54908
rect 18392 54852 18448 54908
rect 26768 54852 26824 54908
rect 26872 54852 26928 54908
rect 26976 54852 27032 54908
rect 27080 54852 27136 54908
rect 27184 54852 27240 54908
rect 27288 54852 27344 54908
rect 27392 54852 27448 54908
rect 35768 54852 35824 54908
rect 35872 54852 35928 54908
rect 35976 54852 36032 54908
rect 36080 54852 36136 54908
rect 36184 54852 36240 54908
rect 36288 54852 36344 54908
rect 36392 54852 36448 54908
rect 44768 54852 44824 54908
rect 44872 54852 44928 54908
rect 44976 54852 45032 54908
rect 45080 54852 45136 54908
rect 45184 54852 45240 54908
rect 45288 54852 45344 54908
rect 45392 54852 45448 54908
rect 53768 54852 53824 54908
rect 53872 54852 53928 54908
rect 53976 54852 54032 54908
rect 54080 54852 54136 54908
rect 54184 54852 54240 54908
rect 54288 54852 54344 54908
rect 54392 54852 54448 54908
rect 62768 54852 62824 54908
rect 62872 54852 62928 54908
rect 62976 54852 63032 54908
rect 63080 54852 63136 54908
rect 63184 54852 63240 54908
rect 63288 54852 63344 54908
rect 63392 54852 63448 54908
rect 71768 54852 71824 54908
rect 71872 54852 71928 54908
rect 71976 54852 72032 54908
rect 72080 54852 72136 54908
rect 72184 54852 72240 54908
rect 72288 54852 72344 54908
rect 72392 54852 72448 54908
rect 80768 54852 80824 54908
rect 80872 54852 80928 54908
rect 80976 54852 81032 54908
rect 81080 54852 81136 54908
rect 81184 54852 81240 54908
rect 81288 54852 81344 54908
rect 81392 54852 81448 54908
rect 89768 54852 89824 54908
rect 89872 54852 89928 54908
rect 89976 54852 90032 54908
rect 90080 54852 90136 54908
rect 90184 54852 90240 54908
rect 90288 54852 90344 54908
rect 90392 54852 90448 54908
rect 4268 54068 4324 54124
rect 4372 54068 4428 54124
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 4788 54068 4844 54124
rect 4892 54068 4948 54124
rect 13268 54068 13324 54124
rect 13372 54068 13428 54124
rect 13476 54068 13532 54124
rect 13580 54068 13636 54124
rect 13684 54068 13740 54124
rect 13788 54068 13844 54124
rect 13892 54068 13948 54124
rect 22268 54068 22324 54124
rect 22372 54068 22428 54124
rect 22476 54068 22532 54124
rect 22580 54068 22636 54124
rect 22684 54068 22740 54124
rect 22788 54068 22844 54124
rect 22892 54068 22948 54124
rect 31268 54068 31324 54124
rect 31372 54068 31428 54124
rect 31476 54068 31532 54124
rect 31580 54068 31636 54124
rect 31684 54068 31740 54124
rect 31788 54068 31844 54124
rect 31892 54068 31948 54124
rect 40268 54068 40324 54124
rect 40372 54068 40428 54124
rect 40476 54068 40532 54124
rect 40580 54068 40636 54124
rect 40684 54068 40740 54124
rect 40788 54068 40844 54124
rect 40892 54068 40948 54124
rect 49268 54068 49324 54124
rect 49372 54068 49428 54124
rect 49476 54068 49532 54124
rect 49580 54068 49636 54124
rect 49684 54068 49740 54124
rect 49788 54068 49844 54124
rect 49892 54068 49948 54124
rect 58268 54068 58324 54124
rect 58372 54068 58428 54124
rect 58476 54068 58532 54124
rect 58580 54068 58636 54124
rect 58684 54068 58740 54124
rect 58788 54068 58844 54124
rect 58892 54068 58948 54124
rect 67268 54068 67324 54124
rect 67372 54068 67428 54124
rect 67476 54068 67532 54124
rect 67580 54068 67636 54124
rect 67684 54068 67740 54124
rect 67788 54068 67844 54124
rect 67892 54068 67948 54124
rect 76268 54068 76324 54124
rect 76372 54068 76428 54124
rect 76476 54068 76532 54124
rect 76580 54068 76636 54124
rect 76684 54068 76740 54124
rect 76788 54068 76844 54124
rect 76892 54068 76948 54124
rect 85268 54068 85324 54124
rect 85372 54068 85428 54124
rect 85476 54068 85532 54124
rect 85580 54068 85636 54124
rect 85684 54068 85740 54124
rect 85788 54068 85844 54124
rect 85892 54068 85948 54124
rect 94268 54068 94324 54124
rect 94372 54068 94428 54124
rect 94476 54068 94532 54124
rect 94580 54068 94636 54124
rect 94684 54068 94740 54124
rect 94788 54068 94844 54124
rect 94892 54068 94948 54124
rect 8768 53284 8824 53340
rect 8872 53284 8928 53340
rect 8976 53284 9032 53340
rect 9080 53284 9136 53340
rect 9184 53284 9240 53340
rect 9288 53284 9344 53340
rect 9392 53284 9448 53340
rect 17768 53284 17824 53340
rect 17872 53284 17928 53340
rect 17976 53284 18032 53340
rect 18080 53284 18136 53340
rect 18184 53284 18240 53340
rect 18288 53284 18344 53340
rect 18392 53284 18448 53340
rect 26768 53284 26824 53340
rect 26872 53284 26928 53340
rect 26976 53284 27032 53340
rect 27080 53284 27136 53340
rect 27184 53284 27240 53340
rect 27288 53284 27344 53340
rect 27392 53284 27448 53340
rect 35768 53284 35824 53340
rect 35872 53284 35928 53340
rect 35976 53284 36032 53340
rect 36080 53284 36136 53340
rect 36184 53284 36240 53340
rect 36288 53284 36344 53340
rect 36392 53284 36448 53340
rect 44768 53284 44824 53340
rect 44872 53284 44928 53340
rect 44976 53284 45032 53340
rect 45080 53284 45136 53340
rect 45184 53284 45240 53340
rect 45288 53284 45344 53340
rect 45392 53284 45448 53340
rect 53768 53284 53824 53340
rect 53872 53284 53928 53340
rect 53976 53284 54032 53340
rect 54080 53284 54136 53340
rect 54184 53284 54240 53340
rect 54288 53284 54344 53340
rect 54392 53284 54448 53340
rect 62768 53284 62824 53340
rect 62872 53284 62928 53340
rect 62976 53284 63032 53340
rect 63080 53284 63136 53340
rect 63184 53284 63240 53340
rect 63288 53284 63344 53340
rect 63392 53284 63448 53340
rect 71768 53284 71824 53340
rect 71872 53284 71928 53340
rect 71976 53284 72032 53340
rect 72080 53284 72136 53340
rect 72184 53284 72240 53340
rect 72288 53284 72344 53340
rect 72392 53284 72448 53340
rect 80768 53284 80824 53340
rect 80872 53284 80928 53340
rect 80976 53284 81032 53340
rect 81080 53284 81136 53340
rect 81184 53284 81240 53340
rect 81288 53284 81344 53340
rect 81392 53284 81448 53340
rect 89768 53284 89824 53340
rect 89872 53284 89928 53340
rect 89976 53284 90032 53340
rect 90080 53284 90136 53340
rect 90184 53284 90240 53340
rect 90288 53284 90344 53340
rect 90392 53284 90448 53340
rect 4268 52500 4324 52556
rect 4372 52500 4428 52556
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 4788 52500 4844 52556
rect 4892 52500 4948 52556
rect 13268 52500 13324 52556
rect 13372 52500 13428 52556
rect 13476 52500 13532 52556
rect 13580 52500 13636 52556
rect 13684 52500 13740 52556
rect 13788 52500 13844 52556
rect 13892 52500 13948 52556
rect 22268 52500 22324 52556
rect 22372 52500 22428 52556
rect 22476 52500 22532 52556
rect 22580 52500 22636 52556
rect 22684 52500 22740 52556
rect 22788 52500 22844 52556
rect 22892 52500 22948 52556
rect 31268 52500 31324 52556
rect 31372 52500 31428 52556
rect 31476 52500 31532 52556
rect 31580 52500 31636 52556
rect 31684 52500 31740 52556
rect 31788 52500 31844 52556
rect 31892 52500 31948 52556
rect 40268 52500 40324 52556
rect 40372 52500 40428 52556
rect 40476 52500 40532 52556
rect 40580 52500 40636 52556
rect 40684 52500 40740 52556
rect 40788 52500 40844 52556
rect 40892 52500 40948 52556
rect 49268 52500 49324 52556
rect 49372 52500 49428 52556
rect 49476 52500 49532 52556
rect 49580 52500 49636 52556
rect 49684 52500 49740 52556
rect 49788 52500 49844 52556
rect 49892 52500 49948 52556
rect 58268 52500 58324 52556
rect 58372 52500 58428 52556
rect 58476 52500 58532 52556
rect 58580 52500 58636 52556
rect 58684 52500 58740 52556
rect 58788 52500 58844 52556
rect 58892 52500 58948 52556
rect 67268 52500 67324 52556
rect 67372 52500 67428 52556
rect 67476 52500 67532 52556
rect 67580 52500 67636 52556
rect 67684 52500 67740 52556
rect 67788 52500 67844 52556
rect 67892 52500 67948 52556
rect 76268 52500 76324 52556
rect 76372 52500 76428 52556
rect 76476 52500 76532 52556
rect 76580 52500 76636 52556
rect 76684 52500 76740 52556
rect 76788 52500 76844 52556
rect 76892 52500 76948 52556
rect 85268 52500 85324 52556
rect 85372 52500 85428 52556
rect 85476 52500 85532 52556
rect 85580 52500 85636 52556
rect 85684 52500 85740 52556
rect 85788 52500 85844 52556
rect 85892 52500 85948 52556
rect 94268 52500 94324 52556
rect 94372 52500 94428 52556
rect 94476 52500 94532 52556
rect 94580 52500 94636 52556
rect 94684 52500 94740 52556
rect 94788 52500 94844 52556
rect 94892 52500 94948 52556
rect 8768 51716 8824 51772
rect 8872 51716 8928 51772
rect 8976 51716 9032 51772
rect 9080 51716 9136 51772
rect 9184 51716 9240 51772
rect 9288 51716 9344 51772
rect 9392 51716 9448 51772
rect 17768 51716 17824 51772
rect 17872 51716 17928 51772
rect 17976 51716 18032 51772
rect 18080 51716 18136 51772
rect 18184 51716 18240 51772
rect 18288 51716 18344 51772
rect 18392 51716 18448 51772
rect 26768 51716 26824 51772
rect 26872 51716 26928 51772
rect 26976 51716 27032 51772
rect 27080 51716 27136 51772
rect 27184 51716 27240 51772
rect 27288 51716 27344 51772
rect 27392 51716 27448 51772
rect 35768 51716 35824 51772
rect 35872 51716 35928 51772
rect 35976 51716 36032 51772
rect 36080 51716 36136 51772
rect 36184 51716 36240 51772
rect 36288 51716 36344 51772
rect 36392 51716 36448 51772
rect 44768 51716 44824 51772
rect 44872 51716 44928 51772
rect 44976 51716 45032 51772
rect 45080 51716 45136 51772
rect 45184 51716 45240 51772
rect 45288 51716 45344 51772
rect 45392 51716 45448 51772
rect 53768 51716 53824 51772
rect 53872 51716 53928 51772
rect 53976 51716 54032 51772
rect 54080 51716 54136 51772
rect 54184 51716 54240 51772
rect 54288 51716 54344 51772
rect 54392 51716 54448 51772
rect 62768 51716 62824 51772
rect 62872 51716 62928 51772
rect 62976 51716 63032 51772
rect 63080 51716 63136 51772
rect 63184 51716 63240 51772
rect 63288 51716 63344 51772
rect 63392 51716 63448 51772
rect 71768 51716 71824 51772
rect 71872 51716 71928 51772
rect 71976 51716 72032 51772
rect 72080 51716 72136 51772
rect 72184 51716 72240 51772
rect 72288 51716 72344 51772
rect 72392 51716 72448 51772
rect 80768 51716 80824 51772
rect 80872 51716 80928 51772
rect 80976 51716 81032 51772
rect 81080 51716 81136 51772
rect 81184 51716 81240 51772
rect 81288 51716 81344 51772
rect 81392 51716 81448 51772
rect 89768 51716 89824 51772
rect 89872 51716 89928 51772
rect 89976 51716 90032 51772
rect 90080 51716 90136 51772
rect 90184 51716 90240 51772
rect 90288 51716 90344 51772
rect 90392 51716 90448 51772
rect 4268 50932 4324 50988
rect 4372 50932 4428 50988
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 4788 50932 4844 50988
rect 4892 50932 4948 50988
rect 13268 50932 13324 50988
rect 13372 50932 13428 50988
rect 13476 50932 13532 50988
rect 13580 50932 13636 50988
rect 13684 50932 13740 50988
rect 13788 50932 13844 50988
rect 13892 50932 13948 50988
rect 22268 50932 22324 50988
rect 22372 50932 22428 50988
rect 22476 50932 22532 50988
rect 22580 50932 22636 50988
rect 22684 50932 22740 50988
rect 22788 50932 22844 50988
rect 22892 50932 22948 50988
rect 31268 50932 31324 50988
rect 31372 50932 31428 50988
rect 31476 50932 31532 50988
rect 31580 50932 31636 50988
rect 31684 50932 31740 50988
rect 31788 50932 31844 50988
rect 31892 50932 31948 50988
rect 40268 50932 40324 50988
rect 40372 50932 40428 50988
rect 40476 50932 40532 50988
rect 40580 50932 40636 50988
rect 40684 50932 40740 50988
rect 40788 50932 40844 50988
rect 40892 50932 40948 50988
rect 49268 50932 49324 50988
rect 49372 50932 49428 50988
rect 49476 50932 49532 50988
rect 49580 50932 49636 50988
rect 49684 50932 49740 50988
rect 49788 50932 49844 50988
rect 49892 50932 49948 50988
rect 58268 50932 58324 50988
rect 58372 50932 58428 50988
rect 58476 50932 58532 50988
rect 58580 50932 58636 50988
rect 58684 50932 58740 50988
rect 58788 50932 58844 50988
rect 58892 50932 58948 50988
rect 67268 50932 67324 50988
rect 67372 50932 67428 50988
rect 67476 50932 67532 50988
rect 67580 50932 67636 50988
rect 67684 50932 67740 50988
rect 67788 50932 67844 50988
rect 67892 50932 67948 50988
rect 76268 50932 76324 50988
rect 76372 50932 76428 50988
rect 76476 50932 76532 50988
rect 76580 50932 76636 50988
rect 76684 50932 76740 50988
rect 76788 50932 76844 50988
rect 76892 50932 76948 50988
rect 85268 50932 85324 50988
rect 85372 50932 85428 50988
rect 85476 50932 85532 50988
rect 85580 50932 85636 50988
rect 85684 50932 85740 50988
rect 85788 50932 85844 50988
rect 85892 50932 85948 50988
rect 94268 50932 94324 50988
rect 94372 50932 94428 50988
rect 94476 50932 94532 50988
rect 94580 50932 94636 50988
rect 94684 50932 94740 50988
rect 94788 50932 94844 50988
rect 94892 50932 94948 50988
rect 8768 50148 8824 50204
rect 8872 50148 8928 50204
rect 8976 50148 9032 50204
rect 9080 50148 9136 50204
rect 9184 50148 9240 50204
rect 9288 50148 9344 50204
rect 9392 50148 9448 50204
rect 17768 50148 17824 50204
rect 17872 50148 17928 50204
rect 17976 50148 18032 50204
rect 18080 50148 18136 50204
rect 18184 50148 18240 50204
rect 18288 50148 18344 50204
rect 18392 50148 18448 50204
rect 26768 50148 26824 50204
rect 26872 50148 26928 50204
rect 26976 50148 27032 50204
rect 27080 50148 27136 50204
rect 27184 50148 27240 50204
rect 27288 50148 27344 50204
rect 27392 50148 27448 50204
rect 35768 50148 35824 50204
rect 35872 50148 35928 50204
rect 35976 50148 36032 50204
rect 36080 50148 36136 50204
rect 36184 50148 36240 50204
rect 36288 50148 36344 50204
rect 36392 50148 36448 50204
rect 44768 50148 44824 50204
rect 44872 50148 44928 50204
rect 44976 50148 45032 50204
rect 45080 50148 45136 50204
rect 45184 50148 45240 50204
rect 45288 50148 45344 50204
rect 45392 50148 45448 50204
rect 53768 50148 53824 50204
rect 53872 50148 53928 50204
rect 53976 50148 54032 50204
rect 54080 50148 54136 50204
rect 54184 50148 54240 50204
rect 54288 50148 54344 50204
rect 54392 50148 54448 50204
rect 62768 50148 62824 50204
rect 62872 50148 62928 50204
rect 62976 50148 63032 50204
rect 63080 50148 63136 50204
rect 63184 50148 63240 50204
rect 63288 50148 63344 50204
rect 63392 50148 63448 50204
rect 71768 50148 71824 50204
rect 71872 50148 71928 50204
rect 71976 50148 72032 50204
rect 72080 50148 72136 50204
rect 72184 50148 72240 50204
rect 72288 50148 72344 50204
rect 72392 50148 72448 50204
rect 80768 50148 80824 50204
rect 80872 50148 80928 50204
rect 80976 50148 81032 50204
rect 81080 50148 81136 50204
rect 81184 50148 81240 50204
rect 81288 50148 81344 50204
rect 81392 50148 81448 50204
rect 89768 50148 89824 50204
rect 89872 50148 89928 50204
rect 89976 50148 90032 50204
rect 90080 50148 90136 50204
rect 90184 50148 90240 50204
rect 90288 50148 90344 50204
rect 90392 50148 90448 50204
rect 4268 49364 4324 49420
rect 4372 49364 4428 49420
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 4788 49364 4844 49420
rect 4892 49364 4948 49420
rect 13268 49364 13324 49420
rect 13372 49364 13428 49420
rect 13476 49364 13532 49420
rect 13580 49364 13636 49420
rect 13684 49364 13740 49420
rect 13788 49364 13844 49420
rect 13892 49364 13948 49420
rect 22268 49364 22324 49420
rect 22372 49364 22428 49420
rect 22476 49364 22532 49420
rect 22580 49364 22636 49420
rect 22684 49364 22740 49420
rect 22788 49364 22844 49420
rect 22892 49364 22948 49420
rect 31268 49364 31324 49420
rect 31372 49364 31428 49420
rect 31476 49364 31532 49420
rect 31580 49364 31636 49420
rect 31684 49364 31740 49420
rect 31788 49364 31844 49420
rect 31892 49364 31948 49420
rect 40268 49364 40324 49420
rect 40372 49364 40428 49420
rect 40476 49364 40532 49420
rect 40580 49364 40636 49420
rect 40684 49364 40740 49420
rect 40788 49364 40844 49420
rect 40892 49364 40948 49420
rect 49268 49364 49324 49420
rect 49372 49364 49428 49420
rect 49476 49364 49532 49420
rect 49580 49364 49636 49420
rect 49684 49364 49740 49420
rect 49788 49364 49844 49420
rect 49892 49364 49948 49420
rect 58268 49364 58324 49420
rect 58372 49364 58428 49420
rect 58476 49364 58532 49420
rect 58580 49364 58636 49420
rect 58684 49364 58740 49420
rect 58788 49364 58844 49420
rect 58892 49364 58948 49420
rect 67268 49364 67324 49420
rect 67372 49364 67428 49420
rect 67476 49364 67532 49420
rect 67580 49364 67636 49420
rect 67684 49364 67740 49420
rect 67788 49364 67844 49420
rect 67892 49364 67948 49420
rect 76268 49364 76324 49420
rect 76372 49364 76428 49420
rect 76476 49364 76532 49420
rect 76580 49364 76636 49420
rect 76684 49364 76740 49420
rect 76788 49364 76844 49420
rect 76892 49364 76948 49420
rect 85268 49364 85324 49420
rect 85372 49364 85428 49420
rect 85476 49364 85532 49420
rect 85580 49364 85636 49420
rect 85684 49364 85740 49420
rect 85788 49364 85844 49420
rect 85892 49364 85948 49420
rect 94268 49364 94324 49420
rect 94372 49364 94428 49420
rect 94476 49364 94532 49420
rect 94580 49364 94636 49420
rect 94684 49364 94740 49420
rect 94788 49364 94844 49420
rect 94892 49364 94948 49420
rect 8768 48580 8824 48636
rect 8872 48580 8928 48636
rect 8976 48580 9032 48636
rect 9080 48580 9136 48636
rect 9184 48580 9240 48636
rect 9288 48580 9344 48636
rect 9392 48580 9448 48636
rect 17768 48580 17824 48636
rect 17872 48580 17928 48636
rect 17976 48580 18032 48636
rect 18080 48580 18136 48636
rect 18184 48580 18240 48636
rect 18288 48580 18344 48636
rect 18392 48580 18448 48636
rect 26768 48580 26824 48636
rect 26872 48580 26928 48636
rect 26976 48580 27032 48636
rect 27080 48580 27136 48636
rect 27184 48580 27240 48636
rect 27288 48580 27344 48636
rect 27392 48580 27448 48636
rect 35768 48580 35824 48636
rect 35872 48580 35928 48636
rect 35976 48580 36032 48636
rect 36080 48580 36136 48636
rect 36184 48580 36240 48636
rect 36288 48580 36344 48636
rect 36392 48580 36448 48636
rect 44768 48580 44824 48636
rect 44872 48580 44928 48636
rect 44976 48580 45032 48636
rect 45080 48580 45136 48636
rect 45184 48580 45240 48636
rect 45288 48580 45344 48636
rect 45392 48580 45448 48636
rect 53768 48580 53824 48636
rect 53872 48580 53928 48636
rect 53976 48580 54032 48636
rect 54080 48580 54136 48636
rect 54184 48580 54240 48636
rect 54288 48580 54344 48636
rect 54392 48580 54448 48636
rect 62768 48580 62824 48636
rect 62872 48580 62928 48636
rect 62976 48580 63032 48636
rect 63080 48580 63136 48636
rect 63184 48580 63240 48636
rect 63288 48580 63344 48636
rect 63392 48580 63448 48636
rect 71768 48580 71824 48636
rect 71872 48580 71928 48636
rect 71976 48580 72032 48636
rect 72080 48580 72136 48636
rect 72184 48580 72240 48636
rect 72288 48580 72344 48636
rect 72392 48580 72448 48636
rect 80768 48580 80824 48636
rect 80872 48580 80928 48636
rect 80976 48580 81032 48636
rect 81080 48580 81136 48636
rect 81184 48580 81240 48636
rect 81288 48580 81344 48636
rect 81392 48580 81448 48636
rect 89768 48580 89824 48636
rect 89872 48580 89928 48636
rect 89976 48580 90032 48636
rect 90080 48580 90136 48636
rect 90184 48580 90240 48636
rect 90288 48580 90344 48636
rect 90392 48580 90448 48636
rect 4268 47796 4324 47852
rect 4372 47796 4428 47852
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 4788 47796 4844 47852
rect 4892 47796 4948 47852
rect 13268 47796 13324 47852
rect 13372 47796 13428 47852
rect 13476 47796 13532 47852
rect 13580 47796 13636 47852
rect 13684 47796 13740 47852
rect 13788 47796 13844 47852
rect 13892 47796 13948 47852
rect 22268 47796 22324 47852
rect 22372 47796 22428 47852
rect 22476 47796 22532 47852
rect 22580 47796 22636 47852
rect 22684 47796 22740 47852
rect 22788 47796 22844 47852
rect 22892 47796 22948 47852
rect 31268 47796 31324 47852
rect 31372 47796 31428 47852
rect 31476 47796 31532 47852
rect 31580 47796 31636 47852
rect 31684 47796 31740 47852
rect 31788 47796 31844 47852
rect 31892 47796 31948 47852
rect 40268 47796 40324 47852
rect 40372 47796 40428 47852
rect 40476 47796 40532 47852
rect 40580 47796 40636 47852
rect 40684 47796 40740 47852
rect 40788 47796 40844 47852
rect 40892 47796 40948 47852
rect 49268 47796 49324 47852
rect 49372 47796 49428 47852
rect 49476 47796 49532 47852
rect 49580 47796 49636 47852
rect 49684 47796 49740 47852
rect 49788 47796 49844 47852
rect 49892 47796 49948 47852
rect 58268 47796 58324 47852
rect 58372 47796 58428 47852
rect 58476 47796 58532 47852
rect 58580 47796 58636 47852
rect 58684 47796 58740 47852
rect 58788 47796 58844 47852
rect 58892 47796 58948 47852
rect 67268 47796 67324 47852
rect 67372 47796 67428 47852
rect 67476 47796 67532 47852
rect 67580 47796 67636 47852
rect 67684 47796 67740 47852
rect 67788 47796 67844 47852
rect 67892 47796 67948 47852
rect 76268 47796 76324 47852
rect 76372 47796 76428 47852
rect 76476 47796 76532 47852
rect 76580 47796 76636 47852
rect 76684 47796 76740 47852
rect 76788 47796 76844 47852
rect 76892 47796 76948 47852
rect 85268 47796 85324 47852
rect 85372 47796 85428 47852
rect 85476 47796 85532 47852
rect 85580 47796 85636 47852
rect 85684 47796 85740 47852
rect 85788 47796 85844 47852
rect 85892 47796 85948 47852
rect 94268 47796 94324 47852
rect 94372 47796 94428 47852
rect 94476 47796 94532 47852
rect 94580 47796 94636 47852
rect 94684 47796 94740 47852
rect 94788 47796 94844 47852
rect 94892 47796 94948 47852
rect 8768 47012 8824 47068
rect 8872 47012 8928 47068
rect 8976 47012 9032 47068
rect 9080 47012 9136 47068
rect 9184 47012 9240 47068
rect 9288 47012 9344 47068
rect 9392 47012 9448 47068
rect 17768 47012 17824 47068
rect 17872 47012 17928 47068
rect 17976 47012 18032 47068
rect 18080 47012 18136 47068
rect 18184 47012 18240 47068
rect 18288 47012 18344 47068
rect 18392 47012 18448 47068
rect 26768 47012 26824 47068
rect 26872 47012 26928 47068
rect 26976 47012 27032 47068
rect 27080 47012 27136 47068
rect 27184 47012 27240 47068
rect 27288 47012 27344 47068
rect 27392 47012 27448 47068
rect 35768 47012 35824 47068
rect 35872 47012 35928 47068
rect 35976 47012 36032 47068
rect 36080 47012 36136 47068
rect 36184 47012 36240 47068
rect 36288 47012 36344 47068
rect 36392 47012 36448 47068
rect 44768 47012 44824 47068
rect 44872 47012 44928 47068
rect 44976 47012 45032 47068
rect 45080 47012 45136 47068
rect 45184 47012 45240 47068
rect 45288 47012 45344 47068
rect 45392 47012 45448 47068
rect 53768 47012 53824 47068
rect 53872 47012 53928 47068
rect 53976 47012 54032 47068
rect 54080 47012 54136 47068
rect 54184 47012 54240 47068
rect 54288 47012 54344 47068
rect 54392 47012 54448 47068
rect 62768 47012 62824 47068
rect 62872 47012 62928 47068
rect 62976 47012 63032 47068
rect 63080 47012 63136 47068
rect 63184 47012 63240 47068
rect 63288 47012 63344 47068
rect 63392 47012 63448 47068
rect 71768 47012 71824 47068
rect 71872 47012 71928 47068
rect 71976 47012 72032 47068
rect 72080 47012 72136 47068
rect 72184 47012 72240 47068
rect 72288 47012 72344 47068
rect 72392 47012 72448 47068
rect 80768 47012 80824 47068
rect 80872 47012 80928 47068
rect 80976 47012 81032 47068
rect 81080 47012 81136 47068
rect 81184 47012 81240 47068
rect 81288 47012 81344 47068
rect 81392 47012 81448 47068
rect 89768 47012 89824 47068
rect 89872 47012 89928 47068
rect 89976 47012 90032 47068
rect 90080 47012 90136 47068
rect 90184 47012 90240 47068
rect 90288 47012 90344 47068
rect 90392 47012 90448 47068
rect 4268 46228 4324 46284
rect 4372 46228 4428 46284
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 4788 46228 4844 46284
rect 4892 46228 4948 46284
rect 13268 46228 13324 46284
rect 13372 46228 13428 46284
rect 13476 46228 13532 46284
rect 13580 46228 13636 46284
rect 13684 46228 13740 46284
rect 13788 46228 13844 46284
rect 13892 46228 13948 46284
rect 22268 46228 22324 46284
rect 22372 46228 22428 46284
rect 22476 46228 22532 46284
rect 22580 46228 22636 46284
rect 22684 46228 22740 46284
rect 22788 46228 22844 46284
rect 22892 46228 22948 46284
rect 31268 46228 31324 46284
rect 31372 46228 31428 46284
rect 31476 46228 31532 46284
rect 31580 46228 31636 46284
rect 31684 46228 31740 46284
rect 31788 46228 31844 46284
rect 31892 46228 31948 46284
rect 40268 46228 40324 46284
rect 40372 46228 40428 46284
rect 40476 46228 40532 46284
rect 40580 46228 40636 46284
rect 40684 46228 40740 46284
rect 40788 46228 40844 46284
rect 40892 46228 40948 46284
rect 49268 46228 49324 46284
rect 49372 46228 49428 46284
rect 49476 46228 49532 46284
rect 49580 46228 49636 46284
rect 49684 46228 49740 46284
rect 49788 46228 49844 46284
rect 49892 46228 49948 46284
rect 58268 46228 58324 46284
rect 58372 46228 58428 46284
rect 58476 46228 58532 46284
rect 58580 46228 58636 46284
rect 58684 46228 58740 46284
rect 58788 46228 58844 46284
rect 58892 46228 58948 46284
rect 67268 46228 67324 46284
rect 67372 46228 67428 46284
rect 67476 46228 67532 46284
rect 67580 46228 67636 46284
rect 67684 46228 67740 46284
rect 67788 46228 67844 46284
rect 67892 46228 67948 46284
rect 76268 46228 76324 46284
rect 76372 46228 76428 46284
rect 76476 46228 76532 46284
rect 76580 46228 76636 46284
rect 76684 46228 76740 46284
rect 76788 46228 76844 46284
rect 76892 46228 76948 46284
rect 85268 46228 85324 46284
rect 85372 46228 85428 46284
rect 85476 46228 85532 46284
rect 85580 46228 85636 46284
rect 85684 46228 85740 46284
rect 85788 46228 85844 46284
rect 85892 46228 85948 46284
rect 94268 46228 94324 46284
rect 94372 46228 94428 46284
rect 94476 46228 94532 46284
rect 94580 46228 94636 46284
rect 94684 46228 94740 46284
rect 94788 46228 94844 46284
rect 94892 46228 94948 46284
rect 8768 45444 8824 45500
rect 8872 45444 8928 45500
rect 8976 45444 9032 45500
rect 9080 45444 9136 45500
rect 9184 45444 9240 45500
rect 9288 45444 9344 45500
rect 9392 45444 9448 45500
rect 17768 45444 17824 45500
rect 17872 45444 17928 45500
rect 17976 45444 18032 45500
rect 18080 45444 18136 45500
rect 18184 45444 18240 45500
rect 18288 45444 18344 45500
rect 18392 45444 18448 45500
rect 26768 45444 26824 45500
rect 26872 45444 26928 45500
rect 26976 45444 27032 45500
rect 27080 45444 27136 45500
rect 27184 45444 27240 45500
rect 27288 45444 27344 45500
rect 27392 45444 27448 45500
rect 35768 45444 35824 45500
rect 35872 45444 35928 45500
rect 35976 45444 36032 45500
rect 36080 45444 36136 45500
rect 36184 45444 36240 45500
rect 36288 45444 36344 45500
rect 36392 45444 36448 45500
rect 44768 45444 44824 45500
rect 44872 45444 44928 45500
rect 44976 45444 45032 45500
rect 45080 45444 45136 45500
rect 45184 45444 45240 45500
rect 45288 45444 45344 45500
rect 45392 45444 45448 45500
rect 53768 45444 53824 45500
rect 53872 45444 53928 45500
rect 53976 45444 54032 45500
rect 54080 45444 54136 45500
rect 54184 45444 54240 45500
rect 54288 45444 54344 45500
rect 54392 45444 54448 45500
rect 62768 45444 62824 45500
rect 62872 45444 62928 45500
rect 62976 45444 63032 45500
rect 63080 45444 63136 45500
rect 63184 45444 63240 45500
rect 63288 45444 63344 45500
rect 63392 45444 63448 45500
rect 71768 45444 71824 45500
rect 71872 45444 71928 45500
rect 71976 45444 72032 45500
rect 72080 45444 72136 45500
rect 72184 45444 72240 45500
rect 72288 45444 72344 45500
rect 72392 45444 72448 45500
rect 80768 45444 80824 45500
rect 80872 45444 80928 45500
rect 80976 45444 81032 45500
rect 81080 45444 81136 45500
rect 81184 45444 81240 45500
rect 81288 45444 81344 45500
rect 81392 45444 81448 45500
rect 89768 45444 89824 45500
rect 89872 45444 89928 45500
rect 89976 45444 90032 45500
rect 90080 45444 90136 45500
rect 90184 45444 90240 45500
rect 90288 45444 90344 45500
rect 90392 45444 90448 45500
rect 4268 44660 4324 44716
rect 4372 44660 4428 44716
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 4788 44660 4844 44716
rect 4892 44660 4948 44716
rect 13268 44660 13324 44716
rect 13372 44660 13428 44716
rect 13476 44660 13532 44716
rect 13580 44660 13636 44716
rect 13684 44660 13740 44716
rect 13788 44660 13844 44716
rect 13892 44660 13948 44716
rect 22268 44660 22324 44716
rect 22372 44660 22428 44716
rect 22476 44660 22532 44716
rect 22580 44660 22636 44716
rect 22684 44660 22740 44716
rect 22788 44660 22844 44716
rect 22892 44660 22948 44716
rect 31268 44660 31324 44716
rect 31372 44660 31428 44716
rect 31476 44660 31532 44716
rect 31580 44660 31636 44716
rect 31684 44660 31740 44716
rect 31788 44660 31844 44716
rect 31892 44660 31948 44716
rect 40268 44660 40324 44716
rect 40372 44660 40428 44716
rect 40476 44660 40532 44716
rect 40580 44660 40636 44716
rect 40684 44660 40740 44716
rect 40788 44660 40844 44716
rect 40892 44660 40948 44716
rect 49268 44660 49324 44716
rect 49372 44660 49428 44716
rect 49476 44660 49532 44716
rect 49580 44660 49636 44716
rect 49684 44660 49740 44716
rect 49788 44660 49844 44716
rect 49892 44660 49948 44716
rect 58268 44660 58324 44716
rect 58372 44660 58428 44716
rect 58476 44660 58532 44716
rect 58580 44660 58636 44716
rect 58684 44660 58740 44716
rect 58788 44660 58844 44716
rect 58892 44660 58948 44716
rect 67268 44660 67324 44716
rect 67372 44660 67428 44716
rect 67476 44660 67532 44716
rect 67580 44660 67636 44716
rect 67684 44660 67740 44716
rect 67788 44660 67844 44716
rect 67892 44660 67948 44716
rect 76268 44660 76324 44716
rect 76372 44660 76428 44716
rect 76476 44660 76532 44716
rect 76580 44660 76636 44716
rect 76684 44660 76740 44716
rect 76788 44660 76844 44716
rect 76892 44660 76948 44716
rect 85268 44660 85324 44716
rect 85372 44660 85428 44716
rect 85476 44660 85532 44716
rect 85580 44660 85636 44716
rect 85684 44660 85740 44716
rect 85788 44660 85844 44716
rect 85892 44660 85948 44716
rect 94268 44660 94324 44716
rect 94372 44660 94428 44716
rect 94476 44660 94532 44716
rect 94580 44660 94636 44716
rect 94684 44660 94740 44716
rect 94788 44660 94844 44716
rect 94892 44660 94948 44716
rect 8768 43876 8824 43932
rect 8872 43876 8928 43932
rect 8976 43876 9032 43932
rect 9080 43876 9136 43932
rect 9184 43876 9240 43932
rect 9288 43876 9344 43932
rect 9392 43876 9448 43932
rect 17768 43876 17824 43932
rect 17872 43876 17928 43932
rect 17976 43876 18032 43932
rect 18080 43876 18136 43932
rect 18184 43876 18240 43932
rect 18288 43876 18344 43932
rect 18392 43876 18448 43932
rect 26768 43876 26824 43932
rect 26872 43876 26928 43932
rect 26976 43876 27032 43932
rect 27080 43876 27136 43932
rect 27184 43876 27240 43932
rect 27288 43876 27344 43932
rect 27392 43876 27448 43932
rect 35768 43876 35824 43932
rect 35872 43876 35928 43932
rect 35976 43876 36032 43932
rect 36080 43876 36136 43932
rect 36184 43876 36240 43932
rect 36288 43876 36344 43932
rect 36392 43876 36448 43932
rect 44768 43876 44824 43932
rect 44872 43876 44928 43932
rect 44976 43876 45032 43932
rect 45080 43876 45136 43932
rect 45184 43876 45240 43932
rect 45288 43876 45344 43932
rect 45392 43876 45448 43932
rect 53768 43876 53824 43932
rect 53872 43876 53928 43932
rect 53976 43876 54032 43932
rect 54080 43876 54136 43932
rect 54184 43876 54240 43932
rect 54288 43876 54344 43932
rect 54392 43876 54448 43932
rect 62768 43876 62824 43932
rect 62872 43876 62928 43932
rect 62976 43876 63032 43932
rect 63080 43876 63136 43932
rect 63184 43876 63240 43932
rect 63288 43876 63344 43932
rect 63392 43876 63448 43932
rect 71768 43876 71824 43932
rect 71872 43876 71928 43932
rect 71976 43876 72032 43932
rect 72080 43876 72136 43932
rect 72184 43876 72240 43932
rect 72288 43876 72344 43932
rect 72392 43876 72448 43932
rect 80768 43876 80824 43932
rect 80872 43876 80928 43932
rect 80976 43876 81032 43932
rect 81080 43876 81136 43932
rect 81184 43876 81240 43932
rect 81288 43876 81344 43932
rect 81392 43876 81448 43932
rect 89768 43876 89824 43932
rect 89872 43876 89928 43932
rect 89976 43876 90032 43932
rect 90080 43876 90136 43932
rect 90184 43876 90240 43932
rect 90288 43876 90344 43932
rect 90392 43876 90448 43932
rect 4268 43092 4324 43148
rect 4372 43092 4428 43148
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 4788 43092 4844 43148
rect 4892 43092 4948 43148
rect 13268 43092 13324 43148
rect 13372 43092 13428 43148
rect 13476 43092 13532 43148
rect 13580 43092 13636 43148
rect 13684 43092 13740 43148
rect 13788 43092 13844 43148
rect 13892 43092 13948 43148
rect 22268 43092 22324 43148
rect 22372 43092 22428 43148
rect 22476 43092 22532 43148
rect 22580 43092 22636 43148
rect 22684 43092 22740 43148
rect 22788 43092 22844 43148
rect 22892 43092 22948 43148
rect 31268 43092 31324 43148
rect 31372 43092 31428 43148
rect 31476 43092 31532 43148
rect 31580 43092 31636 43148
rect 31684 43092 31740 43148
rect 31788 43092 31844 43148
rect 31892 43092 31948 43148
rect 40268 43092 40324 43148
rect 40372 43092 40428 43148
rect 40476 43092 40532 43148
rect 40580 43092 40636 43148
rect 40684 43092 40740 43148
rect 40788 43092 40844 43148
rect 40892 43092 40948 43148
rect 49268 43092 49324 43148
rect 49372 43092 49428 43148
rect 49476 43092 49532 43148
rect 49580 43092 49636 43148
rect 49684 43092 49740 43148
rect 49788 43092 49844 43148
rect 49892 43092 49948 43148
rect 58268 43092 58324 43148
rect 58372 43092 58428 43148
rect 58476 43092 58532 43148
rect 58580 43092 58636 43148
rect 58684 43092 58740 43148
rect 58788 43092 58844 43148
rect 58892 43092 58948 43148
rect 67268 43092 67324 43148
rect 67372 43092 67428 43148
rect 67476 43092 67532 43148
rect 67580 43092 67636 43148
rect 67684 43092 67740 43148
rect 67788 43092 67844 43148
rect 67892 43092 67948 43148
rect 76268 43092 76324 43148
rect 76372 43092 76428 43148
rect 76476 43092 76532 43148
rect 76580 43092 76636 43148
rect 76684 43092 76740 43148
rect 76788 43092 76844 43148
rect 76892 43092 76948 43148
rect 85268 43092 85324 43148
rect 85372 43092 85428 43148
rect 85476 43092 85532 43148
rect 85580 43092 85636 43148
rect 85684 43092 85740 43148
rect 85788 43092 85844 43148
rect 85892 43092 85948 43148
rect 94268 43092 94324 43148
rect 94372 43092 94428 43148
rect 94476 43092 94532 43148
rect 94580 43092 94636 43148
rect 94684 43092 94740 43148
rect 94788 43092 94844 43148
rect 94892 43092 94948 43148
rect 8768 42308 8824 42364
rect 8872 42308 8928 42364
rect 8976 42308 9032 42364
rect 9080 42308 9136 42364
rect 9184 42308 9240 42364
rect 9288 42308 9344 42364
rect 9392 42308 9448 42364
rect 17768 42308 17824 42364
rect 17872 42308 17928 42364
rect 17976 42308 18032 42364
rect 18080 42308 18136 42364
rect 18184 42308 18240 42364
rect 18288 42308 18344 42364
rect 18392 42308 18448 42364
rect 26768 42308 26824 42364
rect 26872 42308 26928 42364
rect 26976 42308 27032 42364
rect 27080 42308 27136 42364
rect 27184 42308 27240 42364
rect 27288 42308 27344 42364
rect 27392 42308 27448 42364
rect 35768 42308 35824 42364
rect 35872 42308 35928 42364
rect 35976 42308 36032 42364
rect 36080 42308 36136 42364
rect 36184 42308 36240 42364
rect 36288 42308 36344 42364
rect 36392 42308 36448 42364
rect 44768 42308 44824 42364
rect 44872 42308 44928 42364
rect 44976 42308 45032 42364
rect 45080 42308 45136 42364
rect 45184 42308 45240 42364
rect 45288 42308 45344 42364
rect 45392 42308 45448 42364
rect 53768 42308 53824 42364
rect 53872 42308 53928 42364
rect 53976 42308 54032 42364
rect 54080 42308 54136 42364
rect 54184 42308 54240 42364
rect 54288 42308 54344 42364
rect 54392 42308 54448 42364
rect 62768 42308 62824 42364
rect 62872 42308 62928 42364
rect 62976 42308 63032 42364
rect 63080 42308 63136 42364
rect 63184 42308 63240 42364
rect 63288 42308 63344 42364
rect 63392 42308 63448 42364
rect 71768 42308 71824 42364
rect 71872 42308 71928 42364
rect 71976 42308 72032 42364
rect 72080 42308 72136 42364
rect 72184 42308 72240 42364
rect 72288 42308 72344 42364
rect 72392 42308 72448 42364
rect 80768 42308 80824 42364
rect 80872 42308 80928 42364
rect 80976 42308 81032 42364
rect 81080 42308 81136 42364
rect 81184 42308 81240 42364
rect 81288 42308 81344 42364
rect 81392 42308 81448 42364
rect 89768 42308 89824 42364
rect 89872 42308 89928 42364
rect 89976 42308 90032 42364
rect 90080 42308 90136 42364
rect 90184 42308 90240 42364
rect 90288 42308 90344 42364
rect 90392 42308 90448 42364
rect 49084 42028 49140 42084
rect 4268 41524 4324 41580
rect 4372 41524 4428 41580
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 4788 41524 4844 41580
rect 4892 41524 4948 41580
rect 13268 41524 13324 41580
rect 13372 41524 13428 41580
rect 13476 41524 13532 41580
rect 13580 41524 13636 41580
rect 13684 41524 13740 41580
rect 13788 41524 13844 41580
rect 13892 41524 13948 41580
rect 22268 41524 22324 41580
rect 22372 41524 22428 41580
rect 22476 41524 22532 41580
rect 22580 41524 22636 41580
rect 22684 41524 22740 41580
rect 22788 41524 22844 41580
rect 22892 41524 22948 41580
rect 31268 41524 31324 41580
rect 31372 41524 31428 41580
rect 31476 41524 31532 41580
rect 31580 41524 31636 41580
rect 31684 41524 31740 41580
rect 31788 41524 31844 41580
rect 31892 41524 31948 41580
rect 40268 41524 40324 41580
rect 40372 41524 40428 41580
rect 40476 41524 40532 41580
rect 40580 41524 40636 41580
rect 40684 41524 40740 41580
rect 40788 41524 40844 41580
rect 40892 41524 40948 41580
rect 49268 41524 49324 41580
rect 49372 41524 49428 41580
rect 49476 41524 49532 41580
rect 49580 41524 49636 41580
rect 49684 41524 49740 41580
rect 49788 41524 49844 41580
rect 49892 41524 49948 41580
rect 58268 41524 58324 41580
rect 58372 41524 58428 41580
rect 58476 41524 58532 41580
rect 58580 41524 58636 41580
rect 58684 41524 58740 41580
rect 58788 41524 58844 41580
rect 58892 41524 58948 41580
rect 67268 41524 67324 41580
rect 67372 41524 67428 41580
rect 67476 41524 67532 41580
rect 67580 41524 67636 41580
rect 67684 41524 67740 41580
rect 67788 41524 67844 41580
rect 67892 41524 67948 41580
rect 76268 41524 76324 41580
rect 76372 41524 76428 41580
rect 76476 41524 76532 41580
rect 76580 41524 76636 41580
rect 76684 41524 76740 41580
rect 76788 41524 76844 41580
rect 76892 41524 76948 41580
rect 85268 41524 85324 41580
rect 85372 41524 85428 41580
rect 85476 41524 85532 41580
rect 85580 41524 85636 41580
rect 85684 41524 85740 41580
rect 85788 41524 85844 41580
rect 85892 41524 85948 41580
rect 94268 41524 94324 41580
rect 94372 41524 94428 41580
rect 94476 41524 94532 41580
rect 94580 41524 94636 41580
rect 94684 41524 94740 41580
rect 94788 41524 94844 41580
rect 94892 41524 94948 41580
rect 8768 40740 8824 40796
rect 8872 40740 8928 40796
rect 8976 40740 9032 40796
rect 9080 40740 9136 40796
rect 9184 40740 9240 40796
rect 9288 40740 9344 40796
rect 9392 40740 9448 40796
rect 17768 40740 17824 40796
rect 17872 40740 17928 40796
rect 17976 40740 18032 40796
rect 18080 40740 18136 40796
rect 18184 40740 18240 40796
rect 18288 40740 18344 40796
rect 18392 40740 18448 40796
rect 26768 40740 26824 40796
rect 26872 40740 26928 40796
rect 26976 40740 27032 40796
rect 27080 40740 27136 40796
rect 27184 40740 27240 40796
rect 27288 40740 27344 40796
rect 27392 40740 27448 40796
rect 35768 40740 35824 40796
rect 35872 40740 35928 40796
rect 35976 40740 36032 40796
rect 36080 40740 36136 40796
rect 36184 40740 36240 40796
rect 36288 40740 36344 40796
rect 36392 40740 36448 40796
rect 44768 40740 44824 40796
rect 44872 40740 44928 40796
rect 44976 40740 45032 40796
rect 45080 40740 45136 40796
rect 45184 40740 45240 40796
rect 45288 40740 45344 40796
rect 45392 40740 45448 40796
rect 53768 40740 53824 40796
rect 53872 40740 53928 40796
rect 53976 40740 54032 40796
rect 54080 40740 54136 40796
rect 54184 40740 54240 40796
rect 54288 40740 54344 40796
rect 54392 40740 54448 40796
rect 62768 40740 62824 40796
rect 62872 40740 62928 40796
rect 62976 40740 63032 40796
rect 63080 40740 63136 40796
rect 63184 40740 63240 40796
rect 63288 40740 63344 40796
rect 63392 40740 63448 40796
rect 71768 40740 71824 40796
rect 71872 40740 71928 40796
rect 71976 40740 72032 40796
rect 72080 40740 72136 40796
rect 72184 40740 72240 40796
rect 72288 40740 72344 40796
rect 72392 40740 72448 40796
rect 80768 40740 80824 40796
rect 80872 40740 80928 40796
rect 80976 40740 81032 40796
rect 81080 40740 81136 40796
rect 81184 40740 81240 40796
rect 81288 40740 81344 40796
rect 81392 40740 81448 40796
rect 89768 40740 89824 40796
rect 89872 40740 89928 40796
rect 89976 40740 90032 40796
rect 90080 40740 90136 40796
rect 90184 40740 90240 40796
rect 90288 40740 90344 40796
rect 90392 40740 90448 40796
rect 49084 40348 49140 40404
rect 4268 39956 4324 40012
rect 4372 39956 4428 40012
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 4788 39956 4844 40012
rect 4892 39956 4948 40012
rect 13268 39956 13324 40012
rect 13372 39956 13428 40012
rect 13476 39956 13532 40012
rect 13580 39956 13636 40012
rect 13684 39956 13740 40012
rect 13788 39956 13844 40012
rect 13892 39956 13948 40012
rect 22268 39956 22324 40012
rect 22372 39956 22428 40012
rect 22476 39956 22532 40012
rect 22580 39956 22636 40012
rect 22684 39956 22740 40012
rect 22788 39956 22844 40012
rect 22892 39956 22948 40012
rect 31268 39956 31324 40012
rect 31372 39956 31428 40012
rect 31476 39956 31532 40012
rect 31580 39956 31636 40012
rect 31684 39956 31740 40012
rect 31788 39956 31844 40012
rect 31892 39956 31948 40012
rect 40268 39956 40324 40012
rect 40372 39956 40428 40012
rect 40476 39956 40532 40012
rect 40580 39956 40636 40012
rect 40684 39956 40740 40012
rect 40788 39956 40844 40012
rect 40892 39956 40948 40012
rect 49268 39956 49324 40012
rect 49372 39956 49428 40012
rect 49476 39956 49532 40012
rect 49580 39956 49636 40012
rect 49684 39956 49740 40012
rect 49788 39956 49844 40012
rect 49892 39956 49948 40012
rect 58268 39956 58324 40012
rect 58372 39956 58428 40012
rect 58476 39956 58532 40012
rect 58580 39956 58636 40012
rect 58684 39956 58740 40012
rect 58788 39956 58844 40012
rect 58892 39956 58948 40012
rect 67268 39956 67324 40012
rect 67372 39956 67428 40012
rect 67476 39956 67532 40012
rect 67580 39956 67636 40012
rect 67684 39956 67740 40012
rect 67788 39956 67844 40012
rect 67892 39956 67948 40012
rect 76268 39956 76324 40012
rect 76372 39956 76428 40012
rect 76476 39956 76532 40012
rect 76580 39956 76636 40012
rect 76684 39956 76740 40012
rect 76788 39956 76844 40012
rect 76892 39956 76948 40012
rect 85268 39956 85324 40012
rect 85372 39956 85428 40012
rect 85476 39956 85532 40012
rect 85580 39956 85636 40012
rect 85684 39956 85740 40012
rect 85788 39956 85844 40012
rect 85892 39956 85948 40012
rect 94268 39956 94324 40012
rect 94372 39956 94428 40012
rect 94476 39956 94532 40012
rect 94580 39956 94636 40012
rect 94684 39956 94740 40012
rect 94788 39956 94844 40012
rect 94892 39956 94948 40012
rect 8768 39172 8824 39228
rect 8872 39172 8928 39228
rect 8976 39172 9032 39228
rect 9080 39172 9136 39228
rect 9184 39172 9240 39228
rect 9288 39172 9344 39228
rect 9392 39172 9448 39228
rect 17768 39172 17824 39228
rect 17872 39172 17928 39228
rect 17976 39172 18032 39228
rect 18080 39172 18136 39228
rect 18184 39172 18240 39228
rect 18288 39172 18344 39228
rect 18392 39172 18448 39228
rect 26768 39172 26824 39228
rect 26872 39172 26928 39228
rect 26976 39172 27032 39228
rect 27080 39172 27136 39228
rect 27184 39172 27240 39228
rect 27288 39172 27344 39228
rect 27392 39172 27448 39228
rect 35768 39172 35824 39228
rect 35872 39172 35928 39228
rect 35976 39172 36032 39228
rect 36080 39172 36136 39228
rect 36184 39172 36240 39228
rect 36288 39172 36344 39228
rect 36392 39172 36448 39228
rect 44768 39172 44824 39228
rect 44872 39172 44928 39228
rect 44976 39172 45032 39228
rect 45080 39172 45136 39228
rect 45184 39172 45240 39228
rect 45288 39172 45344 39228
rect 45392 39172 45448 39228
rect 53768 39172 53824 39228
rect 53872 39172 53928 39228
rect 53976 39172 54032 39228
rect 54080 39172 54136 39228
rect 54184 39172 54240 39228
rect 54288 39172 54344 39228
rect 54392 39172 54448 39228
rect 62768 39172 62824 39228
rect 62872 39172 62928 39228
rect 62976 39172 63032 39228
rect 63080 39172 63136 39228
rect 63184 39172 63240 39228
rect 63288 39172 63344 39228
rect 63392 39172 63448 39228
rect 71768 39172 71824 39228
rect 71872 39172 71928 39228
rect 71976 39172 72032 39228
rect 72080 39172 72136 39228
rect 72184 39172 72240 39228
rect 72288 39172 72344 39228
rect 72392 39172 72448 39228
rect 80768 39172 80824 39228
rect 80872 39172 80928 39228
rect 80976 39172 81032 39228
rect 81080 39172 81136 39228
rect 81184 39172 81240 39228
rect 81288 39172 81344 39228
rect 81392 39172 81448 39228
rect 89768 39172 89824 39228
rect 89872 39172 89928 39228
rect 89976 39172 90032 39228
rect 90080 39172 90136 39228
rect 90184 39172 90240 39228
rect 90288 39172 90344 39228
rect 90392 39172 90448 39228
rect 4268 38388 4324 38444
rect 4372 38388 4428 38444
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 4788 38388 4844 38444
rect 4892 38388 4948 38444
rect 13268 38388 13324 38444
rect 13372 38388 13428 38444
rect 13476 38388 13532 38444
rect 13580 38388 13636 38444
rect 13684 38388 13740 38444
rect 13788 38388 13844 38444
rect 13892 38388 13948 38444
rect 22268 38388 22324 38444
rect 22372 38388 22428 38444
rect 22476 38388 22532 38444
rect 22580 38388 22636 38444
rect 22684 38388 22740 38444
rect 22788 38388 22844 38444
rect 22892 38388 22948 38444
rect 31268 38388 31324 38444
rect 31372 38388 31428 38444
rect 31476 38388 31532 38444
rect 31580 38388 31636 38444
rect 31684 38388 31740 38444
rect 31788 38388 31844 38444
rect 31892 38388 31948 38444
rect 40268 38388 40324 38444
rect 40372 38388 40428 38444
rect 40476 38388 40532 38444
rect 40580 38388 40636 38444
rect 40684 38388 40740 38444
rect 40788 38388 40844 38444
rect 40892 38388 40948 38444
rect 49268 38388 49324 38444
rect 49372 38388 49428 38444
rect 49476 38388 49532 38444
rect 49580 38388 49636 38444
rect 49684 38388 49740 38444
rect 49788 38388 49844 38444
rect 49892 38388 49948 38444
rect 58268 38388 58324 38444
rect 58372 38388 58428 38444
rect 58476 38388 58532 38444
rect 58580 38388 58636 38444
rect 58684 38388 58740 38444
rect 58788 38388 58844 38444
rect 58892 38388 58948 38444
rect 67268 38388 67324 38444
rect 67372 38388 67428 38444
rect 67476 38388 67532 38444
rect 67580 38388 67636 38444
rect 67684 38388 67740 38444
rect 67788 38388 67844 38444
rect 67892 38388 67948 38444
rect 76268 38388 76324 38444
rect 76372 38388 76428 38444
rect 76476 38388 76532 38444
rect 76580 38388 76636 38444
rect 76684 38388 76740 38444
rect 76788 38388 76844 38444
rect 76892 38388 76948 38444
rect 85268 38388 85324 38444
rect 85372 38388 85428 38444
rect 85476 38388 85532 38444
rect 85580 38388 85636 38444
rect 85684 38388 85740 38444
rect 85788 38388 85844 38444
rect 85892 38388 85948 38444
rect 94268 38388 94324 38444
rect 94372 38388 94428 38444
rect 94476 38388 94532 38444
rect 94580 38388 94636 38444
rect 94684 38388 94740 38444
rect 94788 38388 94844 38444
rect 94892 38388 94948 38444
rect 8768 37604 8824 37660
rect 8872 37604 8928 37660
rect 8976 37604 9032 37660
rect 9080 37604 9136 37660
rect 9184 37604 9240 37660
rect 9288 37604 9344 37660
rect 9392 37604 9448 37660
rect 17768 37604 17824 37660
rect 17872 37604 17928 37660
rect 17976 37604 18032 37660
rect 18080 37604 18136 37660
rect 18184 37604 18240 37660
rect 18288 37604 18344 37660
rect 18392 37604 18448 37660
rect 26768 37604 26824 37660
rect 26872 37604 26928 37660
rect 26976 37604 27032 37660
rect 27080 37604 27136 37660
rect 27184 37604 27240 37660
rect 27288 37604 27344 37660
rect 27392 37604 27448 37660
rect 35768 37604 35824 37660
rect 35872 37604 35928 37660
rect 35976 37604 36032 37660
rect 36080 37604 36136 37660
rect 36184 37604 36240 37660
rect 36288 37604 36344 37660
rect 36392 37604 36448 37660
rect 44768 37604 44824 37660
rect 44872 37604 44928 37660
rect 44976 37604 45032 37660
rect 45080 37604 45136 37660
rect 45184 37604 45240 37660
rect 45288 37604 45344 37660
rect 45392 37604 45448 37660
rect 53768 37604 53824 37660
rect 53872 37604 53928 37660
rect 53976 37604 54032 37660
rect 54080 37604 54136 37660
rect 54184 37604 54240 37660
rect 54288 37604 54344 37660
rect 54392 37604 54448 37660
rect 62768 37604 62824 37660
rect 62872 37604 62928 37660
rect 62976 37604 63032 37660
rect 63080 37604 63136 37660
rect 63184 37604 63240 37660
rect 63288 37604 63344 37660
rect 63392 37604 63448 37660
rect 71768 37604 71824 37660
rect 71872 37604 71928 37660
rect 71976 37604 72032 37660
rect 72080 37604 72136 37660
rect 72184 37604 72240 37660
rect 72288 37604 72344 37660
rect 72392 37604 72448 37660
rect 80768 37604 80824 37660
rect 80872 37604 80928 37660
rect 80976 37604 81032 37660
rect 81080 37604 81136 37660
rect 81184 37604 81240 37660
rect 81288 37604 81344 37660
rect 81392 37604 81448 37660
rect 89768 37604 89824 37660
rect 89872 37604 89928 37660
rect 89976 37604 90032 37660
rect 90080 37604 90136 37660
rect 90184 37604 90240 37660
rect 90288 37604 90344 37660
rect 90392 37604 90448 37660
rect 68236 37548 68292 37604
rect 4268 36820 4324 36876
rect 4372 36820 4428 36876
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 4788 36820 4844 36876
rect 4892 36820 4948 36876
rect 13268 36820 13324 36876
rect 13372 36820 13428 36876
rect 13476 36820 13532 36876
rect 13580 36820 13636 36876
rect 13684 36820 13740 36876
rect 13788 36820 13844 36876
rect 13892 36820 13948 36876
rect 22268 36820 22324 36876
rect 22372 36820 22428 36876
rect 22476 36820 22532 36876
rect 22580 36820 22636 36876
rect 22684 36820 22740 36876
rect 22788 36820 22844 36876
rect 22892 36820 22948 36876
rect 31268 36820 31324 36876
rect 31372 36820 31428 36876
rect 31476 36820 31532 36876
rect 31580 36820 31636 36876
rect 31684 36820 31740 36876
rect 31788 36820 31844 36876
rect 31892 36820 31948 36876
rect 40268 36820 40324 36876
rect 40372 36820 40428 36876
rect 40476 36820 40532 36876
rect 40580 36820 40636 36876
rect 40684 36820 40740 36876
rect 40788 36820 40844 36876
rect 40892 36820 40948 36876
rect 49268 36820 49324 36876
rect 49372 36820 49428 36876
rect 49476 36820 49532 36876
rect 49580 36820 49636 36876
rect 49684 36820 49740 36876
rect 49788 36820 49844 36876
rect 49892 36820 49948 36876
rect 58268 36820 58324 36876
rect 58372 36820 58428 36876
rect 58476 36820 58532 36876
rect 58580 36820 58636 36876
rect 58684 36820 58740 36876
rect 58788 36820 58844 36876
rect 58892 36820 58948 36876
rect 67268 36820 67324 36876
rect 67372 36820 67428 36876
rect 67476 36820 67532 36876
rect 67580 36820 67636 36876
rect 67684 36820 67740 36876
rect 67788 36820 67844 36876
rect 67892 36820 67948 36876
rect 76268 36820 76324 36876
rect 76372 36820 76428 36876
rect 76476 36820 76532 36876
rect 76580 36820 76636 36876
rect 76684 36820 76740 36876
rect 76788 36820 76844 36876
rect 76892 36820 76948 36876
rect 85268 36820 85324 36876
rect 85372 36820 85428 36876
rect 85476 36820 85532 36876
rect 85580 36820 85636 36876
rect 85684 36820 85740 36876
rect 85788 36820 85844 36876
rect 85892 36820 85948 36876
rect 94268 36820 94324 36876
rect 94372 36820 94428 36876
rect 94476 36820 94532 36876
rect 94580 36820 94636 36876
rect 94684 36820 94740 36876
rect 94788 36820 94844 36876
rect 94892 36820 94948 36876
rect 8768 36036 8824 36092
rect 8872 36036 8928 36092
rect 8976 36036 9032 36092
rect 9080 36036 9136 36092
rect 9184 36036 9240 36092
rect 9288 36036 9344 36092
rect 9392 36036 9448 36092
rect 17768 36036 17824 36092
rect 17872 36036 17928 36092
rect 17976 36036 18032 36092
rect 18080 36036 18136 36092
rect 18184 36036 18240 36092
rect 18288 36036 18344 36092
rect 18392 36036 18448 36092
rect 26768 36036 26824 36092
rect 26872 36036 26928 36092
rect 26976 36036 27032 36092
rect 27080 36036 27136 36092
rect 27184 36036 27240 36092
rect 27288 36036 27344 36092
rect 27392 36036 27448 36092
rect 35768 36036 35824 36092
rect 35872 36036 35928 36092
rect 35976 36036 36032 36092
rect 36080 36036 36136 36092
rect 36184 36036 36240 36092
rect 36288 36036 36344 36092
rect 36392 36036 36448 36092
rect 44768 36036 44824 36092
rect 44872 36036 44928 36092
rect 44976 36036 45032 36092
rect 45080 36036 45136 36092
rect 45184 36036 45240 36092
rect 45288 36036 45344 36092
rect 45392 36036 45448 36092
rect 53768 36036 53824 36092
rect 53872 36036 53928 36092
rect 53976 36036 54032 36092
rect 54080 36036 54136 36092
rect 54184 36036 54240 36092
rect 54288 36036 54344 36092
rect 54392 36036 54448 36092
rect 62768 36036 62824 36092
rect 62872 36036 62928 36092
rect 62976 36036 63032 36092
rect 63080 36036 63136 36092
rect 63184 36036 63240 36092
rect 63288 36036 63344 36092
rect 63392 36036 63448 36092
rect 71768 36036 71824 36092
rect 71872 36036 71928 36092
rect 71976 36036 72032 36092
rect 72080 36036 72136 36092
rect 72184 36036 72240 36092
rect 72288 36036 72344 36092
rect 72392 36036 72448 36092
rect 80768 36036 80824 36092
rect 80872 36036 80928 36092
rect 80976 36036 81032 36092
rect 81080 36036 81136 36092
rect 81184 36036 81240 36092
rect 81288 36036 81344 36092
rect 81392 36036 81448 36092
rect 89768 36036 89824 36092
rect 89872 36036 89928 36092
rect 89976 36036 90032 36092
rect 90080 36036 90136 36092
rect 90184 36036 90240 36092
rect 90288 36036 90344 36092
rect 90392 36036 90448 36092
rect 68236 35644 68292 35700
rect 4268 35252 4324 35308
rect 4372 35252 4428 35308
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 4788 35252 4844 35308
rect 4892 35252 4948 35308
rect 13268 35252 13324 35308
rect 13372 35252 13428 35308
rect 13476 35252 13532 35308
rect 13580 35252 13636 35308
rect 13684 35252 13740 35308
rect 13788 35252 13844 35308
rect 13892 35252 13948 35308
rect 22268 35252 22324 35308
rect 22372 35252 22428 35308
rect 22476 35252 22532 35308
rect 22580 35252 22636 35308
rect 22684 35252 22740 35308
rect 22788 35252 22844 35308
rect 22892 35252 22948 35308
rect 31268 35252 31324 35308
rect 31372 35252 31428 35308
rect 31476 35252 31532 35308
rect 31580 35252 31636 35308
rect 31684 35252 31740 35308
rect 31788 35252 31844 35308
rect 31892 35252 31948 35308
rect 40268 35252 40324 35308
rect 40372 35252 40428 35308
rect 40476 35252 40532 35308
rect 40580 35252 40636 35308
rect 40684 35252 40740 35308
rect 40788 35252 40844 35308
rect 40892 35252 40948 35308
rect 49268 35252 49324 35308
rect 49372 35252 49428 35308
rect 49476 35252 49532 35308
rect 49580 35252 49636 35308
rect 49684 35252 49740 35308
rect 49788 35252 49844 35308
rect 49892 35252 49948 35308
rect 58268 35252 58324 35308
rect 58372 35252 58428 35308
rect 58476 35252 58532 35308
rect 58580 35252 58636 35308
rect 58684 35252 58740 35308
rect 58788 35252 58844 35308
rect 58892 35252 58948 35308
rect 67268 35252 67324 35308
rect 67372 35252 67428 35308
rect 67476 35252 67532 35308
rect 67580 35252 67636 35308
rect 67684 35252 67740 35308
rect 67788 35252 67844 35308
rect 67892 35252 67948 35308
rect 76268 35252 76324 35308
rect 76372 35252 76428 35308
rect 76476 35252 76532 35308
rect 76580 35252 76636 35308
rect 76684 35252 76740 35308
rect 76788 35252 76844 35308
rect 76892 35252 76948 35308
rect 85268 35252 85324 35308
rect 85372 35252 85428 35308
rect 85476 35252 85532 35308
rect 85580 35252 85636 35308
rect 85684 35252 85740 35308
rect 85788 35252 85844 35308
rect 85892 35252 85948 35308
rect 94268 35252 94324 35308
rect 94372 35252 94428 35308
rect 94476 35252 94532 35308
rect 94580 35252 94636 35308
rect 94684 35252 94740 35308
rect 94788 35252 94844 35308
rect 94892 35252 94948 35308
rect 8768 34468 8824 34524
rect 8872 34468 8928 34524
rect 8976 34468 9032 34524
rect 9080 34468 9136 34524
rect 9184 34468 9240 34524
rect 9288 34468 9344 34524
rect 9392 34468 9448 34524
rect 17768 34468 17824 34524
rect 17872 34468 17928 34524
rect 17976 34468 18032 34524
rect 18080 34468 18136 34524
rect 18184 34468 18240 34524
rect 18288 34468 18344 34524
rect 18392 34468 18448 34524
rect 26768 34468 26824 34524
rect 26872 34468 26928 34524
rect 26976 34468 27032 34524
rect 27080 34468 27136 34524
rect 27184 34468 27240 34524
rect 27288 34468 27344 34524
rect 27392 34468 27448 34524
rect 35768 34468 35824 34524
rect 35872 34468 35928 34524
rect 35976 34468 36032 34524
rect 36080 34468 36136 34524
rect 36184 34468 36240 34524
rect 36288 34468 36344 34524
rect 36392 34468 36448 34524
rect 44768 34468 44824 34524
rect 44872 34468 44928 34524
rect 44976 34468 45032 34524
rect 45080 34468 45136 34524
rect 45184 34468 45240 34524
rect 45288 34468 45344 34524
rect 45392 34468 45448 34524
rect 53768 34468 53824 34524
rect 53872 34468 53928 34524
rect 53976 34468 54032 34524
rect 54080 34468 54136 34524
rect 54184 34468 54240 34524
rect 54288 34468 54344 34524
rect 54392 34468 54448 34524
rect 62768 34468 62824 34524
rect 62872 34468 62928 34524
rect 62976 34468 63032 34524
rect 63080 34468 63136 34524
rect 63184 34468 63240 34524
rect 63288 34468 63344 34524
rect 63392 34468 63448 34524
rect 71768 34468 71824 34524
rect 71872 34468 71928 34524
rect 71976 34468 72032 34524
rect 72080 34468 72136 34524
rect 72184 34468 72240 34524
rect 72288 34468 72344 34524
rect 72392 34468 72448 34524
rect 80768 34468 80824 34524
rect 80872 34468 80928 34524
rect 80976 34468 81032 34524
rect 81080 34468 81136 34524
rect 81184 34468 81240 34524
rect 81288 34468 81344 34524
rect 81392 34468 81448 34524
rect 89768 34468 89824 34524
rect 89872 34468 89928 34524
rect 89976 34468 90032 34524
rect 90080 34468 90136 34524
rect 90184 34468 90240 34524
rect 90288 34468 90344 34524
rect 90392 34468 90448 34524
rect 4268 33684 4324 33740
rect 4372 33684 4428 33740
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 4788 33684 4844 33740
rect 4892 33684 4948 33740
rect 13268 33684 13324 33740
rect 13372 33684 13428 33740
rect 13476 33684 13532 33740
rect 13580 33684 13636 33740
rect 13684 33684 13740 33740
rect 13788 33684 13844 33740
rect 13892 33684 13948 33740
rect 22268 33684 22324 33740
rect 22372 33684 22428 33740
rect 22476 33684 22532 33740
rect 22580 33684 22636 33740
rect 22684 33684 22740 33740
rect 22788 33684 22844 33740
rect 22892 33684 22948 33740
rect 31268 33684 31324 33740
rect 31372 33684 31428 33740
rect 31476 33684 31532 33740
rect 31580 33684 31636 33740
rect 31684 33684 31740 33740
rect 31788 33684 31844 33740
rect 31892 33684 31948 33740
rect 40268 33684 40324 33740
rect 40372 33684 40428 33740
rect 40476 33684 40532 33740
rect 40580 33684 40636 33740
rect 40684 33684 40740 33740
rect 40788 33684 40844 33740
rect 40892 33684 40948 33740
rect 49268 33684 49324 33740
rect 49372 33684 49428 33740
rect 49476 33684 49532 33740
rect 49580 33684 49636 33740
rect 49684 33684 49740 33740
rect 49788 33684 49844 33740
rect 49892 33684 49948 33740
rect 58268 33684 58324 33740
rect 58372 33684 58428 33740
rect 58476 33684 58532 33740
rect 58580 33684 58636 33740
rect 58684 33684 58740 33740
rect 58788 33684 58844 33740
rect 58892 33684 58948 33740
rect 67268 33684 67324 33740
rect 67372 33684 67428 33740
rect 67476 33684 67532 33740
rect 67580 33684 67636 33740
rect 67684 33684 67740 33740
rect 67788 33684 67844 33740
rect 67892 33684 67948 33740
rect 76268 33684 76324 33740
rect 76372 33684 76428 33740
rect 76476 33684 76532 33740
rect 76580 33684 76636 33740
rect 76684 33684 76740 33740
rect 76788 33684 76844 33740
rect 76892 33684 76948 33740
rect 85268 33684 85324 33740
rect 85372 33684 85428 33740
rect 85476 33684 85532 33740
rect 85580 33684 85636 33740
rect 85684 33684 85740 33740
rect 85788 33684 85844 33740
rect 85892 33684 85948 33740
rect 94268 33684 94324 33740
rect 94372 33684 94428 33740
rect 94476 33684 94532 33740
rect 94580 33684 94636 33740
rect 94684 33684 94740 33740
rect 94788 33684 94844 33740
rect 94892 33684 94948 33740
rect 8768 32900 8824 32956
rect 8872 32900 8928 32956
rect 8976 32900 9032 32956
rect 9080 32900 9136 32956
rect 9184 32900 9240 32956
rect 9288 32900 9344 32956
rect 9392 32900 9448 32956
rect 17768 32900 17824 32956
rect 17872 32900 17928 32956
rect 17976 32900 18032 32956
rect 18080 32900 18136 32956
rect 18184 32900 18240 32956
rect 18288 32900 18344 32956
rect 18392 32900 18448 32956
rect 26768 32900 26824 32956
rect 26872 32900 26928 32956
rect 26976 32900 27032 32956
rect 27080 32900 27136 32956
rect 27184 32900 27240 32956
rect 27288 32900 27344 32956
rect 27392 32900 27448 32956
rect 35768 32900 35824 32956
rect 35872 32900 35928 32956
rect 35976 32900 36032 32956
rect 36080 32900 36136 32956
rect 36184 32900 36240 32956
rect 36288 32900 36344 32956
rect 36392 32900 36448 32956
rect 44768 32900 44824 32956
rect 44872 32900 44928 32956
rect 44976 32900 45032 32956
rect 45080 32900 45136 32956
rect 45184 32900 45240 32956
rect 45288 32900 45344 32956
rect 45392 32900 45448 32956
rect 53768 32900 53824 32956
rect 53872 32900 53928 32956
rect 53976 32900 54032 32956
rect 54080 32900 54136 32956
rect 54184 32900 54240 32956
rect 54288 32900 54344 32956
rect 54392 32900 54448 32956
rect 62768 32900 62824 32956
rect 62872 32900 62928 32956
rect 62976 32900 63032 32956
rect 63080 32900 63136 32956
rect 63184 32900 63240 32956
rect 63288 32900 63344 32956
rect 63392 32900 63448 32956
rect 71768 32900 71824 32956
rect 71872 32900 71928 32956
rect 71976 32900 72032 32956
rect 72080 32900 72136 32956
rect 72184 32900 72240 32956
rect 72288 32900 72344 32956
rect 72392 32900 72448 32956
rect 80768 32900 80824 32956
rect 80872 32900 80928 32956
rect 80976 32900 81032 32956
rect 81080 32900 81136 32956
rect 81184 32900 81240 32956
rect 81288 32900 81344 32956
rect 81392 32900 81448 32956
rect 89768 32900 89824 32956
rect 89872 32900 89928 32956
rect 89976 32900 90032 32956
rect 90080 32900 90136 32956
rect 90184 32900 90240 32956
rect 90288 32900 90344 32956
rect 90392 32900 90448 32956
rect 4268 32116 4324 32172
rect 4372 32116 4428 32172
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 4788 32116 4844 32172
rect 4892 32116 4948 32172
rect 13268 32116 13324 32172
rect 13372 32116 13428 32172
rect 13476 32116 13532 32172
rect 13580 32116 13636 32172
rect 13684 32116 13740 32172
rect 13788 32116 13844 32172
rect 13892 32116 13948 32172
rect 22268 32116 22324 32172
rect 22372 32116 22428 32172
rect 22476 32116 22532 32172
rect 22580 32116 22636 32172
rect 22684 32116 22740 32172
rect 22788 32116 22844 32172
rect 22892 32116 22948 32172
rect 31268 32116 31324 32172
rect 31372 32116 31428 32172
rect 31476 32116 31532 32172
rect 31580 32116 31636 32172
rect 31684 32116 31740 32172
rect 31788 32116 31844 32172
rect 31892 32116 31948 32172
rect 40268 32116 40324 32172
rect 40372 32116 40428 32172
rect 40476 32116 40532 32172
rect 40580 32116 40636 32172
rect 40684 32116 40740 32172
rect 40788 32116 40844 32172
rect 40892 32116 40948 32172
rect 49268 32116 49324 32172
rect 49372 32116 49428 32172
rect 49476 32116 49532 32172
rect 49580 32116 49636 32172
rect 49684 32116 49740 32172
rect 49788 32116 49844 32172
rect 49892 32116 49948 32172
rect 58268 32116 58324 32172
rect 58372 32116 58428 32172
rect 58476 32116 58532 32172
rect 58580 32116 58636 32172
rect 58684 32116 58740 32172
rect 58788 32116 58844 32172
rect 58892 32116 58948 32172
rect 67268 32116 67324 32172
rect 67372 32116 67428 32172
rect 67476 32116 67532 32172
rect 67580 32116 67636 32172
rect 67684 32116 67740 32172
rect 67788 32116 67844 32172
rect 67892 32116 67948 32172
rect 76268 32116 76324 32172
rect 76372 32116 76428 32172
rect 76476 32116 76532 32172
rect 76580 32116 76636 32172
rect 76684 32116 76740 32172
rect 76788 32116 76844 32172
rect 76892 32116 76948 32172
rect 85268 32116 85324 32172
rect 85372 32116 85428 32172
rect 85476 32116 85532 32172
rect 85580 32116 85636 32172
rect 85684 32116 85740 32172
rect 85788 32116 85844 32172
rect 85892 32116 85948 32172
rect 94268 32116 94324 32172
rect 94372 32116 94428 32172
rect 94476 32116 94532 32172
rect 94580 32116 94636 32172
rect 94684 32116 94740 32172
rect 94788 32116 94844 32172
rect 94892 32116 94948 32172
rect 8768 31332 8824 31388
rect 8872 31332 8928 31388
rect 8976 31332 9032 31388
rect 9080 31332 9136 31388
rect 9184 31332 9240 31388
rect 9288 31332 9344 31388
rect 9392 31332 9448 31388
rect 17768 31332 17824 31388
rect 17872 31332 17928 31388
rect 17976 31332 18032 31388
rect 18080 31332 18136 31388
rect 18184 31332 18240 31388
rect 18288 31332 18344 31388
rect 18392 31332 18448 31388
rect 26768 31332 26824 31388
rect 26872 31332 26928 31388
rect 26976 31332 27032 31388
rect 27080 31332 27136 31388
rect 27184 31332 27240 31388
rect 27288 31332 27344 31388
rect 27392 31332 27448 31388
rect 35768 31332 35824 31388
rect 35872 31332 35928 31388
rect 35976 31332 36032 31388
rect 36080 31332 36136 31388
rect 36184 31332 36240 31388
rect 36288 31332 36344 31388
rect 36392 31332 36448 31388
rect 44768 31332 44824 31388
rect 44872 31332 44928 31388
rect 44976 31332 45032 31388
rect 45080 31332 45136 31388
rect 45184 31332 45240 31388
rect 45288 31332 45344 31388
rect 45392 31332 45448 31388
rect 53768 31332 53824 31388
rect 53872 31332 53928 31388
rect 53976 31332 54032 31388
rect 54080 31332 54136 31388
rect 54184 31332 54240 31388
rect 54288 31332 54344 31388
rect 54392 31332 54448 31388
rect 62768 31332 62824 31388
rect 62872 31332 62928 31388
rect 62976 31332 63032 31388
rect 63080 31332 63136 31388
rect 63184 31332 63240 31388
rect 63288 31332 63344 31388
rect 63392 31332 63448 31388
rect 71768 31332 71824 31388
rect 71872 31332 71928 31388
rect 71976 31332 72032 31388
rect 72080 31332 72136 31388
rect 72184 31332 72240 31388
rect 72288 31332 72344 31388
rect 72392 31332 72448 31388
rect 80768 31332 80824 31388
rect 80872 31332 80928 31388
rect 80976 31332 81032 31388
rect 81080 31332 81136 31388
rect 81184 31332 81240 31388
rect 81288 31332 81344 31388
rect 81392 31332 81448 31388
rect 89768 31332 89824 31388
rect 89872 31332 89928 31388
rect 89976 31332 90032 31388
rect 90080 31332 90136 31388
rect 90184 31332 90240 31388
rect 90288 31332 90344 31388
rect 90392 31332 90448 31388
rect 4268 30548 4324 30604
rect 4372 30548 4428 30604
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 4788 30548 4844 30604
rect 4892 30548 4948 30604
rect 13268 30548 13324 30604
rect 13372 30548 13428 30604
rect 13476 30548 13532 30604
rect 13580 30548 13636 30604
rect 13684 30548 13740 30604
rect 13788 30548 13844 30604
rect 13892 30548 13948 30604
rect 22268 30548 22324 30604
rect 22372 30548 22428 30604
rect 22476 30548 22532 30604
rect 22580 30548 22636 30604
rect 22684 30548 22740 30604
rect 22788 30548 22844 30604
rect 22892 30548 22948 30604
rect 31268 30548 31324 30604
rect 31372 30548 31428 30604
rect 31476 30548 31532 30604
rect 31580 30548 31636 30604
rect 31684 30548 31740 30604
rect 31788 30548 31844 30604
rect 31892 30548 31948 30604
rect 40268 30548 40324 30604
rect 40372 30548 40428 30604
rect 40476 30548 40532 30604
rect 40580 30548 40636 30604
rect 40684 30548 40740 30604
rect 40788 30548 40844 30604
rect 40892 30548 40948 30604
rect 49268 30548 49324 30604
rect 49372 30548 49428 30604
rect 49476 30548 49532 30604
rect 49580 30548 49636 30604
rect 49684 30548 49740 30604
rect 49788 30548 49844 30604
rect 49892 30548 49948 30604
rect 58268 30548 58324 30604
rect 58372 30548 58428 30604
rect 58476 30548 58532 30604
rect 58580 30548 58636 30604
rect 58684 30548 58740 30604
rect 58788 30548 58844 30604
rect 58892 30548 58948 30604
rect 67268 30548 67324 30604
rect 67372 30548 67428 30604
rect 67476 30548 67532 30604
rect 67580 30548 67636 30604
rect 67684 30548 67740 30604
rect 67788 30548 67844 30604
rect 67892 30548 67948 30604
rect 76268 30548 76324 30604
rect 76372 30548 76428 30604
rect 76476 30548 76532 30604
rect 76580 30548 76636 30604
rect 76684 30548 76740 30604
rect 76788 30548 76844 30604
rect 76892 30548 76948 30604
rect 85268 30548 85324 30604
rect 85372 30548 85428 30604
rect 85476 30548 85532 30604
rect 85580 30548 85636 30604
rect 85684 30548 85740 30604
rect 85788 30548 85844 30604
rect 85892 30548 85948 30604
rect 94268 30548 94324 30604
rect 94372 30548 94428 30604
rect 94476 30548 94532 30604
rect 94580 30548 94636 30604
rect 94684 30548 94740 30604
rect 94788 30548 94844 30604
rect 94892 30548 94948 30604
rect 8768 29764 8824 29820
rect 8872 29764 8928 29820
rect 8976 29764 9032 29820
rect 9080 29764 9136 29820
rect 9184 29764 9240 29820
rect 9288 29764 9344 29820
rect 9392 29764 9448 29820
rect 17768 29764 17824 29820
rect 17872 29764 17928 29820
rect 17976 29764 18032 29820
rect 18080 29764 18136 29820
rect 18184 29764 18240 29820
rect 18288 29764 18344 29820
rect 18392 29764 18448 29820
rect 26768 29764 26824 29820
rect 26872 29764 26928 29820
rect 26976 29764 27032 29820
rect 27080 29764 27136 29820
rect 27184 29764 27240 29820
rect 27288 29764 27344 29820
rect 27392 29764 27448 29820
rect 35768 29764 35824 29820
rect 35872 29764 35928 29820
rect 35976 29764 36032 29820
rect 36080 29764 36136 29820
rect 36184 29764 36240 29820
rect 36288 29764 36344 29820
rect 36392 29764 36448 29820
rect 44768 29764 44824 29820
rect 44872 29764 44928 29820
rect 44976 29764 45032 29820
rect 45080 29764 45136 29820
rect 45184 29764 45240 29820
rect 45288 29764 45344 29820
rect 45392 29764 45448 29820
rect 53768 29764 53824 29820
rect 53872 29764 53928 29820
rect 53976 29764 54032 29820
rect 54080 29764 54136 29820
rect 54184 29764 54240 29820
rect 54288 29764 54344 29820
rect 54392 29764 54448 29820
rect 62768 29764 62824 29820
rect 62872 29764 62928 29820
rect 62976 29764 63032 29820
rect 63080 29764 63136 29820
rect 63184 29764 63240 29820
rect 63288 29764 63344 29820
rect 63392 29764 63448 29820
rect 71768 29764 71824 29820
rect 71872 29764 71928 29820
rect 71976 29764 72032 29820
rect 72080 29764 72136 29820
rect 72184 29764 72240 29820
rect 72288 29764 72344 29820
rect 72392 29764 72448 29820
rect 80768 29764 80824 29820
rect 80872 29764 80928 29820
rect 80976 29764 81032 29820
rect 81080 29764 81136 29820
rect 81184 29764 81240 29820
rect 81288 29764 81344 29820
rect 81392 29764 81448 29820
rect 89768 29764 89824 29820
rect 89872 29764 89928 29820
rect 89976 29764 90032 29820
rect 90080 29764 90136 29820
rect 90184 29764 90240 29820
rect 90288 29764 90344 29820
rect 90392 29764 90448 29820
rect 4268 28980 4324 29036
rect 4372 28980 4428 29036
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 4788 28980 4844 29036
rect 4892 28980 4948 29036
rect 13268 28980 13324 29036
rect 13372 28980 13428 29036
rect 13476 28980 13532 29036
rect 13580 28980 13636 29036
rect 13684 28980 13740 29036
rect 13788 28980 13844 29036
rect 13892 28980 13948 29036
rect 22268 28980 22324 29036
rect 22372 28980 22428 29036
rect 22476 28980 22532 29036
rect 22580 28980 22636 29036
rect 22684 28980 22740 29036
rect 22788 28980 22844 29036
rect 22892 28980 22948 29036
rect 31268 28980 31324 29036
rect 31372 28980 31428 29036
rect 31476 28980 31532 29036
rect 31580 28980 31636 29036
rect 31684 28980 31740 29036
rect 31788 28980 31844 29036
rect 31892 28980 31948 29036
rect 40268 28980 40324 29036
rect 40372 28980 40428 29036
rect 40476 28980 40532 29036
rect 40580 28980 40636 29036
rect 40684 28980 40740 29036
rect 40788 28980 40844 29036
rect 40892 28980 40948 29036
rect 49268 28980 49324 29036
rect 49372 28980 49428 29036
rect 49476 28980 49532 29036
rect 49580 28980 49636 29036
rect 49684 28980 49740 29036
rect 49788 28980 49844 29036
rect 49892 28980 49948 29036
rect 58268 28980 58324 29036
rect 58372 28980 58428 29036
rect 58476 28980 58532 29036
rect 58580 28980 58636 29036
rect 58684 28980 58740 29036
rect 58788 28980 58844 29036
rect 58892 28980 58948 29036
rect 67268 28980 67324 29036
rect 67372 28980 67428 29036
rect 67476 28980 67532 29036
rect 67580 28980 67636 29036
rect 67684 28980 67740 29036
rect 67788 28980 67844 29036
rect 67892 28980 67948 29036
rect 76268 28980 76324 29036
rect 76372 28980 76428 29036
rect 76476 28980 76532 29036
rect 76580 28980 76636 29036
rect 76684 28980 76740 29036
rect 76788 28980 76844 29036
rect 76892 28980 76948 29036
rect 85268 28980 85324 29036
rect 85372 28980 85428 29036
rect 85476 28980 85532 29036
rect 85580 28980 85636 29036
rect 85684 28980 85740 29036
rect 85788 28980 85844 29036
rect 85892 28980 85948 29036
rect 94268 28980 94324 29036
rect 94372 28980 94428 29036
rect 94476 28980 94532 29036
rect 94580 28980 94636 29036
rect 94684 28980 94740 29036
rect 94788 28980 94844 29036
rect 94892 28980 94948 29036
rect 68124 28588 68180 28644
rect 8768 28196 8824 28252
rect 8872 28196 8928 28252
rect 8976 28196 9032 28252
rect 9080 28196 9136 28252
rect 9184 28196 9240 28252
rect 9288 28196 9344 28252
rect 9392 28196 9448 28252
rect 17768 28196 17824 28252
rect 17872 28196 17928 28252
rect 17976 28196 18032 28252
rect 18080 28196 18136 28252
rect 18184 28196 18240 28252
rect 18288 28196 18344 28252
rect 18392 28196 18448 28252
rect 26768 28196 26824 28252
rect 26872 28196 26928 28252
rect 26976 28196 27032 28252
rect 27080 28196 27136 28252
rect 27184 28196 27240 28252
rect 27288 28196 27344 28252
rect 27392 28196 27448 28252
rect 35768 28196 35824 28252
rect 35872 28196 35928 28252
rect 35976 28196 36032 28252
rect 36080 28196 36136 28252
rect 36184 28196 36240 28252
rect 36288 28196 36344 28252
rect 36392 28196 36448 28252
rect 44768 28196 44824 28252
rect 44872 28196 44928 28252
rect 44976 28196 45032 28252
rect 45080 28196 45136 28252
rect 45184 28196 45240 28252
rect 45288 28196 45344 28252
rect 45392 28196 45448 28252
rect 53768 28196 53824 28252
rect 53872 28196 53928 28252
rect 53976 28196 54032 28252
rect 54080 28196 54136 28252
rect 54184 28196 54240 28252
rect 54288 28196 54344 28252
rect 54392 28196 54448 28252
rect 62768 28196 62824 28252
rect 62872 28196 62928 28252
rect 62976 28196 63032 28252
rect 63080 28196 63136 28252
rect 63184 28196 63240 28252
rect 63288 28196 63344 28252
rect 63392 28196 63448 28252
rect 71768 28196 71824 28252
rect 71872 28196 71928 28252
rect 71976 28196 72032 28252
rect 72080 28196 72136 28252
rect 72184 28196 72240 28252
rect 72288 28196 72344 28252
rect 72392 28196 72448 28252
rect 80768 28196 80824 28252
rect 80872 28196 80928 28252
rect 80976 28196 81032 28252
rect 81080 28196 81136 28252
rect 81184 28196 81240 28252
rect 81288 28196 81344 28252
rect 81392 28196 81448 28252
rect 89768 28196 89824 28252
rect 89872 28196 89928 28252
rect 89976 28196 90032 28252
rect 90080 28196 90136 28252
rect 90184 28196 90240 28252
rect 90288 28196 90344 28252
rect 90392 28196 90448 28252
rect 4268 27412 4324 27468
rect 4372 27412 4428 27468
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 4788 27412 4844 27468
rect 4892 27412 4948 27468
rect 13268 27412 13324 27468
rect 13372 27412 13428 27468
rect 13476 27412 13532 27468
rect 13580 27412 13636 27468
rect 13684 27412 13740 27468
rect 13788 27412 13844 27468
rect 13892 27412 13948 27468
rect 22268 27412 22324 27468
rect 22372 27412 22428 27468
rect 22476 27412 22532 27468
rect 22580 27412 22636 27468
rect 22684 27412 22740 27468
rect 22788 27412 22844 27468
rect 22892 27412 22948 27468
rect 31268 27412 31324 27468
rect 31372 27412 31428 27468
rect 31476 27412 31532 27468
rect 31580 27412 31636 27468
rect 31684 27412 31740 27468
rect 31788 27412 31844 27468
rect 31892 27412 31948 27468
rect 40268 27412 40324 27468
rect 40372 27412 40428 27468
rect 40476 27412 40532 27468
rect 40580 27412 40636 27468
rect 40684 27412 40740 27468
rect 40788 27412 40844 27468
rect 40892 27412 40948 27468
rect 49268 27412 49324 27468
rect 49372 27412 49428 27468
rect 49476 27412 49532 27468
rect 49580 27412 49636 27468
rect 49684 27412 49740 27468
rect 49788 27412 49844 27468
rect 49892 27412 49948 27468
rect 58268 27412 58324 27468
rect 58372 27412 58428 27468
rect 58476 27412 58532 27468
rect 58580 27412 58636 27468
rect 58684 27412 58740 27468
rect 58788 27412 58844 27468
rect 58892 27412 58948 27468
rect 67268 27412 67324 27468
rect 67372 27412 67428 27468
rect 67476 27412 67532 27468
rect 67580 27412 67636 27468
rect 67684 27412 67740 27468
rect 67788 27412 67844 27468
rect 67892 27412 67948 27468
rect 76268 27412 76324 27468
rect 76372 27412 76428 27468
rect 76476 27412 76532 27468
rect 76580 27412 76636 27468
rect 76684 27412 76740 27468
rect 76788 27412 76844 27468
rect 76892 27412 76948 27468
rect 85268 27412 85324 27468
rect 85372 27412 85428 27468
rect 85476 27412 85532 27468
rect 85580 27412 85636 27468
rect 85684 27412 85740 27468
rect 85788 27412 85844 27468
rect 85892 27412 85948 27468
rect 94268 27412 94324 27468
rect 94372 27412 94428 27468
rect 94476 27412 94532 27468
rect 94580 27412 94636 27468
rect 94684 27412 94740 27468
rect 94788 27412 94844 27468
rect 94892 27412 94948 27468
rect 8768 26628 8824 26684
rect 8872 26628 8928 26684
rect 8976 26628 9032 26684
rect 9080 26628 9136 26684
rect 9184 26628 9240 26684
rect 9288 26628 9344 26684
rect 9392 26628 9448 26684
rect 17768 26628 17824 26684
rect 17872 26628 17928 26684
rect 17976 26628 18032 26684
rect 18080 26628 18136 26684
rect 18184 26628 18240 26684
rect 18288 26628 18344 26684
rect 18392 26628 18448 26684
rect 26768 26628 26824 26684
rect 26872 26628 26928 26684
rect 26976 26628 27032 26684
rect 27080 26628 27136 26684
rect 27184 26628 27240 26684
rect 27288 26628 27344 26684
rect 27392 26628 27448 26684
rect 35768 26628 35824 26684
rect 35872 26628 35928 26684
rect 35976 26628 36032 26684
rect 36080 26628 36136 26684
rect 36184 26628 36240 26684
rect 36288 26628 36344 26684
rect 36392 26628 36448 26684
rect 44768 26628 44824 26684
rect 44872 26628 44928 26684
rect 44976 26628 45032 26684
rect 45080 26628 45136 26684
rect 45184 26628 45240 26684
rect 45288 26628 45344 26684
rect 45392 26628 45448 26684
rect 53768 26628 53824 26684
rect 53872 26628 53928 26684
rect 53976 26628 54032 26684
rect 54080 26628 54136 26684
rect 54184 26628 54240 26684
rect 54288 26628 54344 26684
rect 54392 26628 54448 26684
rect 62768 26628 62824 26684
rect 62872 26628 62928 26684
rect 62976 26628 63032 26684
rect 63080 26628 63136 26684
rect 63184 26628 63240 26684
rect 63288 26628 63344 26684
rect 63392 26628 63448 26684
rect 71768 26628 71824 26684
rect 71872 26628 71928 26684
rect 71976 26628 72032 26684
rect 72080 26628 72136 26684
rect 72184 26628 72240 26684
rect 72288 26628 72344 26684
rect 72392 26628 72448 26684
rect 80768 26628 80824 26684
rect 80872 26628 80928 26684
rect 80976 26628 81032 26684
rect 81080 26628 81136 26684
rect 81184 26628 81240 26684
rect 81288 26628 81344 26684
rect 81392 26628 81448 26684
rect 89768 26628 89824 26684
rect 89872 26628 89928 26684
rect 89976 26628 90032 26684
rect 90080 26628 90136 26684
rect 90184 26628 90240 26684
rect 90288 26628 90344 26684
rect 90392 26628 90448 26684
rect 67116 26124 67172 26180
rect 4268 25844 4324 25900
rect 4372 25844 4428 25900
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 4788 25844 4844 25900
rect 4892 25844 4948 25900
rect 13268 25844 13324 25900
rect 13372 25844 13428 25900
rect 13476 25844 13532 25900
rect 13580 25844 13636 25900
rect 13684 25844 13740 25900
rect 13788 25844 13844 25900
rect 13892 25844 13948 25900
rect 22268 25844 22324 25900
rect 22372 25844 22428 25900
rect 22476 25844 22532 25900
rect 22580 25844 22636 25900
rect 22684 25844 22740 25900
rect 22788 25844 22844 25900
rect 22892 25844 22948 25900
rect 31268 25844 31324 25900
rect 31372 25844 31428 25900
rect 31476 25844 31532 25900
rect 31580 25844 31636 25900
rect 31684 25844 31740 25900
rect 31788 25844 31844 25900
rect 31892 25844 31948 25900
rect 40268 25844 40324 25900
rect 40372 25844 40428 25900
rect 40476 25844 40532 25900
rect 40580 25844 40636 25900
rect 40684 25844 40740 25900
rect 40788 25844 40844 25900
rect 40892 25844 40948 25900
rect 49268 25844 49324 25900
rect 49372 25844 49428 25900
rect 49476 25844 49532 25900
rect 49580 25844 49636 25900
rect 49684 25844 49740 25900
rect 49788 25844 49844 25900
rect 49892 25844 49948 25900
rect 58268 25844 58324 25900
rect 58372 25844 58428 25900
rect 58476 25844 58532 25900
rect 58580 25844 58636 25900
rect 58684 25844 58740 25900
rect 58788 25844 58844 25900
rect 58892 25844 58948 25900
rect 67268 25844 67324 25900
rect 67372 25844 67428 25900
rect 67476 25844 67532 25900
rect 67580 25844 67636 25900
rect 67684 25844 67740 25900
rect 67788 25844 67844 25900
rect 67892 25844 67948 25900
rect 76268 25844 76324 25900
rect 76372 25844 76428 25900
rect 76476 25844 76532 25900
rect 76580 25844 76636 25900
rect 76684 25844 76740 25900
rect 76788 25844 76844 25900
rect 76892 25844 76948 25900
rect 85268 25844 85324 25900
rect 85372 25844 85428 25900
rect 85476 25844 85532 25900
rect 85580 25844 85636 25900
rect 85684 25844 85740 25900
rect 85788 25844 85844 25900
rect 85892 25844 85948 25900
rect 94268 25844 94324 25900
rect 94372 25844 94428 25900
rect 94476 25844 94532 25900
rect 94580 25844 94636 25900
rect 94684 25844 94740 25900
rect 94788 25844 94844 25900
rect 94892 25844 94948 25900
rect 67116 25228 67172 25284
rect 8768 25060 8824 25116
rect 8872 25060 8928 25116
rect 8976 25060 9032 25116
rect 9080 25060 9136 25116
rect 9184 25060 9240 25116
rect 9288 25060 9344 25116
rect 9392 25060 9448 25116
rect 17768 25060 17824 25116
rect 17872 25060 17928 25116
rect 17976 25060 18032 25116
rect 18080 25060 18136 25116
rect 18184 25060 18240 25116
rect 18288 25060 18344 25116
rect 18392 25060 18448 25116
rect 26768 25060 26824 25116
rect 26872 25060 26928 25116
rect 26976 25060 27032 25116
rect 27080 25060 27136 25116
rect 27184 25060 27240 25116
rect 27288 25060 27344 25116
rect 27392 25060 27448 25116
rect 35768 25060 35824 25116
rect 35872 25060 35928 25116
rect 35976 25060 36032 25116
rect 36080 25060 36136 25116
rect 36184 25060 36240 25116
rect 36288 25060 36344 25116
rect 36392 25060 36448 25116
rect 44768 25060 44824 25116
rect 44872 25060 44928 25116
rect 44976 25060 45032 25116
rect 45080 25060 45136 25116
rect 45184 25060 45240 25116
rect 45288 25060 45344 25116
rect 45392 25060 45448 25116
rect 53768 25060 53824 25116
rect 53872 25060 53928 25116
rect 53976 25060 54032 25116
rect 54080 25060 54136 25116
rect 54184 25060 54240 25116
rect 54288 25060 54344 25116
rect 54392 25060 54448 25116
rect 62768 25060 62824 25116
rect 62872 25060 62928 25116
rect 62976 25060 63032 25116
rect 63080 25060 63136 25116
rect 63184 25060 63240 25116
rect 63288 25060 63344 25116
rect 63392 25060 63448 25116
rect 71768 25060 71824 25116
rect 71872 25060 71928 25116
rect 71976 25060 72032 25116
rect 72080 25060 72136 25116
rect 72184 25060 72240 25116
rect 72288 25060 72344 25116
rect 72392 25060 72448 25116
rect 80768 25060 80824 25116
rect 80872 25060 80928 25116
rect 80976 25060 81032 25116
rect 81080 25060 81136 25116
rect 81184 25060 81240 25116
rect 81288 25060 81344 25116
rect 81392 25060 81448 25116
rect 89768 25060 89824 25116
rect 89872 25060 89928 25116
rect 89976 25060 90032 25116
rect 90080 25060 90136 25116
rect 90184 25060 90240 25116
rect 90288 25060 90344 25116
rect 90392 25060 90448 25116
rect 4268 24276 4324 24332
rect 4372 24276 4428 24332
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 4788 24276 4844 24332
rect 4892 24276 4948 24332
rect 13268 24276 13324 24332
rect 13372 24276 13428 24332
rect 13476 24276 13532 24332
rect 13580 24276 13636 24332
rect 13684 24276 13740 24332
rect 13788 24276 13844 24332
rect 13892 24276 13948 24332
rect 22268 24276 22324 24332
rect 22372 24276 22428 24332
rect 22476 24276 22532 24332
rect 22580 24276 22636 24332
rect 22684 24276 22740 24332
rect 22788 24276 22844 24332
rect 22892 24276 22948 24332
rect 31268 24276 31324 24332
rect 31372 24276 31428 24332
rect 31476 24276 31532 24332
rect 31580 24276 31636 24332
rect 31684 24276 31740 24332
rect 31788 24276 31844 24332
rect 31892 24276 31948 24332
rect 40268 24276 40324 24332
rect 40372 24276 40428 24332
rect 40476 24276 40532 24332
rect 40580 24276 40636 24332
rect 40684 24276 40740 24332
rect 40788 24276 40844 24332
rect 40892 24276 40948 24332
rect 49268 24276 49324 24332
rect 49372 24276 49428 24332
rect 49476 24276 49532 24332
rect 49580 24276 49636 24332
rect 49684 24276 49740 24332
rect 49788 24276 49844 24332
rect 49892 24276 49948 24332
rect 58268 24276 58324 24332
rect 58372 24276 58428 24332
rect 58476 24276 58532 24332
rect 58580 24276 58636 24332
rect 58684 24276 58740 24332
rect 58788 24276 58844 24332
rect 58892 24276 58948 24332
rect 67268 24276 67324 24332
rect 67372 24276 67428 24332
rect 67476 24276 67532 24332
rect 67580 24276 67636 24332
rect 67684 24276 67740 24332
rect 67788 24276 67844 24332
rect 67892 24276 67948 24332
rect 76268 24276 76324 24332
rect 76372 24276 76428 24332
rect 76476 24276 76532 24332
rect 76580 24276 76636 24332
rect 76684 24276 76740 24332
rect 76788 24276 76844 24332
rect 76892 24276 76948 24332
rect 85268 24276 85324 24332
rect 85372 24276 85428 24332
rect 85476 24276 85532 24332
rect 85580 24276 85636 24332
rect 85684 24276 85740 24332
rect 85788 24276 85844 24332
rect 85892 24276 85948 24332
rect 94268 24276 94324 24332
rect 94372 24276 94428 24332
rect 94476 24276 94532 24332
rect 94580 24276 94636 24332
rect 94684 24276 94740 24332
rect 94788 24276 94844 24332
rect 94892 24276 94948 24332
rect 8768 23492 8824 23548
rect 8872 23492 8928 23548
rect 8976 23492 9032 23548
rect 9080 23492 9136 23548
rect 9184 23492 9240 23548
rect 9288 23492 9344 23548
rect 9392 23492 9448 23548
rect 17768 23492 17824 23548
rect 17872 23492 17928 23548
rect 17976 23492 18032 23548
rect 18080 23492 18136 23548
rect 18184 23492 18240 23548
rect 18288 23492 18344 23548
rect 18392 23492 18448 23548
rect 26768 23492 26824 23548
rect 26872 23492 26928 23548
rect 26976 23492 27032 23548
rect 27080 23492 27136 23548
rect 27184 23492 27240 23548
rect 27288 23492 27344 23548
rect 27392 23492 27448 23548
rect 35768 23492 35824 23548
rect 35872 23492 35928 23548
rect 35976 23492 36032 23548
rect 36080 23492 36136 23548
rect 36184 23492 36240 23548
rect 36288 23492 36344 23548
rect 36392 23492 36448 23548
rect 44768 23492 44824 23548
rect 44872 23492 44928 23548
rect 44976 23492 45032 23548
rect 45080 23492 45136 23548
rect 45184 23492 45240 23548
rect 45288 23492 45344 23548
rect 45392 23492 45448 23548
rect 53768 23492 53824 23548
rect 53872 23492 53928 23548
rect 53976 23492 54032 23548
rect 54080 23492 54136 23548
rect 54184 23492 54240 23548
rect 54288 23492 54344 23548
rect 54392 23492 54448 23548
rect 62768 23492 62824 23548
rect 62872 23492 62928 23548
rect 62976 23492 63032 23548
rect 63080 23492 63136 23548
rect 63184 23492 63240 23548
rect 63288 23492 63344 23548
rect 63392 23492 63448 23548
rect 71768 23492 71824 23548
rect 71872 23492 71928 23548
rect 71976 23492 72032 23548
rect 72080 23492 72136 23548
rect 72184 23492 72240 23548
rect 72288 23492 72344 23548
rect 72392 23492 72448 23548
rect 80768 23492 80824 23548
rect 80872 23492 80928 23548
rect 80976 23492 81032 23548
rect 81080 23492 81136 23548
rect 81184 23492 81240 23548
rect 81288 23492 81344 23548
rect 81392 23492 81448 23548
rect 89768 23492 89824 23548
rect 89872 23492 89928 23548
rect 89976 23492 90032 23548
rect 90080 23492 90136 23548
rect 90184 23492 90240 23548
rect 90288 23492 90344 23548
rect 90392 23492 90448 23548
rect 4268 22708 4324 22764
rect 4372 22708 4428 22764
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 4788 22708 4844 22764
rect 4892 22708 4948 22764
rect 13268 22708 13324 22764
rect 13372 22708 13428 22764
rect 13476 22708 13532 22764
rect 13580 22708 13636 22764
rect 13684 22708 13740 22764
rect 13788 22708 13844 22764
rect 13892 22708 13948 22764
rect 22268 22708 22324 22764
rect 22372 22708 22428 22764
rect 22476 22708 22532 22764
rect 22580 22708 22636 22764
rect 22684 22708 22740 22764
rect 22788 22708 22844 22764
rect 22892 22708 22948 22764
rect 31268 22708 31324 22764
rect 31372 22708 31428 22764
rect 31476 22708 31532 22764
rect 31580 22708 31636 22764
rect 31684 22708 31740 22764
rect 31788 22708 31844 22764
rect 31892 22708 31948 22764
rect 40268 22708 40324 22764
rect 40372 22708 40428 22764
rect 40476 22708 40532 22764
rect 40580 22708 40636 22764
rect 40684 22708 40740 22764
rect 40788 22708 40844 22764
rect 40892 22708 40948 22764
rect 49268 22708 49324 22764
rect 49372 22708 49428 22764
rect 49476 22708 49532 22764
rect 49580 22708 49636 22764
rect 49684 22708 49740 22764
rect 49788 22708 49844 22764
rect 49892 22708 49948 22764
rect 58268 22708 58324 22764
rect 58372 22708 58428 22764
rect 58476 22708 58532 22764
rect 58580 22708 58636 22764
rect 58684 22708 58740 22764
rect 58788 22708 58844 22764
rect 58892 22708 58948 22764
rect 67268 22708 67324 22764
rect 67372 22708 67428 22764
rect 67476 22708 67532 22764
rect 67580 22708 67636 22764
rect 67684 22708 67740 22764
rect 67788 22708 67844 22764
rect 67892 22708 67948 22764
rect 76268 22708 76324 22764
rect 76372 22708 76428 22764
rect 76476 22708 76532 22764
rect 76580 22708 76636 22764
rect 76684 22708 76740 22764
rect 76788 22708 76844 22764
rect 76892 22708 76948 22764
rect 85268 22708 85324 22764
rect 85372 22708 85428 22764
rect 85476 22708 85532 22764
rect 85580 22708 85636 22764
rect 85684 22708 85740 22764
rect 85788 22708 85844 22764
rect 85892 22708 85948 22764
rect 94268 22708 94324 22764
rect 94372 22708 94428 22764
rect 94476 22708 94532 22764
rect 94580 22708 94636 22764
rect 94684 22708 94740 22764
rect 94788 22708 94844 22764
rect 94892 22708 94948 22764
rect 67116 22204 67172 22260
rect 8768 21924 8824 21980
rect 8872 21924 8928 21980
rect 8976 21924 9032 21980
rect 9080 21924 9136 21980
rect 9184 21924 9240 21980
rect 9288 21924 9344 21980
rect 9392 21924 9448 21980
rect 17768 21924 17824 21980
rect 17872 21924 17928 21980
rect 17976 21924 18032 21980
rect 18080 21924 18136 21980
rect 18184 21924 18240 21980
rect 18288 21924 18344 21980
rect 18392 21924 18448 21980
rect 26768 21924 26824 21980
rect 26872 21924 26928 21980
rect 26976 21924 27032 21980
rect 27080 21924 27136 21980
rect 27184 21924 27240 21980
rect 27288 21924 27344 21980
rect 27392 21924 27448 21980
rect 35768 21924 35824 21980
rect 35872 21924 35928 21980
rect 35976 21924 36032 21980
rect 36080 21924 36136 21980
rect 36184 21924 36240 21980
rect 36288 21924 36344 21980
rect 36392 21924 36448 21980
rect 44768 21924 44824 21980
rect 44872 21924 44928 21980
rect 44976 21924 45032 21980
rect 45080 21924 45136 21980
rect 45184 21924 45240 21980
rect 45288 21924 45344 21980
rect 45392 21924 45448 21980
rect 53768 21924 53824 21980
rect 53872 21924 53928 21980
rect 53976 21924 54032 21980
rect 54080 21924 54136 21980
rect 54184 21924 54240 21980
rect 54288 21924 54344 21980
rect 54392 21924 54448 21980
rect 62768 21924 62824 21980
rect 62872 21924 62928 21980
rect 62976 21924 63032 21980
rect 63080 21924 63136 21980
rect 63184 21924 63240 21980
rect 63288 21924 63344 21980
rect 63392 21924 63448 21980
rect 71768 21924 71824 21980
rect 71872 21924 71928 21980
rect 71976 21924 72032 21980
rect 72080 21924 72136 21980
rect 72184 21924 72240 21980
rect 72288 21924 72344 21980
rect 72392 21924 72448 21980
rect 80768 21924 80824 21980
rect 80872 21924 80928 21980
rect 80976 21924 81032 21980
rect 81080 21924 81136 21980
rect 81184 21924 81240 21980
rect 81288 21924 81344 21980
rect 81392 21924 81448 21980
rect 89768 21924 89824 21980
rect 89872 21924 89928 21980
rect 89976 21924 90032 21980
rect 90080 21924 90136 21980
rect 90184 21924 90240 21980
rect 90288 21924 90344 21980
rect 90392 21924 90448 21980
rect 68124 21644 68180 21700
rect 4268 21140 4324 21196
rect 4372 21140 4428 21196
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 4788 21140 4844 21196
rect 4892 21140 4948 21196
rect 13268 21140 13324 21196
rect 13372 21140 13428 21196
rect 13476 21140 13532 21196
rect 13580 21140 13636 21196
rect 13684 21140 13740 21196
rect 13788 21140 13844 21196
rect 13892 21140 13948 21196
rect 22268 21140 22324 21196
rect 22372 21140 22428 21196
rect 22476 21140 22532 21196
rect 22580 21140 22636 21196
rect 22684 21140 22740 21196
rect 22788 21140 22844 21196
rect 22892 21140 22948 21196
rect 31268 21140 31324 21196
rect 31372 21140 31428 21196
rect 31476 21140 31532 21196
rect 31580 21140 31636 21196
rect 31684 21140 31740 21196
rect 31788 21140 31844 21196
rect 31892 21140 31948 21196
rect 40268 21140 40324 21196
rect 40372 21140 40428 21196
rect 40476 21140 40532 21196
rect 40580 21140 40636 21196
rect 40684 21140 40740 21196
rect 40788 21140 40844 21196
rect 40892 21140 40948 21196
rect 49268 21140 49324 21196
rect 49372 21140 49428 21196
rect 49476 21140 49532 21196
rect 49580 21140 49636 21196
rect 49684 21140 49740 21196
rect 49788 21140 49844 21196
rect 49892 21140 49948 21196
rect 58268 21140 58324 21196
rect 58372 21140 58428 21196
rect 58476 21140 58532 21196
rect 58580 21140 58636 21196
rect 58684 21140 58740 21196
rect 58788 21140 58844 21196
rect 58892 21140 58948 21196
rect 67268 21140 67324 21196
rect 67372 21140 67428 21196
rect 67476 21140 67532 21196
rect 67580 21140 67636 21196
rect 67684 21140 67740 21196
rect 67788 21140 67844 21196
rect 67892 21140 67948 21196
rect 76268 21140 76324 21196
rect 76372 21140 76428 21196
rect 76476 21140 76532 21196
rect 76580 21140 76636 21196
rect 76684 21140 76740 21196
rect 76788 21140 76844 21196
rect 76892 21140 76948 21196
rect 85268 21140 85324 21196
rect 85372 21140 85428 21196
rect 85476 21140 85532 21196
rect 85580 21140 85636 21196
rect 85684 21140 85740 21196
rect 85788 21140 85844 21196
rect 85892 21140 85948 21196
rect 94268 21140 94324 21196
rect 94372 21140 94428 21196
rect 94476 21140 94532 21196
rect 94580 21140 94636 21196
rect 94684 21140 94740 21196
rect 94788 21140 94844 21196
rect 94892 21140 94948 21196
rect 8768 20356 8824 20412
rect 8872 20356 8928 20412
rect 8976 20356 9032 20412
rect 9080 20356 9136 20412
rect 9184 20356 9240 20412
rect 9288 20356 9344 20412
rect 9392 20356 9448 20412
rect 17768 20356 17824 20412
rect 17872 20356 17928 20412
rect 17976 20356 18032 20412
rect 18080 20356 18136 20412
rect 18184 20356 18240 20412
rect 18288 20356 18344 20412
rect 18392 20356 18448 20412
rect 26768 20356 26824 20412
rect 26872 20356 26928 20412
rect 26976 20356 27032 20412
rect 27080 20356 27136 20412
rect 27184 20356 27240 20412
rect 27288 20356 27344 20412
rect 27392 20356 27448 20412
rect 35768 20356 35824 20412
rect 35872 20356 35928 20412
rect 35976 20356 36032 20412
rect 36080 20356 36136 20412
rect 36184 20356 36240 20412
rect 36288 20356 36344 20412
rect 36392 20356 36448 20412
rect 44768 20356 44824 20412
rect 44872 20356 44928 20412
rect 44976 20356 45032 20412
rect 45080 20356 45136 20412
rect 45184 20356 45240 20412
rect 45288 20356 45344 20412
rect 45392 20356 45448 20412
rect 53768 20356 53824 20412
rect 53872 20356 53928 20412
rect 53976 20356 54032 20412
rect 54080 20356 54136 20412
rect 54184 20356 54240 20412
rect 54288 20356 54344 20412
rect 54392 20356 54448 20412
rect 62768 20356 62824 20412
rect 62872 20356 62928 20412
rect 62976 20356 63032 20412
rect 63080 20356 63136 20412
rect 63184 20356 63240 20412
rect 63288 20356 63344 20412
rect 63392 20356 63448 20412
rect 71768 20356 71824 20412
rect 71872 20356 71928 20412
rect 71976 20356 72032 20412
rect 72080 20356 72136 20412
rect 72184 20356 72240 20412
rect 72288 20356 72344 20412
rect 72392 20356 72448 20412
rect 80768 20356 80824 20412
rect 80872 20356 80928 20412
rect 80976 20356 81032 20412
rect 81080 20356 81136 20412
rect 81184 20356 81240 20412
rect 81288 20356 81344 20412
rect 81392 20356 81448 20412
rect 89768 20356 89824 20412
rect 89872 20356 89928 20412
rect 89976 20356 90032 20412
rect 90080 20356 90136 20412
rect 90184 20356 90240 20412
rect 90288 20356 90344 20412
rect 90392 20356 90448 20412
rect 4268 19572 4324 19628
rect 4372 19572 4428 19628
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 4788 19572 4844 19628
rect 4892 19572 4948 19628
rect 13268 19572 13324 19628
rect 13372 19572 13428 19628
rect 13476 19572 13532 19628
rect 13580 19572 13636 19628
rect 13684 19572 13740 19628
rect 13788 19572 13844 19628
rect 13892 19572 13948 19628
rect 22268 19572 22324 19628
rect 22372 19572 22428 19628
rect 22476 19572 22532 19628
rect 22580 19572 22636 19628
rect 22684 19572 22740 19628
rect 22788 19572 22844 19628
rect 22892 19572 22948 19628
rect 31268 19572 31324 19628
rect 31372 19572 31428 19628
rect 31476 19572 31532 19628
rect 31580 19572 31636 19628
rect 31684 19572 31740 19628
rect 31788 19572 31844 19628
rect 31892 19572 31948 19628
rect 40268 19572 40324 19628
rect 40372 19572 40428 19628
rect 40476 19572 40532 19628
rect 40580 19572 40636 19628
rect 40684 19572 40740 19628
rect 40788 19572 40844 19628
rect 40892 19572 40948 19628
rect 49268 19572 49324 19628
rect 49372 19572 49428 19628
rect 49476 19572 49532 19628
rect 49580 19572 49636 19628
rect 49684 19572 49740 19628
rect 49788 19572 49844 19628
rect 49892 19572 49948 19628
rect 58268 19572 58324 19628
rect 58372 19572 58428 19628
rect 58476 19572 58532 19628
rect 58580 19572 58636 19628
rect 58684 19572 58740 19628
rect 58788 19572 58844 19628
rect 58892 19572 58948 19628
rect 67268 19572 67324 19628
rect 67372 19572 67428 19628
rect 67476 19572 67532 19628
rect 67580 19572 67636 19628
rect 67684 19572 67740 19628
rect 67788 19572 67844 19628
rect 67892 19572 67948 19628
rect 76268 19572 76324 19628
rect 76372 19572 76428 19628
rect 76476 19572 76532 19628
rect 76580 19572 76636 19628
rect 76684 19572 76740 19628
rect 76788 19572 76844 19628
rect 76892 19572 76948 19628
rect 85268 19572 85324 19628
rect 85372 19572 85428 19628
rect 85476 19572 85532 19628
rect 85580 19572 85636 19628
rect 85684 19572 85740 19628
rect 85788 19572 85844 19628
rect 85892 19572 85948 19628
rect 94268 19572 94324 19628
rect 94372 19572 94428 19628
rect 94476 19572 94532 19628
rect 94580 19572 94636 19628
rect 94684 19572 94740 19628
rect 94788 19572 94844 19628
rect 94892 19572 94948 19628
rect 8768 18788 8824 18844
rect 8872 18788 8928 18844
rect 8976 18788 9032 18844
rect 9080 18788 9136 18844
rect 9184 18788 9240 18844
rect 9288 18788 9344 18844
rect 9392 18788 9448 18844
rect 17768 18788 17824 18844
rect 17872 18788 17928 18844
rect 17976 18788 18032 18844
rect 18080 18788 18136 18844
rect 18184 18788 18240 18844
rect 18288 18788 18344 18844
rect 18392 18788 18448 18844
rect 26768 18788 26824 18844
rect 26872 18788 26928 18844
rect 26976 18788 27032 18844
rect 27080 18788 27136 18844
rect 27184 18788 27240 18844
rect 27288 18788 27344 18844
rect 27392 18788 27448 18844
rect 35768 18788 35824 18844
rect 35872 18788 35928 18844
rect 35976 18788 36032 18844
rect 36080 18788 36136 18844
rect 36184 18788 36240 18844
rect 36288 18788 36344 18844
rect 36392 18788 36448 18844
rect 44768 18788 44824 18844
rect 44872 18788 44928 18844
rect 44976 18788 45032 18844
rect 45080 18788 45136 18844
rect 45184 18788 45240 18844
rect 45288 18788 45344 18844
rect 45392 18788 45448 18844
rect 53768 18788 53824 18844
rect 53872 18788 53928 18844
rect 53976 18788 54032 18844
rect 54080 18788 54136 18844
rect 54184 18788 54240 18844
rect 54288 18788 54344 18844
rect 54392 18788 54448 18844
rect 62768 18788 62824 18844
rect 62872 18788 62928 18844
rect 62976 18788 63032 18844
rect 63080 18788 63136 18844
rect 63184 18788 63240 18844
rect 63288 18788 63344 18844
rect 63392 18788 63448 18844
rect 71768 18788 71824 18844
rect 71872 18788 71928 18844
rect 71976 18788 72032 18844
rect 72080 18788 72136 18844
rect 72184 18788 72240 18844
rect 72288 18788 72344 18844
rect 72392 18788 72448 18844
rect 80768 18788 80824 18844
rect 80872 18788 80928 18844
rect 80976 18788 81032 18844
rect 81080 18788 81136 18844
rect 81184 18788 81240 18844
rect 81288 18788 81344 18844
rect 81392 18788 81448 18844
rect 89768 18788 89824 18844
rect 89872 18788 89928 18844
rect 89976 18788 90032 18844
rect 90080 18788 90136 18844
rect 90184 18788 90240 18844
rect 90288 18788 90344 18844
rect 90392 18788 90448 18844
rect 4268 18004 4324 18060
rect 4372 18004 4428 18060
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 4788 18004 4844 18060
rect 4892 18004 4948 18060
rect 13268 18004 13324 18060
rect 13372 18004 13428 18060
rect 13476 18004 13532 18060
rect 13580 18004 13636 18060
rect 13684 18004 13740 18060
rect 13788 18004 13844 18060
rect 13892 18004 13948 18060
rect 22268 18004 22324 18060
rect 22372 18004 22428 18060
rect 22476 18004 22532 18060
rect 22580 18004 22636 18060
rect 22684 18004 22740 18060
rect 22788 18004 22844 18060
rect 22892 18004 22948 18060
rect 31268 18004 31324 18060
rect 31372 18004 31428 18060
rect 31476 18004 31532 18060
rect 31580 18004 31636 18060
rect 31684 18004 31740 18060
rect 31788 18004 31844 18060
rect 31892 18004 31948 18060
rect 40268 18004 40324 18060
rect 40372 18004 40428 18060
rect 40476 18004 40532 18060
rect 40580 18004 40636 18060
rect 40684 18004 40740 18060
rect 40788 18004 40844 18060
rect 40892 18004 40948 18060
rect 49268 18004 49324 18060
rect 49372 18004 49428 18060
rect 49476 18004 49532 18060
rect 49580 18004 49636 18060
rect 49684 18004 49740 18060
rect 49788 18004 49844 18060
rect 49892 18004 49948 18060
rect 58268 18004 58324 18060
rect 58372 18004 58428 18060
rect 58476 18004 58532 18060
rect 58580 18004 58636 18060
rect 58684 18004 58740 18060
rect 58788 18004 58844 18060
rect 58892 18004 58948 18060
rect 67268 18004 67324 18060
rect 67372 18004 67428 18060
rect 67476 18004 67532 18060
rect 67580 18004 67636 18060
rect 67684 18004 67740 18060
rect 67788 18004 67844 18060
rect 67892 18004 67948 18060
rect 76268 18004 76324 18060
rect 76372 18004 76428 18060
rect 76476 18004 76532 18060
rect 76580 18004 76636 18060
rect 76684 18004 76740 18060
rect 76788 18004 76844 18060
rect 76892 18004 76948 18060
rect 85268 18004 85324 18060
rect 85372 18004 85428 18060
rect 85476 18004 85532 18060
rect 85580 18004 85636 18060
rect 85684 18004 85740 18060
rect 85788 18004 85844 18060
rect 85892 18004 85948 18060
rect 94268 18004 94324 18060
rect 94372 18004 94428 18060
rect 94476 18004 94532 18060
rect 94580 18004 94636 18060
rect 94684 18004 94740 18060
rect 94788 18004 94844 18060
rect 94892 18004 94948 18060
rect 8768 17220 8824 17276
rect 8872 17220 8928 17276
rect 8976 17220 9032 17276
rect 9080 17220 9136 17276
rect 9184 17220 9240 17276
rect 9288 17220 9344 17276
rect 9392 17220 9448 17276
rect 17768 17220 17824 17276
rect 17872 17220 17928 17276
rect 17976 17220 18032 17276
rect 18080 17220 18136 17276
rect 18184 17220 18240 17276
rect 18288 17220 18344 17276
rect 18392 17220 18448 17276
rect 26768 17220 26824 17276
rect 26872 17220 26928 17276
rect 26976 17220 27032 17276
rect 27080 17220 27136 17276
rect 27184 17220 27240 17276
rect 27288 17220 27344 17276
rect 27392 17220 27448 17276
rect 35768 17220 35824 17276
rect 35872 17220 35928 17276
rect 35976 17220 36032 17276
rect 36080 17220 36136 17276
rect 36184 17220 36240 17276
rect 36288 17220 36344 17276
rect 36392 17220 36448 17276
rect 44768 17220 44824 17276
rect 44872 17220 44928 17276
rect 44976 17220 45032 17276
rect 45080 17220 45136 17276
rect 45184 17220 45240 17276
rect 45288 17220 45344 17276
rect 45392 17220 45448 17276
rect 53768 17220 53824 17276
rect 53872 17220 53928 17276
rect 53976 17220 54032 17276
rect 54080 17220 54136 17276
rect 54184 17220 54240 17276
rect 54288 17220 54344 17276
rect 54392 17220 54448 17276
rect 62768 17220 62824 17276
rect 62872 17220 62928 17276
rect 62976 17220 63032 17276
rect 63080 17220 63136 17276
rect 63184 17220 63240 17276
rect 63288 17220 63344 17276
rect 63392 17220 63448 17276
rect 71768 17220 71824 17276
rect 71872 17220 71928 17276
rect 71976 17220 72032 17276
rect 72080 17220 72136 17276
rect 72184 17220 72240 17276
rect 72288 17220 72344 17276
rect 72392 17220 72448 17276
rect 80768 17220 80824 17276
rect 80872 17220 80928 17276
rect 80976 17220 81032 17276
rect 81080 17220 81136 17276
rect 81184 17220 81240 17276
rect 81288 17220 81344 17276
rect 81392 17220 81448 17276
rect 89768 17220 89824 17276
rect 89872 17220 89928 17276
rect 89976 17220 90032 17276
rect 90080 17220 90136 17276
rect 90184 17220 90240 17276
rect 90288 17220 90344 17276
rect 90392 17220 90448 17276
rect 4268 16436 4324 16492
rect 4372 16436 4428 16492
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 4788 16436 4844 16492
rect 4892 16436 4948 16492
rect 13268 16436 13324 16492
rect 13372 16436 13428 16492
rect 13476 16436 13532 16492
rect 13580 16436 13636 16492
rect 13684 16436 13740 16492
rect 13788 16436 13844 16492
rect 13892 16436 13948 16492
rect 22268 16436 22324 16492
rect 22372 16436 22428 16492
rect 22476 16436 22532 16492
rect 22580 16436 22636 16492
rect 22684 16436 22740 16492
rect 22788 16436 22844 16492
rect 22892 16436 22948 16492
rect 31268 16436 31324 16492
rect 31372 16436 31428 16492
rect 31476 16436 31532 16492
rect 31580 16436 31636 16492
rect 31684 16436 31740 16492
rect 31788 16436 31844 16492
rect 31892 16436 31948 16492
rect 40268 16436 40324 16492
rect 40372 16436 40428 16492
rect 40476 16436 40532 16492
rect 40580 16436 40636 16492
rect 40684 16436 40740 16492
rect 40788 16436 40844 16492
rect 40892 16436 40948 16492
rect 49268 16436 49324 16492
rect 49372 16436 49428 16492
rect 49476 16436 49532 16492
rect 49580 16436 49636 16492
rect 49684 16436 49740 16492
rect 49788 16436 49844 16492
rect 49892 16436 49948 16492
rect 58268 16436 58324 16492
rect 58372 16436 58428 16492
rect 58476 16436 58532 16492
rect 58580 16436 58636 16492
rect 58684 16436 58740 16492
rect 58788 16436 58844 16492
rect 58892 16436 58948 16492
rect 67268 16436 67324 16492
rect 67372 16436 67428 16492
rect 67476 16436 67532 16492
rect 67580 16436 67636 16492
rect 67684 16436 67740 16492
rect 67788 16436 67844 16492
rect 67892 16436 67948 16492
rect 76268 16436 76324 16492
rect 76372 16436 76428 16492
rect 76476 16436 76532 16492
rect 76580 16436 76636 16492
rect 76684 16436 76740 16492
rect 76788 16436 76844 16492
rect 76892 16436 76948 16492
rect 85268 16436 85324 16492
rect 85372 16436 85428 16492
rect 85476 16436 85532 16492
rect 85580 16436 85636 16492
rect 85684 16436 85740 16492
rect 85788 16436 85844 16492
rect 85892 16436 85948 16492
rect 94268 16436 94324 16492
rect 94372 16436 94428 16492
rect 94476 16436 94532 16492
rect 94580 16436 94636 16492
rect 94684 16436 94740 16492
rect 94788 16436 94844 16492
rect 94892 16436 94948 16492
rect 8768 15652 8824 15708
rect 8872 15652 8928 15708
rect 8976 15652 9032 15708
rect 9080 15652 9136 15708
rect 9184 15652 9240 15708
rect 9288 15652 9344 15708
rect 9392 15652 9448 15708
rect 17768 15652 17824 15708
rect 17872 15652 17928 15708
rect 17976 15652 18032 15708
rect 18080 15652 18136 15708
rect 18184 15652 18240 15708
rect 18288 15652 18344 15708
rect 18392 15652 18448 15708
rect 26768 15652 26824 15708
rect 26872 15652 26928 15708
rect 26976 15652 27032 15708
rect 27080 15652 27136 15708
rect 27184 15652 27240 15708
rect 27288 15652 27344 15708
rect 27392 15652 27448 15708
rect 35768 15652 35824 15708
rect 35872 15652 35928 15708
rect 35976 15652 36032 15708
rect 36080 15652 36136 15708
rect 36184 15652 36240 15708
rect 36288 15652 36344 15708
rect 36392 15652 36448 15708
rect 44768 15652 44824 15708
rect 44872 15652 44928 15708
rect 44976 15652 45032 15708
rect 45080 15652 45136 15708
rect 45184 15652 45240 15708
rect 45288 15652 45344 15708
rect 45392 15652 45448 15708
rect 53768 15652 53824 15708
rect 53872 15652 53928 15708
rect 53976 15652 54032 15708
rect 54080 15652 54136 15708
rect 54184 15652 54240 15708
rect 54288 15652 54344 15708
rect 54392 15652 54448 15708
rect 62768 15652 62824 15708
rect 62872 15652 62928 15708
rect 62976 15652 63032 15708
rect 63080 15652 63136 15708
rect 63184 15652 63240 15708
rect 63288 15652 63344 15708
rect 63392 15652 63448 15708
rect 71768 15652 71824 15708
rect 71872 15652 71928 15708
rect 71976 15652 72032 15708
rect 72080 15652 72136 15708
rect 72184 15652 72240 15708
rect 72288 15652 72344 15708
rect 72392 15652 72448 15708
rect 80768 15652 80824 15708
rect 80872 15652 80928 15708
rect 80976 15652 81032 15708
rect 81080 15652 81136 15708
rect 81184 15652 81240 15708
rect 81288 15652 81344 15708
rect 81392 15652 81448 15708
rect 89768 15652 89824 15708
rect 89872 15652 89928 15708
rect 89976 15652 90032 15708
rect 90080 15652 90136 15708
rect 90184 15652 90240 15708
rect 90288 15652 90344 15708
rect 90392 15652 90448 15708
rect 4268 14868 4324 14924
rect 4372 14868 4428 14924
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 4788 14868 4844 14924
rect 4892 14868 4948 14924
rect 13268 14868 13324 14924
rect 13372 14868 13428 14924
rect 13476 14868 13532 14924
rect 13580 14868 13636 14924
rect 13684 14868 13740 14924
rect 13788 14868 13844 14924
rect 13892 14868 13948 14924
rect 22268 14868 22324 14924
rect 22372 14868 22428 14924
rect 22476 14868 22532 14924
rect 22580 14868 22636 14924
rect 22684 14868 22740 14924
rect 22788 14868 22844 14924
rect 22892 14868 22948 14924
rect 31268 14868 31324 14924
rect 31372 14868 31428 14924
rect 31476 14868 31532 14924
rect 31580 14868 31636 14924
rect 31684 14868 31740 14924
rect 31788 14868 31844 14924
rect 31892 14868 31948 14924
rect 40268 14868 40324 14924
rect 40372 14868 40428 14924
rect 40476 14868 40532 14924
rect 40580 14868 40636 14924
rect 40684 14868 40740 14924
rect 40788 14868 40844 14924
rect 40892 14868 40948 14924
rect 49268 14868 49324 14924
rect 49372 14868 49428 14924
rect 49476 14868 49532 14924
rect 49580 14868 49636 14924
rect 49684 14868 49740 14924
rect 49788 14868 49844 14924
rect 49892 14868 49948 14924
rect 58268 14868 58324 14924
rect 58372 14868 58428 14924
rect 58476 14868 58532 14924
rect 58580 14868 58636 14924
rect 58684 14868 58740 14924
rect 58788 14868 58844 14924
rect 58892 14868 58948 14924
rect 67268 14868 67324 14924
rect 67372 14868 67428 14924
rect 67476 14868 67532 14924
rect 67580 14868 67636 14924
rect 67684 14868 67740 14924
rect 67788 14868 67844 14924
rect 67892 14868 67948 14924
rect 76268 14868 76324 14924
rect 76372 14868 76428 14924
rect 76476 14868 76532 14924
rect 76580 14868 76636 14924
rect 76684 14868 76740 14924
rect 76788 14868 76844 14924
rect 76892 14868 76948 14924
rect 85268 14868 85324 14924
rect 85372 14868 85428 14924
rect 85476 14868 85532 14924
rect 85580 14868 85636 14924
rect 85684 14868 85740 14924
rect 85788 14868 85844 14924
rect 85892 14868 85948 14924
rect 94268 14868 94324 14924
rect 94372 14868 94428 14924
rect 94476 14868 94532 14924
rect 94580 14868 94636 14924
rect 94684 14868 94740 14924
rect 94788 14868 94844 14924
rect 94892 14868 94948 14924
rect 8768 14084 8824 14140
rect 8872 14084 8928 14140
rect 8976 14084 9032 14140
rect 9080 14084 9136 14140
rect 9184 14084 9240 14140
rect 9288 14084 9344 14140
rect 9392 14084 9448 14140
rect 17768 14084 17824 14140
rect 17872 14084 17928 14140
rect 17976 14084 18032 14140
rect 18080 14084 18136 14140
rect 18184 14084 18240 14140
rect 18288 14084 18344 14140
rect 18392 14084 18448 14140
rect 26768 14084 26824 14140
rect 26872 14084 26928 14140
rect 26976 14084 27032 14140
rect 27080 14084 27136 14140
rect 27184 14084 27240 14140
rect 27288 14084 27344 14140
rect 27392 14084 27448 14140
rect 35768 14084 35824 14140
rect 35872 14084 35928 14140
rect 35976 14084 36032 14140
rect 36080 14084 36136 14140
rect 36184 14084 36240 14140
rect 36288 14084 36344 14140
rect 36392 14084 36448 14140
rect 44768 14084 44824 14140
rect 44872 14084 44928 14140
rect 44976 14084 45032 14140
rect 45080 14084 45136 14140
rect 45184 14084 45240 14140
rect 45288 14084 45344 14140
rect 45392 14084 45448 14140
rect 53768 14084 53824 14140
rect 53872 14084 53928 14140
rect 53976 14084 54032 14140
rect 54080 14084 54136 14140
rect 54184 14084 54240 14140
rect 54288 14084 54344 14140
rect 54392 14084 54448 14140
rect 62768 14084 62824 14140
rect 62872 14084 62928 14140
rect 62976 14084 63032 14140
rect 63080 14084 63136 14140
rect 63184 14084 63240 14140
rect 63288 14084 63344 14140
rect 63392 14084 63448 14140
rect 71768 14084 71824 14140
rect 71872 14084 71928 14140
rect 71976 14084 72032 14140
rect 72080 14084 72136 14140
rect 72184 14084 72240 14140
rect 72288 14084 72344 14140
rect 72392 14084 72448 14140
rect 80768 14084 80824 14140
rect 80872 14084 80928 14140
rect 80976 14084 81032 14140
rect 81080 14084 81136 14140
rect 81184 14084 81240 14140
rect 81288 14084 81344 14140
rect 81392 14084 81448 14140
rect 89768 14084 89824 14140
rect 89872 14084 89928 14140
rect 89976 14084 90032 14140
rect 90080 14084 90136 14140
rect 90184 14084 90240 14140
rect 90288 14084 90344 14140
rect 90392 14084 90448 14140
rect 4268 13300 4324 13356
rect 4372 13300 4428 13356
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 4788 13300 4844 13356
rect 4892 13300 4948 13356
rect 13268 13300 13324 13356
rect 13372 13300 13428 13356
rect 13476 13300 13532 13356
rect 13580 13300 13636 13356
rect 13684 13300 13740 13356
rect 13788 13300 13844 13356
rect 13892 13300 13948 13356
rect 22268 13300 22324 13356
rect 22372 13300 22428 13356
rect 22476 13300 22532 13356
rect 22580 13300 22636 13356
rect 22684 13300 22740 13356
rect 22788 13300 22844 13356
rect 22892 13300 22948 13356
rect 31268 13300 31324 13356
rect 31372 13300 31428 13356
rect 31476 13300 31532 13356
rect 31580 13300 31636 13356
rect 31684 13300 31740 13356
rect 31788 13300 31844 13356
rect 31892 13300 31948 13356
rect 40268 13300 40324 13356
rect 40372 13300 40428 13356
rect 40476 13300 40532 13356
rect 40580 13300 40636 13356
rect 40684 13300 40740 13356
rect 40788 13300 40844 13356
rect 40892 13300 40948 13356
rect 49268 13300 49324 13356
rect 49372 13300 49428 13356
rect 49476 13300 49532 13356
rect 49580 13300 49636 13356
rect 49684 13300 49740 13356
rect 49788 13300 49844 13356
rect 49892 13300 49948 13356
rect 58268 13300 58324 13356
rect 58372 13300 58428 13356
rect 58476 13300 58532 13356
rect 58580 13300 58636 13356
rect 58684 13300 58740 13356
rect 58788 13300 58844 13356
rect 58892 13300 58948 13356
rect 67268 13300 67324 13356
rect 67372 13300 67428 13356
rect 67476 13300 67532 13356
rect 67580 13300 67636 13356
rect 67684 13300 67740 13356
rect 67788 13300 67844 13356
rect 67892 13300 67948 13356
rect 76268 13300 76324 13356
rect 76372 13300 76428 13356
rect 76476 13300 76532 13356
rect 76580 13300 76636 13356
rect 76684 13300 76740 13356
rect 76788 13300 76844 13356
rect 76892 13300 76948 13356
rect 85268 13300 85324 13356
rect 85372 13300 85428 13356
rect 85476 13300 85532 13356
rect 85580 13300 85636 13356
rect 85684 13300 85740 13356
rect 85788 13300 85844 13356
rect 85892 13300 85948 13356
rect 94268 13300 94324 13356
rect 94372 13300 94428 13356
rect 94476 13300 94532 13356
rect 94580 13300 94636 13356
rect 94684 13300 94740 13356
rect 94788 13300 94844 13356
rect 94892 13300 94948 13356
rect 8768 12516 8824 12572
rect 8872 12516 8928 12572
rect 8976 12516 9032 12572
rect 9080 12516 9136 12572
rect 9184 12516 9240 12572
rect 9288 12516 9344 12572
rect 9392 12516 9448 12572
rect 17768 12516 17824 12572
rect 17872 12516 17928 12572
rect 17976 12516 18032 12572
rect 18080 12516 18136 12572
rect 18184 12516 18240 12572
rect 18288 12516 18344 12572
rect 18392 12516 18448 12572
rect 26768 12516 26824 12572
rect 26872 12516 26928 12572
rect 26976 12516 27032 12572
rect 27080 12516 27136 12572
rect 27184 12516 27240 12572
rect 27288 12516 27344 12572
rect 27392 12516 27448 12572
rect 35768 12516 35824 12572
rect 35872 12516 35928 12572
rect 35976 12516 36032 12572
rect 36080 12516 36136 12572
rect 36184 12516 36240 12572
rect 36288 12516 36344 12572
rect 36392 12516 36448 12572
rect 44768 12516 44824 12572
rect 44872 12516 44928 12572
rect 44976 12516 45032 12572
rect 45080 12516 45136 12572
rect 45184 12516 45240 12572
rect 45288 12516 45344 12572
rect 45392 12516 45448 12572
rect 53768 12516 53824 12572
rect 53872 12516 53928 12572
rect 53976 12516 54032 12572
rect 54080 12516 54136 12572
rect 54184 12516 54240 12572
rect 54288 12516 54344 12572
rect 54392 12516 54448 12572
rect 62768 12516 62824 12572
rect 62872 12516 62928 12572
rect 62976 12516 63032 12572
rect 63080 12516 63136 12572
rect 63184 12516 63240 12572
rect 63288 12516 63344 12572
rect 63392 12516 63448 12572
rect 71768 12516 71824 12572
rect 71872 12516 71928 12572
rect 71976 12516 72032 12572
rect 72080 12516 72136 12572
rect 72184 12516 72240 12572
rect 72288 12516 72344 12572
rect 72392 12516 72448 12572
rect 80768 12516 80824 12572
rect 80872 12516 80928 12572
rect 80976 12516 81032 12572
rect 81080 12516 81136 12572
rect 81184 12516 81240 12572
rect 81288 12516 81344 12572
rect 81392 12516 81448 12572
rect 89768 12516 89824 12572
rect 89872 12516 89928 12572
rect 89976 12516 90032 12572
rect 90080 12516 90136 12572
rect 90184 12516 90240 12572
rect 90288 12516 90344 12572
rect 90392 12516 90448 12572
rect 4268 11732 4324 11788
rect 4372 11732 4428 11788
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 4788 11732 4844 11788
rect 4892 11732 4948 11788
rect 13268 11732 13324 11788
rect 13372 11732 13428 11788
rect 13476 11732 13532 11788
rect 13580 11732 13636 11788
rect 13684 11732 13740 11788
rect 13788 11732 13844 11788
rect 13892 11732 13948 11788
rect 22268 11732 22324 11788
rect 22372 11732 22428 11788
rect 22476 11732 22532 11788
rect 22580 11732 22636 11788
rect 22684 11732 22740 11788
rect 22788 11732 22844 11788
rect 22892 11732 22948 11788
rect 31268 11732 31324 11788
rect 31372 11732 31428 11788
rect 31476 11732 31532 11788
rect 31580 11732 31636 11788
rect 31684 11732 31740 11788
rect 31788 11732 31844 11788
rect 31892 11732 31948 11788
rect 40268 11732 40324 11788
rect 40372 11732 40428 11788
rect 40476 11732 40532 11788
rect 40580 11732 40636 11788
rect 40684 11732 40740 11788
rect 40788 11732 40844 11788
rect 40892 11732 40948 11788
rect 49268 11732 49324 11788
rect 49372 11732 49428 11788
rect 49476 11732 49532 11788
rect 49580 11732 49636 11788
rect 49684 11732 49740 11788
rect 49788 11732 49844 11788
rect 49892 11732 49948 11788
rect 58268 11732 58324 11788
rect 58372 11732 58428 11788
rect 58476 11732 58532 11788
rect 58580 11732 58636 11788
rect 58684 11732 58740 11788
rect 58788 11732 58844 11788
rect 58892 11732 58948 11788
rect 67268 11732 67324 11788
rect 67372 11732 67428 11788
rect 67476 11732 67532 11788
rect 67580 11732 67636 11788
rect 67684 11732 67740 11788
rect 67788 11732 67844 11788
rect 67892 11732 67948 11788
rect 76268 11732 76324 11788
rect 76372 11732 76428 11788
rect 76476 11732 76532 11788
rect 76580 11732 76636 11788
rect 76684 11732 76740 11788
rect 76788 11732 76844 11788
rect 76892 11732 76948 11788
rect 85268 11732 85324 11788
rect 85372 11732 85428 11788
rect 85476 11732 85532 11788
rect 85580 11732 85636 11788
rect 85684 11732 85740 11788
rect 85788 11732 85844 11788
rect 85892 11732 85948 11788
rect 94268 11732 94324 11788
rect 94372 11732 94428 11788
rect 94476 11732 94532 11788
rect 94580 11732 94636 11788
rect 94684 11732 94740 11788
rect 94788 11732 94844 11788
rect 94892 11732 94948 11788
rect 8768 10948 8824 11004
rect 8872 10948 8928 11004
rect 8976 10948 9032 11004
rect 9080 10948 9136 11004
rect 9184 10948 9240 11004
rect 9288 10948 9344 11004
rect 9392 10948 9448 11004
rect 17768 10948 17824 11004
rect 17872 10948 17928 11004
rect 17976 10948 18032 11004
rect 18080 10948 18136 11004
rect 18184 10948 18240 11004
rect 18288 10948 18344 11004
rect 18392 10948 18448 11004
rect 26768 10948 26824 11004
rect 26872 10948 26928 11004
rect 26976 10948 27032 11004
rect 27080 10948 27136 11004
rect 27184 10948 27240 11004
rect 27288 10948 27344 11004
rect 27392 10948 27448 11004
rect 35768 10948 35824 11004
rect 35872 10948 35928 11004
rect 35976 10948 36032 11004
rect 36080 10948 36136 11004
rect 36184 10948 36240 11004
rect 36288 10948 36344 11004
rect 36392 10948 36448 11004
rect 44768 10948 44824 11004
rect 44872 10948 44928 11004
rect 44976 10948 45032 11004
rect 45080 10948 45136 11004
rect 45184 10948 45240 11004
rect 45288 10948 45344 11004
rect 45392 10948 45448 11004
rect 53768 10948 53824 11004
rect 53872 10948 53928 11004
rect 53976 10948 54032 11004
rect 54080 10948 54136 11004
rect 54184 10948 54240 11004
rect 54288 10948 54344 11004
rect 54392 10948 54448 11004
rect 62768 10948 62824 11004
rect 62872 10948 62928 11004
rect 62976 10948 63032 11004
rect 63080 10948 63136 11004
rect 63184 10948 63240 11004
rect 63288 10948 63344 11004
rect 63392 10948 63448 11004
rect 71768 10948 71824 11004
rect 71872 10948 71928 11004
rect 71976 10948 72032 11004
rect 72080 10948 72136 11004
rect 72184 10948 72240 11004
rect 72288 10948 72344 11004
rect 72392 10948 72448 11004
rect 80768 10948 80824 11004
rect 80872 10948 80928 11004
rect 80976 10948 81032 11004
rect 81080 10948 81136 11004
rect 81184 10948 81240 11004
rect 81288 10948 81344 11004
rect 81392 10948 81448 11004
rect 89768 10948 89824 11004
rect 89872 10948 89928 11004
rect 89976 10948 90032 11004
rect 90080 10948 90136 11004
rect 90184 10948 90240 11004
rect 90288 10948 90344 11004
rect 90392 10948 90448 11004
rect 4268 10164 4324 10220
rect 4372 10164 4428 10220
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 4788 10164 4844 10220
rect 4892 10164 4948 10220
rect 13268 10164 13324 10220
rect 13372 10164 13428 10220
rect 13476 10164 13532 10220
rect 13580 10164 13636 10220
rect 13684 10164 13740 10220
rect 13788 10164 13844 10220
rect 13892 10164 13948 10220
rect 22268 10164 22324 10220
rect 22372 10164 22428 10220
rect 22476 10164 22532 10220
rect 22580 10164 22636 10220
rect 22684 10164 22740 10220
rect 22788 10164 22844 10220
rect 22892 10164 22948 10220
rect 31268 10164 31324 10220
rect 31372 10164 31428 10220
rect 31476 10164 31532 10220
rect 31580 10164 31636 10220
rect 31684 10164 31740 10220
rect 31788 10164 31844 10220
rect 31892 10164 31948 10220
rect 40268 10164 40324 10220
rect 40372 10164 40428 10220
rect 40476 10164 40532 10220
rect 40580 10164 40636 10220
rect 40684 10164 40740 10220
rect 40788 10164 40844 10220
rect 40892 10164 40948 10220
rect 49268 10164 49324 10220
rect 49372 10164 49428 10220
rect 49476 10164 49532 10220
rect 49580 10164 49636 10220
rect 49684 10164 49740 10220
rect 49788 10164 49844 10220
rect 49892 10164 49948 10220
rect 58268 10164 58324 10220
rect 58372 10164 58428 10220
rect 58476 10164 58532 10220
rect 58580 10164 58636 10220
rect 58684 10164 58740 10220
rect 58788 10164 58844 10220
rect 58892 10164 58948 10220
rect 67268 10164 67324 10220
rect 67372 10164 67428 10220
rect 67476 10164 67532 10220
rect 67580 10164 67636 10220
rect 67684 10164 67740 10220
rect 67788 10164 67844 10220
rect 67892 10164 67948 10220
rect 76268 10164 76324 10220
rect 76372 10164 76428 10220
rect 76476 10164 76532 10220
rect 76580 10164 76636 10220
rect 76684 10164 76740 10220
rect 76788 10164 76844 10220
rect 76892 10164 76948 10220
rect 85268 10164 85324 10220
rect 85372 10164 85428 10220
rect 85476 10164 85532 10220
rect 85580 10164 85636 10220
rect 85684 10164 85740 10220
rect 85788 10164 85844 10220
rect 85892 10164 85948 10220
rect 94268 10164 94324 10220
rect 94372 10164 94428 10220
rect 94476 10164 94532 10220
rect 94580 10164 94636 10220
rect 94684 10164 94740 10220
rect 94788 10164 94844 10220
rect 94892 10164 94948 10220
rect 8768 9380 8824 9436
rect 8872 9380 8928 9436
rect 8976 9380 9032 9436
rect 9080 9380 9136 9436
rect 9184 9380 9240 9436
rect 9288 9380 9344 9436
rect 9392 9380 9448 9436
rect 17768 9380 17824 9436
rect 17872 9380 17928 9436
rect 17976 9380 18032 9436
rect 18080 9380 18136 9436
rect 18184 9380 18240 9436
rect 18288 9380 18344 9436
rect 18392 9380 18448 9436
rect 26768 9380 26824 9436
rect 26872 9380 26928 9436
rect 26976 9380 27032 9436
rect 27080 9380 27136 9436
rect 27184 9380 27240 9436
rect 27288 9380 27344 9436
rect 27392 9380 27448 9436
rect 35768 9380 35824 9436
rect 35872 9380 35928 9436
rect 35976 9380 36032 9436
rect 36080 9380 36136 9436
rect 36184 9380 36240 9436
rect 36288 9380 36344 9436
rect 36392 9380 36448 9436
rect 44768 9380 44824 9436
rect 44872 9380 44928 9436
rect 44976 9380 45032 9436
rect 45080 9380 45136 9436
rect 45184 9380 45240 9436
rect 45288 9380 45344 9436
rect 45392 9380 45448 9436
rect 53768 9380 53824 9436
rect 53872 9380 53928 9436
rect 53976 9380 54032 9436
rect 54080 9380 54136 9436
rect 54184 9380 54240 9436
rect 54288 9380 54344 9436
rect 54392 9380 54448 9436
rect 62768 9380 62824 9436
rect 62872 9380 62928 9436
rect 62976 9380 63032 9436
rect 63080 9380 63136 9436
rect 63184 9380 63240 9436
rect 63288 9380 63344 9436
rect 63392 9380 63448 9436
rect 71768 9380 71824 9436
rect 71872 9380 71928 9436
rect 71976 9380 72032 9436
rect 72080 9380 72136 9436
rect 72184 9380 72240 9436
rect 72288 9380 72344 9436
rect 72392 9380 72448 9436
rect 80768 9380 80824 9436
rect 80872 9380 80928 9436
rect 80976 9380 81032 9436
rect 81080 9380 81136 9436
rect 81184 9380 81240 9436
rect 81288 9380 81344 9436
rect 81392 9380 81448 9436
rect 89768 9380 89824 9436
rect 89872 9380 89928 9436
rect 89976 9380 90032 9436
rect 90080 9380 90136 9436
rect 90184 9380 90240 9436
rect 90288 9380 90344 9436
rect 90392 9380 90448 9436
rect 4268 8596 4324 8652
rect 4372 8596 4428 8652
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 4788 8596 4844 8652
rect 4892 8596 4948 8652
rect 13268 8596 13324 8652
rect 13372 8596 13428 8652
rect 13476 8596 13532 8652
rect 13580 8596 13636 8652
rect 13684 8596 13740 8652
rect 13788 8596 13844 8652
rect 13892 8596 13948 8652
rect 22268 8596 22324 8652
rect 22372 8596 22428 8652
rect 22476 8596 22532 8652
rect 22580 8596 22636 8652
rect 22684 8596 22740 8652
rect 22788 8596 22844 8652
rect 22892 8596 22948 8652
rect 31268 8596 31324 8652
rect 31372 8596 31428 8652
rect 31476 8596 31532 8652
rect 31580 8596 31636 8652
rect 31684 8596 31740 8652
rect 31788 8596 31844 8652
rect 31892 8596 31948 8652
rect 40268 8596 40324 8652
rect 40372 8596 40428 8652
rect 40476 8596 40532 8652
rect 40580 8596 40636 8652
rect 40684 8596 40740 8652
rect 40788 8596 40844 8652
rect 40892 8596 40948 8652
rect 49268 8596 49324 8652
rect 49372 8596 49428 8652
rect 49476 8596 49532 8652
rect 49580 8596 49636 8652
rect 49684 8596 49740 8652
rect 49788 8596 49844 8652
rect 49892 8596 49948 8652
rect 58268 8596 58324 8652
rect 58372 8596 58428 8652
rect 58476 8596 58532 8652
rect 58580 8596 58636 8652
rect 58684 8596 58740 8652
rect 58788 8596 58844 8652
rect 58892 8596 58948 8652
rect 67268 8596 67324 8652
rect 67372 8596 67428 8652
rect 67476 8596 67532 8652
rect 67580 8596 67636 8652
rect 67684 8596 67740 8652
rect 67788 8596 67844 8652
rect 67892 8596 67948 8652
rect 76268 8596 76324 8652
rect 76372 8596 76428 8652
rect 76476 8596 76532 8652
rect 76580 8596 76636 8652
rect 76684 8596 76740 8652
rect 76788 8596 76844 8652
rect 76892 8596 76948 8652
rect 85268 8596 85324 8652
rect 85372 8596 85428 8652
rect 85476 8596 85532 8652
rect 85580 8596 85636 8652
rect 85684 8596 85740 8652
rect 85788 8596 85844 8652
rect 85892 8596 85948 8652
rect 94268 8596 94324 8652
rect 94372 8596 94428 8652
rect 94476 8596 94532 8652
rect 94580 8596 94636 8652
rect 94684 8596 94740 8652
rect 94788 8596 94844 8652
rect 94892 8596 94948 8652
rect 8768 7812 8824 7868
rect 8872 7812 8928 7868
rect 8976 7812 9032 7868
rect 9080 7812 9136 7868
rect 9184 7812 9240 7868
rect 9288 7812 9344 7868
rect 9392 7812 9448 7868
rect 17768 7812 17824 7868
rect 17872 7812 17928 7868
rect 17976 7812 18032 7868
rect 18080 7812 18136 7868
rect 18184 7812 18240 7868
rect 18288 7812 18344 7868
rect 18392 7812 18448 7868
rect 26768 7812 26824 7868
rect 26872 7812 26928 7868
rect 26976 7812 27032 7868
rect 27080 7812 27136 7868
rect 27184 7812 27240 7868
rect 27288 7812 27344 7868
rect 27392 7812 27448 7868
rect 35768 7812 35824 7868
rect 35872 7812 35928 7868
rect 35976 7812 36032 7868
rect 36080 7812 36136 7868
rect 36184 7812 36240 7868
rect 36288 7812 36344 7868
rect 36392 7812 36448 7868
rect 44768 7812 44824 7868
rect 44872 7812 44928 7868
rect 44976 7812 45032 7868
rect 45080 7812 45136 7868
rect 45184 7812 45240 7868
rect 45288 7812 45344 7868
rect 45392 7812 45448 7868
rect 53768 7812 53824 7868
rect 53872 7812 53928 7868
rect 53976 7812 54032 7868
rect 54080 7812 54136 7868
rect 54184 7812 54240 7868
rect 54288 7812 54344 7868
rect 54392 7812 54448 7868
rect 62768 7812 62824 7868
rect 62872 7812 62928 7868
rect 62976 7812 63032 7868
rect 63080 7812 63136 7868
rect 63184 7812 63240 7868
rect 63288 7812 63344 7868
rect 63392 7812 63448 7868
rect 71768 7812 71824 7868
rect 71872 7812 71928 7868
rect 71976 7812 72032 7868
rect 72080 7812 72136 7868
rect 72184 7812 72240 7868
rect 72288 7812 72344 7868
rect 72392 7812 72448 7868
rect 80768 7812 80824 7868
rect 80872 7812 80928 7868
rect 80976 7812 81032 7868
rect 81080 7812 81136 7868
rect 81184 7812 81240 7868
rect 81288 7812 81344 7868
rect 81392 7812 81448 7868
rect 89768 7812 89824 7868
rect 89872 7812 89928 7868
rect 89976 7812 90032 7868
rect 90080 7812 90136 7868
rect 90184 7812 90240 7868
rect 90288 7812 90344 7868
rect 90392 7812 90448 7868
rect 48860 7644 48916 7700
rect 4268 7028 4324 7084
rect 4372 7028 4428 7084
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 4788 7028 4844 7084
rect 4892 7028 4948 7084
rect 13268 7028 13324 7084
rect 13372 7028 13428 7084
rect 13476 7028 13532 7084
rect 13580 7028 13636 7084
rect 13684 7028 13740 7084
rect 13788 7028 13844 7084
rect 13892 7028 13948 7084
rect 22268 7028 22324 7084
rect 22372 7028 22428 7084
rect 22476 7028 22532 7084
rect 22580 7028 22636 7084
rect 22684 7028 22740 7084
rect 22788 7028 22844 7084
rect 22892 7028 22948 7084
rect 31268 7028 31324 7084
rect 31372 7028 31428 7084
rect 31476 7028 31532 7084
rect 31580 7028 31636 7084
rect 31684 7028 31740 7084
rect 31788 7028 31844 7084
rect 31892 7028 31948 7084
rect 40268 7028 40324 7084
rect 40372 7028 40428 7084
rect 40476 7028 40532 7084
rect 40580 7028 40636 7084
rect 40684 7028 40740 7084
rect 40788 7028 40844 7084
rect 40892 7028 40948 7084
rect 49268 7028 49324 7084
rect 49372 7028 49428 7084
rect 49476 7028 49532 7084
rect 49580 7028 49636 7084
rect 49684 7028 49740 7084
rect 49788 7028 49844 7084
rect 49892 7028 49948 7084
rect 58268 7028 58324 7084
rect 58372 7028 58428 7084
rect 58476 7028 58532 7084
rect 58580 7028 58636 7084
rect 58684 7028 58740 7084
rect 58788 7028 58844 7084
rect 58892 7028 58948 7084
rect 67268 7028 67324 7084
rect 67372 7028 67428 7084
rect 67476 7028 67532 7084
rect 67580 7028 67636 7084
rect 67684 7028 67740 7084
rect 67788 7028 67844 7084
rect 67892 7028 67948 7084
rect 76268 7028 76324 7084
rect 76372 7028 76428 7084
rect 76476 7028 76532 7084
rect 76580 7028 76636 7084
rect 76684 7028 76740 7084
rect 76788 7028 76844 7084
rect 76892 7028 76948 7084
rect 85268 7028 85324 7084
rect 85372 7028 85428 7084
rect 85476 7028 85532 7084
rect 85580 7028 85636 7084
rect 85684 7028 85740 7084
rect 85788 7028 85844 7084
rect 85892 7028 85948 7084
rect 94268 7028 94324 7084
rect 94372 7028 94428 7084
rect 94476 7028 94532 7084
rect 94580 7028 94636 7084
rect 94684 7028 94740 7084
rect 94788 7028 94844 7084
rect 94892 7028 94948 7084
rect 8768 6244 8824 6300
rect 8872 6244 8928 6300
rect 8976 6244 9032 6300
rect 9080 6244 9136 6300
rect 9184 6244 9240 6300
rect 9288 6244 9344 6300
rect 9392 6244 9448 6300
rect 17768 6244 17824 6300
rect 17872 6244 17928 6300
rect 17976 6244 18032 6300
rect 18080 6244 18136 6300
rect 18184 6244 18240 6300
rect 18288 6244 18344 6300
rect 18392 6244 18448 6300
rect 26768 6244 26824 6300
rect 26872 6244 26928 6300
rect 26976 6244 27032 6300
rect 27080 6244 27136 6300
rect 27184 6244 27240 6300
rect 27288 6244 27344 6300
rect 27392 6244 27448 6300
rect 35768 6244 35824 6300
rect 35872 6244 35928 6300
rect 35976 6244 36032 6300
rect 36080 6244 36136 6300
rect 36184 6244 36240 6300
rect 36288 6244 36344 6300
rect 36392 6244 36448 6300
rect 44768 6244 44824 6300
rect 44872 6244 44928 6300
rect 44976 6244 45032 6300
rect 45080 6244 45136 6300
rect 45184 6244 45240 6300
rect 45288 6244 45344 6300
rect 45392 6244 45448 6300
rect 53768 6244 53824 6300
rect 53872 6244 53928 6300
rect 53976 6244 54032 6300
rect 54080 6244 54136 6300
rect 54184 6244 54240 6300
rect 54288 6244 54344 6300
rect 54392 6244 54448 6300
rect 62768 6244 62824 6300
rect 62872 6244 62928 6300
rect 62976 6244 63032 6300
rect 63080 6244 63136 6300
rect 63184 6244 63240 6300
rect 63288 6244 63344 6300
rect 63392 6244 63448 6300
rect 71768 6244 71824 6300
rect 71872 6244 71928 6300
rect 71976 6244 72032 6300
rect 72080 6244 72136 6300
rect 72184 6244 72240 6300
rect 72288 6244 72344 6300
rect 72392 6244 72448 6300
rect 80768 6244 80824 6300
rect 80872 6244 80928 6300
rect 80976 6244 81032 6300
rect 81080 6244 81136 6300
rect 81184 6244 81240 6300
rect 81288 6244 81344 6300
rect 81392 6244 81448 6300
rect 89768 6244 89824 6300
rect 89872 6244 89928 6300
rect 89976 6244 90032 6300
rect 90080 6244 90136 6300
rect 90184 6244 90240 6300
rect 90288 6244 90344 6300
rect 90392 6244 90448 6300
rect 48860 6076 48916 6132
rect 4268 5460 4324 5516
rect 4372 5460 4428 5516
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 4788 5460 4844 5516
rect 4892 5460 4948 5516
rect 13268 5460 13324 5516
rect 13372 5460 13428 5516
rect 13476 5460 13532 5516
rect 13580 5460 13636 5516
rect 13684 5460 13740 5516
rect 13788 5460 13844 5516
rect 13892 5460 13948 5516
rect 22268 5460 22324 5516
rect 22372 5460 22428 5516
rect 22476 5460 22532 5516
rect 22580 5460 22636 5516
rect 22684 5460 22740 5516
rect 22788 5460 22844 5516
rect 22892 5460 22948 5516
rect 31268 5460 31324 5516
rect 31372 5460 31428 5516
rect 31476 5460 31532 5516
rect 31580 5460 31636 5516
rect 31684 5460 31740 5516
rect 31788 5460 31844 5516
rect 31892 5460 31948 5516
rect 40268 5460 40324 5516
rect 40372 5460 40428 5516
rect 40476 5460 40532 5516
rect 40580 5460 40636 5516
rect 40684 5460 40740 5516
rect 40788 5460 40844 5516
rect 40892 5460 40948 5516
rect 49268 5460 49324 5516
rect 49372 5460 49428 5516
rect 49476 5460 49532 5516
rect 49580 5460 49636 5516
rect 49684 5460 49740 5516
rect 49788 5460 49844 5516
rect 49892 5460 49948 5516
rect 58268 5460 58324 5516
rect 58372 5460 58428 5516
rect 58476 5460 58532 5516
rect 58580 5460 58636 5516
rect 58684 5460 58740 5516
rect 58788 5460 58844 5516
rect 58892 5460 58948 5516
rect 67268 5460 67324 5516
rect 67372 5460 67428 5516
rect 67476 5460 67532 5516
rect 67580 5460 67636 5516
rect 67684 5460 67740 5516
rect 67788 5460 67844 5516
rect 67892 5460 67948 5516
rect 76268 5460 76324 5516
rect 76372 5460 76428 5516
rect 76476 5460 76532 5516
rect 76580 5460 76636 5516
rect 76684 5460 76740 5516
rect 76788 5460 76844 5516
rect 76892 5460 76948 5516
rect 85268 5460 85324 5516
rect 85372 5460 85428 5516
rect 85476 5460 85532 5516
rect 85580 5460 85636 5516
rect 85684 5460 85740 5516
rect 85788 5460 85844 5516
rect 85892 5460 85948 5516
rect 94268 5460 94324 5516
rect 94372 5460 94428 5516
rect 94476 5460 94532 5516
rect 94580 5460 94636 5516
rect 94684 5460 94740 5516
rect 94788 5460 94844 5516
rect 94892 5460 94948 5516
rect 59612 4956 59668 5012
rect 8768 4676 8824 4732
rect 8872 4676 8928 4732
rect 8976 4676 9032 4732
rect 9080 4676 9136 4732
rect 9184 4676 9240 4732
rect 9288 4676 9344 4732
rect 9392 4676 9448 4732
rect 17768 4676 17824 4732
rect 17872 4676 17928 4732
rect 17976 4676 18032 4732
rect 18080 4676 18136 4732
rect 18184 4676 18240 4732
rect 18288 4676 18344 4732
rect 18392 4676 18448 4732
rect 26768 4676 26824 4732
rect 26872 4676 26928 4732
rect 26976 4676 27032 4732
rect 27080 4676 27136 4732
rect 27184 4676 27240 4732
rect 27288 4676 27344 4732
rect 27392 4676 27448 4732
rect 35768 4676 35824 4732
rect 35872 4676 35928 4732
rect 35976 4676 36032 4732
rect 36080 4676 36136 4732
rect 36184 4676 36240 4732
rect 36288 4676 36344 4732
rect 36392 4676 36448 4732
rect 44768 4676 44824 4732
rect 44872 4676 44928 4732
rect 44976 4676 45032 4732
rect 45080 4676 45136 4732
rect 45184 4676 45240 4732
rect 45288 4676 45344 4732
rect 45392 4676 45448 4732
rect 53768 4676 53824 4732
rect 53872 4676 53928 4732
rect 53976 4676 54032 4732
rect 54080 4676 54136 4732
rect 54184 4676 54240 4732
rect 54288 4676 54344 4732
rect 54392 4676 54448 4732
rect 62768 4676 62824 4732
rect 62872 4676 62928 4732
rect 62976 4676 63032 4732
rect 63080 4676 63136 4732
rect 63184 4676 63240 4732
rect 63288 4676 63344 4732
rect 63392 4676 63448 4732
rect 71768 4676 71824 4732
rect 71872 4676 71928 4732
rect 71976 4676 72032 4732
rect 72080 4676 72136 4732
rect 72184 4676 72240 4732
rect 72288 4676 72344 4732
rect 72392 4676 72448 4732
rect 80768 4676 80824 4732
rect 80872 4676 80928 4732
rect 80976 4676 81032 4732
rect 81080 4676 81136 4732
rect 81184 4676 81240 4732
rect 81288 4676 81344 4732
rect 81392 4676 81448 4732
rect 89768 4676 89824 4732
rect 89872 4676 89928 4732
rect 89976 4676 90032 4732
rect 90080 4676 90136 4732
rect 90184 4676 90240 4732
rect 90288 4676 90344 4732
rect 90392 4676 90448 4732
rect 75628 4396 75684 4452
rect 4268 3892 4324 3948
rect 4372 3892 4428 3948
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 4788 3892 4844 3948
rect 4892 3892 4948 3948
rect 13268 3892 13324 3948
rect 13372 3892 13428 3948
rect 13476 3892 13532 3948
rect 13580 3892 13636 3948
rect 13684 3892 13740 3948
rect 13788 3892 13844 3948
rect 13892 3892 13948 3948
rect 22268 3892 22324 3948
rect 22372 3892 22428 3948
rect 22476 3892 22532 3948
rect 22580 3892 22636 3948
rect 22684 3892 22740 3948
rect 22788 3892 22844 3948
rect 22892 3892 22948 3948
rect 31268 3892 31324 3948
rect 31372 3892 31428 3948
rect 31476 3892 31532 3948
rect 31580 3892 31636 3948
rect 31684 3892 31740 3948
rect 31788 3892 31844 3948
rect 31892 3892 31948 3948
rect 40268 3892 40324 3948
rect 40372 3892 40428 3948
rect 40476 3892 40532 3948
rect 40580 3892 40636 3948
rect 40684 3892 40740 3948
rect 40788 3892 40844 3948
rect 40892 3892 40948 3948
rect 49268 3892 49324 3948
rect 49372 3892 49428 3948
rect 49476 3892 49532 3948
rect 49580 3892 49636 3948
rect 49684 3892 49740 3948
rect 49788 3892 49844 3948
rect 49892 3892 49948 3948
rect 58268 3892 58324 3948
rect 58372 3892 58428 3948
rect 58476 3892 58532 3948
rect 58580 3892 58636 3948
rect 58684 3892 58740 3948
rect 58788 3892 58844 3948
rect 58892 3892 58948 3948
rect 67268 3892 67324 3948
rect 67372 3892 67428 3948
rect 67476 3892 67532 3948
rect 67580 3892 67636 3948
rect 67684 3892 67740 3948
rect 67788 3892 67844 3948
rect 67892 3892 67948 3948
rect 76268 3892 76324 3948
rect 76372 3892 76428 3948
rect 76476 3892 76532 3948
rect 76580 3892 76636 3948
rect 76684 3892 76740 3948
rect 76788 3892 76844 3948
rect 76892 3892 76948 3948
rect 85268 3892 85324 3948
rect 85372 3892 85428 3948
rect 85476 3892 85532 3948
rect 85580 3892 85636 3948
rect 85684 3892 85740 3948
rect 85788 3892 85844 3948
rect 85892 3892 85948 3948
rect 94268 3892 94324 3948
rect 94372 3892 94428 3948
rect 94476 3892 94532 3948
rect 94580 3892 94636 3948
rect 94684 3892 94740 3948
rect 94788 3892 94844 3948
rect 94892 3892 94948 3948
rect 8768 3108 8824 3164
rect 8872 3108 8928 3164
rect 8976 3108 9032 3164
rect 9080 3108 9136 3164
rect 9184 3108 9240 3164
rect 9288 3108 9344 3164
rect 9392 3108 9448 3164
rect 17768 3108 17824 3164
rect 17872 3108 17928 3164
rect 17976 3108 18032 3164
rect 18080 3108 18136 3164
rect 18184 3108 18240 3164
rect 18288 3108 18344 3164
rect 18392 3108 18448 3164
rect 26768 3108 26824 3164
rect 26872 3108 26928 3164
rect 26976 3108 27032 3164
rect 27080 3108 27136 3164
rect 27184 3108 27240 3164
rect 27288 3108 27344 3164
rect 27392 3108 27448 3164
rect 35768 3108 35824 3164
rect 35872 3108 35928 3164
rect 35976 3108 36032 3164
rect 36080 3108 36136 3164
rect 36184 3108 36240 3164
rect 36288 3108 36344 3164
rect 36392 3108 36448 3164
rect 44768 3108 44824 3164
rect 44872 3108 44928 3164
rect 44976 3108 45032 3164
rect 45080 3108 45136 3164
rect 45184 3108 45240 3164
rect 45288 3108 45344 3164
rect 45392 3108 45448 3164
rect 53768 3108 53824 3164
rect 53872 3108 53928 3164
rect 53976 3108 54032 3164
rect 54080 3108 54136 3164
rect 54184 3108 54240 3164
rect 54288 3108 54344 3164
rect 54392 3108 54448 3164
rect 62768 3108 62824 3164
rect 62872 3108 62928 3164
rect 62976 3108 63032 3164
rect 63080 3108 63136 3164
rect 63184 3108 63240 3164
rect 63288 3108 63344 3164
rect 63392 3108 63448 3164
rect 71768 3108 71824 3164
rect 71872 3108 71928 3164
rect 71976 3108 72032 3164
rect 72080 3108 72136 3164
rect 72184 3108 72240 3164
rect 72288 3108 72344 3164
rect 72392 3108 72448 3164
rect 80768 3108 80824 3164
rect 80872 3108 80928 3164
rect 80976 3108 81032 3164
rect 81080 3108 81136 3164
rect 81184 3108 81240 3164
rect 81288 3108 81344 3164
rect 81392 3108 81448 3164
rect 89768 3108 89824 3164
rect 89872 3108 89928 3164
rect 89976 3108 90032 3164
rect 90080 3108 90136 3164
rect 90184 3108 90240 3164
rect 90288 3108 90344 3164
rect 90392 3108 90448 3164
<< metal4 >>
rect 4258 55692 4958 56508
rect 4258 55636 4268 55692
rect 4324 55636 4372 55692
rect 4428 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4788 55692
rect 4844 55636 4892 55692
rect 4948 55636 4958 55692
rect 4258 54124 4958 55636
rect 4258 54068 4268 54124
rect 4324 54068 4372 54124
rect 4428 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4788 54124
rect 4844 54068 4892 54124
rect 4948 54068 4958 54124
rect 4258 52556 4958 54068
rect 4258 52500 4268 52556
rect 4324 52500 4372 52556
rect 4428 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4788 52556
rect 4844 52500 4892 52556
rect 4948 52500 4958 52556
rect 4258 50988 4958 52500
rect 4258 50932 4268 50988
rect 4324 50932 4372 50988
rect 4428 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4788 50988
rect 4844 50932 4892 50988
rect 4948 50932 4958 50988
rect 4258 49420 4958 50932
rect 4258 49364 4268 49420
rect 4324 49364 4372 49420
rect 4428 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4788 49420
rect 4844 49364 4892 49420
rect 4948 49364 4958 49420
rect 4258 47852 4958 49364
rect 4258 47796 4268 47852
rect 4324 47796 4372 47852
rect 4428 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4788 47852
rect 4844 47796 4892 47852
rect 4948 47796 4958 47852
rect 4258 46284 4958 47796
rect 4258 46228 4268 46284
rect 4324 46228 4372 46284
rect 4428 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4788 46284
rect 4844 46228 4892 46284
rect 4948 46228 4958 46284
rect 4258 44716 4958 46228
rect 4258 44660 4268 44716
rect 4324 44660 4372 44716
rect 4428 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4788 44716
rect 4844 44660 4892 44716
rect 4948 44660 4958 44716
rect 4258 43148 4958 44660
rect 4258 43092 4268 43148
rect 4324 43092 4372 43148
rect 4428 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4788 43148
rect 4844 43092 4892 43148
rect 4948 43092 4958 43148
rect 4258 41580 4958 43092
rect 4258 41524 4268 41580
rect 4324 41524 4372 41580
rect 4428 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4788 41580
rect 4844 41524 4892 41580
rect 4948 41524 4958 41580
rect 4258 40012 4958 41524
rect 4258 39956 4268 40012
rect 4324 39956 4372 40012
rect 4428 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4788 40012
rect 4844 39956 4892 40012
rect 4948 39956 4958 40012
rect 4258 38444 4958 39956
rect 4258 38388 4268 38444
rect 4324 38388 4372 38444
rect 4428 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4788 38444
rect 4844 38388 4892 38444
rect 4948 38388 4958 38444
rect 4258 36876 4958 38388
rect 4258 36820 4268 36876
rect 4324 36820 4372 36876
rect 4428 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4788 36876
rect 4844 36820 4892 36876
rect 4948 36820 4958 36876
rect 4258 35308 4958 36820
rect 4258 35252 4268 35308
rect 4324 35252 4372 35308
rect 4428 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4788 35308
rect 4844 35252 4892 35308
rect 4948 35252 4958 35308
rect 4258 33740 4958 35252
rect 4258 33684 4268 33740
rect 4324 33684 4372 33740
rect 4428 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4788 33740
rect 4844 33684 4892 33740
rect 4948 33684 4958 33740
rect 4258 32172 4958 33684
rect 4258 32116 4268 32172
rect 4324 32116 4372 32172
rect 4428 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4788 32172
rect 4844 32116 4892 32172
rect 4948 32116 4958 32172
rect 4258 30604 4958 32116
rect 4258 30548 4268 30604
rect 4324 30548 4372 30604
rect 4428 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4788 30604
rect 4844 30548 4892 30604
rect 4948 30548 4958 30604
rect 4258 29036 4958 30548
rect 4258 28980 4268 29036
rect 4324 28980 4372 29036
rect 4428 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4788 29036
rect 4844 28980 4892 29036
rect 4948 28980 4958 29036
rect 4258 27468 4958 28980
rect 4258 27412 4268 27468
rect 4324 27412 4372 27468
rect 4428 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4788 27468
rect 4844 27412 4892 27468
rect 4948 27412 4958 27468
rect 4258 25900 4958 27412
rect 4258 25844 4268 25900
rect 4324 25844 4372 25900
rect 4428 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4788 25900
rect 4844 25844 4892 25900
rect 4948 25844 4958 25900
rect 4258 24332 4958 25844
rect 4258 24276 4268 24332
rect 4324 24276 4372 24332
rect 4428 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4788 24332
rect 4844 24276 4892 24332
rect 4948 24276 4958 24332
rect 4258 22764 4958 24276
rect 4258 22708 4268 22764
rect 4324 22708 4372 22764
rect 4428 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4788 22764
rect 4844 22708 4892 22764
rect 4948 22708 4958 22764
rect 4258 21196 4958 22708
rect 4258 21140 4268 21196
rect 4324 21140 4372 21196
rect 4428 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4788 21196
rect 4844 21140 4892 21196
rect 4948 21140 4958 21196
rect 4258 19628 4958 21140
rect 4258 19572 4268 19628
rect 4324 19572 4372 19628
rect 4428 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4788 19628
rect 4844 19572 4892 19628
rect 4948 19572 4958 19628
rect 4258 18060 4958 19572
rect 4258 18004 4268 18060
rect 4324 18004 4372 18060
rect 4428 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4788 18060
rect 4844 18004 4892 18060
rect 4948 18004 4958 18060
rect 4258 16492 4958 18004
rect 4258 16436 4268 16492
rect 4324 16436 4372 16492
rect 4428 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4788 16492
rect 4844 16436 4892 16492
rect 4948 16436 4958 16492
rect 4258 14924 4958 16436
rect 4258 14868 4268 14924
rect 4324 14868 4372 14924
rect 4428 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4788 14924
rect 4844 14868 4892 14924
rect 4948 14868 4958 14924
rect 4258 13356 4958 14868
rect 4258 13300 4268 13356
rect 4324 13300 4372 13356
rect 4428 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4788 13356
rect 4844 13300 4892 13356
rect 4948 13300 4958 13356
rect 4258 11788 4958 13300
rect 4258 11732 4268 11788
rect 4324 11732 4372 11788
rect 4428 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4788 11788
rect 4844 11732 4892 11788
rect 4948 11732 4958 11788
rect 4258 10220 4958 11732
rect 4258 10164 4268 10220
rect 4324 10164 4372 10220
rect 4428 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4788 10220
rect 4844 10164 4892 10220
rect 4948 10164 4958 10220
rect 4258 8652 4958 10164
rect 4258 8596 4268 8652
rect 4324 8596 4372 8652
rect 4428 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4788 8652
rect 4844 8596 4892 8652
rect 4948 8596 4958 8652
rect 4258 7084 4958 8596
rect 4258 7028 4268 7084
rect 4324 7028 4372 7084
rect 4428 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4788 7084
rect 4844 7028 4892 7084
rect 4948 7028 4958 7084
rect 4258 5516 4958 7028
rect 4258 5460 4268 5516
rect 4324 5460 4372 5516
rect 4428 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4788 5516
rect 4844 5460 4892 5516
rect 4948 5460 4958 5516
rect 4258 3948 4958 5460
rect 4258 3892 4268 3948
rect 4324 3892 4372 3948
rect 4428 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4788 3948
rect 4844 3892 4892 3948
rect 4948 3892 4958 3948
rect 4258 3076 4958 3892
rect 8758 56476 9458 56508
rect 8758 56420 8768 56476
rect 8824 56420 8872 56476
rect 8928 56420 8976 56476
rect 9032 56420 9080 56476
rect 9136 56420 9184 56476
rect 9240 56420 9288 56476
rect 9344 56420 9392 56476
rect 9448 56420 9458 56476
rect 8758 54908 9458 56420
rect 8758 54852 8768 54908
rect 8824 54852 8872 54908
rect 8928 54852 8976 54908
rect 9032 54852 9080 54908
rect 9136 54852 9184 54908
rect 9240 54852 9288 54908
rect 9344 54852 9392 54908
rect 9448 54852 9458 54908
rect 8758 53340 9458 54852
rect 8758 53284 8768 53340
rect 8824 53284 8872 53340
rect 8928 53284 8976 53340
rect 9032 53284 9080 53340
rect 9136 53284 9184 53340
rect 9240 53284 9288 53340
rect 9344 53284 9392 53340
rect 9448 53284 9458 53340
rect 8758 51772 9458 53284
rect 8758 51716 8768 51772
rect 8824 51716 8872 51772
rect 8928 51716 8976 51772
rect 9032 51716 9080 51772
rect 9136 51716 9184 51772
rect 9240 51716 9288 51772
rect 9344 51716 9392 51772
rect 9448 51716 9458 51772
rect 8758 50204 9458 51716
rect 8758 50148 8768 50204
rect 8824 50148 8872 50204
rect 8928 50148 8976 50204
rect 9032 50148 9080 50204
rect 9136 50148 9184 50204
rect 9240 50148 9288 50204
rect 9344 50148 9392 50204
rect 9448 50148 9458 50204
rect 8758 48636 9458 50148
rect 8758 48580 8768 48636
rect 8824 48580 8872 48636
rect 8928 48580 8976 48636
rect 9032 48580 9080 48636
rect 9136 48580 9184 48636
rect 9240 48580 9288 48636
rect 9344 48580 9392 48636
rect 9448 48580 9458 48636
rect 8758 47068 9458 48580
rect 8758 47012 8768 47068
rect 8824 47012 8872 47068
rect 8928 47012 8976 47068
rect 9032 47012 9080 47068
rect 9136 47012 9184 47068
rect 9240 47012 9288 47068
rect 9344 47012 9392 47068
rect 9448 47012 9458 47068
rect 8758 45500 9458 47012
rect 8758 45444 8768 45500
rect 8824 45444 8872 45500
rect 8928 45444 8976 45500
rect 9032 45444 9080 45500
rect 9136 45444 9184 45500
rect 9240 45444 9288 45500
rect 9344 45444 9392 45500
rect 9448 45444 9458 45500
rect 8758 43932 9458 45444
rect 8758 43876 8768 43932
rect 8824 43876 8872 43932
rect 8928 43876 8976 43932
rect 9032 43876 9080 43932
rect 9136 43876 9184 43932
rect 9240 43876 9288 43932
rect 9344 43876 9392 43932
rect 9448 43876 9458 43932
rect 8758 42364 9458 43876
rect 8758 42308 8768 42364
rect 8824 42308 8872 42364
rect 8928 42308 8976 42364
rect 9032 42308 9080 42364
rect 9136 42308 9184 42364
rect 9240 42308 9288 42364
rect 9344 42308 9392 42364
rect 9448 42308 9458 42364
rect 8758 40796 9458 42308
rect 8758 40740 8768 40796
rect 8824 40740 8872 40796
rect 8928 40740 8976 40796
rect 9032 40740 9080 40796
rect 9136 40740 9184 40796
rect 9240 40740 9288 40796
rect 9344 40740 9392 40796
rect 9448 40740 9458 40796
rect 8758 39228 9458 40740
rect 8758 39172 8768 39228
rect 8824 39172 8872 39228
rect 8928 39172 8976 39228
rect 9032 39172 9080 39228
rect 9136 39172 9184 39228
rect 9240 39172 9288 39228
rect 9344 39172 9392 39228
rect 9448 39172 9458 39228
rect 8758 37660 9458 39172
rect 8758 37604 8768 37660
rect 8824 37604 8872 37660
rect 8928 37604 8976 37660
rect 9032 37604 9080 37660
rect 9136 37604 9184 37660
rect 9240 37604 9288 37660
rect 9344 37604 9392 37660
rect 9448 37604 9458 37660
rect 8758 36092 9458 37604
rect 8758 36036 8768 36092
rect 8824 36036 8872 36092
rect 8928 36036 8976 36092
rect 9032 36036 9080 36092
rect 9136 36036 9184 36092
rect 9240 36036 9288 36092
rect 9344 36036 9392 36092
rect 9448 36036 9458 36092
rect 8758 34524 9458 36036
rect 8758 34468 8768 34524
rect 8824 34468 8872 34524
rect 8928 34468 8976 34524
rect 9032 34468 9080 34524
rect 9136 34468 9184 34524
rect 9240 34468 9288 34524
rect 9344 34468 9392 34524
rect 9448 34468 9458 34524
rect 8758 32956 9458 34468
rect 8758 32900 8768 32956
rect 8824 32900 8872 32956
rect 8928 32900 8976 32956
rect 9032 32900 9080 32956
rect 9136 32900 9184 32956
rect 9240 32900 9288 32956
rect 9344 32900 9392 32956
rect 9448 32900 9458 32956
rect 8758 31388 9458 32900
rect 8758 31332 8768 31388
rect 8824 31332 8872 31388
rect 8928 31332 8976 31388
rect 9032 31332 9080 31388
rect 9136 31332 9184 31388
rect 9240 31332 9288 31388
rect 9344 31332 9392 31388
rect 9448 31332 9458 31388
rect 8758 29820 9458 31332
rect 8758 29764 8768 29820
rect 8824 29764 8872 29820
rect 8928 29764 8976 29820
rect 9032 29764 9080 29820
rect 9136 29764 9184 29820
rect 9240 29764 9288 29820
rect 9344 29764 9392 29820
rect 9448 29764 9458 29820
rect 8758 28252 9458 29764
rect 8758 28196 8768 28252
rect 8824 28196 8872 28252
rect 8928 28196 8976 28252
rect 9032 28196 9080 28252
rect 9136 28196 9184 28252
rect 9240 28196 9288 28252
rect 9344 28196 9392 28252
rect 9448 28196 9458 28252
rect 8758 26684 9458 28196
rect 8758 26628 8768 26684
rect 8824 26628 8872 26684
rect 8928 26628 8976 26684
rect 9032 26628 9080 26684
rect 9136 26628 9184 26684
rect 9240 26628 9288 26684
rect 9344 26628 9392 26684
rect 9448 26628 9458 26684
rect 8758 25116 9458 26628
rect 8758 25060 8768 25116
rect 8824 25060 8872 25116
rect 8928 25060 8976 25116
rect 9032 25060 9080 25116
rect 9136 25060 9184 25116
rect 9240 25060 9288 25116
rect 9344 25060 9392 25116
rect 9448 25060 9458 25116
rect 8758 23548 9458 25060
rect 8758 23492 8768 23548
rect 8824 23492 8872 23548
rect 8928 23492 8976 23548
rect 9032 23492 9080 23548
rect 9136 23492 9184 23548
rect 9240 23492 9288 23548
rect 9344 23492 9392 23548
rect 9448 23492 9458 23548
rect 8758 21980 9458 23492
rect 8758 21924 8768 21980
rect 8824 21924 8872 21980
rect 8928 21924 8976 21980
rect 9032 21924 9080 21980
rect 9136 21924 9184 21980
rect 9240 21924 9288 21980
rect 9344 21924 9392 21980
rect 9448 21924 9458 21980
rect 8758 20412 9458 21924
rect 8758 20356 8768 20412
rect 8824 20356 8872 20412
rect 8928 20356 8976 20412
rect 9032 20356 9080 20412
rect 9136 20356 9184 20412
rect 9240 20356 9288 20412
rect 9344 20356 9392 20412
rect 9448 20356 9458 20412
rect 8758 18844 9458 20356
rect 8758 18788 8768 18844
rect 8824 18788 8872 18844
rect 8928 18788 8976 18844
rect 9032 18788 9080 18844
rect 9136 18788 9184 18844
rect 9240 18788 9288 18844
rect 9344 18788 9392 18844
rect 9448 18788 9458 18844
rect 8758 17276 9458 18788
rect 8758 17220 8768 17276
rect 8824 17220 8872 17276
rect 8928 17220 8976 17276
rect 9032 17220 9080 17276
rect 9136 17220 9184 17276
rect 9240 17220 9288 17276
rect 9344 17220 9392 17276
rect 9448 17220 9458 17276
rect 8758 15708 9458 17220
rect 8758 15652 8768 15708
rect 8824 15652 8872 15708
rect 8928 15652 8976 15708
rect 9032 15652 9080 15708
rect 9136 15652 9184 15708
rect 9240 15652 9288 15708
rect 9344 15652 9392 15708
rect 9448 15652 9458 15708
rect 8758 14140 9458 15652
rect 8758 14084 8768 14140
rect 8824 14084 8872 14140
rect 8928 14084 8976 14140
rect 9032 14084 9080 14140
rect 9136 14084 9184 14140
rect 9240 14084 9288 14140
rect 9344 14084 9392 14140
rect 9448 14084 9458 14140
rect 8758 12572 9458 14084
rect 8758 12516 8768 12572
rect 8824 12516 8872 12572
rect 8928 12516 8976 12572
rect 9032 12516 9080 12572
rect 9136 12516 9184 12572
rect 9240 12516 9288 12572
rect 9344 12516 9392 12572
rect 9448 12516 9458 12572
rect 8758 11004 9458 12516
rect 8758 10948 8768 11004
rect 8824 10948 8872 11004
rect 8928 10948 8976 11004
rect 9032 10948 9080 11004
rect 9136 10948 9184 11004
rect 9240 10948 9288 11004
rect 9344 10948 9392 11004
rect 9448 10948 9458 11004
rect 8758 9436 9458 10948
rect 8758 9380 8768 9436
rect 8824 9380 8872 9436
rect 8928 9380 8976 9436
rect 9032 9380 9080 9436
rect 9136 9380 9184 9436
rect 9240 9380 9288 9436
rect 9344 9380 9392 9436
rect 9448 9380 9458 9436
rect 8758 7868 9458 9380
rect 8758 7812 8768 7868
rect 8824 7812 8872 7868
rect 8928 7812 8976 7868
rect 9032 7812 9080 7868
rect 9136 7812 9184 7868
rect 9240 7812 9288 7868
rect 9344 7812 9392 7868
rect 9448 7812 9458 7868
rect 8758 6300 9458 7812
rect 8758 6244 8768 6300
rect 8824 6244 8872 6300
rect 8928 6244 8976 6300
rect 9032 6244 9080 6300
rect 9136 6244 9184 6300
rect 9240 6244 9288 6300
rect 9344 6244 9392 6300
rect 9448 6244 9458 6300
rect 8758 4732 9458 6244
rect 8758 4676 8768 4732
rect 8824 4676 8872 4732
rect 8928 4676 8976 4732
rect 9032 4676 9080 4732
rect 9136 4676 9184 4732
rect 9240 4676 9288 4732
rect 9344 4676 9392 4732
rect 9448 4676 9458 4732
rect 8758 3164 9458 4676
rect 8758 3108 8768 3164
rect 8824 3108 8872 3164
rect 8928 3108 8976 3164
rect 9032 3108 9080 3164
rect 9136 3108 9184 3164
rect 9240 3108 9288 3164
rect 9344 3108 9392 3164
rect 9448 3108 9458 3164
rect 8758 3076 9458 3108
rect 13258 55692 13958 56508
rect 13258 55636 13268 55692
rect 13324 55636 13372 55692
rect 13428 55636 13476 55692
rect 13532 55636 13580 55692
rect 13636 55636 13684 55692
rect 13740 55636 13788 55692
rect 13844 55636 13892 55692
rect 13948 55636 13958 55692
rect 13258 54124 13958 55636
rect 13258 54068 13268 54124
rect 13324 54068 13372 54124
rect 13428 54068 13476 54124
rect 13532 54068 13580 54124
rect 13636 54068 13684 54124
rect 13740 54068 13788 54124
rect 13844 54068 13892 54124
rect 13948 54068 13958 54124
rect 13258 52556 13958 54068
rect 13258 52500 13268 52556
rect 13324 52500 13372 52556
rect 13428 52500 13476 52556
rect 13532 52500 13580 52556
rect 13636 52500 13684 52556
rect 13740 52500 13788 52556
rect 13844 52500 13892 52556
rect 13948 52500 13958 52556
rect 13258 50988 13958 52500
rect 13258 50932 13268 50988
rect 13324 50932 13372 50988
rect 13428 50932 13476 50988
rect 13532 50932 13580 50988
rect 13636 50932 13684 50988
rect 13740 50932 13788 50988
rect 13844 50932 13892 50988
rect 13948 50932 13958 50988
rect 13258 49420 13958 50932
rect 13258 49364 13268 49420
rect 13324 49364 13372 49420
rect 13428 49364 13476 49420
rect 13532 49364 13580 49420
rect 13636 49364 13684 49420
rect 13740 49364 13788 49420
rect 13844 49364 13892 49420
rect 13948 49364 13958 49420
rect 13258 47852 13958 49364
rect 13258 47796 13268 47852
rect 13324 47796 13372 47852
rect 13428 47796 13476 47852
rect 13532 47796 13580 47852
rect 13636 47796 13684 47852
rect 13740 47796 13788 47852
rect 13844 47796 13892 47852
rect 13948 47796 13958 47852
rect 13258 46284 13958 47796
rect 13258 46228 13268 46284
rect 13324 46228 13372 46284
rect 13428 46228 13476 46284
rect 13532 46228 13580 46284
rect 13636 46228 13684 46284
rect 13740 46228 13788 46284
rect 13844 46228 13892 46284
rect 13948 46228 13958 46284
rect 13258 44716 13958 46228
rect 13258 44660 13268 44716
rect 13324 44660 13372 44716
rect 13428 44660 13476 44716
rect 13532 44660 13580 44716
rect 13636 44660 13684 44716
rect 13740 44660 13788 44716
rect 13844 44660 13892 44716
rect 13948 44660 13958 44716
rect 13258 43148 13958 44660
rect 13258 43092 13268 43148
rect 13324 43092 13372 43148
rect 13428 43092 13476 43148
rect 13532 43092 13580 43148
rect 13636 43092 13684 43148
rect 13740 43092 13788 43148
rect 13844 43092 13892 43148
rect 13948 43092 13958 43148
rect 13258 41580 13958 43092
rect 13258 41524 13268 41580
rect 13324 41524 13372 41580
rect 13428 41524 13476 41580
rect 13532 41524 13580 41580
rect 13636 41524 13684 41580
rect 13740 41524 13788 41580
rect 13844 41524 13892 41580
rect 13948 41524 13958 41580
rect 13258 40012 13958 41524
rect 13258 39956 13268 40012
rect 13324 39956 13372 40012
rect 13428 39956 13476 40012
rect 13532 39956 13580 40012
rect 13636 39956 13684 40012
rect 13740 39956 13788 40012
rect 13844 39956 13892 40012
rect 13948 39956 13958 40012
rect 13258 38444 13958 39956
rect 13258 38388 13268 38444
rect 13324 38388 13372 38444
rect 13428 38388 13476 38444
rect 13532 38388 13580 38444
rect 13636 38388 13684 38444
rect 13740 38388 13788 38444
rect 13844 38388 13892 38444
rect 13948 38388 13958 38444
rect 13258 36876 13958 38388
rect 13258 36820 13268 36876
rect 13324 36820 13372 36876
rect 13428 36820 13476 36876
rect 13532 36820 13580 36876
rect 13636 36820 13684 36876
rect 13740 36820 13788 36876
rect 13844 36820 13892 36876
rect 13948 36820 13958 36876
rect 13258 35308 13958 36820
rect 13258 35252 13268 35308
rect 13324 35252 13372 35308
rect 13428 35252 13476 35308
rect 13532 35252 13580 35308
rect 13636 35252 13684 35308
rect 13740 35252 13788 35308
rect 13844 35252 13892 35308
rect 13948 35252 13958 35308
rect 13258 33740 13958 35252
rect 13258 33684 13268 33740
rect 13324 33684 13372 33740
rect 13428 33684 13476 33740
rect 13532 33684 13580 33740
rect 13636 33684 13684 33740
rect 13740 33684 13788 33740
rect 13844 33684 13892 33740
rect 13948 33684 13958 33740
rect 13258 32172 13958 33684
rect 13258 32116 13268 32172
rect 13324 32116 13372 32172
rect 13428 32116 13476 32172
rect 13532 32116 13580 32172
rect 13636 32116 13684 32172
rect 13740 32116 13788 32172
rect 13844 32116 13892 32172
rect 13948 32116 13958 32172
rect 13258 30604 13958 32116
rect 13258 30548 13268 30604
rect 13324 30548 13372 30604
rect 13428 30548 13476 30604
rect 13532 30548 13580 30604
rect 13636 30548 13684 30604
rect 13740 30548 13788 30604
rect 13844 30548 13892 30604
rect 13948 30548 13958 30604
rect 13258 29036 13958 30548
rect 13258 28980 13268 29036
rect 13324 28980 13372 29036
rect 13428 28980 13476 29036
rect 13532 28980 13580 29036
rect 13636 28980 13684 29036
rect 13740 28980 13788 29036
rect 13844 28980 13892 29036
rect 13948 28980 13958 29036
rect 13258 27468 13958 28980
rect 13258 27412 13268 27468
rect 13324 27412 13372 27468
rect 13428 27412 13476 27468
rect 13532 27412 13580 27468
rect 13636 27412 13684 27468
rect 13740 27412 13788 27468
rect 13844 27412 13892 27468
rect 13948 27412 13958 27468
rect 13258 25900 13958 27412
rect 13258 25844 13268 25900
rect 13324 25844 13372 25900
rect 13428 25844 13476 25900
rect 13532 25844 13580 25900
rect 13636 25844 13684 25900
rect 13740 25844 13788 25900
rect 13844 25844 13892 25900
rect 13948 25844 13958 25900
rect 13258 24332 13958 25844
rect 13258 24276 13268 24332
rect 13324 24276 13372 24332
rect 13428 24276 13476 24332
rect 13532 24276 13580 24332
rect 13636 24276 13684 24332
rect 13740 24276 13788 24332
rect 13844 24276 13892 24332
rect 13948 24276 13958 24332
rect 13258 22764 13958 24276
rect 13258 22708 13268 22764
rect 13324 22708 13372 22764
rect 13428 22708 13476 22764
rect 13532 22708 13580 22764
rect 13636 22708 13684 22764
rect 13740 22708 13788 22764
rect 13844 22708 13892 22764
rect 13948 22708 13958 22764
rect 13258 21196 13958 22708
rect 13258 21140 13268 21196
rect 13324 21140 13372 21196
rect 13428 21140 13476 21196
rect 13532 21140 13580 21196
rect 13636 21140 13684 21196
rect 13740 21140 13788 21196
rect 13844 21140 13892 21196
rect 13948 21140 13958 21196
rect 13258 19628 13958 21140
rect 13258 19572 13268 19628
rect 13324 19572 13372 19628
rect 13428 19572 13476 19628
rect 13532 19572 13580 19628
rect 13636 19572 13684 19628
rect 13740 19572 13788 19628
rect 13844 19572 13892 19628
rect 13948 19572 13958 19628
rect 13258 18060 13958 19572
rect 13258 18004 13268 18060
rect 13324 18004 13372 18060
rect 13428 18004 13476 18060
rect 13532 18004 13580 18060
rect 13636 18004 13684 18060
rect 13740 18004 13788 18060
rect 13844 18004 13892 18060
rect 13948 18004 13958 18060
rect 13258 16492 13958 18004
rect 13258 16436 13268 16492
rect 13324 16436 13372 16492
rect 13428 16436 13476 16492
rect 13532 16436 13580 16492
rect 13636 16436 13684 16492
rect 13740 16436 13788 16492
rect 13844 16436 13892 16492
rect 13948 16436 13958 16492
rect 13258 14924 13958 16436
rect 13258 14868 13268 14924
rect 13324 14868 13372 14924
rect 13428 14868 13476 14924
rect 13532 14868 13580 14924
rect 13636 14868 13684 14924
rect 13740 14868 13788 14924
rect 13844 14868 13892 14924
rect 13948 14868 13958 14924
rect 13258 13356 13958 14868
rect 13258 13300 13268 13356
rect 13324 13300 13372 13356
rect 13428 13300 13476 13356
rect 13532 13300 13580 13356
rect 13636 13300 13684 13356
rect 13740 13300 13788 13356
rect 13844 13300 13892 13356
rect 13948 13300 13958 13356
rect 13258 11788 13958 13300
rect 13258 11732 13268 11788
rect 13324 11732 13372 11788
rect 13428 11732 13476 11788
rect 13532 11732 13580 11788
rect 13636 11732 13684 11788
rect 13740 11732 13788 11788
rect 13844 11732 13892 11788
rect 13948 11732 13958 11788
rect 13258 10220 13958 11732
rect 13258 10164 13268 10220
rect 13324 10164 13372 10220
rect 13428 10164 13476 10220
rect 13532 10164 13580 10220
rect 13636 10164 13684 10220
rect 13740 10164 13788 10220
rect 13844 10164 13892 10220
rect 13948 10164 13958 10220
rect 13258 8652 13958 10164
rect 13258 8596 13268 8652
rect 13324 8596 13372 8652
rect 13428 8596 13476 8652
rect 13532 8596 13580 8652
rect 13636 8596 13684 8652
rect 13740 8596 13788 8652
rect 13844 8596 13892 8652
rect 13948 8596 13958 8652
rect 13258 7084 13958 8596
rect 13258 7028 13268 7084
rect 13324 7028 13372 7084
rect 13428 7028 13476 7084
rect 13532 7028 13580 7084
rect 13636 7028 13684 7084
rect 13740 7028 13788 7084
rect 13844 7028 13892 7084
rect 13948 7028 13958 7084
rect 13258 5516 13958 7028
rect 13258 5460 13268 5516
rect 13324 5460 13372 5516
rect 13428 5460 13476 5516
rect 13532 5460 13580 5516
rect 13636 5460 13684 5516
rect 13740 5460 13788 5516
rect 13844 5460 13892 5516
rect 13948 5460 13958 5516
rect 13258 3948 13958 5460
rect 13258 3892 13268 3948
rect 13324 3892 13372 3948
rect 13428 3892 13476 3948
rect 13532 3892 13580 3948
rect 13636 3892 13684 3948
rect 13740 3892 13788 3948
rect 13844 3892 13892 3948
rect 13948 3892 13958 3948
rect 13258 3076 13958 3892
rect 17758 56476 18458 56508
rect 17758 56420 17768 56476
rect 17824 56420 17872 56476
rect 17928 56420 17976 56476
rect 18032 56420 18080 56476
rect 18136 56420 18184 56476
rect 18240 56420 18288 56476
rect 18344 56420 18392 56476
rect 18448 56420 18458 56476
rect 17758 54908 18458 56420
rect 17758 54852 17768 54908
rect 17824 54852 17872 54908
rect 17928 54852 17976 54908
rect 18032 54852 18080 54908
rect 18136 54852 18184 54908
rect 18240 54852 18288 54908
rect 18344 54852 18392 54908
rect 18448 54852 18458 54908
rect 17758 53340 18458 54852
rect 17758 53284 17768 53340
rect 17824 53284 17872 53340
rect 17928 53284 17976 53340
rect 18032 53284 18080 53340
rect 18136 53284 18184 53340
rect 18240 53284 18288 53340
rect 18344 53284 18392 53340
rect 18448 53284 18458 53340
rect 17758 51772 18458 53284
rect 17758 51716 17768 51772
rect 17824 51716 17872 51772
rect 17928 51716 17976 51772
rect 18032 51716 18080 51772
rect 18136 51716 18184 51772
rect 18240 51716 18288 51772
rect 18344 51716 18392 51772
rect 18448 51716 18458 51772
rect 17758 50204 18458 51716
rect 17758 50148 17768 50204
rect 17824 50148 17872 50204
rect 17928 50148 17976 50204
rect 18032 50148 18080 50204
rect 18136 50148 18184 50204
rect 18240 50148 18288 50204
rect 18344 50148 18392 50204
rect 18448 50148 18458 50204
rect 17758 48636 18458 50148
rect 17758 48580 17768 48636
rect 17824 48580 17872 48636
rect 17928 48580 17976 48636
rect 18032 48580 18080 48636
rect 18136 48580 18184 48636
rect 18240 48580 18288 48636
rect 18344 48580 18392 48636
rect 18448 48580 18458 48636
rect 17758 47068 18458 48580
rect 17758 47012 17768 47068
rect 17824 47012 17872 47068
rect 17928 47012 17976 47068
rect 18032 47012 18080 47068
rect 18136 47012 18184 47068
rect 18240 47012 18288 47068
rect 18344 47012 18392 47068
rect 18448 47012 18458 47068
rect 17758 45500 18458 47012
rect 17758 45444 17768 45500
rect 17824 45444 17872 45500
rect 17928 45444 17976 45500
rect 18032 45444 18080 45500
rect 18136 45444 18184 45500
rect 18240 45444 18288 45500
rect 18344 45444 18392 45500
rect 18448 45444 18458 45500
rect 17758 43932 18458 45444
rect 17758 43876 17768 43932
rect 17824 43876 17872 43932
rect 17928 43876 17976 43932
rect 18032 43876 18080 43932
rect 18136 43876 18184 43932
rect 18240 43876 18288 43932
rect 18344 43876 18392 43932
rect 18448 43876 18458 43932
rect 17758 42364 18458 43876
rect 17758 42308 17768 42364
rect 17824 42308 17872 42364
rect 17928 42308 17976 42364
rect 18032 42308 18080 42364
rect 18136 42308 18184 42364
rect 18240 42308 18288 42364
rect 18344 42308 18392 42364
rect 18448 42308 18458 42364
rect 17758 40796 18458 42308
rect 17758 40740 17768 40796
rect 17824 40740 17872 40796
rect 17928 40740 17976 40796
rect 18032 40740 18080 40796
rect 18136 40740 18184 40796
rect 18240 40740 18288 40796
rect 18344 40740 18392 40796
rect 18448 40740 18458 40796
rect 17758 39228 18458 40740
rect 17758 39172 17768 39228
rect 17824 39172 17872 39228
rect 17928 39172 17976 39228
rect 18032 39172 18080 39228
rect 18136 39172 18184 39228
rect 18240 39172 18288 39228
rect 18344 39172 18392 39228
rect 18448 39172 18458 39228
rect 17758 37660 18458 39172
rect 17758 37604 17768 37660
rect 17824 37604 17872 37660
rect 17928 37604 17976 37660
rect 18032 37604 18080 37660
rect 18136 37604 18184 37660
rect 18240 37604 18288 37660
rect 18344 37604 18392 37660
rect 18448 37604 18458 37660
rect 17758 36092 18458 37604
rect 17758 36036 17768 36092
rect 17824 36036 17872 36092
rect 17928 36036 17976 36092
rect 18032 36036 18080 36092
rect 18136 36036 18184 36092
rect 18240 36036 18288 36092
rect 18344 36036 18392 36092
rect 18448 36036 18458 36092
rect 17758 34524 18458 36036
rect 17758 34468 17768 34524
rect 17824 34468 17872 34524
rect 17928 34468 17976 34524
rect 18032 34468 18080 34524
rect 18136 34468 18184 34524
rect 18240 34468 18288 34524
rect 18344 34468 18392 34524
rect 18448 34468 18458 34524
rect 17758 32956 18458 34468
rect 17758 32900 17768 32956
rect 17824 32900 17872 32956
rect 17928 32900 17976 32956
rect 18032 32900 18080 32956
rect 18136 32900 18184 32956
rect 18240 32900 18288 32956
rect 18344 32900 18392 32956
rect 18448 32900 18458 32956
rect 17758 31388 18458 32900
rect 17758 31332 17768 31388
rect 17824 31332 17872 31388
rect 17928 31332 17976 31388
rect 18032 31332 18080 31388
rect 18136 31332 18184 31388
rect 18240 31332 18288 31388
rect 18344 31332 18392 31388
rect 18448 31332 18458 31388
rect 17758 29820 18458 31332
rect 17758 29764 17768 29820
rect 17824 29764 17872 29820
rect 17928 29764 17976 29820
rect 18032 29764 18080 29820
rect 18136 29764 18184 29820
rect 18240 29764 18288 29820
rect 18344 29764 18392 29820
rect 18448 29764 18458 29820
rect 17758 28252 18458 29764
rect 17758 28196 17768 28252
rect 17824 28196 17872 28252
rect 17928 28196 17976 28252
rect 18032 28196 18080 28252
rect 18136 28196 18184 28252
rect 18240 28196 18288 28252
rect 18344 28196 18392 28252
rect 18448 28196 18458 28252
rect 17758 26684 18458 28196
rect 17758 26628 17768 26684
rect 17824 26628 17872 26684
rect 17928 26628 17976 26684
rect 18032 26628 18080 26684
rect 18136 26628 18184 26684
rect 18240 26628 18288 26684
rect 18344 26628 18392 26684
rect 18448 26628 18458 26684
rect 17758 25116 18458 26628
rect 17758 25060 17768 25116
rect 17824 25060 17872 25116
rect 17928 25060 17976 25116
rect 18032 25060 18080 25116
rect 18136 25060 18184 25116
rect 18240 25060 18288 25116
rect 18344 25060 18392 25116
rect 18448 25060 18458 25116
rect 17758 23548 18458 25060
rect 17758 23492 17768 23548
rect 17824 23492 17872 23548
rect 17928 23492 17976 23548
rect 18032 23492 18080 23548
rect 18136 23492 18184 23548
rect 18240 23492 18288 23548
rect 18344 23492 18392 23548
rect 18448 23492 18458 23548
rect 17758 21980 18458 23492
rect 17758 21924 17768 21980
rect 17824 21924 17872 21980
rect 17928 21924 17976 21980
rect 18032 21924 18080 21980
rect 18136 21924 18184 21980
rect 18240 21924 18288 21980
rect 18344 21924 18392 21980
rect 18448 21924 18458 21980
rect 17758 20412 18458 21924
rect 17758 20356 17768 20412
rect 17824 20356 17872 20412
rect 17928 20356 17976 20412
rect 18032 20356 18080 20412
rect 18136 20356 18184 20412
rect 18240 20356 18288 20412
rect 18344 20356 18392 20412
rect 18448 20356 18458 20412
rect 17758 18844 18458 20356
rect 17758 18788 17768 18844
rect 17824 18788 17872 18844
rect 17928 18788 17976 18844
rect 18032 18788 18080 18844
rect 18136 18788 18184 18844
rect 18240 18788 18288 18844
rect 18344 18788 18392 18844
rect 18448 18788 18458 18844
rect 17758 17276 18458 18788
rect 17758 17220 17768 17276
rect 17824 17220 17872 17276
rect 17928 17220 17976 17276
rect 18032 17220 18080 17276
rect 18136 17220 18184 17276
rect 18240 17220 18288 17276
rect 18344 17220 18392 17276
rect 18448 17220 18458 17276
rect 17758 15708 18458 17220
rect 17758 15652 17768 15708
rect 17824 15652 17872 15708
rect 17928 15652 17976 15708
rect 18032 15652 18080 15708
rect 18136 15652 18184 15708
rect 18240 15652 18288 15708
rect 18344 15652 18392 15708
rect 18448 15652 18458 15708
rect 17758 14140 18458 15652
rect 17758 14084 17768 14140
rect 17824 14084 17872 14140
rect 17928 14084 17976 14140
rect 18032 14084 18080 14140
rect 18136 14084 18184 14140
rect 18240 14084 18288 14140
rect 18344 14084 18392 14140
rect 18448 14084 18458 14140
rect 17758 12572 18458 14084
rect 17758 12516 17768 12572
rect 17824 12516 17872 12572
rect 17928 12516 17976 12572
rect 18032 12516 18080 12572
rect 18136 12516 18184 12572
rect 18240 12516 18288 12572
rect 18344 12516 18392 12572
rect 18448 12516 18458 12572
rect 17758 11004 18458 12516
rect 17758 10948 17768 11004
rect 17824 10948 17872 11004
rect 17928 10948 17976 11004
rect 18032 10948 18080 11004
rect 18136 10948 18184 11004
rect 18240 10948 18288 11004
rect 18344 10948 18392 11004
rect 18448 10948 18458 11004
rect 17758 9436 18458 10948
rect 17758 9380 17768 9436
rect 17824 9380 17872 9436
rect 17928 9380 17976 9436
rect 18032 9380 18080 9436
rect 18136 9380 18184 9436
rect 18240 9380 18288 9436
rect 18344 9380 18392 9436
rect 18448 9380 18458 9436
rect 17758 7868 18458 9380
rect 17758 7812 17768 7868
rect 17824 7812 17872 7868
rect 17928 7812 17976 7868
rect 18032 7812 18080 7868
rect 18136 7812 18184 7868
rect 18240 7812 18288 7868
rect 18344 7812 18392 7868
rect 18448 7812 18458 7868
rect 17758 6300 18458 7812
rect 17758 6244 17768 6300
rect 17824 6244 17872 6300
rect 17928 6244 17976 6300
rect 18032 6244 18080 6300
rect 18136 6244 18184 6300
rect 18240 6244 18288 6300
rect 18344 6244 18392 6300
rect 18448 6244 18458 6300
rect 17758 4732 18458 6244
rect 17758 4676 17768 4732
rect 17824 4676 17872 4732
rect 17928 4676 17976 4732
rect 18032 4676 18080 4732
rect 18136 4676 18184 4732
rect 18240 4676 18288 4732
rect 18344 4676 18392 4732
rect 18448 4676 18458 4732
rect 17758 3164 18458 4676
rect 17758 3108 17768 3164
rect 17824 3108 17872 3164
rect 17928 3108 17976 3164
rect 18032 3108 18080 3164
rect 18136 3108 18184 3164
rect 18240 3108 18288 3164
rect 18344 3108 18392 3164
rect 18448 3108 18458 3164
rect 17758 3076 18458 3108
rect 22258 55692 22958 56508
rect 22258 55636 22268 55692
rect 22324 55636 22372 55692
rect 22428 55636 22476 55692
rect 22532 55636 22580 55692
rect 22636 55636 22684 55692
rect 22740 55636 22788 55692
rect 22844 55636 22892 55692
rect 22948 55636 22958 55692
rect 22258 54124 22958 55636
rect 22258 54068 22268 54124
rect 22324 54068 22372 54124
rect 22428 54068 22476 54124
rect 22532 54068 22580 54124
rect 22636 54068 22684 54124
rect 22740 54068 22788 54124
rect 22844 54068 22892 54124
rect 22948 54068 22958 54124
rect 22258 52556 22958 54068
rect 22258 52500 22268 52556
rect 22324 52500 22372 52556
rect 22428 52500 22476 52556
rect 22532 52500 22580 52556
rect 22636 52500 22684 52556
rect 22740 52500 22788 52556
rect 22844 52500 22892 52556
rect 22948 52500 22958 52556
rect 22258 50988 22958 52500
rect 22258 50932 22268 50988
rect 22324 50932 22372 50988
rect 22428 50932 22476 50988
rect 22532 50932 22580 50988
rect 22636 50932 22684 50988
rect 22740 50932 22788 50988
rect 22844 50932 22892 50988
rect 22948 50932 22958 50988
rect 22258 49420 22958 50932
rect 22258 49364 22268 49420
rect 22324 49364 22372 49420
rect 22428 49364 22476 49420
rect 22532 49364 22580 49420
rect 22636 49364 22684 49420
rect 22740 49364 22788 49420
rect 22844 49364 22892 49420
rect 22948 49364 22958 49420
rect 22258 47852 22958 49364
rect 22258 47796 22268 47852
rect 22324 47796 22372 47852
rect 22428 47796 22476 47852
rect 22532 47796 22580 47852
rect 22636 47796 22684 47852
rect 22740 47796 22788 47852
rect 22844 47796 22892 47852
rect 22948 47796 22958 47852
rect 22258 46284 22958 47796
rect 22258 46228 22268 46284
rect 22324 46228 22372 46284
rect 22428 46228 22476 46284
rect 22532 46228 22580 46284
rect 22636 46228 22684 46284
rect 22740 46228 22788 46284
rect 22844 46228 22892 46284
rect 22948 46228 22958 46284
rect 22258 44716 22958 46228
rect 22258 44660 22268 44716
rect 22324 44660 22372 44716
rect 22428 44660 22476 44716
rect 22532 44660 22580 44716
rect 22636 44660 22684 44716
rect 22740 44660 22788 44716
rect 22844 44660 22892 44716
rect 22948 44660 22958 44716
rect 22258 43148 22958 44660
rect 22258 43092 22268 43148
rect 22324 43092 22372 43148
rect 22428 43092 22476 43148
rect 22532 43092 22580 43148
rect 22636 43092 22684 43148
rect 22740 43092 22788 43148
rect 22844 43092 22892 43148
rect 22948 43092 22958 43148
rect 22258 41580 22958 43092
rect 22258 41524 22268 41580
rect 22324 41524 22372 41580
rect 22428 41524 22476 41580
rect 22532 41524 22580 41580
rect 22636 41524 22684 41580
rect 22740 41524 22788 41580
rect 22844 41524 22892 41580
rect 22948 41524 22958 41580
rect 22258 40012 22958 41524
rect 22258 39956 22268 40012
rect 22324 39956 22372 40012
rect 22428 39956 22476 40012
rect 22532 39956 22580 40012
rect 22636 39956 22684 40012
rect 22740 39956 22788 40012
rect 22844 39956 22892 40012
rect 22948 39956 22958 40012
rect 22258 38444 22958 39956
rect 22258 38388 22268 38444
rect 22324 38388 22372 38444
rect 22428 38388 22476 38444
rect 22532 38388 22580 38444
rect 22636 38388 22684 38444
rect 22740 38388 22788 38444
rect 22844 38388 22892 38444
rect 22948 38388 22958 38444
rect 22258 36876 22958 38388
rect 22258 36820 22268 36876
rect 22324 36820 22372 36876
rect 22428 36820 22476 36876
rect 22532 36820 22580 36876
rect 22636 36820 22684 36876
rect 22740 36820 22788 36876
rect 22844 36820 22892 36876
rect 22948 36820 22958 36876
rect 22258 35308 22958 36820
rect 22258 35252 22268 35308
rect 22324 35252 22372 35308
rect 22428 35252 22476 35308
rect 22532 35252 22580 35308
rect 22636 35252 22684 35308
rect 22740 35252 22788 35308
rect 22844 35252 22892 35308
rect 22948 35252 22958 35308
rect 22258 33740 22958 35252
rect 22258 33684 22268 33740
rect 22324 33684 22372 33740
rect 22428 33684 22476 33740
rect 22532 33684 22580 33740
rect 22636 33684 22684 33740
rect 22740 33684 22788 33740
rect 22844 33684 22892 33740
rect 22948 33684 22958 33740
rect 22258 32172 22958 33684
rect 22258 32116 22268 32172
rect 22324 32116 22372 32172
rect 22428 32116 22476 32172
rect 22532 32116 22580 32172
rect 22636 32116 22684 32172
rect 22740 32116 22788 32172
rect 22844 32116 22892 32172
rect 22948 32116 22958 32172
rect 22258 30604 22958 32116
rect 22258 30548 22268 30604
rect 22324 30548 22372 30604
rect 22428 30548 22476 30604
rect 22532 30548 22580 30604
rect 22636 30548 22684 30604
rect 22740 30548 22788 30604
rect 22844 30548 22892 30604
rect 22948 30548 22958 30604
rect 22258 29036 22958 30548
rect 22258 28980 22268 29036
rect 22324 28980 22372 29036
rect 22428 28980 22476 29036
rect 22532 28980 22580 29036
rect 22636 28980 22684 29036
rect 22740 28980 22788 29036
rect 22844 28980 22892 29036
rect 22948 28980 22958 29036
rect 22258 27468 22958 28980
rect 22258 27412 22268 27468
rect 22324 27412 22372 27468
rect 22428 27412 22476 27468
rect 22532 27412 22580 27468
rect 22636 27412 22684 27468
rect 22740 27412 22788 27468
rect 22844 27412 22892 27468
rect 22948 27412 22958 27468
rect 22258 25900 22958 27412
rect 22258 25844 22268 25900
rect 22324 25844 22372 25900
rect 22428 25844 22476 25900
rect 22532 25844 22580 25900
rect 22636 25844 22684 25900
rect 22740 25844 22788 25900
rect 22844 25844 22892 25900
rect 22948 25844 22958 25900
rect 22258 24332 22958 25844
rect 22258 24276 22268 24332
rect 22324 24276 22372 24332
rect 22428 24276 22476 24332
rect 22532 24276 22580 24332
rect 22636 24276 22684 24332
rect 22740 24276 22788 24332
rect 22844 24276 22892 24332
rect 22948 24276 22958 24332
rect 22258 22764 22958 24276
rect 22258 22708 22268 22764
rect 22324 22708 22372 22764
rect 22428 22708 22476 22764
rect 22532 22708 22580 22764
rect 22636 22708 22684 22764
rect 22740 22708 22788 22764
rect 22844 22708 22892 22764
rect 22948 22708 22958 22764
rect 22258 21196 22958 22708
rect 22258 21140 22268 21196
rect 22324 21140 22372 21196
rect 22428 21140 22476 21196
rect 22532 21140 22580 21196
rect 22636 21140 22684 21196
rect 22740 21140 22788 21196
rect 22844 21140 22892 21196
rect 22948 21140 22958 21196
rect 22258 19628 22958 21140
rect 22258 19572 22268 19628
rect 22324 19572 22372 19628
rect 22428 19572 22476 19628
rect 22532 19572 22580 19628
rect 22636 19572 22684 19628
rect 22740 19572 22788 19628
rect 22844 19572 22892 19628
rect 22948 19572 22958 19628
rect 22258 18060 22958 19572
rect 22258 18004 22268 18060
rect 22324 18004 22372 18060
rect 22428 18004 22476 18060
rect 22532 18004 22580 18060
rect 22636 18004 22684 18060
rect 22740 18004 22788 18060
rect 22844 18004 22892 18060
rect 22948 18004 22958 18060
rect 22258 16492 22958 18004
rect 22258 16436 22268 16492
rect 22324 16436 22372 16492
rect 22428 16436 22476 16492
rect 22532 16436 22580 16492
rect 22636 16436 22684 16492
rect 22740 16436 22788 16492
rect 22844 16436 22892 16492
rect 22948 16436 22958 16492
rect 22258 14924 22958 16436
rect 22258 14868 22268 14924
rect 22324 14868 22372 14924
rect 22428 14868 22476 14924
rect 22532 14868 22580 14924
rect 22636 14868 22684 14924
rect 22740 14868 22788 14924
rect 22844 14868 22892 14924
rect 22948 14868 22958 14924
rect 22258 13356 22958 14868
rect 22258 13300 22268 13356
rect 22324 13300 22372 13356
rect 22428 13300 22476 13356
rect 22532 13300 22580 13356
rect 22636 13300 22684 13356
rect 22740 13300 22788 13356
rect 22844 13300 22892 13356
rect 22948 13300 22958 13356
rect 22258 11788 22958 13300
rect 22258 11732 22268 11788
rect 22324 11732 22372 11788
rect 22428 11732 22476 11788
rect 22532 11732 22580 11788
rect 22636 11732 22684 11788
rect 22740 11732 22788 11788
rect 22844 11732 22892 11788
rect 22948 11732 22958 11788
rect 22258 10220 22958 11732
rect 22258 10164 22268 10220
rect 22324 10164 22372 10220
rect 22428 10164 22476 10220
rect 22532 10164 22580 10220
rect 22636 10164 22684 10220
rect 22740 10164 22788 10220
rect 22844 10164 22892 10220
rect 22948 10164 22958 10220
rect 22258 8652 22958 10164
rect 22258 8596 22268 8652
rect 22324 8596 22372 8652
rect 22428 8596 22476 8652
rect 22532 8596 22580 8652
rect 22636 8596 22684 8652
rect 22740 8596 22788 8652
rect 22844 8596 22892 8652
rect 22948 8596 22958 8652
rect 22258 7084 22958 8596
rect 22258 7028 22268 7084
rect 22324 7028 22372 7084
rect 22428 7028 22476 7084
rect 22532 7028 22580 7084
rect 22636 7028 22684 7084
rect 22740 7028 22788 7084
rect 22844 7028 22892 7084
rect 22948 7028 22958 7084
rect 22258 5516 22958 7028
rect 22258 5460 22268 5516
rect 22324 5460 22372 5516
rect 22428 5460 22476 5516
rect 22532 5460 22580 5516
rect 22636 5460 22684 5516
rect 22740 5460 22788 5516
rect 22844 5460 22892 5516
rect 22948 5460 22958 5516
rect 22258 3948 22958 5460
rect 22258 3892 22268 3948
rect 22324 3892 22372 3948
rect 22428 3892 22476 3948
rect 22532 3892 22580 3948
rect 22636 3892 22684 3948
rect 22740 3892 22788 3948
rect 22844 3892 22892 3948
rect 22948 3892 22958 3948
rect 22258 3076 22958 3892
rect 26758 56476 27458 56508
rect 26758 56420 26768 56476
rect 26824 56420 26872 56476
rect 26928 56420 26976 56476
rect 27032 56420 27080 56476
rect 27136 56420 27184 56476
rect 27240 56420 27288 56476
rect 27344 56420 27392 56476
rect 27448 56420 27458 56476
rect 26758 54908 27458 56420
rect 26758 54852 26768 54908
rect 26824 54852 26872 54908
rect 26928 54852 26976 54908
rect 27032 54852 27080 54908
rect 27136 54852 27184 54908
rect 27240 54852 27288 54908
rect 27344 54852 27392 54908
rect 27448 54852 27458 54908
rect 26758 53340 27458 54852
rect 26758 53284 26768 53340
rect 26824 53284 26872 53340
rect 26928 53284 26976 53340
rect 27032 53284 27080 53340
rect 27136 53284 27184 53340
rect 27240 53284 27288 53340
rect 27344 53284 27392 53340
rect 27448 53284 27458 53340
rect 26758 51772 27458 53284
rect 26758 51716 26768 51772
rect 26824 51716 26872 51772
rect 26928 51716 26976 51772
rect 27032 51716 27080 51772
rect 27136 51716 27184 51772
rect 27240 51716 27288 51772
rect 27344 51716 27392 51772
rect 27448 51716 27458 51772
rect 26758 50204 27458 51716
rect 26758 50148 26768 50204
rect 26824 50148 26872 50204
rect 26928 50148 26976 50204
rect 27032 50148 27080 50204
rect 27136 50148 27184 50204
rect 27240 50148 27288 50204
rect 27344 50148 27392 50204
rect 27448 50148 27458 50204
rect 26758 48636 27458 50148
rect 26758 48580 26768 48636
rect 26824 48580 26872 48636
rect 26928 48580 26976 48636
rect 27032 48580 27080 48636
rect 27136 48580 27184 48636
rect 27240 48580 27288 48636
rect 27344 48580 27392 48636
rect 27448 48580 27458 48636
rect 26758 47068 27458 48580
rect 26758 47012 26768 47068
rect 26824 47012 26872 47068
rect 26928 47012 26976 47068
rect 27032 47012 27080 47068
rect 27136 47012 27184 47068
rect 27240 47012 27288 47068
rect 27344 47012 27392 47068
rect 27448 47012 27458 47068
rect 26758 45500 27458 47012
rect 26758 45444 26768 45500
rect 26824 45444 26872 45500
rect 26928 45444 26976 45500
rect 27032 45444 27080 45500
rect 27136 45444 27184 45500
rect 27240 45444 27288 45500
rect 27344 45444 27392 45500
rect 27448 45444 27458 45500
rect 26758 43932 27458 45444
rect 26758 43876 26768 43932
rect 26824 43876 26872 43932
rect 26928 43876 26976 43932
rect 27032 43876 27080 43932
rect 27136 43876 27184 43932
rect 27240 43876 27288 43932
rect 27344 43876 27392 43932
rect 27448 43876 27458 43932
rect 26758 42364 27458 43876
rect 26758 42308 26768 42364
rect 26824 42308 26872 42364
rect 26928 42308 26976 42364
rect 27032 42308 27080 42364
rect 27136 42308 27184 42364
rect 27240 42308 27288 42364
rect 27344 42308 27392 42364
rect 27448 42308 27458 42364
rect 26758 40796 27458 42308
rect 26758 40740 26768 40796
rect 26824 40740 26872 40796
rect 26928 40740 26976 40796
rect 27032 40740 27080 40796
rect 27136 40740 27184 40796
rect 27240 40740 27288 40796
rect 27344 40740 27392 40796
rect 27448 40740 27458 40796
rect 26758 39228 27458 40740
rect 26758 39172 26768 39228
rect 26824 39172 26872 39228
rect 26928 39172 26976 39228
rect 27032 39172 27080 39228
rect 27136 39172 27184 39228
rect 27240 39172 27288 39228
rect 27344 39172 27392 39228
rect 27448 39172 27458 39228
rect 26758 37660 27458 39172
rect 26758 37604 26768 37660
rect 26824 37604 26872 37660
rect 26928 37604 26976 37660
rect 27032 37604 27080 37660
rect 27136 37604 27184 37660
rect 27240 37604 27288 37660
rect 27344 37604 27392 37660
rect 27448 37604 27458 37660
rect 26758 36092 27458 37604
rect 26758 36036 26768 36092
rect 26824 36036 26872 36092
rect 26928 36036 26976 36092
rect 27032 36036 27080 36092
rect 27136 36036 27184 36092
rect 27240 36036 27288 36092
rect 27344 36036 27392 36092
rect 27448 36036 27458 36092
rect 26758 34524 27458 36036
rect 26758 34468 26768 34524
rect 26824 34468 26872 34524
rect 26928 34468 26976 34524
rect 27032 34468 27080 34524
rect 27136 34468 27184 34524
rect 27240 34468 27288 34524
rect 27344 34468 27392 34524
rect 27448 34468 27458 34524
rect 26758 32956 27458 34468
rect 26758 32900 26768 32956
rect 26824 32900 26872 32956
rect 26928 32900 26976 32956
rect 27032 32900 27080 32956
rect 27136 32900 27184 32956
rect 27240 32900 27288 32956
rect 27344 32900 27392 32956
rect 27448 32900 27458 32956
rect 26758 31388 27458 32900
rect 26758 31332 26768 31388
rect 26824 31332 26872 31388
rect 26928 31332 26976 31388
rect 27032 31332 27080 31388
rect 27136 31332 27184 31388
rect 27240 31332 27288 31388
rect 27344 31332 27392 31388
rect 27448 31332 27458 31388
rect 26758 29820 27458 31332
rect 26758 29764 26768 29820
rect 26824 29764 26872 29820
rect 26928 29764 26976 29820
rect 27032 29764 27080 29820
rect 27136 29764 27184 29820
rect 27240 29764 27288 29820
rect 27344 29764 27392 29820
rect 27448 29764 27458 29820
rect 26758 28252 27458 29764
rect 26758 28196 26768 28252
rect 26824 28196 26872 28252
rect 26928 28196 26976 28252
rect 27032 28196 27080 28252
rect 27136 28196 27184 28252
rect 27240 28196 27288 28252
rect 27344 28196 27392 28252
rect 27448 28196 27458 28252
rect 26758 26684 27458 28196
rect 26758 26628 26768 26684
rect 26824 26628 26872 26684
rect 26928 26628 26976 26684
rect 27032 26628 27080 26684
rect 27136 26628 27184 26684
rect 27240 26628 27288 26684
rect 27344 26628 27392 26684
rect 27448 26628 27458 26684
rect 26758 25116 27458 26628
rect 26758 25060 26768 25116
rect 26824 25060 26872 25116
rect 26928 25060 26976 25116
rect 27032 25060 27080 25116
rect 27136 25060 27184 25116
rect 27240 25060 27288 25116
rect 27344 25060 27392 25116
rect 27448 25060 27458 25116
rect 26758 23548 27458 25060
rect 26758 23492 26768 23548
rect 26824 23492 26872 23548
rect 26928 23492 26976 23548
rect 27032 23492 27080 23548
rect 27136 23492 27184 23548
rect 27240 23492 27288 23548
rect 27344 23492 27392 23548
rect 27448 23492 27458 23548
rect 26758 21980 27458 23492
rect 26758 21924 26768 21980
rect 26824 21924 26872 21980
rect 26928 21924 26976 21980
rect 27032 21924 27080 21980
rect 27136 21924 27184 21980
rect 27240 21924 27288 21980
rect 27344 21924 27392 21980
rect 27448 21924 27458 21980
rect 26758 20412 27458 21924
rect 26758 20356 26768 20412
rect 26824 20356 26872 20412
rect 26928 20356 26976 20412
rect 27032 20356 27080 20412
rect 27136 20356 27184 20412
rect 27240 20356 27288 20412
rect 27344 20356 27392 20412
rect 27448 20356 27458 20412
rect 26758 18844 27458 20356
rect 26758 18788 26768 18844
rect 26824 18788 26872 18844
rect 26928 18788 26976 18844
rect 27032 18788 27080 18844
rect 27136 18788 27184 18844
rect 27240 18788 27288 18844
rect 27344 18788 27392 18844
rect 27448 18788 27458 18844
rect 26758 17276 27458 18788
rect 26758 17220 26768 17276
rect 26824 17220 26872 17276
rect 26928 17220 26976 17276
rect 27032 17220 27080 17276
rect 27136 17220 27184 17276
rect 27240 17220 27288 17276
rect 27344 17220 27392 17276
rect 27448 17220 27458 17276
rect 26758 15708 27458 17220
rect 26758 15652 26768 15708
rect 26824 15652 26872 15708
rect 26928 15652 26976 15708
rect 27032 15652 27080 15708
rect 27136 15652 27184 15708
rect 27240 15652 27288 15708
rect 27344 15652 27392 15708
rect 27448 15652 27458 15708
rect 26758 14140 27458 15652
rect 26758 14084 26768 14140
rect 26824 14084 26872 14140
rect 26928 14084 26976 14140
rect 27032 14084 27080 14140
rect 27136 14084 27184 14140
rect 27240 14084 27288 14140
rect 27344 14084 27392 14140
rect 27448 14084 27458 14140
rect 26758 12572 27458 14084
rect 26758 12516 26768 12572
rect 26824 12516 26872 12572
rect 26928 12516 26976 12572
rect 27032 12516 27080 12572
rect 27136 12516 27184 12572
rect 27240 12516 27288 12572
rect 27344 12516 27392 12572
rect 27448 12516 27458 12572
rect 26758 11004 27458 12516
rect 26758 10948 26768 11004
rect 26824 10948 26872 11004
rect 26928 10948 26976 11004
rect 27032 10948 27080 11004
rect 27136 10948 27184 11004
rect 27240 10948 27288 11004
rect 27344 10948 27392 11004
rect 27448 10948 27458 11004
rect 26758 9436 27458 10948
rect 26758 9380 26768 9436
rect 26824 9380 26872 9436
rect 26928 9380 26976 9436
rect 27032 9380 27080 9436
rect 27136 9380 27184 9436
rect 27240 9380 27288 9436
rect 27344 9380 27392 9436
rect 27448 9380 27458 9436
rect 26758 7868 27458 9380
rect 26758 7812 26768 7868
rect 26824 7812 26872 7868
rect 26928 7812 26976 7868
rect 27032 7812 27080 7868
rect 27136 7812 27184 7868
rect 27240 7812 27288 7868
rect 27344 7812 27392 7868
rect 27448 7812 27458 7868
rect 26758 6300 27458 7812
rect 26758 6244 26768 6300
rect 26824 6244 26872 6300
rect 26928 6244 26976 6300
rect 27032 6244 27080 6300
rect 27136 6244 27184 6300
rect 27240 6244 27288 6300
rect 27344 6244 27392 6300
rect 27448 6244 27458 6300
rect 26758 4732 27458 6244
rect 26758 4676 26768 4732
rect 26824 4676 26872 4732
rect 26928 4676 26976 4732
rect 27032 4676 27080 4732
rect 27136 4676 27184 4732
rect 27240 4676 27288 4732
rect 27344 4676 27392 4732
rect 27448 4676 27458 4732
rect 26758 3164 27458 4676
rect 26758 3108 26768 3164
rect 26824 3108 26872 3164
rect 26928 3108 26976 3164
rect 27032 3108 27080 3164
rect 27136 3108 27184 3164
rect 27240 3108 27288 3164
rect 27344 3108 27392 3164
rect 27448 3108 27458 3164
rect 26758 3076 27458 3108
rect 31258 55692 31958 56508
rect 31258 55636 31268 55692
rect 31324 55636 31372 55692
rect 31428 55636 31476 55692
rect 31532 55636 31580 55692
rect 31636 55636 31684 55692
rect 31740 55636 31788 55692
rect 31844 55636 31892 55692
rect 31948 55636 31958 55692
rect 31258 54124 31958 55636
rect 31258 54068 31268 54124
rect 31324 54068 31372 54124
rect 31428 54068 31476 54124
rect 31532 54068 31580 54124
rect 31636 54068 31684 54124
rect 31740 54068 31788 54124
rect 31844 54068 31892 54124
rect 31948 54068 31958 54124
rect 31258 52556 31958 54068
rect 31258 52500 31268 52556
rect 31324 52500 31372 52556
rect 31428 52500 31476 52556
rect 31532 52500 31580 52556
rect 31636 52500 31684 52556
rect 31740 52500 31788 52556
rect 31844 52500 31892 52556
rect 31948 52500 31958 52556
rect 31258 50988 31958 52500
rect 31258 50932 31268 50988
rect 31324 50932 31372 50988
rect 31428 50932 31476 50988
rect 31532 50932 31580 50988
rect 31636 50932 31684 50988
rect 31740 50932 31788 50988
rect 31844 50932 31892 50988
rect 31948 50932 31958 50988
rect 31258 49420 31958 50932
rect 31258 49364 31268 49420
rect 31324 49364 31372 49420
rect 31428 49364 31476 49420
rect 31532 49364 31580 49420
rect 31636 49364 31684 49420
rect 31740 49364 31788 49420
rect 31844 49364 31892 49420
rect 31948 49364 31958 49420
rect 31258 47852 31958 49364
rect 31258 47796 31268 47852
rect 31324 47796 31372 47852
rect 31428 47796 31476 47852
rect 31532 47796 31580 47852
rect 31636 47796 31684 47852
rect 31740 47796 31788 47852
rect 31844 47796 31892 47852
rect 31948 47796 31958 47852
rect 31258 46284 31958 47796
rect 31258 46228 31268 46284
rect 31324 46228 31372 46284
rect 31428 46228 31476 46284
rect 31532 46228 31580 46284
rect 31636 46228 31684 46284
rect 31740 46228 31788 46284
rect 31844 46228 31892 46284
rect 31948 46228 31958 46284
rect 31258 44716 31958 46228
rect 31258 44660 31268 44716
rect 31324 44660 31372 44716
rect 31428 44660 31476 44716
rect 31532 44660 31580 44716
rect 31636 44660 31684 44716
rect 31740 44660 31788 44716
rect 31844 44660 31892 44716
rect 31948 44660 31958 44716
rect 31258 43148 31958 44660
rect 31258 43092 31268 43148
rect 31324 43092 31372 43148
rect 31428 43092 31476 43148
rect 31532 43092 31580 43148
rect 31636 43092 31684 43148
rect 31740 43092 31788 43148
rect 31844 43092 31892 43148
rect 31948 43092 31958 43148
rect 31258 41580 31958 43092
rect 31258 41524 31268 41580
rect 31324 41524 31372 41580
rect 31428 41524 31476 41580
rect 31532 41524 31580 41580
rect 31636 41524 31684 41580
rect 31740 41524 31788 41580
rect 31844 41524 31892 41580
rect 31948 41524 31958 41580
rect 31258 40012 31958 41524
rect 31258 39956 31268 40012
rect 31324 39956 31372 40012
rect 31428 39956 31476 40012
rect 31532 39956 31580 40012
rect 31636 39956 31684 40012
rect 31740 39956 31788 40012
rect 31844 39956 31892 40012
rect 31948 39956 31958 40012
rect 31258 38444 31958 39956
rect 31258 38388 31268 38444
rect 31324 38388 31372 38444
rect 31428 38388 31476 38444
rect 31532 38388 31580 38444
rect 31636 38388 31684 38444
rect 31740 38388 31788 38444
rect 31844 38388 31892 38444
rect 31948 38388 31958 38444
rect 31258 36876 31958 38388
rect 31258 36820 31268 36876
rect 31324 36820 31372 36876
rect 31428 36820 31476 36876
rect 31532 36820 31580 36876
rect 31636 36820 31684 36876
rect 31740 36820 31788 36876
rect 31844 36820 31892 36876
rect 31948 36820 31958 36876
rect 31258 35308 31958 36820
rect 31258 35252 31268 35308
rect 31324 35252 31372 35308
rect 31428 35252 31476 35308
rect 31532 35252 31580 35308
rect 31636 35252 31684 35308
rect 31740 35252 31788 35308
rect 31844 35252 31892 35308
rect 31948 35252 31958 35308
rect 31258 33740 31958 35252
rect 31258 33684 31268 33740
rect 31324 33684 31372 33740
rect 31428 33684 31476 33740
rect 31532 33684 31580 33740
rect 31636 33684 31684 33740
rect 31740 33684 31788 33740
rect 31844 33684 31892 33740
rect 31948 33684 31958 33740
rect 31258 32172 31958 33684
rect 31258 32116 31268 32172
rect 31324 32116 31372 32172
rect 31428 32116 31476 32172
rect 31532 32116 31580 32172
rect 31636 32116 31684 32172
rect 31740 32116 31788 32172
rect 31844 32116 31892 32172
rect 31948 32116 31958 32172
rect 31258 30604 31958 32116
rect 31258 30548 31268 30604
rect 31324 30548 31372 30604
rect 31428 30548 31476 30604
rect 31532 30548 31580 30604
rect 31636 30548 31684 30604
rect 31740 30548 31788 30604
rect 31844 30548 31892 30604
rect 31948 30548 31958 30604
rect 31258 29036 31958 30548
rect 31258 28980 31268 29036
rect 31324 28980 31372 29036
rect 31428 28980 31476 29036
rect 31532 28980 31580 29036
rect 31636 28980 31684 29036
rect 31740 28980 31788 29036
rect 31844 28980 31892 29036
rect 31948 28980 31958 29036
rect 31258 27468 31958 28980
rect 31258 27412 31268 27468
rect 31324 27412 31372 27468
rect 31428 27412 31476 27468
rect 31532 27412 31580 27468
rect 31636 27412 31684 27468
rect 31740 27412 31788 27468
rect 31844 27412 31892 27468
rect 31948 27412 31958 27468
rect 31258 25900 31958 27412
rect 31258 25844 31268 25900
rect 31324 25844 31372 25900
rect 31428 25844 31476 25900
rect 31532 25844 31580 25900
rect 31636 25844 31684 25900
rect 31740 25844 31788 25900
rect 31844 25844 31892 25900
rect 31948 25844 31958 25900
rect 31258 24332 31958 25844
rect 31258 24276 31268 24332
rect 31324 24276 31372 24332
rect 31428 24276 31476 24332
rect 31532 24276 31580 24332
rect 31636 24276 31684 24332
rect 31740 24276 31788 24332
rect 31844 24276 31892 24332
rect 31948 24276 31958 24332
rect 31258 22764 31958 24276
rect 31258 22708 31268 22764
rect 31324 22708 31372 22764
rect 31428 22708 31476 22764
rect 31532 22708 31580 22764
rect 31636 22708 31684 22764
rect 31740 22708 31788 22764
rect 31844 22708 31892 22764
rect 31948 22708 31958 22764
rect 31258 21196 31958 22708
rect 31258 21140 31268 21196
rect 31324 21140 31372 21196
rect 31428 21140 31476 21196
rect 31532 21140 31580 21196
rect 31636 21140 31684 21196
rect 31740 21140 31788 21196
rect 31844 21140 31892 21196
rect 31948 21140 31958 21196
rect 31258 19628 31958 21140
rect 31258 19572 31268 19628
rect 31324 19572 31372 19628
rect 31428 19572 31476 19628
rect 31532 19572 31580 19628
rect 31636 19572 31684 19628
rect 31740 19572 31788 19628
rect 31844 19572 31892 19628
rect 31948 19572 31958 19628
rect 31258 18060 31958 19572
rect 31258 18004 31268 18060
rect 31324 18004 31372 18060
rect 31428 18004 31476 18060
rect 31532 18004 31580 18060
rect 31636 18004 31684 18060
rect 31740 18004 31788 18060
rect 31844 18004 31892 18060
rect 31948 18004 31958 18060
rect 31258 16492 31958 18004
rect 31258 16436 31268 16492
rect 31324 16436 31372 16492
rect 31428 16436 31476 16492
rect 31532 16436 31580 16492
rect 31636 16436 31684 16492
rect 31740 16436 31788 16492
rect 31844 16436 31892 16492
rect 31948 16436 31958 16492
rect 31258 14924 31958 16436
rect 31258 14868 31268 14924
rect 31324 14868 31372 14924
rect 31428 14868 31476 14924
rect 31532 14868 31580 14924
rect 31636 14868 31684 14924
rect 31740 14868 31788 14924
rect 31844 14868 31892 14924
rect 31948 14868 31958 14924
rect 31258 13356 31958 14868
rect 31258 13300 31268 13356
rect 31324 13300 31372 13356
rect 31428 13300 31476 13356
rect 31532 13300 31580 13356
rect 31636 13300 31684 13356
rect 31740 13300 31788 13356
rect 31844 13300 31892 13356
rect 31948 13300 31958 13356
rect 31258 11788 31958 13300
rect 31258 11732 31268 11788
rect 31324 11732 31372 11788
rect 31428 11732 31476 11788
rect 31532 11732 31580 11788
rect 31636 11732 31684 11788
rect 31740 11732 31788 11788
rect 31844 11732 31892 11788
rect 31948 11732 31958 11788
rect 31258 10220 31958 11732
rect 31258 10164 31268 10220
rect 31324 10164 31372 10220
rect 31428 10164 31476 10220
rect 31532 10164 31580 10220
rect 31636 10164 31684 10220
rect 31740 10164 31788 10220
rect 31844 10164 31892 10220
rect 31948 10164 31958 10220
rect 31258 8652 31958 10164
rect 31258 8596 31268 8652
rect 31324 8596 31372 8652
rect 31428 8596 31476 8652
rect 31532 8596 31580 8652
rect 31636 8596 31684 8652
rect 31740 8596 31788 8652
rect 31844 8596 31892 8652
rect 31948 8596 31958 8652
rect 31258 7084 31958 8596
rect 31258 7028 31268 7084
rect 31324 7028 31372 7084
rect 31428 7028 31476 7084
rect 31532 7028 31580 7084
rect 31636 7028 31684 7084
rect 31740 7028 31788 7084
rect 31844 7028 31892 7084
rect 31948 7028 31958 7084
rect 31258 5516 31958 7028
rect 31258 5460 31268 5516
rect 31324 5460 31372 5516
rect 31428 5460 31476 5516
rect 31532 5460 31580 5516
rect 31636 5460 31684 5516
rect 31740 5460 31788 5516
rect 31844 5460 31892 5516
rect 31948 5460 31958 5516
rect 31258 3948 31958 5460
rect 31258 3892 31268 3948
rect 31324 3892 31372 3948
rect 31428 3892 31476 3948
rect 31532 3892 31580 3948
rect 31636 3892 31684 3948
rect 31740 3892 31788 3948
rect 31844 3892 31892 3948
rect 31948 3892 31958 3948
rect 31258 3076 31958 3892
rect 35758 56476 36458 56508
rect 35758 56420 35768 56476
rect 35824 56420 35872 56476
rect 35928 56420 35976 56476
rect 36032 56420 36080 56476
rect 36136 56420 36184 56476
rect 36240 56420 36288 56476
rect 36344 56420 36392 56476
rect 36448 56420 36458 56476
rect 35758 54908 36458 56420
rect 35758 54852 35768 54908
rect 35824 54852 35872 54908
rect 35928 54852 35976 54908
rect 36032 54852 36080 54908
rect 36136 54852 36184 54908
rect 36240 54852 36288 54908
rect 36344 54852 36392 54908
rect 36448 54852 36458 54908
rect 35758 53340 36458 54852
rect 35758 53284 35768 53340
rect 35824 53284 35872 53340
rect 35928 53284 35976 53340
rect 36032 53284 36080 53340
rect 36136 53284 36184 53340
rect 36240 53284 36288 53340
rect 36344 53284 36392 53340
rect 36448 53284 36458 53340
rect 35758 51772 36458 53284
rect 35758 51716 35768 51772
rect 35824 51716 35872 51772
rect 35928 51716 35976 51772
rect 36032 51716 36080 51772
rect 36136 51716 36184 51772
rect 36240 51716 36288 51772
rect 36344 51716 36392 51772
rect 36448 51716 36458 51772
rect 35758 50204 36458 51716
rect 35758 50148 35768 50204
rect 35824 50148 35872 50204
rect 35928 50148 35976 50204
rect 36032 50148 36080 50204
rect 36136 50148 36184 50204
rect 36240 50148 36288 50204
rect 36344 50148 36392 50204
rect 36448 50148 36458 50204
rect 35758 48636 36458 50148
rect 35758 48580 35768 48636
rect 35824 48580 35872 48636
rect 35928 48580 35976 48636
rect 36032 48580 36080 48636
rect 36136 48580 36184 48636
rect 36240 48580 36288 48636
rect 36344 48580 36392 48636
rect 36448 48580 36458 48636
rect 35758 47068 36458 48580
rect 35758 47012 35768 47068
rect 35824 47012 35872 47068
rect 35928 47012 35976 47068
rect 36032 47012 36080 47068
rect 36136 47012 36184 47068
rect 36240 47012 36288 47068
rect 36344 47012 36392 47068
rect 36448 47012 36458 47068
rect 35758 45500 36458 47012
rect 35758 45444 35768 45500
rect 35824 45444 35872 45500
rect 35928 45444 35976 45500
rect 36032 45444 36080 45500
rect 36136 45444 36184 45500
rect 36240 45444 36288 45500
rect 36344 45444 36392 45500
rect 36448 45444 36458 45500
rect 35758 43932 36458 45444
rect 35758 43876 35768 43932
rect 35824 43876 35872 43932
rect 35928 43876 35976 43932
rect 36032 43876 36080 43932
rect 36136 43876 36184 43932
rect 36240 43876 36288 43932
rect 36344 43876 36392 43932
rect 36448 43876 36458 43932
rect 35758 42364 36458 43876
rect 35758 42308 35768 42364
rect 35824 42308 35872 42364
rect 35928 42308 35976 42364
rect 36032 42308 36080 42364
rect 36136 42308 36184 42364
rect 36240 42308 36288 42364
rect 36344 42308 36392 42364
rect 36448 42308 36458 42364
rect 35758 40796 36458 42308
rect 35758 40740 35768 40796
rect 35824 40740 35872 40796
rect 35928 40740 35976 40796
rect 36032 40740 36080 40796
rect 36136 40740 36184 40796
rect 36240 40740 36288 40796
rect 36344 40740 36392 40796
rect 36448 40740 36458 40796
rect 35758 39228 36458 40740
rect 35758 39172 35768 39228
rect 35824 39172 35872 39228
rect 35928 39172 35976 39228
rect 36032 39172 36080 39228
rect 36136 39172 36184 39228
rect 36240 39172 36288 39228
rect 36344 39172 36392 39228
rect 36448 39172 36458 39228
rect 35758 37660 36458 39172
rect 35758 37604 35768 37660
rect 35824 37604 35872 37660
rect 35928 37604 35976 37660
rect 36032 37604 36080 37660
rect 36136 37604 36184 37660
rect 36240 37604 36288 37660
rect 36344 37604 36392 37660
rect 36448 37604 36458 37660
rect 35758 36092 36458 37604
rect 35758 36036 35768 36092
rect 35824 36036 35872 36092
rect 35928 36036 35976 36092
rect 36032 36036 36080 36092
rect 36136 36036 36184 36092
rect 36240 36036 36288 36092
rect 36344 36036 36392 36092
rect 36448 36036 36458 36092
rect 35758 34524 36458 36036
rect 35758 34468 35768 34524
rect 35824 34468 35872 34524
rect 35928 34468 35976 34524
rect 36032 34468 36080 34524
rect 36136 34468 36184 34524
rect 36240 34468 36288 34524
rect 36344 34468 36392 34524
rect 36448 34468 36458 34524
rect 35758 32956 36458 34468
rect 35758 32900 35768 32956
rect 35824 32900 35872 32956
rect 35928 32900 35976 32956
rect 36032 32900 36080 32956
rect 36136 32900 36184 32956
rect 36240 32900 36288 32956
rect 36344 32900 36392 32956
rect 36448 32900 36458 32956
rect 35758 31388 36458 32900
rect 35758 31332 35768 31388
rect 35824 31332 35872 31388
rect 35928 31332 35976 31388
rect 36032 31332 36080 31388
rect 36136 31332 36184 31388
rect 36240 31332 36288 31388
rect 36344 31332 36392 31388
rect 36448 31332 36458 31388
rect 35758 29820 36458 31332
rect 35758 29764 35768 29820
rect 35824 29764 35872 29820
rect 35928 29764 35976 29820
rect 36032 29764 36080 29820
rect 36136 29764 36184 29820
rect 36240 29764 36288 29820
rect 36344 29764 36392 29820
rect 36448 29764 36458 29820
rect 35758 28252 36458 29764
rect 35758 28196 35768 28252
rect 35824 28196 35872 28252
rect 35928 28196 35976 28252
rect 36032 28196 36080 28252
rect 36136 28196 36184 28252
rect 36240 28196 36288 28252
rect 36344 28196 36392 28252
rect 36448 28196 36458 28252
rect 35758 26684 36458 28196
rect 35758 26628 35768 26684
rect 35824 26628 35872 26684
rect 35928 26628 35976 26684
rect 36032 26628 36080 26684
rect 36136 26628 36184 26684
rect 36240 26628 36288 26684
rect 36344 26628 36392 26684
rect 36448 26628 36458 26684
rect 35758 25116 36458 26628
rect 35758 25060 35768 25116
rect 35824 25060 35872 25116
rect 35928 25060 35976 25116
rect 36032 25060 36080 25116
rect 36136 25060 36184 25116
rect 36240 25060 36288 25116
rect 36344 25060 36392 25116
rect 36448 25060 36458 25116
rect 35758 23548 36458 25060
rect 35758 23492 35768 23548
rect 35824 23492 35872 23548
rect 35928 23492 35976 23548
rect 36032 23492 36080 23548
rect 36136 23492 36184 23548
rect 36240 23492 36288 23548
rect 36344 23492 36392 23548
rect 36448 23492 36458 23548
rect 35758 21980 36458 23492
rect 35758 21924 35768 21980
rect 35824 21924 35872 21980
rect 35928 21924 35976 21980
rect 36032 21924 36080 21980
rect 36136 21924 36184 21980
rect 36240 21924 36288 21980
rect 36344 21924 36392 21980
rect 36448 21924 36458 21980
rect 35758 20412 36458 21924
rect 35758 20356 35768 20412
rect 35824 20356 35872 20412
rect 35928 20356 35976 20412
rect 36032 20356 36080 20412
rect 36136 20356 36184 20412
rect 36240 20356 36288 20412
rect 36344 20356 36392 20412
rect 36448 20356 36458 20412
rect 35758 18844 36458 20356
rect 35758 18788 35768 18844
rect 35824 18788 35872 18844
rect 35928 18788 35976 18844
rect 36032 18788 36080 18844
rect 36136 18788 36184 18844
rect 36240 18788 36288 18844
rect 36344 18788 36392 18844
rect 36448 18788 36458 18844
rect 35758 17276 36458 18788
rect 35758 17220 35768 17276
rect 35824 17220 35872 17276
rect 35928 17220 35976 17276
rect 36032 17220 36080 17276
rect 36136 17220 36184 17276
rect 36240 17220 36288 17276
rect 36344 17220 36392 17276
rect 36448 17220 36458 17276
rect 35758 15708 36458 17220
rect 35758 15652 35768 15708
rect 35824 15652 35872 15708
rect 35928 15652 35976 15708
rect 36032 15652 36080 15708
rect 36136 15652 36184 15708
rect 36240 15652 36288 15708
rect 36344 15652 36392 15708
rect 36448 15652 36458 15708
rect 35758 14140 36458 15652
rect 35758 14084 35768 14140
rect 35824 14084 35872 14140
rect 35928 14084 35976 14140
rect 36032 14084 36080 14140
rect 36136 14084 36184 14140
rect 36240 14084 36288 14140
rect 36344 14084 36392 14140
rect 36448 14084 36458 14140
rect 35758 12572 36458 14084
rect 35758 12516 35768 12572
rect 35824 12516 35872 12572
rect 35928 12516 35976 12572
rect 36032 12516 36080 12572
rect 36136 12516 36184 12572
rect 36240 12516 36288 12572
rect 36344 12516 36392 12572
rect 36448 12516 36458 12572
rect 35758 11004 36458 12516
rect 35758 10948 35768 11004
rect 35824 10948 35872 11004
rect 35928 10948 35976 11004
rect 36032 10948 36080 11004
rect 36136 10948 36184 11004
rect 36240 10948 36288 11004
rect 36344 10948 36392 11004
rect 36448 10948 36458 11004
rect 35758 9436 36458 10948
rect 35758 9380 35768 9436
rect 35824 9380 35872 9436
rect 35928 9380 35976 9436
rect 36032 9380 36080 9436
rect 36136 9380 36184 9436
rect 36240 9380 36288 9436
rect 36344 9380 36392 9436
rect 36448 9380 36458 9436
rect 35758 7868 36458 9380
rect 35758 7812 35768 7868
rect 35824 7812 35872 7868
rect 35928 7812 35976 7868
rect 36032 7812 36080 7868
rect 36136 7812 36184 7868
rect 36240 7812 36288 7868
rect 36344 7812 36392 7868
rect 36448 7812 36458 7868
rect 35758 6300 36458 7812
rect 35758 6244 35768 6300
rect 35824 6244 35872 6300
rect 35928 6244 35976 6300
rect 36032 6244 36080 6300
rect 36136 6244 36184 6300
rect 36240 6244 36288 6300
rect 36344 6244 36392 6300
rect 36448 6244 36458 6300
rect 35758 4732 36458 6244
rect 35758 4676 35768 4732
rect 35824 4676 35872 4732
rect 35928 4676 35976 4732
rect 36032 4676 36080 4732
rect 36136 4676 36184 4732
rect 36240 4676 36288 4732
rect 36344 4676 36392 4732
rect 36448 4676 36458 4732
rect 35758 3164 36458 4676
rect 35758 3108 35768 3164
rect 35824 3108 35872 3164
rect 35928 3108 35976 3164
rect 36032 3108 36080 3164
rect 36136 3108 36184 3164
rect 36240 3108 36288 3164
rect 36344 3108 36392 3164
rect 36448 3108 36458 3164
rect 35758 3076 36458 3108
rect 40258 55692 40958 56508
rect 40258 55636 40268 55692
rect 40324 55636 40372 55692
rect 40428 55636 40476 55692
rect 40532 55636 40580 55692
rect 40636 55636 40684 55692
rect 40740 55636 40788 55692
rect 40844 55636 40892 55692
rect 40948 55636 40958 55692
rect 40258 54124 40958 55636
rect 40258 54068 40268 54124
rect 40324 54068 40372 54124
rect 40428 54068 40476 54124
rect 40532 54068 40580 54124
rect 40636 54068 40684 54124
rect 40740 54068 40788 54124
rect 40844 54068 40892 54124
rect 40948 54068 40958 54124
rect 40258 52556 40958 54068
rect 40258 52500 40268 52556
rect 40324 52500 40372 52556
rect 40428 52500 40476 52556
rect 40532 52500 40580 52556
rect 40636 52500 40684 52556
rect 40740 52500 40788 52556
rect 40844 52500 40892 52556
rect 40948 52500 40958 52556
rect 40258 50988 40958 52500
rect 40258 50932 40268 50988
rect 40324 50932 40372 50988
rect 40428 50932 40476 50988
rect 40532 50932 40580 50988
rect 40636 50932 40684 50988
rect 40740 50932 40788 50988
rect 40844 50932 40892 50988
rect 40948 50932 40958 50988
rect 40258 49420 40958 50932
rect 40258 49364 40268 49420
rect 40324 49364 40372 49420
rect 40428 49364 40476 49420
rect 40532 49364 40580 49420
rect 40636 49364 40684 49420
rect 40740 49364 40788 49420
rect 40844 49364 40892 49420
rect 40948 49364 40958 49420
rect 40258 47852 40958 49364
rect 40258 47796 40268 47852
rect 40324 47796 40372 47852
rect 40428 47796 40476 47852
rect 40532 47796 40580 47852
rect 40636 47796 40684 47852
rect 40740 47796 40788 47852
rect 40844 47796 40892 47852
rect 40948 47796 40958 47852
rect 40258 46284 40958 47796
rect 40258 46228 40268 46284
rect 40324 46228 40372 46284
rect 40428 46228 40476 46284
rect 40532 46228 40580 46284
rect 40636 46228 40684 46284
rect 40740 46228 40788 46284
rect 40844 46228 40892 46284
rect 40948 46228 40958 46284
rect 40258 44716 40958 46228
rect 40258 44660 40268 44716
rect 40324 44660 40372 44716
rect 40428 44660 40476 44716
rect 40532 44660 40580 44716
rect 40636 44660 40684 44716
rect 40740 44660 40788 44716
rect 40844 44660 40892 44716
rect 40948 44660 40958 44716
rect 40258 43148 40958 44660
rect 40258 43092 40268 43148
rect 40324 43092 40372 43148
rect 40428 43092 40476 43148
rect 40532 43092 40580 43148
rect 40636 43092 40684 43148
rect 40740 43092 40788 43148
rect 40844 43092 40892 43148
rect 40948 43092 40958 43148
rect 40258 41580 40958 43092
rect 40258 41524 40268 41580
rect 40324 41524 40372 41580
rect 40428 41524 40476 41580
rect 40532 41524 40580 41580
rect 40636 41524 40684 41580
rect 40740 41524 40788 41580
rect 40844 41524 40892 41580
rect 40948 41524 40958 41580
rect 40258 40012 40958 41524
rect 40258 39956 40268 40012
rect 40324 39956 40372 40012
rect 40428 39956 40476 40012
rect 40532 39956 40580 40012
rect 40636 39956 40684 40012
rect 40740 39956 40788 40012
rect 40844 39956 40892 40012
rect 40948 39956 40958 40012
rect 40258 38444 40958 39956
rect 40258 38388 40268 38444
rect 40324 38388 40372 38444
rect 40428 38388 40476 38444
rect 40532 38388 40580 38444
rect 40636 38388 40684 38444
rect 40740 38388 40788 38444
rect 40844 38388 40892 38444
rect 40948 38388 40958 38444
rect 40258 36876 40958 38388
rect 40258 36820 40268 36876
rect 40324 36820 40372 36876
rect 40428 36820 40476 36876
rect 40532 36820 40580 36876
rect 40636 36820 40684 36876
rect 40740 36820 40788 36876
rect 40844 36820 40892 36876
rect 40948 36820 40958 36876
rect 40258 35308 40958 36820
rect 40258 35252 40268 35308
rect 40324 35252 40372 35308
rect 40428 35252 40476 35308
rect 40532 35252 40580 35308
rect 40636 35252 40684 35308
rect 40740 35252 40788 35308
rect 40844 35252 40892 35308
rect 40948 35252 40958 35308
rect 40258 33740 40958 35252
rect 40258 33684 40268 33740
rect 40324 33684 40372 33740
rect 40428 33684 40476 33740
rect 40532 33684 40580 33740
rect 40636 33684 40684 33740
rect 40740 33684 40788 33740
rect 40844 33684 40892 33740
rect 40948 33684 40958 33740
rect 40258 32172 40958 33684
rect 40258 32116 40268 32172
rect 40324 32116 40372 32172
rect 40428 32116 40476 32172
rect 40532 32116 40580 32172
rect 40636 32116 40684 32172
rect 40740 32116 40788 32172
rect 40844 32116 40892 32172
rect 40948 32116 40958 32172
rect 40258 30604 40958 32116
rect 40258 30548 40268 30604
rect 40324 30548 40372 30604
rect 40428 30548 40476 30604
rect 40532 30548 40580 30604
rect 40636 30548 40684 30604
rect 40740 30548 40788 30604
rect 40844 30548 40892 30604
rect 40948 30548 40958 30604
rect 40258 29036 40958 30548
rect 40258 28980 40268 29036
rect 40324 28980 40372 29036
rect 40428 28980 40476 29036
rect 40532 28980 40580 29036
rect 40636 28980 40684 29036
rect 40740 28980 40788 29036
rect 40844 28980 40892 29036
rect 40948 28980 40958 29036
rect 40258 27468 40958 28980
rect 40258 27412 40268 27468
rect 40324 27412 40372 27468
rect 40428 27412 40476 27468
rect 40532 27412 40580 27468
rect 40636 27412 40684 27468
rect 40740 27412 40788 27468
rect 40844 27412 40892 27468
rect 40948 27412 40958 27468
rect 40258 25900 40958 27412
rect 40258 25844 40268 25900
rect 40324 25844 40372 25900
rect 40428 25844 40476 25900
rect 40532 25844 40580 25900
rect 40636 25844 40684 25900
rect 40740 25844 40788 25900
rect 40844 25844 40892 25900
rect 40948 25844 40958 25900
rect 40258 24332 40958 25844
rect 40258 24276 40268 24332
rect 40324 24276 40372 24332
rect 40428 24276 40476 24332
rect 40532 24276 40580 24332
rect 40636 24276 40684 24332
rect 40740 24276 40788 24332
rect 40844 24276 40892 24332
rect 40948 24276 40958 24332
rect 40258 22764 40958 24276
rect 40258 22708 40268 22764
rect 40324 22708 40372 22764
rect 40428 22708 40476 22764
rect 40532 22708 40580 22764
rect 40636 22708 40684 22764
rect 40740 22708 40788 22764
rect 40844 22708 40892 22764
rect 40948 22708 40958 22764
rect 40258 21196 40958 22708
rect 40258 21140 40268 21196
rect 40324 21140 40372 21196
rect 40428 21140 40476 21196
rect 40532 21140 40580 21196
rect 40636 21140 40684 21196
rect 40740 21140 40788 21196
rect 40844 21140 40892 21196
rect 40948 21140 40958 21196
rect 40258 19628 40958 21140
rect 40258 19572 40268 19628
rect 40324 19572 40372 19628
rect 40428 19572 40476 19628
rect 40532 19572 40580 19628
rect 40636 19572 40684 19628
rect 40740 19572 40788 19628
rect 40844 19572 40892 19628
rect 40948 19572 40958 19628
rect 40258 18060 40958 19572
rect 40258 18004 40268 18060
rect 40324 18004 40372 18060
rect 40428 18004 40476 18060
rect 40532 18004 40580 18060
rect 40636 18004 40684 18060
rect 40740 18004 40788 18060
rect 40844 18004 40892 18060
rect 40948 18004 40958 18060
rect 40258 16492 40958 18004
rect 40258 16436 40268 16492
rect 40324 16436 40372 16492
rect 40428 16436 40476 16492
rect 40532 16436 40580 16492
rect 40636 16436 40684 16492
rect 40740 16436 40788 16492
rect 40844 16436 40892 16492
rect 40948 16436 40958 16492
rect 40258 14924 40958 16436
rect 40258 14868 40268 14924
rect 40324 14868 40372 14924
rect 40428 14868 40476 14924
rect 40532 14868 40580 14924
rect 40636 14868 40684 14924
rect 40740 14868 40788 14924
rect 40844 14868 40892 14924
rect 40948 14868 40958 14924
rect 40258 13356 40958 14868
rect 40258 13300 40268 13356
rect 40324 13300 40372 13356
rect 40428 13300 40476 13356
rect 40532 13300 40580 13356
rect 40636 13300 40684 13356
rect 40740 13300 40788 13356
rect 40844 13300 40892 13356
rect 40948 13300 40958 13356
rect 40258 11788 40958 13300
rect 40258 11732 40268 11788
rect 40324 11732 40372 11788
rect 40428 11732 40476 11788
rect 40532 11732 40580 11788
rect 40636 11732 40684 11788
rect 40740 11732 40788 11788
rect 40844 11732 40892 11788
rect 40948 11732 40958 11788
rect 40258 10220 40958 11732
rect 40258 10164 40268 10220
rect 40324 10164 40372 10220
rect 40428 10164 40476 10220
rect 40532 10164 40580 10220
rect 40636 10164 40684 10220
rect 40740 10164 40788 10220
rect 40844 10164 40892 10220
rect 40948 10164 40958 10220
rect 40258 8652 40958 10164
rect 40258 8596 40268 8652
rect 40324 8596 40372 8652
rect 40428 8596 40476 8652
rect 40532 8596 40580 8652
rect 40636 8596 40684 8652
rect 40740 8596 40788 8652
rect 40844 8596 40892 8652
rect 40948 8596 40958 8652
rect 40258 7084 40958 8596
rect 40258 7028 40268 7084
rect 40324 7028 40372 7084
rect 40428 7028 40476 7084
rect 40532 7028 40580 7084
rect 40636 7028 40684 7084
rect 40740 7028 40788 7084
rect 40844 7028 40892 7084
rect 40948 7028 40958 7084
rect 40258 5516 40958 7028
rect 40258 5460 40268 5516
rect 40324 5460 40372 5516
rect 40428 5460 40476 5516
rect 40532 5460 40580 5516
rect 40636 5460 40684 5516
rect 40740 5460 40788 5516
rect 40844 5460 40892 5516
rect 40948 5460 40958 5516
rect 40258 3948 40958 5460
rect 40258 3892 40268 3948
rect 40324 3892 40372 3948
rect 40428 3892 40476 3948
rect 40532 3892 40580 3948
rect 40636 3892 40684 3948
rect 40740 3892 40788 3948
rect 40844 3892 40892 3948
rect 40948 3892 40958 3948
rect 40258 3076 40958 3892
rect 44758 56476 45458 56508
rect 44758 56420 44768 56476
rect 44824 56420 44872 56476
rect 44928 56420 44976 56476
rect 45032 56420 45080 56476
rect 45136 56420 45184 56476
rect 45240 56420 45288 56476
rect 45344 56420 45392 56476
rect 45448 56420 45458 56476
rect 44758 54908 45458 56420
rect 44758 54852 44768 54908
rect 44824 54852 44872 54908
rect 44928 54852 44976 54908
rect 45032 54852 45080 54908
rect 45136 54852 45184 54908
rect 45240 54852 45288 54908
rect 45344 54852 45392 54908
rect 45448 54852 45458 54908
rect 44758 53340 45458 54852
rect 44758 53284 44768 53340
rect 44824 53284 44872 53340
rect 44928 53284 44976 53340
rect 45032 53284 45080 53340
rect 45136 53284 45184 53340
rect 45240 53284 45288 53340
rect 45344 53284 45392 53340
rect 45448 53284 45458 53340
rect 44758 51772 45458 53284
rect 44758 51716 44768 51772
rect 44824 51716 44872 51772
rect 44928 51716 44976 51772
rect 45032 51716 45080 51772
rect 45136 51716 45184 51772
rect 45240 51716 45288 51772
rect 45344 51716 45392 51772
rect 45448 51716 45458 51772
rect 44758 50204 45458 51716
rect 44758 50148 44768 50204
rect 44824 50148 44872 50204
rect 44928 50148 44976 50204
rect 45032 50148 45080 50204
rect 45136 50148 45184 50204
rect 45240 50148 45288 50204
rect 45344 50148 45392 50204
rect 45448 50148 45458 50204
rect 44758 48636 45458 50148
rect 44758 48580 44768 48636
rect 44824 48580 44872 48636
rect 44928 48580 44976 48636
rect 45032 48580 45080 48636
rect 45136 48580 45184 48636
rect 45240 48580 45288 48636
rect 45344 48580 45392 48636
rect 45448 48580 45458 48636
rect 44758 47068 45458 48580
rect 44758 47012 44768 47068
rect 44824 47012 44872 47068
rect 44928 47012 44976 47068
rect 45032 47012 45080 47068
rect 45136 47012 45184 47068
rect 45240 47012 45288 47068
rect 45344 47012 45392 47068
rect 45448 47012 45458 47068
rect 44758 45500 45458 47012
rect 44758 45444 44768 45500
rect 44824 45444 44872 45500
rect 44928 45444 44976 45500
rect 45032 45444 45080 45500
rect 45136 45444 45184 45500
rect 45240 45444 45288 45500
rect 45344 45444 45392 45500
rect 45448 45444 45458 45500
rect 44758 43932 45458 45444
rect 44758 43876 44768 43932
rect 44824 43876 44872 43932
rect 44928 43876 44976 43932
rect 45032 43876 45080 43932
rect 45136 43876 45184 43932
rect 45240 43876 45288 43932
rect 45344 43876 45392 43932
rect 45448 43876 45458 43932
rect 44758 42364 45458 43876
rect 44758 42308 44768 42364
rect 44824 42308 44872 42364
rect 44928 42308 44976 42364
rect 45032 42308 45080 42364
rect 45136 42308 45184 42364
rect 45240 42308 45288 42364
rect 45344 42308 45392 42364
rect 45448 42308 45458 42364
rect 44758 40796 45458 42308
rect 49258 55692 49958 56508
rect 49258 55636 49268 55692
rect 49324 55636 49372 55692
rect 49428 55636 49476 55692
rect 49532 55636 49580 55692
rect 49636 55636 49684 55692
rect 49740 55636 49788 55692
rect 49844 55636 49892 55692
rect 49948 55636 49958 55692
rect 49258 54124 49958 55636
rect 49258 54068 49268 54124
rect 49324 54068 49372 54124
rect 49428 54068 49476 54124
rect 49532 54068 49580 54124
rect 49636 54068 49684 54124
rect 49740 54068 49788 54124
rect 49844 54068 49892 54124
rect 49948 54068 49958 54124
rect 49258 52556 49958 54068
rect 49258 52500 49268 52556
rect 49324 52500 49372 52556
rect 49428 52500 49476 52556
rect 49532 52500 49580 52556
rect 49636 52500 49684 52556
rect 49740 52500 49788 52556
rect 49844 52500 49892 52556
rect 49948 52500 49958 52556
rect 49258 50988 49958 52500
rect 49258 50932 49268 50988
rect 49324 50932 49372 50988
rect 49428 50932 49476 50988
rect 49532 50932 49580 50988
rect 49636 50932 49684 50988
rect 49740 50932 49788 50988
rect 49844 50932 49892 50988
rect 49948 50932 49958 50988
rect 49258 49420 49958 50932
rect 49258 49364 49268 49420
rect 49324 49364 49372 49420
rect 49428 49364 49476 49420
rect 49532 49364 49580 49420
rect 49636 49364 49684 49420
rect 49740 49364 49788 49420
rect 49844 49364 49892 49420
rect 49948 49364 49958 49420
rect 49258 47852 49958 49364
rect 49258 47796 49268 47852
rect 49324 47796 49372 47852
rect 49428 47796 49476 47852
rect 49532 47796 49580 47852
rect 49636 47796 49684 47852
rect 49740 47796 49788 47852
rect 49844 47796 49892 47852
rect 49948 47796 49958 47852
rect 49258 46284 49958 47796
rect 49258 46228 49268 46284
rect 49324 46228 49372 46284
rect 49428 46228 49476 46284
rect 49532 46228 49580 46284
rect 49636 46228 49684 46284
rect 49740 46228 49788 46284
rect 49844 46228 49892 46284
rect 49948 46228 49958 46284
rect 49258 44716 49958 46228
rect 49258 44660 49268 44716
rect 49324 44660 49372 44716
rect 49428 44660 49476 44716
rect 49532 44660 49580 44716
rect 49636 44660 49684 44716
rect 49740 44660 49788 44716
rect 49844 44660 49892 44716
rect 49948 44660 49958 44716
rect 49258 43148 49958 44660
rect 49258 43092 49268 43148
rect 49324 43092 49372 43148
rect 49428 43092 49476 43148
rect 49532 43092 49580 43148
rect 49636 43092 49684 43148
rect 49740 43092 49788 43148
rect 49844 43092 49892 43148
rect 49948 43092 49958 43148
rect 44758 40740 44768 40796
rect 44824 40740 44872 40796
rect 44928 40740 44976 40796
rect 45032 40740 45080 40796
rect 45136 40740 45184 40796
rect 45240 40740 45288 40796
rect 45344 40740 45392 40796
rect 45448 40740 45458 40796
rect 44758 39228 45458 40740
rect 49084 42084 49140 42094
rect 49084 40404 49140 42028
rect 49084 40338 49140 40348
rect 49258 41580 49958 43092
rect 49258 41524 49268 41580
rect 49324 41524 49372 41580
rect 49428 41524 49476 41580
rect 49532 41524 49580 41580
rect 49636 41524 49684 41580
rect 49740 41524 49788 41580
rect 49844 41524 49892 41580
rect 49948 41524 49958 41580
rect 44758 39172 44768 39228
rect 44824 39172 44872 39228
rect 44928 39172 44976 39228
rect 45032 39172 45080 39228
rect 45136 39172 45184 39228
rect 45240 39172 45288 39228
rect 45344 39172 45392 39228
rect 45448 39172 45458 39228
rect 44758 37660 45458 39172
rect 44758 37604 44768 37660
rect 44824 37604 44872 37660
rect 44928 37604 44976 37660
rect 45032 37604 45080 37660
rect 45136 37604 45184 37660
rect 45240 37604 45288 37660
rect 45344 37604 45392 37660
rect 45448 37604 45458 37660
rect 44758 36092 45458 37604
rect 44758 36036 44768 36092
rect 44824 36036 44872 36092
rect 44928 36036 44976 36092
rect 45032 36036 45080 36092
rect 45136 36036 45184 36092
rect 45240 36036 45288 36092
rect 45344 36036 45392 36092
rect 45448 36036 45458 36092
rect 44758 34524 45458 36036
rect 44758 34468 44768 34524
rect 44824 34468 44872 34524
rect 44928 34468 44976 34524
rect 45032 34468 45080 34524
rect 45136 34468 45184 34524
rect 45240 34468 45288 34524
rect 45344 34468 45392 34524
rect 45448 34468 45458 34524
rect 44758 32956 45458 34468
rect 44758 32900 44768 32956
rect 44824 32900 44872 32956
rect 44928 32900 44976 32956
rect 45032 32900 45080 32956
rect 45136 32900 45184 32956
rect 45240 32900 45288 32956
rect 45344 32900 45392 32956
rect 45448 32900 45458 32956
rect 44758 31388 45458 32900
rect 44758 31332 44768 31388
rect 44824 31332 44872 31388
rect 44928 31332 44976 31388
rect 45032 31332 45080 31388
rect 45136 31332 45184 31388
rect 45240 31332 45288 31388
rect 45344 31332 45392 31388
rect 45448 31332 45458 31388
rect 44758 29820 45458 31332
rect 44758 29764 44768 29820
rect 44824 29764 44872 29820
rect 44928 29764 44976 29820
rect 45032 29764 45080 29820
rect 45136 29764 45184 29820
rect 45240 29764 45288 29820
rect 45344 29764 45392 29820
rect 45448 29764 45458 29820
rect 44758 28252 45458 29764
rect 44758 28196 44768 28252
rect 44824 28196 44872 28252
rect 44928 28196 44976 28252
rect 45032 28196 45080 28252
rect 45136 28196 45184 28252
rect 45240 28196 45288 28252
rect 45344 28196 45392 28252
rect 45448 28196 45458 28252
rect 44758 26684 45458 28196
rect 44758 26628 44768 26684
rect 44824 26628 44872 26684
rect 44928 26628 44976 26684
rect 45032 26628 45080 26684
rect 45136 26628 45184 26684
rect 45240 26628 45288 26684
rect 45344 26628 45392 26684
rect 45448 26628 45458 26684
rect 44758 25116 45458 26628
rect 44758 25060 44768 25116
rect 44824 25060 44872 25116
rect 44928 25060 44976 25116
rect 45032 25060 45080 25116
rect 45136 25060 45184 25116
rect 45240 25060 45288 25116
rect 45344 25060 45392 25116
rect 45448 25060 45458 25116
rect 44758 23548 45458 25060
rect 44758 23492 44768 23548
rect 44824 23492 44872 23548
rect 44928 23492 44976 23548
rect 45032 23492 45080 23548
rect 45136 23492 45184 23548
rect 45240 23492 45288 23548
rect 45344 23492 45392 23548
rect 45448 23492 45458 23548
rect 44758 21980 45458 23492
rect 44758 21924 44768 21980
rect 44824 21924 44872 21980
rect 44928 21924 44976 21980
rect 45032 21924 45080 21980
rect 45136 21924 45184 21980
rect 45240 21924 45288 21980
rect 45344 21924 45392 21980
rect 45448 21924 45458 21980
rect 44758 20412 45458 21924
rect 44758 20356 44768 20412
rect 44824 20356 44872 20412
rect 44928 20356 44976 20412
rect 45032 20356 45080 20412
rect 45136 20356 45184 20412
rect 45240 20356 45288 20412
rect 45344 20356 45392 20412
rect 45448 20356 45458 20412
rect 44758 18844 45458 20356
rect 44758 18788 44768 18844
rect 44824 18788 44872 18844
rect 44928 18788 44976 18844
rect 45032 18788 45080 18844
rect 45136 18788 45184 18844
rect 45240 18788 45288 18844
rect 45344 18788 45392 18844
rect 45448 18788 45458 18844
rect 44758 17276 45458 18788
rect 44758 17220 44768 17276
rect 44824 17220 44872 17276
rect 44928 17220 44976 17276
rect 45032 17220 45080 17276
rect 45136 17220 45184 17276
rect 45240 17220 45288 17276
rect 45344 17220 45392 17276
rect 45448 17220 45458 17276
rect 44758 15708 45458 17220
rect 44758 15652 44768 15708
rect 44824 15652 44872 15708
rect 44928 15652 44976 15708
rect 45032 15652 45080 15708
rect 45136 15652 45184 15708
rect 45240 15652 45288 15708
rect 45344 15652 45392 15708
rect 45448 15652 45458 15708
rect 44758 14140 45458 15652
rect 44758 14084 44768 14140
rect 44824 14084 44872 14140
rect 44928 14084 44976 14140
rect 45032 14084 45080 14140
rect 45136 14084 45184 14140
rect 45240 14084 45288 14140
rect 45344 14084 45392 14140
rect 45448 14084 45458 14140
rect 44758 12572 45458 14084
rect 44758 12516 44768 12572
rect 44824 12516 44872 12572
rect 44928 12516 44976 12572
rect 45032 12516 45080 12572
rect 45136 12516 45184 12572
rect 45240 12516 45288 12572
rect 45344 12516 45392 12572
rect 45448 12516 45458 12572
rect 44758 11004 45458 12516
rect 44758 10948 44768 11004
rect 44824 10948 44872 11004
rect 44928 10948 44976 11004
rect 45032 10948 45080 11004
rect 45136 10948 45184 11004
rect 45240 10948 45288 11004
rect 45344 10948 45392 11004
rect 45448 10948 45458 11004
rect 44758 9436 45458 10948
rect 44758 9380 44768 9436
rect 44824 9380 44872 9436
rect 44928 9380 44976 9436
rect 45032 9380 45080 9436
rect 45136 9380 45184 9436
rect 45240 9380 45288 9436
rect 45344 9380 45392 9436
rect 45448 9380 45458 9436
rect 44758 7868 45458 9380
rect 44758 7812 44768 7868
rect 44824 7812 44872 7868
rect 44928 7812 44976 7868
rect 45032 7812 45080 7868
rect 45136 7812 45184 7868
rect 45240 7812 45288 7868
rect 45344 7812 45392 7868
rect 45448 7812 45458 7868
rect 44758 6300 45458 7812
rect 49258 40012 49958 41524
rect 49258 39956 49268 40012
rect 49324 39956 49372 40012
rect 49428 39956 49476 40012
rect 49532 39956 49580 40012
rect 49636 39956 49684 40012
rect 49740 39956 49788 40012
rect 49844 39956 49892 40012
rect 49948 39956 49958 40012
rect 49258 38444 49958 39956
rect 49258 38388 49268 38444
rect 49324 38388 49372 38444
rect 49428 38388 49476 38444
rect 49532 38388 49580 38444
rect 49636 38388 49684 38444
rect 49740 38388 49788 38444
rect 49844 38388 49892 38444
rect 49948 38388 49958 38444
rect 49258 36876 49958 38388
rect 49258 36820 49268 36876
rect 49324 36820 49372 36876
rect 49428 36820 49476 36876
rect 49532 36820 49580 36876
rect 49636 36820 49684 36876
rect 49740 36820 49788 36876
rect 49844 36820 49892 36876
rect 49948 36820 49958 36876
rect 49258 35308 49958 36820
rect 49258 35252 49268 35308
rect 49324 35252 49372 35308
rect 49428 35252 49476 35308
rect 49532 35252 49580 35308
rect 49636 35252 49684 35308
rect 49740 35252 49788 35308
rect 49844 35252 49892 35308
rect 49948 35252 49958 35308
rect 49258 33740 49958 35252
rect 49258 33684 49268 33740
rect 49324 33684 49372 33740
rect 49428 33684 49476 33740
rect 49532 33684 49580 33740
rect 49636 33684 49684 33740
rect 49740 33684 49788 33740
rect 49844 33684 49892 33740
rect 49948 33684 49958 33740
rect 49258 32172 49958 33684
rect 49258 32116 49268 32172
rect 49324 32116 49372 32172
rect 49428 32116 49476 32172
rect 49532 32116 49580 32172
rect 49636 32116 49684 32172
rect 49740 32116 49788 32172
rect 49844 32116 49892 32172
rect 49948 32116 49958 32172
rect 49258 30604 49958 32116
rect 49258 30548 49268 30604
rect 49324 30548 49372 30604
rect 49428 30548 49476 30604
rect 49532 30548 49580 30604
rect 49636 30548 49684 30604
rect 49740 30548 49788 30604
rect 49844 30548 49892 30604
rect 49948 30548 49958 30604
rect 49258 29036 49958 30548
rect 49258 28980 49268 29036
rect 49324 28980 49372 29036
rect 49428 28980 49476 29036
rect 49532 28980 49580 29036
rect 49636 28980 49684 29036
rect 49740 28980 49788 29036
rect 49844 28980 49892 29036
rect 49948 28980 49958 29036
rect 49258 27468 49958 28980
rect 49258 27412 49268 27468
rect 49324 27412 49372 27468
rect 49428 27412 49476 27468
rect 49532 27412 49580 27468
rect 49636 27412 49684 27468
rect 49740 27412 49788 27468
rect 49844 27412 49892 27468
rect 49948 27412 49958 27468
rect 49258 25900 49958 27412
rect 49258 25844 49268 25900
rect 49324 25844 49372 25900
rect 49428 25844 49476 25900
rect 49532 25844 49580 25900
rect 49636 25844 49684 25900
rect 49740 25844 49788 25900
rect 49844 25844 49892 25900
rect 49948 25844 49958 25900
rect 49258 24332 49958 25844
rect 49258 24276 49268 24332
rect 49324 24276 49372 24332
rect 49428 24276 49476 24332
rect 49532 24276 49580 24332
rect 49636 24276 49684 24332
rect 49740 24276 49788 24332
rect 49844 24276 49892 24332
rect 49948 24276 49958 24332
rect 49258 22764 49958 24276
rect 49258 22708 49268 22764
rect 49324 22708 49372 22764
rect 49428 22708 49476 22764
rect 49532 22708 49580 22764
rect 49636 22708 49684 22764
rect 49740 22708 49788 22764
rect 49844 22708 49892 22764
rect 49948 22708 49958 22764
rect 49258 21196 49958 22708
rect 49258 21140 49268 21196
rect 49324 21140 49372 21196
rect 49428 21140 49476 21196
rect 49532 21140 49580 21196
rect 49636 21140 49684 21196
rect 49740 21140 49788 21196
rect 49844 21140 49892 21196
rect 49948 21140 49958 21196
rect 49258 19628 49958 21140
rect 49258 19572 49268 19628
rect 49324 19572 49372 19628
rect 49428 19572 49476 19628
rect 49532 19572 49580 19628
rect 49636 19572 49684 19628
rect 49740 19572 49788 19628
rect 49844 19572 49892 19628
rect 49948 19572 49958 19628
rect 49258 18060 49958 19572
rect 49258 18004 49268 18060
rect 49324 18004 49372 18060
rect 49428 18004 49476 18060
rect 49532 18004 49580 18060
rect 49636 18004 49684 18060
rect 49740 18004 49788 18060
rect 49844 18004 49892 18060
rect 49948 18004 49958 18060
rect 49258 16492 49958 18004
rect 49258 16436 49268 16492
rect 49324 16436 49372 16492
rect 49428 16436 49476 16492
rect 49532 16436 49580 16492
rect 49636 16436 49684 16492
rect 49740 16436 49788 16492
rect 49844 16436 49892 16492
rect 49948 16436 49958 16492
rect 49258 14924 49958 16436
rect 49258 14868 49268 14924
rect 49324 14868 49372 14924
rect 49428 14868 49476 14924
rect 49532 14868 49580 14924
rect 49636 14868 49684 14924
rect 49740 14868 49788 14924
rect 49844 14868 49892 14924
rect 49948 14868 49958 14924
rect 49258 13356 49958 14868
rect 49258 13300 49268 13356
rect 49324 13300 49372 13356
rect 49428 13300 49476 13356
rect 49532 13300 49580 13356
rect 49636 13300 49684 13356
rect 49740 13300 49788 13356
rect 49844 13300 49892 13356
rect 49948 13300 49958 13356
rect 49258 11788 49958 13300
rect 49258 11732 49268 11788
rect 49324 11732 49372 11788
rect 49428 11732 49476 11788
rect 49532 11732 49580 11788
rect 49636 11732 49684 11788
rect 49740 11732 49788 11788
rect 49844 11732 49892 11788
rect 49948 11732 49958 11788
rect 49258 10220 49958 11732
rect 49258 10164 49268 10220
rect 49324 10164 49372 10220
rect 49428 10164 49476 10220
rect 49532 10164 49580 10220
rect 49636 10164 49684 10220
rect 49740 10164 49788 10220
rect 49844 10164 49892 10220
rect 49948 10164 49958 10220
rect 49258 8652 49958 10164
rect 49258 8596 49268 8652
rect 49324 8596 49372 8652
rect 49428 8596 49476 8652
rect 49532 8596 49580 8652
rect 49636 8596 49684 8652
rect 49740 8596 49788 8652
rect 49844 8596 49892 8652
rect 49948 8596 49958 8652
rect 44758 6244 44768 6300
rect 44824 6244 44872 6300
rect 44928 6244 44976 6300
rect 45032 6244 45080 6300
rect 45136 6244 45184 6300
rect 45240 6244 45288 6300
rect 45344 6244 45392 6300
rect 45448 6244 45458 6300
rect 44758 4732 45458 6244
rect 48860 7700 48916 7710
rect 48860 6132 48916 7644
rect 48860 6066 48916 6076
rect 49258 7084 49958 8596
rect 49258 7028 49268 7084
rect 49324 7028 49372 7084
rect 49428 7028 49476 7084
rect 49532 7028 49580 7084
rect 49636 7028 49684 7084
rect 49740 7028 49788 7084
rect 49844 7028 49892 7084
rect 49948 7028 49958 7084
rect 44758 4676 44768 4732
rect 44824 4676 44872 4732
rect 44928 4676 44976 4732
rect 45032 4676 45080 4732
rect 45136 4676 45184 4732
rect 45240 4676 45288 4732
rect 45344 4676 45392 4732
rect 45448 4676 45458 4732
rect 44758 3164 45458 4676
rect 44758 3108 44768 3164
rect 44824 3108 44872 3164
rect 44928 3108 44976 3164
rect 45032 3108 45080 3164
rect 45136 3108 45184 3164
rect 45240 3108 45288 3164
rect 45344 3108 45392 3164
rect 45448 3108 45458 3164
rect 44758 3076 45458 3108
rect 49258 5516 49958 7028
rect 49258 5460 49268 5516
rect 49324 5460 49372 5516
rect 49428 5460 49476 5516
rect 49532 5460 49580 5516
rect 49636 5460 49684 5516
rect 49740 5460 49788 5516
rect 49844 5460 49892 5516
rect 49948 5460 49958 5516
rect 49258 3948 49958 5460
rect 49258 3892 49268 3948
rect 49324 3892 49372 3948
rect 49428 3892 49476 3948
rect 49532 3892 49580 3948
rect 49636 3892 49684 3948
rect 49740 3892 49788 3948
rect 49844 3892 49892 3948
rect 49948 3892 49958 3948
rect 49258 3076 49958 3892
rect 53758 56476 54458 56508
rect 53758 56420 53768 56476
rect 53824 56420 53872 56476
rect 53928 56420 53976 56476
rect 54032 56420 54080 56476
rect 54136 56420 54184 56476
rect 54240 56420 54288 56476
rect 54344 56420 54392 56476
rect 54448 56420 54458 56476
rect 53758 54908 54458 56420
rect 53758 54852 53768 54908
rect 53824 54852 53872 54908
rect 53928 54852 53976 54908
rect 54032 54852 54080 54908
rect 54136 54852 54184 54908
rect 54240 54852 54288 54908
rect 54344 54852 54392 54908
rect 54448 54852 54458 54908
rect 53758 53340 54458 54852
rect 53758 53284 53768 53340
rect 53824 53284 53872 53340
rect 53928 53284 53976 53340
rect 54032 53284 54080 53340
rect 54136 53284 54184 53340
rect 54240 53284 54288 53340
rect 54344 53284 54392 53340
rect 54448 53284 54458 53340
rect 53758 51772 54458 53284
rect 53758 51716 53768 51772
rect 53824 51716 53872 51772
rect 53928 51716 53976 51772
rect 54032 51716 54080 51772
rect 54136 51716 54184 51772
rect 54240 51716 54288 51772
rect 54344 51716 54392 51772
rect 54448 51716 54458 51772
rect 53758 50204 54458 51716
rect 53758 50148 53768 50204
rect 53824 50148 53872 50204
rect 53928 50148 53976 50204
rect 54032 50148 54080 50204
rect 54136 50148 54184 50204
rect 54240 50148 54288 50204
rect 54344 50148 54392 50204
rect 54448 50148 54458 50204
rect 53758 48636 54458 50148
rect 53758 48580 53768 48636
rect 53824 48580 53872 48636
rect 53928 48580 53976 48636
rect 54032 48580 54080 48636
rect 54136 48580 54184 48636
rect 54240 48580 54288 48636
rect 54344 48580 54392 48636
rect 54448 48580 54458 48636
rect 53758 47068 54458 48580
rect 53758 47012 53768 47068
rect 53824 47012 53872 47068
rect 53928 47012 53976 47068
rect 54032 47012 54080 47068
rect 54136 47012 54184 47068
rect 54240 47012 54288 47068
rect 54344 47012 54392 47068
rect 54448 47012 54458 47068
rect 53758 45500 54458 47012
rect 53758 45444 53768 45500
rect 53824 45444 53872 45500
rect 53928 45444 53976 45500
rect 54032 45444 54080 45500
rect 54136 45444 54184 45500
rect 54240 45444 54288 45500
rect 54344 45444 54392 45500
rect 54448 45444 54458 45500
rect 53758 43932 54458 45444
rect 53758 43876 53768 43932
rect 53824 43876 53872 43932
rect 53928 43876 53976 43932
rect 54032 43876 54080 43932
rect 54136 43876 54184 43932
rect 54240 43876 54288 43932
rect 54344 43876 54392 43932
rect 54448 43876 54458 43932
rect 53758 42364 54458 43876
rect 53758 42308 53768 42364
rect 53824 42308 53872 42364
rect 53928 42308 53976 42364
rect 54032 42308 54080 42364
rect 54136 42308 54184 42364
rect 54240 42308 54288 42364
rect 54344 42308 54392 42364
rect 54448 42308 54458 42364
rect 53758 40796 54458 42308
rect 53758 40740 53768 40796
rect 53824 40740 53872 40796
rect 53928 40740 53976 40796
rect 54032 40740 54080 40796
rect 54136 40740 54184 40796
rect 54240 40740 54288 40796
rect 54344 40740 54392 40796
rect 54448 40740 54458 40796
rect 53758 39228 54458 40740
rect 53758 39172 53768 39228
rect 53824 39172 53872 39228
rect 53928 39172 53976 39228
rect 54032 39172 54080 39228
rect 54136 39172 54184 39228
rect 54240 39172 54288 39228
rect 54344 39172 54392 39228
rect 54448 39172 54458 39228
rect 53758 37660 54458 39172
rect 53758 37604 53768 37660
rect 53824 37604 53872 37660
rect 53928 37604 53976 37660
rect 54032 37604 54080 37660
rect 54136 37604 54184 37660
rect 54240 37604 54288 37660
rect 54344 37604 54392 37660
rect 54448 37604 54458 37660
rect 53758 36092 54458 37604
rect 53758 36036 53768 36092
rect 53824 36036 53872 36092
rect 53928 36036 53976 36092
rect 54032 36036 54080 36092
rect 54136 36036 54184 36092
rect 54240 36036 54288 36092
rect 54344 36036 54392 36092
rect 54448 36036 54458 36092
rect 53758 34524 54458 36036
rect 53758 34468 53768 34524
rect 53824 34468 53872 34524
rect 53928 34468 53976 34524
rect 54032 34468 54080 34524
rect 54136 34468 54184 34524
rect 54240 34468 54288 34524
rect 54344 34468 54392 34524
rect 54448 34468 54458 34524
rect 53758 32956 54458 34468
rect 53758 32900 53768 32956
rect 53824 32900 53872 32956
rect 53928 32900 53976 32956
rect 54032 32900 54080 32956
rect 54136 32900 54184 32956
rect 54240 32900 54288 32956
rect 54344 32900 54392 32956
rect 54448 32900 54458 32956
rect 53758 31388 54458 32900
rect 53758 31332 53768 31388
rect 53824 31332 53872 31388
rect 53928 31332 53976 31388
rect 54032 31332 54080 31388
rect 54136 31332 54184 31388
rect 54240 31332 54288 31388
rect 54344 31332 54392 31388
rect 54448 31332 54458 31388
rect 53758 29820 54458 31332
rect 53758 29764 53768 29820
rect 53824 29764 53872 29820
rect 53928 29764 53976 29820
rect 54032 29764 54080 29820
rect 54136 29764 54184 29820
rect 54240 29764 54288 29820
rect 54344 29764 54392 29820
rect 54448 29764 54458 29820
rect 53758 28252 54458 29764
rect 53758 28196 53768 28252
rect 53824 28196 53872 28252
rect 53928 28196 53976 28252
rect 54032 28196 54080 28252
rect 54136 28196 54184 28252
rect 54240 28196 54288 28252
rect 54344 28196 54392 28252
rect 54448 28196 54458 28252
rect 53758 26684 54458 28196
rect 53758 26628 53768 26684
rect 53824 26628 53872 26684
rect 53928 26628 53976 26684
rect 54032 26628 54080 26684
rect 54136 26628 54184 26684
rect 54240 26628 54288 26684
rect 54344 26628 54392 26684
rect 54448 26628 54458 26684
rect 53758 25116 54458 26628
rect 53758 25060 53768 25116
rect 53824 25060 53872 25116
rect 53928 25060 53976 25116
rect 54032 25060 54080 25116
rect 54136 25060 54184 25116
rect 54240 25060 54288 25116
rect 54344 25060 54392 25116
rect 54448 25060 54458 25116
rect 53758 23548 54458 25060
rect 53758 23492 53768 23548
rect 53824 23492 53872 23548
rect 53928 23492 53976 23548
rect 54032 23492 54080 23548
rect 54136 23492 54184 23548
rect 54240 23492 54288 23548
rect 54344 23492 54392 23548
rect 54448 23492 54458 23548
rect 53758 21980 54458 23492
rect 53758 21924 53768 21980
rect 53824 21924 53872 21980
rect 53928 21924 53976 21980
rect 54032 21924 54080 21980
rect 54136 21924 54184 21980
rect 54240 21924 54288 21980
rect 54344 21924 54392 21980
rect 54448 21924 54458 21980
rect 53758 20412 54458 21924
rect 53758 20356 53768 20412
rect 53824 20356 53872 20412
rect 53928 20356 53976 20412
rect 54032 20356 54080 20412
rect 54136 20356 54184 20412
rect 54240 20356 54288 20412
rect 54344 20356 54392 20412
rect 54448 20356 54458 20412
rect 53758 18844 54458 20356
rect 53758 18788 53768 18844
rect 53824 18788 53872 18844
rect 53928 18788 53976 18844
rect 54032 18788 54080 18844
rect 54136 18788 54184 18844
rect 54240 18788 54288 18844
rect 54344 18788 54392 18844
rect 54448 18788 54458 18844
rect 53758 17276 54458 18788
rect 53758 17220 53768 17276
rect 53824 17220 53872 17276
rect 53928 17220 53976 17276
rect 54032 17220 54080 17276
rect 54136 17220 54184 17276
rect 54240 17220 54288 17276
rect 54344 17220 54392 17276
rect 54448 17220 54458 17276
rect 53758 15708 54458 17220
rect 53758 15652 53768 15708
rect 53824 15652 53872 15708
rect 53928 15652 53976 15708
rect 54032 15652 54080 15708
rect 54136 15652 54184 15708
rect 54240 15652 54288 15708
rect 54344 15652 54392 15708
rect 54448 15652 54458 15708
rect 53758 14140 54458 15652
rect 53758 14084 53768 14140
rect 53824 14084 53872 14140
rect 53928 14084 53976 14140
rect 54032 14084 54080 14140
rect 54136 14084 54184 14140
rect 54240 14084 54288 14140
rect 54344 14084 54392 14140
rect 54448 14084 54458 14140
rect 53758 12572 54458 14084
rect 53758 12516 53768 12572
rect 53824 12516 53872 12572
rect 53928 12516 53976 12572
rect 54032 12516 54080 12572
rect 54136 12516 54184 12572
rect 54240 12516 54288 12572
rect 54344 12516 54392 12572
rect 54448 12516 54458 12572
rect 53758 11004 54458 12516
rect 53758 10948 53768 11004
rect 53824 10948 53872 11004
rect 53928 10948 53976 11004
rect 54032 10948 54080 11004
rect 54136 10948 54184 11004
rect 54240 10948 54288 11004
rect 54344 10948 54392 11004
rect 54448 10948 54458 11004
rect 53758 9436 54458 10948
rect 53758 9380 53768 9436
rect 53824 9380 53872 9436
rect 53928 9380 53976 9436
rect 54032 9380 54080 9436
rect 54136 9380 54184 9436
rect 54240 9380 54288 9436
rect 54344 9380 54392 9436
rect 54448 9380 54458 9436
rect 53758 7868 54458 9380
rect 53758 7812 53768 7868
rect 53824 7812 53872 7868
rect 53928 7812 53976 7868
rect 54032 7812 54080 7868
rect 54136 7812 54184 7868
rect 54240 7812 54288 7868
rect 54344 7812 54392 7868
rect 54448 7812 54458 7868
rect 53758 6300 54458 7812
rect 53758 6244 53768 6300
rect 53824 6244 53872 6300
rect 53928 6244 53976 6300
rect 54032 6244 54080 6300
rect 54136 6244 54184 6300
rect 54240 6244 54288 6300
rect 54344 6244 54392 6300
rect 54448 6244 54458 6300
rect 53758 4732 54458 6244
rect 53758 4676 53768 4732
rect 53824 4676 53872 4732
rect 53928 4676 53976 4732
rect 54032 4676 54080 4732
rect 54136 4676 54184 4732
rect 54240 4676 54288 4732
rect 54344 4676 54392 4732
rect 54448 4676 54458 4732
rect 53758 3164 54458 4676
rect 53758 3108 53768 3164
rect 53824 3108 53872 3164
rect 53928 3108 53976 3164
rect 54032 3108 54080 3164
rect 54136 3108 54184 3164
rect 54240 3108 54288 3164
rect 54344 3108 54392 3164
rect 54448 3108 54458 3164
rect 53758 3076 54458 3108
rect 58258 55692 58958 56508
rect 58258 55636 58268 55692
rect 58324 55636 58372 55692
rect 58428 55636 58476 55692
rect 58532 55636 58580 55692
rect 58636 55636 58684 55692
rect 58740 55636 58788 55692
rect 58844 55636 58892 55692
rect 58948 55636 58958 55692
rect 58258 54124 58958 55636
rect 58258 54068 58268 54124
rect 58324 54068 58372 54124
rect 58428 54068 58476 54124
rect 58532 54068 58580 54124
rect 58636 54068 58684 54124
rect 58740 54068 58788 54124
rect 58844 54068 58892 54124
rect 58948 54068 58958 54124
rect 58258 52556 58958 54068
rect 58258 52500 58268 52556
rect 58324 52500 58372 52556
rect 58428 52500 58476 52556
rect 58532 52500 58580 52556
rect 58636 52500 58684 52556
rect 58740 52500 58788 52556
rect 58844 52500 58892 52556
rect 58948 52500 58958 52556
rect 58258 50988 58958 52500
rect 58258 50932 58268 50988
rect 58324 50932 58372 50988
rect 58428 50932 58476 50988
rect 58532 50932 58580 50988
rect 58636 50932 58684 50988
rect 58740 50932 58788 50988
rect 58844 50932 58892 50988
rect 58948 50932 58958 50988
rect 58258 49420 58958 50932
rect 58258 49364 58268 49420
rect 58324 49364 58372 49420
rect 58428 49364 58476 49420
rect 58532 49364 58580 49420
rect 58636 49364 58684 49420
rect 58740 49364 58788 49420
rect 58844 49364 58892 49420
rect 58948 49364 58958 49420
rect 58258 47852 58958 49364
rect 58258 47796 58268 47852
rect 58324 47796 58372 47852
rect 58428 47796 58476 47852
rect 58532 47796 58580 47852
rect 58636 47796 58684 47852
rect 58740 47796 58788 47852
rect 58844 47796 58892 47852
rect 58948 47796 58958 47852
rect 58258 46284 58958 47796
rect 58258 46228 58268 46284
rect 58324 46228 58372 46284
rect 58428 46228 58476 46284
rect 58532 46228 58580 46284
rect 58636 46228 58684 46284
rect 58740 46228 58788 46284
rect 58844 46228 58892 46284
rect 58948 46228 58958 46284
rect 58258 44716 58958 46228
rect 58258 44660 58268 44716
rect 58324 44660 58372 44716
rect 58428 44660 58476 44716
rect 58532 44660 58580 44716
rect 58636 44660 58684 44716
rect 58740 44660 58788 44716
rect 58844 44660 58892 44716
rect 58948 44660 58958 44716
rect 58258 43148 58958 44660
rect 58258 43092 58268 43148
rect 58324 43092 58372 43148
rect 58428 43092 58476 43148
rect 58532 43092 58580 43148
rect 58636 43092 58684 43148
rect 58740 43092 58788 43148
rect 58844 43092 58892 43148
rect 58948 43092 58958 43148
rect 58258 41580 58958 43092
rect 58258 41524 58268 41580
rect 58324 41524 58372 41580
rect 58428 41524 58476 41580
rect 58532 41524 58580 41580
rect 58636 41524 58684 41580
rect 58740 41524 58788 41580
rect 58844 41524 58892 41580
rect 58948 41524 58958 41580
rect 58258 40012 58958 41524
rect 58258 39956 58268 40012
rect 58324 39956 58372 40012
rect 58428 39956 58476 40012
rect 58532 39956 58580 40012
rect 58636 39956 58684 40012
rect 58740 39956 58788 40012
rect 58844 39956 58892 40012
rect 58948 39956 58958 40012
rect 58258 38444 58958 39956
rect 58258 38388 58268 38444
rect 58324 38388 58372 38444
rect 58428 38388 58476 38444
rect 58532 38388 58580 38444
rect 58636 38388 58684 38444
rect 58740 38388 58788 38444
rect 58844 38388 58892 38444
rect 58948 38388 58958 38444
rect 58258 36876 58958 38388
rect 58258 36820 58268 36876
rect 58324 36820 58372 36876
rect 58428 36820 58476 36876
rect 58532 36820 58580 36876
rect 58636 36820 58684 36876
rect 58740 36820 58788 36876
rect 58844 36820 58892 36876
rect 58948 36820 58958 36876
rect 58258 35308 58958 36820
rect 58258 35252 58268 35308
rect 58324 35252 58372 35308
rect 58428 35252 58476 35308
rect 58532 35252 58580 35308
rect 58636 35252 58684 35308
rect 58740 35252 58788 35308
rect 58844 35252 58892 35308
rect 58948 35252 58958 35308
rect 58258 33740 58958 35252
rect 58258 33684 58268 33740
rect 58324 33684 58372 33740
rect 58428 33684 58476 33740
rect 58532 33684 58580 33740
rect 58636 33684 58684 33740
rect 58740 33684 58788 33740
rect 58844 33684 58892 33740
rect 58948 33684 58958 33740
rect 58258 32172 58958 33684
rect 58258 32116 58268 32172
rect 58324 32116 58372 32172
rect 58428 32116 58476 32172
rect 58532 32116 58580 32172
rect 58636 32116 58684 32172
rect 58740 32116 58788 32172
rect 58844 32116 58892 32172
rect 58948 32116 58958 32172
rect 58258 30604 58958 32116
rect 58258 30548 58268 30604
rect 58324 30548 58372 30604
rect 58428 30548 58476 30604
rect 58532 30548 58580 30604
rect 58636 30548 58684 30604
rect 58740 30548 58788 30604
rect 58844 30548 58892 30604
rect 58948 30548 58958 30604
rect 58258 29036 58958 30548
rect 58258 28980 58268 29036
rect 58324 28980 58372 29036
rect 58428 28980 58476 29036
rect 58532 28980 58580 29036
rect 58636 28980 58684 29036
rect 58740 28980 58788 29036
rect 58844 28980 58892 29036
rect 58948 28980 58958 29036
rect 58258 27468 58958 28980
rect 58258 27412 58268 27468
rect 58324 27412 58372 27468
rect 58428 27412 58476 27468
rect 58532 27412 58580 27468
rect 58636 27412 58684 27468
rect 58740 27412 58788 27468
rect 58844 27412 58892 27468
rect 58948 27412 58958 27468
rect 58258 25900 58958 27412
rect 58258 25844 58268 25900
rect 58324 25844 58372 25900
rect 58428 25844 58476 25900
rect 58532 25844 58580 25900
rect 58636 25844 58684 25900
rect 58740 25844 58788 25900
rect 58844 25844 58892 25900
rect 58948 25844 58958 25900
rect 58258 24332 58958 25844
rect 58258 24276 58268 24332
rect 58324 24276 58372 24332
rect 58428 24276 58476 24332
rect 58532 24276 58580 24332
rect 58636 24276 58684 24332
rect 58740 24276 58788 24332
rect 58844 24276 58892 24332
rect 58948 24276 58958 24332
rect 58258 22764 58958 24276
rect 58258 22708 58268 22764
rect 58324 22708 58372 22764
rect 58428 22708 58476 22764
rect 58532 22708 58580 22764
rect 58636 22708 58684 22764
rect 58740 22708 58788 22764
rect 58844 22708 58892 22764
rect 58948 22708 58958 22764
rect 58258 21196 58958 22708
rect 58258 21140 58268 21196
rect 58324 21140 58372 21196
rect 58428 21140 58476 21196
rect 58532 21140 58580 21196
rect 58636 21140 58684 21196
rect 58740 21140 58788 21196
rect 58844 21140 58892 21196
rect 58948 21140 58958 21196
rect 58258 19628 58958 21140
rect 58258 19572 58268 19628
rect 58324 19572 58372 19628
rect 58428 19572 58476 19628
rect 58532 19572 58580 19628
rect 58636 19572 58684 19628
rect 58740 19572 58788 19628
rect 58844 19572 58892 19628
rect 58948 19572 58958 19628
rect 58258 18060 58958 19572
rect 58258 18004 58268 18060
rect 58324 18004 58372 18060
rect 58428 18004 58476 18060
rect 58532 18004 58580 18060
rect 58636 18004 58684 18060
rect 58740 18004 58788 18060
rect 58844 18004 58892 18060
rect 58948 18004 58958 18060
rect 58258 16492 58958 18004
rect 58258 16436 58268 16492
rect 58324 16436 58372 16492
rect 58428 16436 58476 16492
rect 58532 16436 58580 16492
rect 58636 16436 58684 16492
rect 58740 16436 58788 16492
rect 58844 16436 58892 16492
rect 58948 16436 58958 16492
rect 58258 14924 58958 16436
rect 58258 14868 58268 14924
rect 58324 14868 58372 14924
rect 58428 14868 58476 14924
rect 58532 14868 58580 14924
rect 58636 14868 58684 14924
rect 58740 14868 58788 14924
rect 58844 14868 58892 14924
rect 58948 14868 58958 14924
rect 58258 13356 58958 14868
rect 58258 13300 58268 13356
rect 58324 13300 58372 13356
rect 58428 13300 58476 13356
rect 58532 13300 58580 13356
rect 58636 13300 58684 13356
rect 58740 13300 58788 13356
rect 58844 13300 58892 13356
rect 58948 13300 58958 13356
rect 58258 11788 58958 13300
rect 58258 11732 58268 11788
rect 58324 11732 58372 11788
rect 58428 11732 58476 11788
rect 58532 11732 58580 11788
rect 58636 11732 58684 11788
rect 58740 11732 58788 11788
rect 58844 11732 58892 11788
rect 58948 11732 58958 11788
rect 58258 10220 58958 11732
rect 58258 10164 58268 10220
rect 58324 10164 58372 10220
rect 58428 10164 58476 10220
rect 58532 10164 58580 10220
rect 58636 10164 58684 10220
rect 58740 10164 58788 10220
rect 58844 10164 58892 10220
rect 58948 10164 58958 10220
rect 58258 8652 58958 10164
rect 58258 8596 58268 8652
rect 58324 8596 58372 8652
rect 58428 8596 58476 8652
rect 58532 8596 58580 8652
rect 58636 8596 58684 8652
rect 58740 8596 58788 8652
rect 58844 8596 58892 8652
rect 58948 8596 58958 8652
rect 58258 7084 58958 8596
rect 58258 7028 58268 7084
rect 58324 7028 58372 7084
rect 58428 7028 58476 7084
rect 58532 7028 58580 7084
rect 58636 7028 58684 7084
rect 58740 7028 58788 7084
rect 58844 7028 58892 7084
rect 58948 7028 58958 7084
rect 58258 5516 58958 7028
rect 58258 5460 58268 5516
rect 58324 5460 58372 5516
rect 58428 5460 58476 5516
rect 58532 5460 58580 5516
rect 58636 5460 58684 5516
rect 58740 5460 58788 5516
rect 58844 5460 58892 5516
rect 58948 5460 58958 5516
rect 58258 3948 58958 5460
rect 62758 56476 63458 56508
rect 62758 56420 62768 56476
rect 62824 56420 62872 56476
rect 62928 56420 62976 56476
rect 63032 56420 63080 56476
rect 63136 56420 63184 56476
rect 63240 56420 63288 56476
rect 63344 56420 63392 56476
rect 63448 56420 63458 56476
rect 62758 54908 63458 56420
rect 62758 54852 62768 54908
rect 62824 54852 62872 54908
rect 62928 54852 62976 54908
rect 63032 54852 63080 54908
rect 63136 54852 63184 54908
rect 63240 54852 63288 54908
rect 63344 54852 63392 54908
rect 63448 54852 63458 54908
rect 62758 53340 63458 54852
rect 62758 53284 62768 53340
rect 62824 53284 62872 53340
rect 62928 53284 62976 53340
rect 63032 53284 63080 53340
rect 63136 53284 63184 53340
rect 63240 53284 63288 53340
rect 63344 53284 63392 53340
rect 63448 53284 63458 53340
rect 62758 51772 63458 53284
rect 62758 51716 62768 51772
rect 62824 51716 62872 51772
rect 62928 51716 62976 51772
rect 63032 51716 63080 51772
rect 63136 51716 63184 51772
rect 63240 51716 63288 51772
rect 63344 51716 63392 51772
rect 63448 51716 63458 51772
rect 62758 50204 63458 51716
rect 62758 50148 62768 50204
rect 62824 50148 62872 50204
rect 62928 50148 62976 50204
rect 63032 50148 63080 50204
rect 63136 50148 63184 50204
rect 63240 50148 63288 50204
rect 63344 50148 63392 50204
rect 63448 50148 63458 50204
rect 62758 48636 63458 50148
rect 62758 48580 62768 48636
rect 62824 48580 62872 48636
rect 62928 48580 62976 48636
rect 63032 48580 63080 48636
rect 63136 48580 63184 48636
rect 63240 48580 63288 48636
rect 63344 48580 63392 48636
rect 63448 48580 63458 48636
rect 62758 47068 63458 48580
rect 62758 47012 62768 47068
rect 62824 47012 62872 47068
rect 62928 47012 62976 47068
rect 63032 47012 63080 47068
rect 63136 47012 63184 47068
rect 63240 47012 63288 47068
rect 63344 47012 63392 47068
rect 63448 47012 63458 47068
rect 62758 45500 63458 47012
rect 62758 45444 62768 45500
rect 62824 45444 62872 45500
rect 62928 45444 62976 45500
rect 63032 45444 63080 45500
rect 63136 45444 63184 45500
rect 63240 45444 63288 45500
rect 63344 45444 63392 45500
rect 63448 45444 63458 45500
rect 62758 43932 63458 45444
rect 62758 43876 62768 43932
rect 62824 43876 62872 43932
rect 62928 43876 62976 43932
rect 63032 43876 63080 43932
rect 63136 43876 63184 43932
rect 63240 43876 63288 43932
rect 63344 43876 63392 43932
rect 63448 43876 63458 43932
rect 62758 42364 63458 43876
rect 62758 42308 62768 42364
rect 62824 42308 62872 42364
rect 62928 42308 62976 42364
rect 63032 42308 63080 42364
rect 63136 42308 63184 42364
rect 63240 42308 63288 42364
rect 63344 42308 63392 42364
rect 63448 42308 63458 42364
rect 62758 40796 63458 42308
rect 62758 40740 62768 40796
rect 62824 40740 62872 40796
rect 62928 40740 62976 40796
rect 63032 40740 63080 40796
rect 63136 40740 63184 40796
rect 63240 40740 63288 40796
rect 63344 40740 63392 40796
rect 63448 40740 63458 40796
rect 62758 39228 63458 40740
rect 62758 39172 62768 39228
rect 62824 39172 62872 39228
rect 62928 39172 62976 39228
rect 63032 39172 63080 39228
rect 63136 39172 63184 39228
rect 63240 39172 63288 39228
rect 63344 39172 63392 39228
rect 63448 39172 63458 39228
rect 62758 37660 63458 39172
rect 62758 37604 62768 37660
rect 62824 37604 62872 37660
rect 62928 37604 62976 37660
rect 63032 37604 63080 37660
rect 63136 37604 63184 37660
rect 63240 37604 63288 37660
rect 63344 37604 63392 37660
rect 63448 37604 63458 37660
rect 62758 36092 63458 37604
rect 62758 36036 62768 36092
rect 62824 36036 62872 36092
rect 62928 36036 62976 36092
rect 63032 36036 63080 36092
rect 63136 36036 63184 36092
rect 63240 36036 63288 36092
rect 63344 36036 63392 36092
rect 63448 36036 63458 36092
rect 62758 34524 63458 36036
rect 62758 34468 62768 34524
rect 62824 34468 62872 34524
rect 62928 34468 62976 34524
rect 63032 34468 63080 34524
rect 63136 34468 63184 34524
rect 63240 34468 63288 34524
rect 63344 34468 63392 34524
rect 63448 34468 63458 34524
rect 62758 32956 63458 34468
rect 62758 32900 62768 32956
rect 62824 32900 62872 32956
rect 62928 32900 62976 32956
rect 63032 32900 63080 32956
rect 63136 32900 63184 32956
rect 63240 32900 63288 32956
rect 63344 32900 63392 32956
rect 63448 32900 63458 32956
rect 62758 31388 63458 32900
rect 62758 31332 62768 31388
rect 62824 31332 62872 31388
rect 62928 31332 62976 31388
rect 63032 31332 63080 31388
rect 63136 31332 63184 31388
rect 63240 31332 63288 31388
rect 63344 31332 63392 31388
rect 63448 31332 63458 31388
rect 62758 29820 63458 31332
rect 62758 29764 62768 29820
rect 62824 29764 62872 29820
rect 62928 29764 62976 29820
rect 63032 29764 63080 29820
rect 63136 29764 63184 29820
rect 63240 29764 63288 29820
rect 63344 29764 63392 29820
rect 63448 29764 63458 29820
rect 62758 28252 63458 29764
rect 62758 28196 62768 28252
rect 62824 28196 62872 28252
rect 62928 28196 62976 28252
rect 63032 28196 63080 28252
rect 63136 28196 63184 28252
rect 63240 28196 63288 28252
rect 63344 28196 63392 28252
rect 63448 28196 63458 28252
rect 62758 26684 63458 28196
rect 62758 26628 62768 26684
rect 62824 26628 62872 26684
rect 62928 26628 62976 26684
rect 63032 26628 63080 26684
rect 63136 26628 63184 26684
rect 63240 26628 63288 26684
rect 63344 26628 63392 26684
rect 63448 26628 63458 26684
rect 62758 25116 63458 26628
rect 67258 55692 67958 56508
rect 67258 55636 67268 55692
rect 67324 55636 67372 55692
rect 67428 55636 67476 55692
rect 67532 55636 67580 55692
rect 67636 55636 67684 55692
rect 67740 55636 67788 55692
rect 67844 55636 67892 55692
rect 67948 55636 67958 55692
rect 67258 54124 67958 55636
rect 67258 54068 67268 54124
rect 67324 54068 67372 54124
rect 67428 54068 67476 54124
rect 67532 54068 67580 54124
rect 67636 54068 67684 54124
rect 67740 54068 67788 54124
rect 67844 54068 67892 54124
rect 67948 54068 67958 54124
rect 67258 52556 67958 54068
rect 67258 52500 67268 52556
rect 67324 52500 67372 52556
rect 67428 52500 67476 52556
rect 67532 52500 67580 52556
rect 67636 52500 67684 52556
rect 67740 52500 67788 52556
rect 67844 52500 67892 52556
rect 67948 52500 67958 52556
rect 67258 50988 67958 52500
rect 67258 50932 67268 50988
rect 67324 50932 67372 50988
rect 67428 50932 67476 50988
rect 67532 50932 67580 50988
rect 67636 50932 67684 50988
rect 67740 50932 67788 50988
rect 67844 50932 67892 50988
rect 67948 50932 67958 50988
rect 67258 49420 67958 50932
rect 67258 49364 67268 49420
rect 67324 49364 67372 49420
rect 67428 49364 67476 49420
rect 67532 49364 67580 49420
rect 67636 49364 67684 49420
rect 67740 49364 67788 49420
rect 67844 49364 67892 49420
rect 67948 49364 67958 49420
rect 67258 47852 67958 49364
rect 67258 47796 67268 47852
rect 67324 47796 67372 47852
rect 67428 47796 67476 47852
rect 67532 47796 67580 47852
rect 67636 47796 67684 47852
rect 67740 47796 67788 47852
rect 67844 47796 67892 47852
rect 67948 47796 67958 47852
rect 67258 46284 67958 47796
rect 67258 46228 67268 46284
rect 67324 46228 67372 46284
rect 67428 46228 67476 46284
rect 67532 46228 67580 46284
rect 67636 46228 67684 46284
rect 67740 46228 67788 46284
rect 67844 46228 67892 46284
rect 67948 46228 67958 46284
rect 67258 44716 67958 46228
rect 67258 44660 67268 44716
rect 67324 44660 67372 44716
rect 67428 44660 67476 44716
rect 67532 44660 67580 44716
rect 67636 44660 67684 44716
rect 67740 44660 67788 44716
rect 67844 44660 67892 44716
rect 67948 44660 67958 44716
rect 67258 43148 67958 44660
rect 67258 43092 67268 43148
rect 67324 43092 67372 43148
rect 67428 43092 67476 43148
rect 67532 43092 67580 43148
rect 67636 43092 67684 43148
rect 67740 43092 67788 43148
rect 67844 43092 67892 43148
rect 67948 43092 67958 43148
rect 67258 41580 67958 43092
rect 67258 41524 67268 41580
rect 67324 41524 67372 41580
rect 67428 41524 67476 41580
rect 67532 41524 67580 41580
rect 67636 41524 67684 41580
rect 67740 41524 67788 41580
rect 67844 41524 67892 41580
rect 67948 41524 67958 41580
rect 67258 40012 67958 41524
rect 67258 39956 67268 40012
rect 67324 39956 67372 40012
rect 67428 39956 67476 40012
rect 67532 39956 67580 40012
rect 67636 39956 67684 40012
rect 67740 39956 67788 40012
rect 67844 39956 67892 40012
rect 67948 39956 67958 40012
rect 67258 38444 67958 39956
rect 67258 38388 67268 38444
rect 67324 38388 67372 38444
rect 67428 38388 67476 38444
rect 67532 38388 67580 38444
rect 67636 38388 67684 38444
rect 67740 38388 67788 38444
rect 67844 38388 67892 38444
rect 67948 38388 67958 38444
rect 67258 36876 67958 38388
rect 71758 56476 72458 56508
rect 71758 56420 71768 56476
rect 71824 56420 71872 56476
rect 71928 56420 71976 56476
rect 72032 56420 72080 56476
rect 72136 56420 72184 56476
rect 72240 56420 72288 56476
rect 72344 56420 72392 56476
rect 72448 56420 72458 56476
rect 71758 54908 72458 56420
rect 71758 54852 71768 54908
rect 71824 54852 71872 54908
rect 71928 54852 71976 54908
rect 72032 54852 72080 54908
rect 72136 54852 72184 54908
rect 72240 54852 72288 54908
rect 72344 54852 72392 54908
rect 72448 54852 72458 54908
rect 71758 53340 72458 54852
rect 71758 53284 71768 53340
rect 71824 53284 71872 53340
rect 71928 53284 71976 53340
rect 72032 53284 72080 53340
rect 72136 53284 72184 53340
rect 72240 53284 72288 53340
rect 72344 53284 72392 53340
rect 72448 53284 72458 53340
rect 71758 51772 72458 53284
rect 71758 51716 71768 51772
rect 71824 51716 71872 51772
rect 71928 51716 71976 51772
rect 72032 51716 72080 51772
rect 72136 51716 72184 51772
rect 72240 51716 72288 51772
rect 72344 51716 72392 51772
rect 72448 51716 72458 51772
rect 71758 50204 72458 51716
rect 71758 50148 71768 50204
rect 71824 50148 71872 50204
rect 71928 50148 71976 50204
rect 72032 50148 72080 50204
rect 72136 50148 72184 50204
rect 72240 50148 72288 50204
rect 72344 50148 72392 50204
rect 72448 50148 72458 50204
rect 71758 48636 72458 50148
rect 71758 48580 71768 48636
rect 71824 48580 71872 48636
rect 71928 48580 71976 48636
rect 72032 48580 72080 48636
rect 72136 48580 72184 48636
rect 72240 48580 72288 48636
rect 72344 48580 72392 48636
rect 72448 48580 72458 48636
rect 71758 47068 72458 48580
rect 71758 47012 71768 47068
rect 71824 47012 71872 47068
rect 71928 47012 71976 47068
rect 72032 47012 72080 47068
rect 72136 47012 72184 47068
rect 72240 47012 72288 47068
rect 72344 47012 72392 47068
rect 72448 47012 72458 47068
rect 71758 45500 72458 47012
rect 71758 45444 71768 45500
rect 71824 45444 71872 45500
rect 71928 45444 71976 45500
rect 72032 45444 72080 45500
rect 72136 45444 72184 45500
rect 72240 45444 72288 45500
rect 72344 45444 72392 45500
rect 72448 45444 72458 45500
rect 71758 43932 72458 45444
rect 71758 43876 71768 43932
rect 71824 43876 71872 43932
rect 71928 43876 71976 43932
rect 72032 43876 72080 43932
rect 72136 43876 72184 43932
rect 72240 43876 72288 43932
rect 72344 43876 72392 43932
rect 72448 43876 72458 43932
rect 71758 42364 72458 43876
rect 71758 42308 71768 42364
rect 71824 42308 71872 42364
rect 71928 42308 71976 42364
rect 72032 42308 72080 42364
rect 72136 42308 72184 42364
rect 72240 42308 72288 42364
rect 72344 42308 72392 42364
rect 72448 42308 72458 42364
rect 71758 40796 72458 42308
rect 71758 40740 71768 40796
rect 71824 40740 71872 40796
rect 71928 40740 71976 40796
rect 72032 40740 72080 40796
rect 72136 40740 72184 40796
rect 72240 40740 72288 40796
rect 72344 40740 72392 40796
rect 72448 40740 72458 40796
rect 71758 39228 72458 40740
rect 71758 39172 71768 39228
rect 71824 39172 71872 39228
rect 71928 39172 71976 39228
rect 72032 39172 72080 39228
rect 72136 39172 72184 39228
rect 72240 39172 72288 39228
rect 72344 39172 72392 39228
rect 72448 39172 72458 39228
rect 71758 37660 72458 39172
rect 67258 36820 67268 36876
rect 67324 36820 67372 36876
rect 67428 36820 67476 36876
rect 67532 36820 67580 36876
rect 67636 36820 67684 36876
rect 67740 36820 67788 36876
rect 67844 36820 67892 36876
rect 67948 36820 67958 36876
rect 67258 35308 67958 36820
rect 68236 37604 68292 37614
rect 68236 35700 68292 37548
rect 68236 35634 68292 35644
rect 71758 37604 71768 37660
rect 71824 37604 71872 37660
rect 71928 37604 71976 37660
rect 72032 37604 72080 37660
rect 72136 37604 72184 37660
rect 72240 37604 72288 37660
rect 72344 37604 72392 37660
rect 72448 37604 72458 37660
rect 71758 36092 72458 37604
rect 71758 36036 71768 36092
rect 71824 36036 71872 36092
rect 71928 36036 71976 36092
rect 72032 36036 72080 36092
rect 72136 36036 72184 36092
rect 72240 36036 72288 36092
rect 72344 36036 72392 36092
rect 72448 36036 72458 36092
rect 67258 35252 67268 35308
rect 67324 35252 67372 35308
rect 67428 35252 67476 35308
rect 67532 35252 67580 35308
rect 67636 35252 67684 35308
rect 67740 35252 67788 35308
rect 67844 35252 67892 35308
rect 67948 35252 67958 35308
rect 67258 33740 67958 35252
rect 67258 33684 67268 33740
rect 67324 33684 67372 33740
rect 67428 33684 67476 33740
rect 67532 33684 67580 33740
rect 67636 33684 67684 33740
rect 67740 33684 67788 33740
rect 67844 33684 67892 33740
rect 67948 33684 67958 33740
rect 67258 32172 67958 33684
rect 67258 32116 67268 32172
rect 67324 32116 67372 32172
rect 67428 32116 67476 32172
rect 67532 32116 67580 32172
rect 67636 32116 67684 32172
rect 67740 32116 67788 32172
rect 67844 32116 67892 32172
rect 67948 32116 67958 32172
rect 67258 30604 67958 32116
rect 67258 30548 67268 30604
rect 67324 30548 67372 30604
rect 67428 30548 67476 30604
rect 67532 30548 67580 30604
rect 67636 30548 67684 30604
rect 67740 30548 67788 30604
rect 67844 30548 67892 30604
rect 67948 30548 67958 30604
rect 67258 29036 67958 30548
rect 67258 28980 67268 29036
rect 67324 28980 67372 29036
rect 67428 28980 67476 29036
rect 67532 28980 67580 29036
rect 67636 28980 67684 29036
rect 67740 28980 67788 29036
rect 67844 28980 67892 29036
rect 67948 28980 67958 29036
rect 67258 27468 67958 28980
rect 71758 34524 72458 36036
rect 71758 34468 71768 34524
rect 71824 34468 71872 34524
rect 71928 34468 71976 34524
rect 72032 34468 72080 34524
rect 72136 34468 72184 34524
rect 72240 34468 72288 34524
rect 72344 34468 72392 34524
rect 72448 34468 72458 34524
rect 71758 32956 72458 34468
rect 71758 32900 71768 32956
rect 71824 32900 71872 32956
rect 71928 32900 71976 32956
rect 72032 32900 72080 32956
rect 72136 32900 72184 32956
rect 72240 32900 72288 32956
rect 72344 32900 72392 32956
rect 72448 32900 72458 32956
rect 71758 31388 72458 32900
rect 71758 31332 71768 31388
rect 71824 31332 71872 31388
rect 71928 31332 71976 31388
rect 72032 31332 72080 31388
rect 72136 31332 72184 31388
rect 72240 31332 72288 31388
rect 72344 31332 72392 31388
rect 72448 31332 72458 31388
rect 71758 29820 72458 31332
rect 71758 29764 71768 29820
rect 71824 29764 71872 29820
rect 71928 29764 71976 29820
rect 72032 29764 72080 29820
rect 72136 29764 72184 29820
rect 72240 29764 72288 29820
rect 72344 29764 72392 29820
rect 72448 29764 72458 29820
rect 67258 27412 67268 27468
rect 67324 27412 67372 27468
rect 67428 27412 67476 27468
rect 67532 27412 67580 27468
rect 67636 27412 67684 27468
rect 67740 27412 67788 27468
rect 67844 27412 67892 27468
rect 67948 27412 67958 27468
rect 62758 25060 62768 25116
rect 62824 25060 62872 25116
rect 62928 25060 62976 25116
rect 63032 25060 63080 25116
rect 63136 25060 63184 25116
rect 63240 25060 63288 25116
rect 63344 25060 63392 25116
rect 63448 25060 63458 25116
rect 62758 23548 63458 25060
rect 62758 23492 62768 23548
rect 62824 23492 62872 23548
rect 62928 23492 62976 23548
rect 63032 23492 63080 23548
rect 63136 23492 63184 23548
rect 63240 23492 63288 23548
rect 63344 23492 63392 23548
rect 63448 23492 63458 23548
rect 62758 21980 63458 23492
rect 67116 26180 67172 26190
rect 67116 25284 67172 26124
rect 67116 22260 67172 25228
rect 67116 22194 67172 22204
rect 67258 25900 67958 27412
rect 67258 25844 67268 25900
rect 67324 25844 67372 25900
rect 67428 25844 67476 25900
rect 67532 25844 67580 25900
rect 67636 25844 67684 25900
rect 67740 25844 67788 25900
rect 67844 25844 67892 25900
rect 67948 25844 67958 25900
rect 67258 24332 67958 25844
rect 67258 24276 67268 24332
rect 67324 24276 67372 24332
rect 67428 24276 67476 24332
rect 67532 24276 67580 24332
rect 67636 24276 67684 24332
rect 67740 24276 67788 24332
rect 67844 24276 67892 24332
rect 67948 24276 67958 24332
rect 67258 22764 67958 24276
rect 67258 22708 67268 22764
rect 67324 22708 67372 22764
rect 67428 22708 67476 22764
rect 67532 22708 67580 22764
rect 67636 22708 67684 22764
rect 67740 22708 67788 22764
rect 67844 22708 67892 22764
rect 67948 22708 67958 22764
rect 62758 21924 62768 21980
rect 62824 21924 62872 21980
rect 62928 21924 62976 21980
rect 63032 21924 63080 21980
rect 63136 21924 63184 21980
rect 63240 21924 63288 21980
rect 63344 21924 63392 21980
rect 63448 21924 63458 21980
rect 62758 20412 63458 21924
rect 62758 20356 62768 20412
rect 62824 20356 62872 20412
rect 62928 20356 62976 20412
rect 63032 20356 63080 20412
rect 63136 20356 63184 20412
rect 63240 20356 63288 20412
rect 63344 20356 63392 20412
rect 63448 20356 63458 20412
rect 62758 18844 63458 20356
rect 62758 18788 62768 18844
rect 62824 18788 62872 18844
rect 62928 18788 62976 18844
rect 63032 18788 63080 18844
rect 63136 18788 63184 18844
rect 63240 18788 63288 18844
rect 63344 18788 63392 18844
rect 63448 18788 63458 18844
rect 62758 17276 63458 18788
rect 62758 17220 62768 17276
rect 62824 17220 62872 17276
rect 62928 17220 62976 17276
rect 63032 17220 63080 17276
rect 63136 17220 63184 17276
rect 63240 17220 63288 17276
rect 63344 17220 63392 17276
rect 63448 17220 63458 17276
rect 62758 15708 63458 17220
rect 62758 15652 62768 15708
rect 62824 15652 62872 15708
rect 62928 15652 62976 15708
rect 63032 15652 63080 15708
rect 63136 15652 63184 15708
rect 63240 15652 63288 15708
rect 63344 15652 63392 15708
rect 63448 15652 63458 15708
rect 62758 14140 63458 15652
rect 62758 14084 62768 14140
rect 62824 14084 62872 14140
rect 62928 14084 62976 14140
rect 63032 14084 63080 14140
rect 63136 14084 63184 14140
rect 63240 14084 63288 14140
rect 63344 14084 63392 14140
rect 63448 14084 63458 14140
rect 62758 12572 63458 14084
rect 62758 12516 62768 12572
rect 62824 12516 62872 12572
rect 62928 12516 62976 12572
rect 63032 12516 63080 12572
rect 63136 12516 63184 12572
rect 63240 12516 63288 12572
rect 63344 12516 63392 12572
rect 63448 12516 63458 12572
rect 62758 11004 63458 12516
rect 62758 10948 62768 11004
rect 62824 10948 62872 11004
rect 62928 10948 62976 11004
rect 63032 10948 63080 11004
rect 63136 10948 63184 11004
rect 63240 10948 63288 11004
rect 63344 10948 63392 11004
rect 63448 10948 63458 11004
rect 62758 9436 63458 10948
rect 62758 9380 62768 9436
rect 62824 9380 62872 9436
rect 62928 9380 62976 9436
rect 63032 9380 63080 9436
rect 63136 9380 63184 9436
rect 63240 9380 63288 9436
rect 63344 9380 63392 9436
rect 63448 9380 63458 9436
rect 62758 7868 63458 9380
rect 62758 7812 62768 7868
rect 62824 7812 62872 7868
rect 62928 7812 62976 7868
rect 63032 7812 63080 7868
rect 63136 7812 63184 7868
rect 63240 7812 63288 7868
rect 63344 7812 63392 7868
rect 63448 7812 63458 7868
rect 62758 6300 63458 7812
rect 62758 6244 62768 6300
rect 62824 6244 62872 6300
rect 62928 6244 62976 6300
rect 63032 6244 63080 6300
rect 63136 6244 63184 6300
rect 63240 6244 63288 6300
rect 63344 6244 63392 6300
rect 63448 6244 63458 6300
rect 59612 5012 59668 5022
rect 59612 4912 59668 4922
rect 58258 3892 58268 3948
rect 58324 3892 58372 3948
rect 58428 3892 58476 3948
rect 58532 3892 58580 3948
rect 58636 3892 58684 3948
rect 58740 3892 58788 3948
rect 58844 3892 58892 3948
rect 58948 3892 58958 3948
rect 58258 3076 58958 3892
rect 62758 4732 63458 6244
rect 62758 4676 62768 4732
rect 62824 4676 62872 4732
rect 62928 4676 62976 4732
rect 63032 4676 63080 4732
rect 63136 4676 63184 4732
rect 63240 4676 63288 4732
rect 63344 4676 63392 4732
rect 63448 4676 63458 4732
rect 62758 3164 63458 4676
rect 62758 3108 62768 3164
rect 62824 3108 62872 3164
rect 62928 3108 62976 3164
rect 63032 3108 63080 3164
rect 63136 3108 63184 3164
rect 63240 3108 63288 3164
rect 63344 3108 63392 3164
rect 63448 3108 63458 3164
rect 62758 3076 63458 3108
rect 67258 21196 67958 22708
rect 68124 28644 68180 28654
rect 68124 21700 68180 28588
rect 68124 21634 68180 21644
rect 71758 28252 72458 29764
rect 71758 28196 71768 28252
rect 71824 28196 71872 28252
rect 71928 28196 71976 28252
rect 72032 28196 72080 28252
rect 72136 28196 72184 28252
rect 72240 28196 72288 28252
rect 72344 28196 72392 28252
rect 72448 28196 72458 28252
rect 71758 26684 72458 28196
rect 71758 26628 71768 26684
rect 71824 26628 71872 26684
rect 71928 26628 71976 26684
rect 72032 26628 72080 26684
rect 72136 26628 72184 26684
rect 72240 26628 72288 26684
rect 72344 26628 72392 26684
rect 72448 26628 72458 26684
rect 71758 25116 72458 26628
rect 71758 25060 71768 25116
rect 71824 25060 71872 25116
rect 71928 25060 71976 25116
rect 72032 25060 72080 25116
rect 72136 25060 72184 25116
rect 72240 25060 72288 25116
rect 72344 25060 72392 25116
rect 72448 25060 72458 25116
rect 71758 23548 72458 25060
rect 71758 23492 71768 23548
rect 71824 23492 71872 23548
rect 71928 23492 71976 23548
rect 72032 23492 72080 23548
rect 72136 23492 72184 23548
rect 72240 23492 72288 23548
rect 72344 23492 72392 23548
rect 72448 23492 72458 23548
rect 71758 21980 72458 23492
rect 71758 21924 71768 21980
rect 71824 21924 71872 21980
rect 71928 21924 71976 21980
rect 72032 21924 72080 21980
rect 72136 21924 72184 21980
rect 72240 21924 72288 21980
rect 72344 21924 72392 21980
rect 72448 21924 72458 21980
rect 67258 21140 67268 21196
rect 67324 21140 67372 21196
rect 67428 21140 67476 21196
rect 67532 21140 67580 21196
rect 67636 21140 67684 21196
rect 67740 21140 67788 21196
rect 67844 21140 67892 21196
rect 67948 21140 67958 21196
rect 67258 19628 67958 21140
rect 67258 19572 67268 19628
rect 67324 19572 67372 19628
rect 67428 19572 67476 19628
rect 67532 19572 67580 19628
rect 67636 19572 67684 19628
rect 67740 19572 67788 19628
rect 67844 19572 67892 19628
rect 67948 19572 67958 19628
rect 67258 18060 67958 19572
rect 67258 18004 67268 18060
rect 67324 18004 67372 18060
rect 67428 18004 67476 18060
rect 67532 18004 67580 18060
rect 67636 18004 67684 18060
rect 67740 18004 67788 18060
rect 67844 18004 67892 18060
rect 67948 18004 67958 18060
rect 67258 16492 67958 18004
rect 67258 16436 67268 16492
rect 67324 16436 67372 16492
rect 67428 16436 67476 16492
rect 67532 16436 67580 16492
rect 67636 16436 67684 16492
rect 67740 16436 67788 16492
rect 67844 16436 67892 16492
rect 67948 16436 67958 16492
rect 67258 14924 67958 16436
rect 67258 14868 67268 14924
rect 67324 14868 67372 14924
rect 67428 14868 67476 14924
rect 67532 14868 67580 14924
rect 67636 14868 67684 14924
rect 67740 14868 67788 14924
rect 67844 14868 67892 14924
rect 67948 14868 67958 14924
rect 67258 13356 67958 14868
rect 67258 13300 67268 13356
rect 67324 13300 67372 13356
rect 67428 13300 67476 13356
rect 67532 13300 67580 13356
rect 67636 13300 67684 13356
rect 67740 13300 67788 13356
rect 67844 13300 67892 13356
rect 67948 13300 67958 13356
rect 67258 11788 67958 13300
rect 67258 11732 67268 11788
rect 67324 11732 67372 11788
rect 67428 11732 67476 11788
rect 67532 11732 67580 11788
rect 67636 11732 67684 11788
rect 67740 11732 67788 11788
rect 67844 11732 67892 11788
rect 67948 11732 67958 11788
rect 67258 10220 67958 11732
rect 67258 10164 67268 10220
rect 67324 10164 67372 10220
rect 67428 10164 67476 10220
rect 67532 10164 67580 10220
rect 67636 10164 67684 10220
rect 67740 10164 67788 10220
rect 67844 10164 67892 10220
rect 67948 10164 67958 10220
rect 67258 8652 67958 10164
rect 67258 8596 67268 8652
rect 67324 8596 67372 8652
rect 67428 8596 67476 8652
rect 67532 8596 67580 8652
rect 67636 8596 67684 8652
rect 67740 8596 67788 8652
rect 67844 8596 67892 8652
rect 67948 8596 67958 8652
rect 67258 7084 67958 8596
rect 67258 7028 67268 7084
rect 67324 7028 67372 7084
rect 67428 7028 67476 7084
rect 67532 7028 67580 7084
rect 67636 7028 67684 7084
rect 67740 7028 67788 7084
rect 67844 7028 67892 7084
rect 67948 7028 67958 7084
rect 67258 5516 67958 7028
rect 67258 5460 67268 5516
rect 67324 5460 67372 5516
rect 67428 5460 67476 5516
rect 67532 5460 67580 5516
rect 67636 5460 67684 5516
rect 67740 5460 67788 5516
rect 67844 5460 67892 5516
rect 67948 5460 67958 5516
rect 67258 3948 67958 5460
rect 67258 3892 67268 3948
rect 67324 3892 67372 3948
rect 67428 3892 67476 3948
rect 67532 3892 67580 3948
rect 67636 3892 67684 3948
rect 67740 3892 67788 3948
rect 67844 3892 67892 3948
rect 67948 3892 67958 3948
rect 67258 3076 67958 3892
rect 71758 20412 72458 21924
rect 71758 20356 71768 20412
rect 71824 20356 71872 20412
rect 71928 20356 71976 20412
rect 72032 20356 72080 20412
rect 72136 20356 72184 20412
rect 72240 20356 72288 20412
rect 72344 20356 72392 20412
rect 72448 20356 72458 20412
rect 71758 18844 72458 20356
rect 71758 18788 71768 18844
rect 71824 18788 71872 18844
rect 71928 18788 71976 18844
rect 72032 18788 72080 18844
rect 72136 18788 72184 18844
rect 72240 18788 72288 18844
rect 72344 18788 72392 18844
rect 72448 18788 72458 18844
rect 71758 17276 72458 18788
rect 71758 17220 71768 17276
rect 71824 17220 71872 17276
rect 71928 17220 71976 17276
rect 72032 17220 72080 17276
rect 72136 17220 72184 17276
rect 72240 17220 72288 17276
rect 72344 17220 72392 17276
rect 72448 17220 72458 17276
rect 71758 15708 72458 17220
rect 71758 15652 71768 15708
rect 71824 15652 71872 15708
rect 71928 15652 71976 15708
rect 72032 15652 72080 15708
rect 72136 15652 72184 15708
rect 72240 15652 72288 15708
rect 72344 15652 72392 15708
rect 72448 15652 72458 15708
rect 71758 14140 72458 15652
rect 71758 14084 71768 14140
rect 71824 14084 71872 14140
rect 71928 14084 71976 14140
rect 72032 14084 72080 14140
rect 72136 14084 72184 14140
rect 72240 14084 72288 14140
rect 72344 14084 72392 14140
rect 72448 14084 72458 14140
rect 71758 12572 72458 14084
rect 71758 12516 71768 12572
rect 71824 12516 71872 12572
rect 71928 12516 71976 12572
rect 72032 12516 72080 12572
rect 72136 12516 72184 12572
rect 72240 12516 72288 12572
rect 72344 12516 72392 12572
rect 72448 12516 72458 12572
rect 71758 11004 72458 12516
rect 71758 10948 71768 11004
rect 71824 10948 71872 11004
rect 71928 10948 71976 11004
rect 72032 10948 72080 11004
rect 72136 10948 72184 11004
rect 72240 10948 72288 11004
rect 72344 10948 72392 11004
rect 72448 10948 72458 11004
rect 71758 9436 72458 10948
rect 71758 9380 71768 9436
rect 71824 9380 71872 9436
rect 71928 9380 71976 9436
rect 72032 9380 72080 9436
rect 72136 9380 72184 9436
rect 72240 9380 72288 9436
rect 72344 9380 72392 9436
rect 72448 9380 72458 9436
rect 71758 7868 72458 9380
rect 71758 7812 71768 7868
rect 71824 7812 71872 7868
rect 71928 7812 71976 7868
rect 72032 7812 72080 7868
rect 72136 7812 72184 7868
rect 72240 7812 72288 7868
rect 72344 7812 72392 7868
rect 72448 7812 72458 7868
rect 71758 6300 72458 7812
rect 71758 6244 71768 6300
rect 71824 6244 71872 6300
rect 71928 6244 71976 6300
rect 72032 6244 72080 6300
rect 72136 6244 72184 6300
rect 72240 6244 72288 6300
rect 72344 6244 72392 6300
rect 72448 6244 72458 6300
rect 71758 4732 72458 6244
rect 76258 55692 76958 56508
rect 76258 55636 76268 55692
rect 76324 55636 76372 55692
rect 76428 55636 76476 55692
rect 76532 55636 76580 55692
rect 76636 55636 76684 55692
rect 76740 55636 76788 55692
rect 76844 55636 76892 55692
rect 76948 55636 76958 55692
rect 76258 54124 76958 55636
rect 76258 54068 76268 54124
rect 76324 54068 76372 54124
rect 76428 54068 76476 54124
rect 76532 54068 76580 54124
rect 76636 54068 76684 54124
rect 76740 54068 76788 54124
rect 76844 54068 76892 54124
rect 76948 54068 76958 54124
rect 76258 52556 76958 54068
rect 76258 52500 76268 52556
rect 76324 52500 76372 52556
rect 76428 52500 76476 52556
rect 76532 52500 76580 52556
rect 76636 52500 76684 52556
rect 76740 52500 76788 52556
rect 76844 52500 76892 52556
rect 76948 52500 76958 52556
rect 76258 50988 76958 52500
rect 76258 50932 76268 50988
rect 76324 50932 76372 50988
rect 76428 50932 76476 50988
rect 76532 50932 76580 50988
rect 76636 50932 76684 50988
rect 76740 50932 76788 50988
rect 76844 50932 76892 50988
rect 76948 50932 76958 50988
rect 76258 49420 76958 50932
rect 76258 49364 76268 49420
rect 76324 49364 76372 49420
rect 76428 49364 76476 49420
rect 76532 49364 76580 49420
rect 76636 49364 76684 49420
rect 76740 49364 76788 49420
rect 76844 49364 76892 49420
rect 76948 49364 76958 49420
rect 76258 47852 76958 49364
rect 76258 47796 76268 47852
rect 76324 47796 76372 47852
rect 76428 47796 76476 47852
rect 76532 47796 76580 47852
rect 76636 47796 76684 47852
rect 76740 47796 76788 47852
rect 76844 47796 76892 47852
rect 76948 47796 76958 47852
rect 76258 46284 76958 47796
rect 76258 46228 76268 46284
rect 76324 46228 76372 46284
rect 76428 46228 76476 46284
rect 76532 46228 76580 46284
rect 76636 46228 76684 46284
rect 76740 46228 76788 46284
rect 76844 46228 76892 46284
rect 76948 46228 76958 46284
rect 76258 44716 76958 46228
rect 76258 44660 76268 44716
rect 76324 44660 76372 44716
rect 76428 44660 76476 44716
rect 76532 44660 76580 44716
rect 76636 44660 76684 44716
rect 76740 44660 76788 44716
rect 76844 44660 76892 44716
rect 76948 44660 76958 44716
rect 76258 43148 76958 44660
rect 76258 43092 76268 43148
rect 76324 43092 76372 43148
rect 76428 43092 76476 43148
rect 76532 43092 76580 43148
rect 76636 43092 76684 43148
rect 76740 43092 76788 43148
rect 76844 43092 76892 43148
rect 76948 43092 76958 43148
rect 76258 41580 76958 43092
rect 76258 41524 76268 41580
rect 76324 41524 76372 41580
rect 76428 41524 76476 41580
rect 76532 41524 76580 41580
rect 76636 41524 76684 41580
rect 76740 41524 76788 41580
rect 76844 41524 76892 41580
rect 76948 41524 76958 41580
rect 76258 40012 76958 41524
rect 76258 39956 76268 40012
rect 76324 39956 76372 40012
rect 76428 39956 76476 40012
rect 76532 39956 76580 40012
rect 76636 39956 76684 40012
rect 76740 39956 76788 40012
rect 76844 39956 76892 40012
rect 76948 39956 76958 40012
rect 76258 38444 76958 39956
rect 76258 38388 76268 38444
rect 76324 38388 76372 38444
rect 76428 38388 76476 38444
rect 76532 38388 76580 38444
rect 76636 38388 76684 38444
rect 76740 38388 76788 38444
rect 76844 38388 76892 38444
rect 76948 38388 76958 38444
rect 76258 36876 76958 38388
rect 76258 36820 76268 36876
rect 76324 36820 76372 36876
rect 76428 36820 76476 36876
rect 76532 36820 76580 36876
rect 76636 36820 76684 36876
rect 76740 36820 76788 36876
rect 76844 36820 76892 36876
rect 76948 36820 76958 36876
rect 76258 35308 76958 36820
rect 76258 35252 76268 35308
rect 76324 35252 76372 35308
rect 76428 35252 76476 35308
rect 76532 35252 76580 35308
rect 76636 35252 76684 35308
rect 76740 35252 76788 35308
rect 76844 35252 76892 35308
rect 76948 35252 76958 35308
rect 76258 33740 76958 35252
rect 76258 33684 76268 33740
rect 76324 33684 76372 33740
rect 76428 33684 76476 33740
rect 76532 33684 76580 33740
rect 76636 33684 76684 33740
rect 76740 33684 76788 33740
rect 76844 33684 76892 33740
rect 76948 33684 76958 33740
rect 76258 32172 76958 33684
rect 76258 32116 76268 32172
rect 76324 32116 76372 32172
rect 76428 32116 76476 32172
rect 76532 32116 76580 32172
rect 76636 32116 76684 32172
rect 76740 32116 76788 32172
rect 76844 32116 76892 32172
rect 76948 32116 76958 32172
rect 76258 30604 76958 32116
rect 76258 30548 76268 30604
rect 76324 30548 76372 30604
rect 76428 30548 76476 30604
rect 76532 30548 76580 30604
rect 76636 30548 76684 30604
rect 76740 30548 76788 30604
rect 76844 30548 76892 30604
rect 76948 30548 76958 30604
rect 76258 29036 76958 30548
rect 76258 28980 76268 29036
rect 76324 28980 76372 29036
rect 76428 28980 76476 29036
rect 76532 28980 76580 29036
rect 76636 28980 76684 29036
rect 76740 28980 76788 29036
rect 76844 28980 76892 29036
rect 76948 28980 76958 29036
rect 76258 27468 76958 28980
rect 76258 27412 76268 27468
rect 76324 27412 76372 27468
rect 76428 27412 76476 27468
rect 76532 27412 76580 27468
rect 76636 27412 76684 27468
rect 76740 27412 76788 27468
rect 76844 27412 76892 27468
rect 76948 27412 76958 27468
rect 76258 25900 76958 27412
rect 76258 25844 76268 25900
rect 76324 25844 76372 25900
rect 76428 25844 76476 25900
rect 76532 25844 76580 25900
rect 76636 25844 76684 25900
rect 76740 25844 76788 25900
rect 76844 25844 76892 25900
rect 76948 25844 76958 25900
rect 76258 24332 76958 25844
rect 76258 24276 76268 24332
rect 76324 24276 76372 24332
rect 76428 24276 76476 24332
rect 76532 24276 76580 24332
rect 76636 24276 76684 24332
rect 76740 24276 76788 24332
rect 76844 24276 76892 24332
rect 76948 24276 76958 24332
rect 76258 22764 76958 24276
rect 76258 22708 76268 22764
rect 76324 22708 76372 22764
rect 76428 22708 76476 22764
rect 76532 22708 76580 22764
rect 76636 22708 76684 22764
rect 76740 22708 76788 22764
rect 76844 22708 76892 22764
rect 76948 22708 76958 22764
rect 76258 21196 76958 22708
rect 76258 21140 76268 21196
rect 76324 21140 76372 21196
rect 76428 21140 76476 21196
rect 76532 21140 76580 21196
rect 76636 21140 76684 21196
rect 76740 21140 76788 21196
rect 76844 21140 76892 21196
rect 76948 21140 76958 21196
rect 76258 19628 76958 21140
rect 76258 19572 76268 19628
rect 76324 19572 76372 19628
rect 76428 19572 76476 19628
rect 76532 19572 76580 19628
rect 76636 19572 76684 19628
rect 76740 19572 76788 19628
rect 76844 19572 76892 19628
rect 76948 19572 76958 19628
rect 76258 18060 76958 19572
rect 76258 18004 76268 18060
rect 76324 18004 76372 18060
rect 76428 18004 76476 18060
rect 76532 18004 76580 18060
rect 76636 18004 76684 18060
rect 76740 18004 76788 18060
rect 76844 18004 76892 18060
rect 76948 18004 76958 18060
rect 76258 16492 76958 18004
rect 76258 16436 76268 16492
rect 76324 16436 76372 16492
rect 76428 16436 76476 16492
rect 76532 16436 76580 16492
rect 76636 16436 76684 16492
rect 76740 16436 76788 16492
rect 76844 16436 76892 16492
rect 76948 16436 76958 16492
rect 76258 14924 76958 16436
rect 76258 14868 76268 14924
rect 76324 14868 76372 14924
rect 76428 14868 76476 14924
rect 76532 14868 76580 14924
rect 76636 14868 76684 14924
rect 76740 14868 76788 14924
rect 76844 14868 76892 14924
rect 76948 14868 76958 14924
rect 76258 13356 76958 14868
rect 76258 13300 76268 13356
rect 76324 13300 76372 13356
rect 76428 13300 76476 13356
rect 76532 13300 76580 13356
rect 76636 13300 76684 13356
rect 76740 13300 76788 13356
rect 76844 13300 76892 13356
rect 76948 13300 76958 13356
rect 76258 11788 76958 13300
rect 76258 11732 76268 11788
rect 76324 11732 76372 11788
rect 76428 11732 76476 11788
rect 76532 11732 76580 11788
rect 76636 11732 76684 11788
rect 76740 11732 76788 11788
rect 76844 11732 76892 11788
rect 76948 11732 76958 11788
rect 76258 10220 76958 11732
rect 76258 10164 76268 10220
rect 76324 10164 76372 10220
rect 76428 10164 76476 10220
rect 76532 10164 76580 10220
rect 76636 10164 76684 10220
rect 76740 10164 76788 10220
rect 76844 10164 76892 10220
rect 76948 10164 76958 10220
rect 76258 8652 76958 10164
rect 76258 8596 76268 8652
rect 76324 8596 76372 8652
rect 76428 8596 76476 8652
rect 76532 8596 76580 8652
rect 76636 8596 76684 8652
rect 76740 8596 76788 8652
rect 76844 8596 76892 8652
rect 76948 8596 76958 8652
rect 76258 7084 76958 8596
rect 76258 7028 76268 7084
rect 76324 7028 76372 7084
rect 76428 7028 76476 7084
rect 76532 7028 76580 7084
rect 76636 7028 76684 7084
rect 76740 7028 76788 7084
rect 76844 7028 76892 7084
rect 76948 7028 76958 7084
rect 76258 5516 76958 7028
rect 76258 5460 76268 5516
rect 76324 5460 76372 5516
rect 76428 5460 76476 5516
rect 76532 5460 76580 5516
rect 76636 5460 76684 5516
rect 76740 5460 76788 5516
rect 76844 5460 76892 5516
rect 76948 5460 76958 5516
rect 71758 4676 71768 4732
rect 71824 4676 71872 4732
rect 71928 4676 71976 4732
rect 72032 4676 72080 4732
rect 72136 4676 72184 4732
rect 72240 4676 72288 4732
rect 72344 4676 72392 4732
rect 72448 4676 72458 4732
rect 71758 3164 72458 4676
rect 75628 4978 75684 4988
rect 75628 4452 75684 4922
rect 75628 4386 75684 4396
rect 71758 3108 71768 3164
rect 71824 3108 71872 3164
rect 71928 3108 71976 3164
rect 72032 3108 72080 3164
rect 72136 3108 72184 3164
rect 72240 3108 72288 3164
rect 72344 3108 72392 3164
rect 72448 3108 72458 3164
rect 71758 3076 72458 3108
rect 76258 3948 76958 5460
rect 76258 3892 76268 3948
rect 76324 3892 76372 3948
rect 76428 3892 76476 3948
rect 76532 3892 76580 3948
rect 76636 3892 76684 3948
rect 76740 3892 76788 3948
rect 76844 3892 76892 3948
rect 76948 3892 76958 3948
rect 76258 3076 76958 3892
rect 80758 56476 81458 56508
rect 80758 56420 80768 56476
rect 80824 56420 80872 56476
rect 80928 56420 80976 56476
rect 81032 56420 81080 56476
rect 81136 56420 81184 56476
rect 81240 56420 81288 56476
rect 81344 56420 81392 56476
rect 81448 56420 81458 56476
rect 80758 54908 81458 56420
rect 80758 54852 80768 54908
rect 80824 54852 80872 54908
rect 80928 54852 80976 54908
rect 81032 54852 81080 54908
rect 81136 54852 81184 54908
rect 81240 54852 81288 54908
rect 81344 54852 81392 54908
rect 81448 54852 81458 54908
rect 80758 53340 81458 54852
rect 80758 53284 80768 53340
rect 80824 53284 80872 53340
rect 80928 53284 80976 53340
rect 81032 53284 81080 53340
rect 81136 53284 81184 53340
rect 81240 53284 81288 53340
rect 81344 53284 81392 53340
rect 81448 53284 81458 53340
rect 80758 51772 81458 53284
rect 80758 51716 80768 51772
rect 80824 51716 80872 51772
rect 80928 51716 80976 51772
rect 81032 51716 81080 51772
rect 81136 51716 81184 51772
rect 81240 51716 81288 51772
rect 81344 51716 81392 51772
rect 81448 51716 81458 51772
rect 80758 50204 81458 51716
rect 80758 50148 80768 50204
rect 80824 50148 80872 50204
rect 80928 50148 80976 50204
rect 81032 50148 81080 50204
rect 81136 50148 81184 50204
rect 81240 50148 81288 50204
rect 81344 50148 81392 50204
rect 81448 50148 81458 50204
rect 80758 48636 81458 50148
rect 80758 48580 80768 48636
rect 80824 48580 80872 48636
rect 80928 48580 80976 48636
rect 81032 48580 81080 48636
rect 81136 48580 81184 48636
rect 81240 48580 81288 48636
rect 81344 48580 81392 48636
rect 81448 48580 81458 48636
rect 80758 47068 81458 48580
rect 80758 47012 80768 47068
rect 80824 47012 80872 47068
rect 80928 47012 80976 47068
rect 81032 47012 81080 47068
rect 81136 47012 81184 47068
rect 81240 47012 81288 47068
rect 81344 47012 81392 47068
rect 81448 47012 81458 47068
rect 80758 45500 81458 47012
rect 80758 45444 80768 45500
rect 80824 45444 80872 45500
rect 80928 45444 80976 45500
rect 81032 45444 81080 45500
rect 81136 45444 81184 45500
rect 81240 45444 81288 45500
rect 81344 45444 81392 45500
rect 81448 45444 81458 45500
rect 80758 43932 81458 45444
rect 80758 43876 80768 43932
rect 80824 43876 80872 43932
rect 80928 43876 80976 43932
rect 81032 43876 81080 43932
rect 81136 43876 81184 43932
rect 81240 43876 81288 43932
rect 81344 43876 81392 43932
rect 81448 43876 81458 43932
rect 80758 42364 81458 43876
rect 80758 42308 80768 42364
rect 80824 42308 80872 42364
rect 80928 42308 80976 42364
rect 81032 42308 81080 42364
rect 81136 42308 81184 42364
rect 81240 42308 81288 42364
rect 81344 42308 81392 42364
rect 81448 42308 81458 42364
rect 80758 40796 81458 42308
rect 80758 40740 80768 40796
rect 80824 40740 80872 40796
rect 80928 40740 80976 40796
rect 81032 40740 81080 40796
rect 81136 40740 81184 40796
rect 81240 40740 81288 40796
rect 81344 40740 81392 40796
rect 81448 40740 81458 40796
rect 80758 39228 81458 40740
rect 80758 39172 80768 39228
rect 80824 39172 80872 39228
rect 80928 39172 80976 39228
rect 81032 39172 81080 39228
rect 81136 39172 81184 39228
rect 81240 39172 81288 39228
rect 81344 39172 81392 39228
rect 81448 39172 81458 39228
rect 80758 37660 81458 39172
rect 80758 37604 80768 37660
rect 80824 37604 80872 37660
rect 80928 37604 80976 37660
rect 81032 37604 81080 37660
rect 81136 37604 81184 37660
rect 81240 37604 81288 37660
rect 81344 37604 81392 37660
rect 81448 37604 81458 37660
rect 80758 36092 81458 37604
rect 80758 36036 80768 36092
rect 80824 36036 80872 36092
rect 80928 36036 80976 36092
rect 81032 36036 81080 36092
rect 81136 36036 81184 36092
rect 81240 36036 81288 36092
rect 81344 36036 81392 36092
rect 81448 36036 81458 36092
rect 80758 34524 81458 36036
rect 80758 34468 80768 34524
rect 80824 34468 80872 34524
rect 80928 34468 80976 34524
rect 81032 34468 81080 34524
rect 81136 34468 81184 34524
rect 81240 34468 81288 34524
rect 81344 34468 81392 34524
rect 81448 34468 81458 34524
rect 80758 32956 81458 34468
rect 80758 32900 80768 32956
rect 80824 32900 80872 32956
rect 80928 32900 80976 32956
rect 81032 32900 81080 32956
rect 81136 32900 81184 32956
rect 81240 32900 81288 32956
rect 81344 32900 81392 32956
rect 81448 32900 81458 32956
rect 80758 31388 81458 32900
rect 80758 31332 80768 31388
rect 80824 31332 80872 31388
rect 80928 31332 80976 31388
rect 81032 31332 81080 31388
rect 81136 31332 81184 31388
rect 81240 31332 81288 31388
rect 81344 31332 81392 31388
rect 81448 31332 81458 31388
rect 80758 29820 81458 31332
rect 80758 29764 80768 29820
rect 80824 29764 80872 29820
rect 80928 29764 80976 29820
rect 81032 29764 81080 29820
rect 81136 29764 81184 29820
rect 81240 29764 81288 29820
rect 81344 29764 81392 29820
rect 81448 29764 81458 29820
rect 80758 28252 81458 29764
rect 80758 28196 80768 28252
rect 80824 28196 80872 28252
rect 80928 28196 80976 28252
rect 81032 28196 81080 28252
rect 81136 28196 81184 28252
rect 81240 28196 81288 28252
rect 81344 28196 81392 28252
rect 81448 28196 81458 28252
rect 80758 26684 81458 28196
rect 80758 26628 80768 26684
rect 80824 26628 80872 26684
rect 80928 26628 80976 26684
rect 81032 26628 81080 26684
rect 81136 26628 81184 26684
rect 81240 26628 81288 26684
rect 81344 26628 81392 26684
rect 81448 26628 81458 26684
rect 80758 25116 81458 26628
rect 80758 25060 80768 25116
rect 80824 25060 80872 25116
rect 80928 25060 80976 25116
rect 81032 25060 81080 25116
rect 81136 25060 81184 25116
rect 81240 25060 81288 25116
rect 81344 25060 81392 25116
rect 81448 25060 81458 25116
rect 80758 23548 81458 25060
rect 80758 23492 80768 23548
rect 80824 23492 80872 23548
rect 80928 23492 80976 23548
rect 81032 23492 81080 23548
rect 81136 23492 81184 23548
rect 81240 23492 81288 23548
rect 81344 23492 81392 23548
rect 81448 23492 81458 23548
rect 80758 21980 81458 23492
rect 80758 21924 80768 21980
rect 80824 21924 80872 21980
rect 80928 21924 80976 21980
rect 81032 21924 81080 21980
rect 81136 21924 81184 21980
rect 81240 21924 81288 21980
rect 81344 21924 81392 21980
rect 81448 21924 81458 21980
rect 80758 20412 81458 21924
rect 80758 20356 80768 20412
rect 80824 20356 80872 20412
rect 80928 20356 80976 20412
rect 81032 20356 81080 20412
rect 81136 20356 81184 20412
rect 81240 20356 81288 20412
rect 81344 20356 81392 20412
rect 81448 20356 81458 20412
rect 80758 18844 81458 20356
rect 80758 18788 80768 18844
rect 80824 18788 80872 18844
rect 80928 18788 80976 18844
rect 81032 18788 81080 18844
rect 81136 18788 81184 18844
rect 81240 18788 81288 18844
rect 81344 18788 81392 18844
rect 81448 18788 81458 18844
rect 80758 17276 81458 18788
rect 80758 17220 80768 17276
rect 80824 17220 80872 17276
rect 80928 17220 80976 17276
rect 81032 17220 81080 17276
rect 81136 17220 81184 17276
rect 81240 17220 81288 17276
rect 81344 17220 81392 17276
rect 81448 17220 81458 17276
rect 80758 15708 81458 17220
rect 80758 15652 80768 15708
rect 80824 15652 80872 15708
rect 80928 15652 80976 15708
rect 81032 15652 81080 15708
rect 81136 15652 81184 15708
rect 81240 15652 81288 15708
rect 81344 15652 81392 15708
rect 81448 15652 81458 15708
rect 80758 14140 81458 15652
rect 80758 14084 80768 14140
rect 80824 14084 80872 14140
rect 80928 14084 80976 14140
rect 81032 14084 81080 14140
rect 81136 14084 81184 14140
rect 81240 14084 81288 14140
rect 81344 14084 81392 14140
rect 81448 14084 81458 14140
rect 80758 12572 81458 14084
rect 80758 12516 80768 12572
rect 80824 12516 80872 12572
rect 80928 12516 80976 12572
rect 81032 12516 81080 12572
rect 81136 12516 81184 12572
rect 81240 12516 81288 12572
rect 81344 12516 81392 12572
rect 81448 12516 81458 12572
rect 80758 11004 81458 12516
rect 80758 10948 80768 11004
rect 80824 10948 80872 11004
rect 80928 10948 80976 11004
rect 81032 10948 81080 11004
rect 81136 10948 81184 11004
rect 81240 10948 81288 11004
rect 81344 10948 81392 11004
rect 81448 10948 81458 11004
rect 80758 9436 81458 10948
rect 80758 9380 80768 9436
rect 80824 9380 80872 9436
rect 80928 9380 80976 9436
rect 81032 9380 81080 9436
rect 81136 9380 81184 9436
rect 81240 9380 81288 9436
rect 81344 9380 81392 9436
rect 81448 9380 81458 9436
rect 80758 7868 81458 9380
rect 80758 7812 80768 7868
rect 80824 7812 80872 7868
rect 80928 7812 80976 7868
rect 81032 7812 81080 7868
rect 81136 7812 81184 7868
rect 81240 7812 81288 7868
rect 81344 7812 81392 7868
rect 81448 7812 81458 7868
rect 80758 6300 81458 7812
rect 80758 6244 80768 6300
rect 80824 6244 80872 6300
rect 80928 6244 80976 6300
rect 81032 6244 81080 6300
rect 81136 6244 81184 6300
rect 81240 6244 81288 6300
rect 81344 6244 81392 6300
rect 81448 6244 81458 6300
rect 80758 4732 81458 6244
rect 80758 4676 80768 4732
rect 80824 4676 80872 4732
rect 80928 4676 80976 4732
rect 81032 4676 81080 4732
rect 81136 4676 81184 4732
rect 81240 4676 81288 4732
rect 81344 4676 81392 4732
rect 81448 4676 81458 4732
rect 80758 3164 81458 4676
rect 80758 3108 80768 3164
rect 80824 3108 80872 3164
rect 80928 3108 80976 3164
rect 81032 3108 81080 3164
rect 81136 3108 81184 3164
rect 81240 3108 81288 3164
rect 81344 3108 81392 3164
rect 81448 3108 81458 3164
rect 80758 3076 81458 3108
rect 85258 55692 85958 56508
rect 85258 55636 85268 55692
rect 85324 55636 85372 55692
rect 85428 55636 85476 55692
rect 85532 55636 85580 55692
rect 85636 55636 85684 55692
rect 85740 55636 85788 55692
rect 85844 55636 85892 55692
rect 85948 55636 85958 55692
rect 85258 54124 85958 55636
rect 85258 54068 85268 54124
rect 85324 54068 85372 54124
rect 85428 54068 85476 54124
rect 85532 54068 85580 54124
rect 85636 54068 85684 54124
rect 85740 54068 85788 54124
rect 85844 54068 85892 54124
rect 85948 54068 85958 54124
rect 85258 52556 85958 54068
rect 85258 52500 85268 52556
rect 85324 52500 85372 52556
rect 85428 52500 85476 52556
rect 85532 52500 85580 52556
rect 85636 52500 85684 52556
rect 85740 52500 85788 52556
rect 85844 52500 85892 52556
rect 85948 52500 85958 52556
rect 85258 50988 85958 52500
rect 85258 50932 85268 50988
rect 85324 50932 85372 50988
rect 85428 50932 85476 50988
rect 85532 50932 85580 50988
rect 85636 50932 85684 50988
rect 85740 50932 85788 50988
rect 85844 50932 85892 50988
rect 85948 50932 85958 50988
rect 85258 49420 85958 50932
rect 85258 49364 85268 49420
rect 85324 49364 85372 49420
rect 85428 49364 85476 49420
rect 85532 49364 85580 49420
rect 85636 49364 85684 49420
rect 85740 49364 85788 49420
rect 85844 49364 85892 49420
rect 85948 49364 85958 49420
rect 85258 47852 85958 49364
rect 85258 47796 85268 47852
rect 85324 47796 85372 47852
rect 85428 47796 85476 47852
rect 85532 47796 85580 47852
rect 85636 47796 85684 47852
rect 85740 47796 85788 47852
rect 85844 47796 85892 47852
rect 85948 47796 85958 47852
rect 85258 46284 85958 47796
rect 85258 46228 85268 46284
rect 85324 46228 85372 46284
rect 85428 46228 85476 46284
rect 85532 46228 85580 46284
rect 85636 46228 85684 46284
rect 85740 46228 85788 46284
rect 85844 46228 85892 46284
rect 85948 46228 85958 46284
rect 85258 44716 85958 46228
rect 85258 44660 85268 44716
rect 85324 44660 85372 44716
rect 85428 44660 85476 44716
rect 85532 44660 85580 44716
rect 85636 44660 85684 44716
rect 85740 44660 85788 44716
rect 85844 44660 85892 44716
rect 85948 44660 85958 44716
rect 85258 43148 85958 44660
rect 85258 43092 85268 43148
rect 85324 43092 85372 43148
rect 85428 43092 85476 43148
rect 85532 43092 85580 43148
rect 85636 43092 85684 43148
rect 85740 43092 85788 43148
rect 85844 43092 85892 43148
rect 85948 43092 85958 43148
rect 85258 41580 85958 43092
rect 85258 41524 85268 41580
rect 85324 41524 85372 41580
rect 85428 41524 85476 41580
rect 85532 41524 85580 41580
rect 85636 41524 85684 41580
rect 85740 41524 85788 41580
rect 85844 41524 85892 41580
rect 85948 41524 85958 41580
rect 85258 40012 85958 41524
rect 85258 39956 85268 40012
rect 85324 39956 85372 40012
rect 85428 39956 85476 40012
rect 85532 39956 85580 40012
rect 85636 39956 85684 40012
rect 85740 39956 85788 40012
rect 85844 39956 85892 40012
rect 85948 39956 85958 40012
rect 85258 38444 85958 39956
rect 85258 38388 85268 38444
rect 85324 38388 85372 38444
rect 85428 38388 85476 38444
rect 85532 38388 85580 38444
rect 85636 38388 85684 38444
rect 85740 38388 85788 38444
rect 85844 38388 85892 38444
rect 85948 38388 85958 38444
rect 85258 36876 85958 38388
rect 85258 36820 85268 36876
rect 85324 36820 85372 36876
rect 85428 36820 85476 36876
rect 85532 36820 85580 36876
rect 85636 36820 85684 36876
rect 85740 36820 85788 36876
rect 85844 36820 85892 36876
rect 85948 36820 85958 36876
rect 85258 35308 85958 36820
rect 85258 35252 85268 35308
rect 85324 35252 85372 35308
rect 85428 35252 85476 35308
rect 85532 35252 85580 35308
rect 85636 35252 85684 35308
rect 85740 35252 85788 35308
rect 85844 35252 85892 35308
rect 85948 35252 85958 35308
rect 85258 33740 85958 35252
rect 85258 33684 85268 33740
rect 85324 33684 85372 33740
rect 85428 33684 85476 33740
rect 85532 33684 85580 33740
rect 85636 33684 85684 33740
rect 85740 33684 85788 33740
rect 85844 33684 85892 33740
rect 85948 33684 85958 33740
rect 85258 32172 85958 33684
rect 85258 32116 85268 32172
rect 85324 32116 85372 32172
rect 85428 32116 85476 32172
rect 85532 32116 85580 32172
rect 85636 32116 85684 32172
rect 85740 32116 85788 32172
rect 85844 32116 85892 32172
rect 85948 32116 85958 32172
rect 85258 30604 85958 32116
rect 85258 30548 85268 30604
rect 85324 30548 85372 30604
rect 85428 30548 85476 30604
rect 85532 30548 85580 30604
rect 85636 30548 85684 30604
rect 85740 30548 85788 30604
rect 85844 30548 85892 30604
rect 85948 30548 85958 30604
rect 85258 29036 85958 30548
rect 85258 28980 85268 29036
rect 85324 28980 85372 29036
rect 85428 28980 85476 29036
rect 85532 28980 85580 29036
rect 85636 28980 85684 29036
rect 85740 28980 85788 29036
rect 85844 28980 85892 29036
rect 85948 28980 85958 29036
rect 85258 27468 85958 28980
rect 85258 27412 85268 27468
rect 85324 27412 85372 27468
rect 85428 27412 85476 27468
rect 85532 27412 85580 27468
rect 85636 27412 85684 27468
rect 85740 27412 85788 27468
rect 85844 27412 85892 27468
rect 85948 27412 85958 27468
rect 85258 25900 85958 27412
rect 85258 25844 85268 25900
rect 85324 25844 85372 25900
rect 85428 25844 85476 25900
rect 85532 25844 85580 25900
rect 85636 25844 85684 25900
rect 85740 25844 85788 25900
rect 85844 25844 85892 25900
rect 85948 25844 85958 25900
rect 85258 24332 85958 25844
rect 85258 24276 85268 24332
rect 85324 24276 85372 24332
rect 85428 24276 85476 24332
rect 85532 24276 85580 24332
rect 85636 24276 85684 24332
rect 85740 24276 85788 24332
rect 85844 24276 85892 24332
rect 85948 24276 85958 24332
rect 85258 22764 85958 24276
rect 85258 22708 85268 22764
rect 85324 22708 85372 22764
rect 85428 22708 85476 22764
rect 85532 22708 85580 22764
rect 85636 22708 85684 22764
rect 85740 22708 85788 22764
rect 85844 22708 85892 22764
rect 85948 22708 85958 22764
rect 85258 21196 85958 22708
rect 85258 21140 85268 21196
rect 85324 21140 85372 21196
rect 85428 21140 85476 21196
rect 85532 21140 85580 21196
rect 85636 21140 85684 21196
rect 85740 21140 85788 21196
rect 85844 21140 85892 21196
rect 85948 21140 85958 21196
rect 85258 19628 85958 21140
rect 85258 19572 85268 19628
rect 85324 19572 85372 19628
rect 85428 19572 85476 19628
rect 85532 19572 85580 19628
rect 85636 19572 85684 19628
rect 85740 19572 85788 19628
rect 85844 19572 85892 19628
rect 85948 19572 85958 19628
rect 85258 18060 85958 19572
rect 85258 18004 85268 18060
rect 85324 18004 85372 18060
rect 85428 18004 85476 18060
rect 85532 18004 85580 18060
rect 85636 18004 85684 18060
rect 85740 18004 85788 18060
rect 85844 18004 85892 18060
rect 85948 18004 85958 18060
rect 85258 16492 85958 18004
rect 85258 16436 85268 16492
rect 85324 16436 85372 16492
rect 85428 16436 85476 16492
rect 85532 16436 85580 16492
rect 85636 16436 85684 16492
rect 85740 16436 85788 16492
rect 85844 16436 85892 16492
rect 85948 16436 85958 16492
rect 85258 14924 85958 16436
rect 85258 14868 85268 14924
rect 85324 14868 85372 14924
rect 85428 14868 85476 14924
rect 85532 14868 85580 14924
rect 85636 14868 85684 14924
rect 85740 14868 85788 14924
rect 85844 14868 85892 14924
rect 85948 14868 85958 14924
rect 85258 13356 85958 14868
rect 85258 13300 85268 13356
rect 85324 13300 85372 13356
rect 85428 13300 85476 13356
rect 85532 13300 85580 13356
rect 85636 13300 85684 13356
rect 85740 13300 85788 13356
rect 85844 13300 85892 13356
rect 85948 13300 85958 13356
rect 85258 11788 85958 13300
rect 85258 11732 85268 11788
rect 85324 11732 85372 11788
rect 85428 11732 85476 11788
rect 85532 11732 85580 11788
rect 85636 11732 85684 11788
rect 85740 11732 85788 11788
rect 85844 11732 85892 11788
rect 85948 11732 85958 11788
rect 85258 10220 85958 11732
rect 85258 10164 85268 10220
rect 85324 10164 85372 10220
rect 85428 10164 85476 10220
rect 85532 10164 85580 10220
rect 85636 10164 85684 10220
rect 85740 10164 85788 10220
rect 85844 10164 85892 10220
rect 85948 10164 85958 10220
rect 85258 8652 85958 10164
rect 85258 8596 85268 8652
rect 85324 8596 85372 8652
rect 85428 8596 85476 8652
rect 85532 8596 85580 8652
rect 85636 8596 85684 8652
rect 85740 8596 85788 8652
rect 85844 8596 85892 8652
rect 85948 8596 85958 8652
rect 85258 7084 85958 8596
rect 85258 7028 85268 7084
rect 85324 7028 85372 7084
rect 85428 7028 85476 7084
rect 85532 7028 85580 7084
rect 85636 7028 85684 7084
rect 85740 7028 85788 7084
rect 85844 7028 85892 7084
rect 85948 7028 85958 7084
rect 85258 5516 85958 7028
rect 85258 5460 85268 5516
rect 85324 5460 85372 5516
rect 85428 5460 85476 5516
rect 85532 5460 85580 5516
rect 85636 5460 85684 5516
rect 85740 5460 85788 5516
rect 85844 5460 85892 5516
rect 85948 5460 85958 5516
rect 85258 3948 85958 5460
rect 85258 3892 85268 3948
rect 85324 3892 85372 3948
rect 85428 3892 85476 3948
rect 85532 3892 85580 3948
rect 85636 3892 85684 3948
rect 85740 3892 85788 3948
rect 85844 3892 85892 3948
rect 85948 3892 85958 3948
rect 85258 3076 85958 3892
rect 89758 56476 90458 56508
rect 89758 56420 89768 56476
rect 89824 56420 89872 56476
rect 89928 56420 89976 56476
rect 90032 56420 90080 56476
rect 90136 56420 90184 56476
rect 90240 56420 90288 56476
rect 90344 56420 90392 56476
rect 90448 56420 90458 56476
rect 89758 54908 90458 56420
rect 89758 54852 89768 54908
rect 89824 54852 89872 54908
rect 89928 54852 89976 54908
rect 90032 54852 90080 54908
rect 90136 54852 90184 54908
rect 90240 54852 90288 54908
rect 90344 54852 90392 54908
rect 90448 54852 90458 54908
rect 89758 53340 90458 54852
rect 89758 53284 89768 53340
rect 89824 53284 89872 53340
rect 89928 53284 89976 53340
rect 90032 53284 90080 53340
rect 90136 53284 90184 53340
rect 90240 53284 90288 53340
rect 90344 53284 90392 53340
rect 90448 53284 90458 53340
rect 89758 51772 90458 53284
rect 89758 51716 89768 51772
rect 89824 51716 89872 51772
rect 89928 51716 89976 51772
rect 90032 51716 90080 51772
rect 90136 51716 90184 51772
rect 90240 51716 90288 51772
rect 90344 51716 90392 51772
rect 90448 51716 90458 51772
rect 89758 50204 90458 51716
rect 89758 50148 89768 50204
rect 89824 50148 89872 50204
rect 89928 50148 89976 50204
rect 90032 50148 90080 50204
rect 90136 50148 90184 50204
rect 90240 50148 90288 50204
rect 90344 50148 90392 50204
rect 90448 50148 90458 50204
rect 89758 48636 90458 50148
rect 89758 48580 89768 48636
rect 89824 48580 89872 48636
rect 89928 48580 89976 48636
rect 90032 48580 90080 48636
rect 90136 48580 90184 48636
rect 90240 48580 90288 48636
rect 90344 48580 90392 48636
rect 90448 48580 90458 48636
rect 89758 47068 90458 48580
rect 89758 47012 89768 47068
rect 89824 47012 89872 47068
rect 89928 47012 89976 47068
rect 90032 47012 90080 47068
rect 90136 47012 90184 47068
rect 90240 47012 90288 47068
rect 90344 47012 90392 47068
rect 90448 47012 90458 47068
rect 89758 45500 90458 47012
rect 89758 45444 89768 45500
rect 89824 45444 89872 45500
rect 89928 45444 89976 45500
rect 90032 45444 90080 45500
rect 90136 45444 90184 45500
rect 90240 45444 90288 45500
rect 90344 45444 90392 45500
rect 90448 45444 90458 45500
rect 89758 43932 90458 45444
rect 89758 43876 89768 43932
rect 89824 43876 89872 43932
rect 89928 43876 89976 43932
rect 90032 43876 90080 43932
rect 90136 43876 90184 43932
rect 90240 43876 90288 43932
rect 90344 43876 90392 43932
rect 90448 43876 90458 43932
rect 89758 42364 90458 43876
rect 89758 42308 89768 42364
rect 89824 42308 89872 42364
rect 89928 42308 89976 42364
rect 90032 42308 90080 42364
rect 90136 42308 90184 42364
rect 90240 42308 90288 42364
rect 90344 42308 90392 42364
rect 90448 42308 90458 42364
rect 89758 40796 90458 42308
rect 89758 40740 89768 40796
rect 89824 40740 89872 40796
rect 89928 40740 89976 40796
rect 90032 40740 90080 40796
rect 90136 40740 90184 40796
rect 90240 40740 90288 40796
rect 90344 40740 90392 40796
rect 90448 40740 90458 40796
rect 89758 39228 90458 40740
rect 89758 39172 89768 39228
rect 89824 39172 89872 39228
rect 89928 39172 89976 39228
rect 90032 39172 90080 39228
rect 90136 39172 90184 39228
rect 90240 39172 90288 39228
rect 90344 39172 90392 39228
rect 90448 39172 90458 39228
rect 89758 37660 90458 39172
rect 89758 37604 89768 37660
rect 89824 37604 89872 37660
rect 89928 37604 89976 37660
rect 90032 37604 90080 37660
rect 90136 37604 90184 37660
rect 90240 37604 90288 37660
rect 90344 37604 90392 37660
rect 90448 37604 90458 37660
rect 89758 36092 90458 37604
rect 89758 36036 89768 36092
rect 89824 36036 89872 36092
rect 89928 36036 89976 36092
rect 90032 36036 90080 36092
rect 90136 36036 90184 36092
rect 90240 36036 90288 36092
rect 90344 36036 90392 36092
rect 90448 36036 90458 36092
rect 89758 34524 90458 36036
rect 89758 34468 89768 34524
rect 89824 34468 89872 34524
rect 89928 34468 89976 34524
rect 90032 34468 90080 34524
rect 90136 34468 90184 34524
rect 90240 34468 90288 34524
rect 90344 34468 90392 34524
rect 90448 34468 90458 34524
rect 89758 32956 90458 34468
rect 89758 32900 89768 32956
rect 89824 32900 89872 32956
rect 89928 32900 89976 32956
rect 90032 32900 90080 32956
rect 90136 32900 90184 32956
rect 90240 32900 90288 32956
rect 90344 32900 90392 32956
rect 90448 32900 90458 32956
rect 89758 31388 90458 32900
rect 89758 31332 89768 31388
rect 89824 31332 89872 31388
rect 89928 31332 89976 31388
rect 90032 31332 90080 31388
rect 90136 31332 90184 31388
rect 90240 31332 90288 31388
rect 90344 31332 90392 31388
rect 90448 31332 90458 31388
rect 89758 29820 90458 31332
rect 89758 29764 89768 29820
rect 89824 29764 89872 29820
rect 89928 29764 89976 29820
rect 90032 29764 90080 29820
rect 90136 29764 90184 29820
rect 90240 29764 90288 29820
rect 90344 29764 90392 29820
rect 90448 29764 90458 29820
rect 89758 28252 90458 29764
rect 89758 28196 89768 28252
rect 89824 28196 89872 28252
rect 89928 28196 89976 28252
rect 90032 28196 90080 28252
rect 90136 28196 90184 28252
rect 90240 28196 90288 28252
rect 90344 28196 90392 28252
rect 90448 28196 90458 28252
rect 89758 26684 90458 28196
rect 89758 26628 89768 26684
rect 89824 26628 89872 26684
rect 89928 26628 89976 26684
rect 90032 26628 90080 26684
rect 90136 26628 90184 26684
rect 90240 26628 90288 26684
rect 90344 26628 90392 26684
rect 90448 26628 90458 26684
rect 89758 25116 90458 26628
rect 89758 25060 89768 25116
rect 89824 25060 89872 25116
rect 89928 25060 89976 25116
rect 90032 25060 90080 25116
rect 90136 25060 90184 25116
rect 90240 25060 90288 25116
rect 90344 25060 90392 25116
rect 90448 25060 90458 25116
rect 89758 23548 90458 25060
rect 89758 23492 89768 23548
rect 89824 23492 89872 23548
rect 89928 23492 89976 23548
rect 90032 23492 90080 23548
rect 90136 23492 90184 23548
rect 90240 23492 90288 23548
rect 90344 23492 90392 23548
rect 90448 23492 90458 23548
rect 89758 21980 90458 23492
rect 89758 21924 89768 21980
rect 89824 21924 89872 21980
rect 89928 21924 89976 21980
rect 90032 21924 90080 21980
rect 90136 21924 90184 21980
rect 90240 21924 90288 21980
rect 90344 21924 90392 21980
rect 90448 21924 90458 21980
rect 89758 20412 90458 21924
rect 89758 20356 89768 20412
rect 89824 20356 89872 20412
rect 89928 20356 89976 20412
rect 90032 20356 90080 20412
rect 90136 20356 90184 20412
rect 90240 20356 90288 20412
rect 90344 20356 90392 20412
rect 90448 20356 90458 20412
rect 89758 18844 90458 20356
rect 89758 18788 89768 18844
rect 89824 18788 89872 18844
rect 89928 18788 89976 18844
rect 90032 18788 90080 18844
rect 90136 18788 90184 18844
rect 90240 18788 90288 18844
rect 90344 18788 90392 18844
rect 90448 18788 90458 18844
rect 89758 17276 90458 18788
rect 89758 17220 89768 17276
rect 89824 17220 89872 17276
rect 89928 17220 89976 17276
rect 90032 17220 90080 17276
rect 90136 17220 90184 17276
rect 90240 17220 90288 17276
rect 90344 17220 90392 17276
rect 90448 17220 90458 17276
rect 89758 15708 90458 17220
rect 89758 15652 89768 15708
rect 89824 15652 89872 15708
rect 89928 15652 89976 15708
rect 90032 15652 90080 15708
rect 90136 15652 90184 15708
rect 90240 15652 90288 15708
rect 90344 15652 90392 15708
rect 90448 15652 90458 15708
rect 89758 14140 90458 15652
rect 89758 14084 89768 14140
rect 89824 14084 89872 14140
rect 89928 14084 89976 14140
rect 90032 14084 90080 14140
rect 90136 14084 90184 14140
rect 90240 14084 90288 14140
rect 90344 14084 90392 14140
rect 90448 14084 90458 14140
rect 89758 12572 90458 14084
rect 89758 12516 89768 12572
rect 89824 12516 89872 12572
rect 89928 12516 89976 12572
rect 90032 12516 90080 12572
rect 90136 12516 90184 12572
rect 90240 12516 90288 12572
rect 90344 12516 90392 12572
rect 90448 12516 90458 12572
rect 89758 11004 90458 12516
rect 89758 10948 89768 11004
rect 89824 10948 89872 11004
rect 89928 10948 89976 11004
rect 90032 10948 90080 11004
rect 90136 10948 90184 11004
rect 90240 10948 90288 11004
rect 90344 10948 90392 11004
rect 90448 10948 90458 11004
rect 89758 9436 90458 10948
rect 89758 9380 89768 9436
rect 89824 9380 89872 9436
rect 89928 9380 89976 9436
rect 90032 9380 90080 9436
rect 90136 9380 90184 9436
rect 90240 9380 90288 9436
rect 90344 9380 90392 9436
rect 90448 9380 90458 9436
rect 89758 7868 90458 9380
rect 89758 7812 89768 7868
rect 89824 7812 89872 7868
rect 89928 7812 89976 7868
rect 90032 7812 90080 7868
rect 90136 7812 90184 7868
rect 90240 7812 90288 7868
rect 90344 7812 90392 7868
rect 90448 7812 90458 7868
rect 89758 6300 90458 7812
rect 89758 6244 89768 6300
rect 89824 6244 89872 6300
rect 89928 6244 89976 6300
rect 90032 6244 90080 6300
rect 90136 6244 90184 6300
rect 90240 6244 90288 6300
rect 90344 6244 90392 6300
rect 90448 6244 90458 6300
rect 89758 4732 90458 6244
rect 89758 4676 89768 4732
rect 89824 4676 89872 4732
rect 89928 4676 89976 4732
rect 90032 4676 90080 4732
rect 90136 4676 90184 4732
rect 90240 4676 90288 4732
rect 90344 4676 90392 4732
rect 90448 4676 90458 4732
rect 89758 3164 90458 4676
rect 89758 3108 89768 3164
rect 89824 3108 89872 3164
rect 89928 3108 89976 3164
rect 90032 3108 90080 3164
rect 90136 3108 90184 3164
rect 90240 3108 90288 3164
rect 90344 3108 90392 3164
rect 90448 3108 90458 3164
rect 89758 3076 90458 3108
rect 94258 55692 94958 56508
rect 94258 55636 94268 55692
rect 94324 55636 94372 55692
rect 94428 55636 94476 55692
rect 94532 55636 94580 55692
rect 94636 55636 94684 55692
rect 94740 55636 94788 55692
rect 94844 55636 94892 55692
rect 94948 55636 94958 55692
rect 94258 54124 94958 55636
rect 94258 54068 94268 54124
rect 94324 54068 94372 54124
rect 94428 54068 94476 54124
rect 94532 54068 94580 54124
rect 94636 54068 94684 54124
rect 94740 54068 94788 54124
rect 94844 54068 94892 54124
rect 94948 54068 94958 54124
rect 94258 52556 94958 54068
rect 94258 52500 94268 52556
rect 94324 52500 94372 52556
rect 94428 52500 94476 52556
rect 94532 52500 94580 52556
rect 94636 52500 94684 52556
rect 94740 52500 94788 52556
rect 94844 52500 94892 52556
rect 94948 52500 94958 52556
rect 94258 50988 94958 52500
rect 94258 50932 94268 50988
rect 94324 50932 94372 50988
rect 94428 50932 94476 50988
rect 94532 50932 94580 50988
rect 94636 50932 94684 50988
rect 94740 50932 94788 50988
rect 94844 50932 94892 50988
rect 94948 50932 94958 50988
rect 94258 49420 94958 50932
rect 94258 49364 94268 49420
rect 94324 49364 94372 49420
rect 94428 49364 94476 49420
rect 94532 49364 94580 49420
rect 94636 49364 94684 49420
rect 94740 49364 94788 49420
rect 94844 49364 94892 49420
rect 94948 49364 94958 49420
rect 94258 47852 94958 49364
rect 94258 47796 94268 47852
rect 94324 47796 94372 47852
rect 94428 47796 94476 47852
rect 94532 47796 94580 47852
rect 94636 47796 94684 47852
rect 94740 47796 94788 47852
rect 94844 47796 94892 47852
rect 94948 47796 94958 47852
rect 94258 46284 94958 47796
rect 94258 46228 94268 46284
rect 94324 46228 94372 46284
rect 94428 46228 94476 46284
rect 94532 46228 94580 46284
rect 94636 46228 94684 46284
rect 94740 46228 94788 46284
rect 94844 46228 94892 46284
rect 94948 46228 94958 46284
rect 94258 44716 94958 46228
rect 94258 44660 94268 44716
rect 94324 44660 94372 44716
rect 94428 44660 94476 44716
rect 94532 44660 94580 44716
rect 94636 44660 94684 44716
rect 94740 44660 94788 44716
rect 94844 44660 94892 44716
rect 94948 44660 94958 44716
rect 94258 43148 94958 44660
rect 94258 43092 94268 43148
rect 94324 43092 94372 43148
rect 94428 43092 94476 43148
rect 94532 43092 94580 43148
rect 94636 43092 94684 43148
rect 94740 43092 94788 43148
rect 94844 43092 94892 43148
rect 94948 43092 94958 43148
rect 94258 41580 94958 43092
rect 94258 41524 94268 41580
rect 94324 41524 94372 41580
rect 94428 41524 94476 41580
rect 94532 41524 94580 41580
rect 94636 41524 94684 41580
rect 94740 41524 94788 41580
rect 94844 41524 94892 41580
rect 94948 41524 94958 41580
rect 94258 40012 94958 41524
rect 94258 39956 94268 40012
rect 94324 39956 94372 40012
rect 94428 39956 94476 40012
rect 94532 39956 94580 40012
rect 94636 39956 94684 40012
rect 94740 39956 94788 40012
rect 94844 39956 94892 40012
rect 94948 39956 94958 40012
rect 94258 38444 94958 39956
rect 94258 38388 94268 38444
rect 94324 38388 94372 38444
rect 94428 38388 94476 38444
rect 94532 38388 94580 38444
rect 94636 38388 94684 38444
rect 94740 38388 94788 38444
rect 94844 38388 94892 38444
rect 94948 38388 94958 38444
rect 94258 36876 94958 38388
rect 94258 36820 94268 36876
rect 94324 36820 94372 36876
rect 94428 36820 94476 36876
rect 94532 36820 94580 36876
rect 94636 36820 94684 36876
rect 94740 36820 94788 36876
rect 94844 36820 94892 36876
rect 94948 36820 94958 36876
rect 94258 35308 94958 36820
rect 94258 35252 94268 35308
rect 94324 35252 94372 35308
rect 94428 35252 94476 35308
rect 94532 35252 94580 35308
rect 94636 35252 94684 35308
rect 94740 35252 94788 35308
rect 94844 35252 94892 35308
rect 94948 35252 94958 35308
rect 94258 33740 94958 35252
rect 94258 33684 94268 33740
rect 94324 33684 94372 33740
rect 94428 33684 94476 33740
rect 94532 33684 94580 33740
rect 94636 33684 94684 33740
rect 94740 33684 94788 33740
rect 94844 33684 94892 33740
rect 94948 33684 94958 33740
rect 94258 32172 94958 33684
rect 94258 32116 94268 32172
rect 94324 32116 94372 32172
rect 94428 32116 94476 32172
rect 94532 32116 94580 32172
rect 94636 32116 94684 32172
rect 94740 32116 94788 32172
rect 94844 32116 94892 32172
rect 94948 32116 94958 32172
rect 94258 30604 94958 32116
rect 94258 30548 94268 30604
rect 94324 30548 94372 30604
rect 94428 30548 94476 30604
rect 94532 30548 94580 30604
rect 94636 30548 94684 30604
rect 94740 30548 94788 30604
rect 94844 30548 94892 30604
rect 94948 30548 94958 30604
rect 94258 29036 94958 30548
rect 94258 28980 94268 29036
rect 94324 28980 94372 29036
rect 94428 28980 94476 29036
rect 94532 28980 94580 29036
rect 94636 28980 94684 29036
rect 94740 28980 94788 29036
rect 94844 28980 94892 29036
rect 94948 28980 94958 29036
rect 94258 27468 94958 28980
rect 94258 27412 94268 27468
rect 94324 27412 94372 27468
rect 94428 27412 94476 27468
rect 94532 27412 94580 27468
rect 94636 27412 94684 27468
rect 94740 27412 94788 27468
rect 94844 27412 94892 27468
rect 94948 27412 94958 27468
rect 94258 25900 94958 27412
rect 94258 25844 94268 25900
rect 94324 25844 94372 25900
rect 94428 25844 94476 25900
rect 94532 25844 94580 25900
rect 94636 25844 94684 25900
rect 94740 25844 94788 25900
rect 94844 25844 94892 25900
rect 94948 25844 94958 25900
rect 94258 24332 94958 25844
rect 94258 24276 94268 24332
rect 94324 24276 94372 24332
rect 94428 24276 94476 24332
rect 94532 24276 94580 24332
rect 94636 24276 94684 24332
rect 94740 24276 94788 24332
rect 94844 24276 94892 24332
rect 94948 24276 94958 24332
rect 94258 22764 94958 24276
rect 94258 22708 94268 22764
rect 94324 22708 94372 22764
rect 94428 22708 94476 22764
rect 94532 22708 94580 22764
rect 94636 22708 94684 22764
rect 94740 22708 94788 22764
rect 94844 22708 94892 22764
rect 94948 22708 94958 22764
rect 94258 21196 94958 22708
rect 94258 21140 94268 21196
rect 94324 21140 94372 21196
rect 94428 21140 94476 21196
rect 94532 21140 94580 21196
rect 94636 21140 94684 21196
rect 94740 21140 94788 21196
rect 94844 21140 94892 21196
rect 94948 21140 94958 21196
rect 94258 19628 94958 21140
rect 94258 19572 94268 19628
rect 94324 19572 94372 19628
rect 94428 19572 94476 19628
rect 94532 19572 94580 19628
rect 94636 19572 94684 19628
rect 94740 19572 94788 19628
rect 94844 19572 94892 19628
rect 94948 19572 94958 19628
rect 94258 18060 94958 19572
rect 94258 18004 94268 18060
rect 94324 18004 94372 18060
rect 94428 18004 94476 18060
rect 94532 18004 94580 18060
rect 94636 18004 94684 18060
rect 94740 18004 94788 18060
rect 94844 18004 94892 18060
rect 94948 18004 94958 18060
rect 94258 16492 94958 18004
rect 94258 16436 94268 16492
rect 94324 16436 94372 16492
rect 94428 16436 94476 16492
rect 94532 16436 94580 16492
rect 94636 16436 94684 16492
rect 94740 16436 94788 16492
rect 94844 16436 94892 16492
rect 94948 16436 94958 16492
rect 94258 14924 94958 16436
rect 94258 14868 94268 14924
rect 94324 14868 94372 14924
rect 94428 14868 94476 14924
rect 94532 14868 94580 14924
rect 94636 14868 94684 14924
rect 94740 14868 94788 14924
rect 94844 14868 94892 14924
rect 94948 14868 94958 14924
rect 94258 13356 94958 14868
rect 94258 13300 94268 13356
rect 94324 13300 94372 13356
rect 94428 13300 94476 13356
rect 94532 13300 94580 13356
rect 94636 13300 94684 13356
rect 94740 13300 94788 13356
rect 94844 13300 94892 13356
rect 94948 13300 94958 13356
rect 94258 11788 94958 13300
rect 94258 11732 94268 11788
rect 94324 11732 94372 11788
rect 94428 11732 94476 11788
rect 94532 11732 94580 11788
rect 94636 11732 94684 11788
rect 94740 11732 94788 11788
rect 94844 11732 94892 11788
rect 94948 11732 94958 11788
rect 94258 10220 94958 11732
rect 94258 10164 94268 10220
rect 94324 10164 94372 10220
rect 94428 10164 94476 10220
rect 94532 10164 94580 10220
rect 94636 10164 94684 10220
rect 94740 10164 94788 10220
rect 94844 10164 94892 10220
rect 94948 10164 94958 10220
rect 94258 8652 94958 10164
rect 94258 8596 94268 8652
rect 94324 8596 94372 8652
rect 94428 8596 94476 8652
rect 94532 8596 94580 8652
rect 94636 8596 94684 8652
rect 94740 8596 94788 8652
rect 94844 8596 94892 8652
rect 94948 8596 94958 8652
rect 94258 7084 94958 8596
rect 94258 7028 94268 7084
rect 94324 7028 94372 7084
rect 94428 7028 94476 7084
rect 94532 7028 94580 7084
rect 94636 7028 94684 7084
rect 94740 7028 94788 7084
rect 94844 7028 94892 7084
rect 94948 7028 94958 7084
rect 94258 5516 94958 7028
rect 94258 5460 94268 5516
rect 94324 5460 94372 5516
rect 94428 5460 94476 5516
rect 94532 5460 94580 5516
rect 94636 5460 94684 5516
rect 94740 5460 94788 5516
rect 94844 5460 94892 5516
rect 94948 5460 94958 5516
rect 94258 3948 94958 5460
rect 94258 3892 94268 3948
rect 94324 3892 94372 3948
rect 94428 3892 94476 3948
rect 94532 3892 94580 3948
rect 94636 3892 94684 3948
rect 94740 3892 94788 3948
rect 94844 3892 94892 3948
rect 94948 3892 94958 3948
rect 94258 3076 94958 3892
<< via4 >>
rect 59612 4956 59668 4978
rect 59612 4922 59668 4956
rect 75628 4922 75684 4978
<< metal5 >>
rect 59596 4978 75700 4994
rect 59596 4922 59612 4978
rect 59668 4922 75628 4978
rect 75684 4922 75700 4978
rect 59596 4906 75700 4922
use gf180mcu_fd_sc_mcu7t5v0__mux4_2  _07_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 51072 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _08__25 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 46256 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _09_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 46592 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _10_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 44912 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _11_
timestamp 1698175906
transform -1 0 49056 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _12_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 44688 0 1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_4  _13_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 44800 0 1 14112
box -86 -86 4006 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _15_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 95984 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _16_
timestamp 1698175906
transform 1 0 90496 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _17_
timestamp 1698175906
transform 1 0 96096 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _18_
timestamp 1698175906
transform 1 0 96096 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _19_
timestamp 1698175906
transform 1 0 96096 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _20_
timestamp 1698175906
transform 1 0 96096 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _21_
timestamp 1698175906
transform 1 0 95424 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _22_
timestamp 1698175906
transform 1 0 96096 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _23_
timestamp 1698175906
transform 1 0 96096 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _24_
timestamp 1698175906
transform 1 0 96096 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _25_
timestamp 1698175906
transform 1 0 96096 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _26_
timestamp 1698175906
transform 1 0 96096 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _27_
timestamp 1698175906
transform 1 0 96096 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _28_
timestamp 1698175906
transform 1 0 76048 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _29_
timestamp 1698175906
transform 1 0 73920 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _30_
timestamp 1698175906
transform 1 0 72352 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _31_
timestamp 1698175906
transform 1 0 72240 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _32_
timestamp 1698175906
transform 1 0 67088 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _33_
timestamp 1698175906
transform 1 0 83776 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _34_
timestamp 1698175906
transform 1 0 76160 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _35_
timestamp 1698175906
transform 1 0 66192 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _36_
timestamp 1698175906
transform 1 0 71008 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _37_
timestamp 1698175906
transform 1 0 82992 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _38_
timestamp 1698175906
transform 1 0 65744 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _39_
timestamp 1698175906
transform 1 0 82656 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _40_
timestamp 1698175906
transform 1 0 72128 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _41_
timestamp 1698175906
transform 1 0 77728 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _42_
timestamp 1698175906
transform 1 0 86912 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _43_
timestamp 1698175906
transform 1 0 89824 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _44_
timestamp 1698175906
transform 1 0 80080 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _45_
timestamp 1698175906
transform 1 0 75040 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _46_
timestamp 1698175906
transform 1 0 85568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _47_
timestamp 1698175906
transform 1 0 81648 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _48_
timestamp 1698175906
transform 1 0 68208 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _49_
timestamp 1698175906
transform 1 0 66640 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _50_
timestamp 1698175906
transform 1 0 55552 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _51_
timestamp 1698175906
transform 1 0 42784 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _52_
timestamp 1698175906
transform -1 0 32928 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _53_
timestamp 1698175906
transform -1 0 25984 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _54_
timestamp 1698175906
transform -1 0 26656 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__07__S0 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 55104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__07__S1
timestamp 1698175906
transform 1 0 55552 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__09__A1
timestamp 1698175906
transform -1 0 45472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__10__I
timestamp 1698175906
transform 1 0 45360 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__11__I
timestamp 1698175906
transform -1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__12__B
timestamp 1698175906
transform -1 0 42784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__13__A1
timestamp 1698175906
transform 1 0 44240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__47__I
timestamp 1698175906
transform 1 0 81424 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 52080 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_COMP_1.net2_I
timestamp 1698175906
transform 1 0 82320 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_CTRL.cmp_I
timestamp 1698175906
transform 1 0 49616 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_0__f_COMP_1.net2_I
timestamp 1698175906
transform 1 0 74256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_0__f_COMP_2.net4_I
timestamp 1698175906
transform 1 0 66528 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_0__f_COMP_4.net2_I
timestamp 1698175906
transform -1 0 31360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_1__f_COMP_1.net2_I
timestamp 1698175906
transform 1 0 81872 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_1__f_COMP_2.net4_I
timestamp 1698175906
transform 1 0 66192 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_1__f_COMP_4.net2_I
timestamp 1698175906
transform 1 0 48160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_clk_I
timestamp 1698175906
transform 1 0 44240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_clk_I
timestamp 1698175906
transform 1 0 43680 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_clk_I
timestamp 1698175906
transform 1 0 62160 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_clk_I
timestamp 1698175906
transform 1 0 61600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clone1_I
timestamp 1698175906
transform -1 0 66080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_0.x6_B1
timestamp 1698175906
transform 1 0 78848 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_0.x7_C
timestamp 1698175906
transform -1 0 82880 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_0.x8_A1
timestamp 1698175906
transform -1 0 79744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_0.x8_A2
timestamp 1698175906
transform -1 0 80416 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_0.x9_A1
timestamp 1698175906
transform 1 0 79296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_0.x9_A2
timestamp 1698175906
transform 1 0 79296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_0.x9_B1
timestamp 1698175906
transform 1 0 74032 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_0.x15_1_I
timestamp 1698175906
transform 1 0 79408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_1.x6_B1
timestamp 1698175906
transform 1 0 70336 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_1.x8_A1
timestamp 1698175906
transform 1 0 75040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_1.x8_A2
timestamp 1698175906
transform 1 0 74592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_1.x9_A1
timestamp 1698175906
transform 1 0 74480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_1.x9_A2
timestamp 1698175906
transform 1 0 75376 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_1.x9_B1
timestamp 1698175906
transform -1 0 74368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_1.x15_3_I
timestamp 1698175906
transform 1 0 67312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_1.x15_4_I
timestamp 1698175906
transform 1 0 73248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_2.x6_B1
timestamp 1698175906
transform 1 0 62720 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_2.x8_A1
timestamp 1698175906
transform 1 0 61040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_2.x8_A2
timestamp 1698175906
transform 1 0 60592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_2.x9_A1
timestamp 1698175906
transform 1 0 62720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_2.x9_A2
timestamp 1698175906
transform 1 0 59360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_2.x9_B1
timestamp 1698175906
transform 1 0 63168 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_2.x15_5_I
timestamp 1698175906
transform -1 0 57568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_2.x15_6_I
timestamp 1698175906
transform 1 0 57792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_3.x6_B1
timestamp 1698175906
transform 1 0 52640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_3.x8_A1
timestamp 1698175906
transform 1 0 50848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_3.x8_A2
timestamp 1698175906
transform 1 0 51296 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_3.x9_A1
timestamp 1698175906
transform -1 0 52416 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_3.x9_A2
timestamp 1698175906
transform -1 0 51968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_3.x9_B1
timestamp 1698175906
transform -1 0 51520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_3.x15_7_I
timestamp 1698175906
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_3.x15_8_I
timestamp 1698175906
transform 1 0 48832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_4.x6_B1
timestamp 1698175906
transform 1 0 37856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_4.x7_C
timestamp 1698175906
transform -1 0 41216 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_4.x8_A1
timestamp 1698175906
transform 1 0 44912 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_4.x8_A2
timestamp 1698175906
transform 1 0 42560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_4.x9_A1
timestamp 1698175906
transform 1 0 41664 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_4.x9_A2
timestamp 1698175906
transform 1 0 38752 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_4.x9_B1
timestamp 1698175906
transform 1 0 42112 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_4.x15_9_I
timestamp 1698175906
transform 1 0 38304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_4.x15_10_I
timestamp 1698175906
transform 1 0 37408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_5.x6_B1
timestamp 1698175906
transform -1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_5.x7_C
timestamp 1698175906
transform -1 0 29456 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_5.x8_A1
timestamp 1698175906
transform 1 0 35168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_5.x8_A2
timestamp 1698175906
transform 1 0 37968 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_5.x9_A1
timestamp 1698175906
transform 1 0 36512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_5.x9_A2
timestamp 1698175906
transform -1 0 33152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_5.x9_B1
timestamp 1698175906
transform 1 0 36064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_5.x15_11_I
timestamp 1698175906
transform 1 0 34496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_COMP_5.x15_12_I
timestamp 1698175906
transform 1 0 32480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._053__I
timestamp 1698175906
transform 1 0 44912 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._055__A1
timestamp 1698175906
transform 1 0 40096 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._055__A2
timestamp 1698175906
transform -1 0 40432 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._057__I
timestamp 1698175906
transform 1 0 45584 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._062__A1
timestamp 1698175906
transform -1 0 39200 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._062__A2
timestamp 1698175906
transform 1 0 38528 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._063__A1
timestamp 1698175906
transform 1 0 40320 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._063__A2
timestamp 1698175906
transform -1 0 39648 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._064__A1
timestamp 1698175906
transform 1 0 43680 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._064__A2
timestamp 1698175906
transform 1 0 43232 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._065__A1
timestamp 1698175906
transform 1 0 48720 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._065__A2
timestamp 1698175906
transform 1 0 48272 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._066__A1
timestamp 1698175906
transform 1 0 47824 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._068__I
timestamp 1698175906
transform 1 0 61712 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._069__I
timestamp 1698175906
transform 1 0 67648 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._070__I
timestamp 1698175906
transform 1 0 66528 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._071__I
timestamp 1698175906
transform -1 0 55552 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._072__I
timestamp 1698175906
transform 1 0 42336 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._073__I
timestamp 1698175906
transform 1 0 32816 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._074__I
timestamp 1698175906
transform 1 0 29904 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._075__I
timestamp 1698175906
transform 1 0 28448 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._077__A2
timestamp 1698175906
transform 1 0 50736 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._077__A3
timestamp 1698175906
transform 1 0 51184 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._080__A1
timestamp 1698175906
transform 1 0 51632 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._080__B2
timestamp 1698175906
transform 1 0 48160 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._080__C
timestamp 1698175906
transform 1 0 49168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._081__A2
timestamp 1698175906
transform 1 0 55552 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._081__A3
timestamp 1698175906
transform 1 0 56000 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._082__A2
timestamp 1698175906
transform 1 0 52416 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._082__A3
timestamp 1698175906
transform 1 0 52080 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._083__C
timestamp 1698175906
transform -1 0 65856 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._084__A2
timestamp 1698175906
transform -1 0 57792 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._084__A3
timestamp 1698175906
transform 1 0 57120 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._086__A2
timestamp 1698175906
transform 1 0 55104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._086__A3
timestamp 1698175906
transform 1 0 55552 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._087__C
timestamp 1698175906
transform 1 0 64512 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._088__A2
timestamp 1698175906
transform 1 0 45920 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._088__A3
timestamp 1698175906
transform 1 0 45472 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._090__A2
timestamp 1698175906
transform 1 0 53312 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._090__A3
timestamp 1698175906
transform 1 0 53760 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._091__C
timestamp 1698175906
transform 1 0 56000 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._092__A2
timestamp 1698175906
transform 1 0 39872 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._092__A3
timestamp 1698175906
transform 1 0 38416 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._094__A2
timestamp 1698175906
transform 1 0 44240 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._094__A3
timestamp 1698175906
transform 1 0 43792 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._095__C
timestamp 1698175906
transform 1 0 38864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._096__A2
timestamp 1698175906
transform 1 0 36736 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._096__A3
timestamp 1698175906
transform 1 0 36288 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._098__A2
timestamp 1698175906
transform 1 0 36176 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._098__A3
timestamp 1698175906
transform 1 0 35728 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._099__C
timestamp 1698175906
transform 1 0 34160 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._100__A2
timestamp 1698175906
transform 1 0 36960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._100__A3
timestamp 1698175906
transform 1 0 36512 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._102__A2
timestamp 1698175906
transform 1 0 32144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._102__A3
timestamp 1698175906
transform 1 0 31696 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._103__C
timestamp 1698175906
transform 1 0 30800 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._105__A2
timestamp 1698175906
transform 1 0 28784 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._105__A3
timestamp 1698175906
transform 1 0 29232 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._106__A1
timestamp 1698175906
transform 1 0 29232 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._106__A2
timestamp 1698175906
transform 1 0 31248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._108__A2
timestamp 1698175906
transform -1 0 48720 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._109__A2
timestamp 1698175906
transform -1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._110__A2
timestamp 1698175906
transform -1 0 57344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._111__A2
timestamp 1698175906
transform 1 0 57904 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._112__A2
timestamp 1698175906
transform 1 0 41888 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._113__A2
timestamp 1698175906
transform 1 0 35168 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._114__A2
timestamp 1698175906
transform 1 0 31248 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._115__A2
timestamp 1698175906
transform -1 0 28560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._116__CLK
timestamp 1698175906
transform 1 0 50400 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._117__CLK
timestamp 1698175906
transform 1 0 69552 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._118__CLK
timestamp 1698175906
transform 1 0 68768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._119__CLK
timestamp 1698175906
transform 1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._120__CLK
timestamp 1698175906
transform -1 0 39088 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._121__CLK
timestamp 1698175906
transform 1 0 35728 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._122__CLK
timestamp 1698175906
transform 1 0 32480 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._123__CLK
timestamp 1698175906
transform 1 0 29232 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._124__CLK
timestamp 1698175906
transform 1 0 44240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._125__CLK
timestamp 1698175906
transform 1 0 50624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._126__CLK
timestamp 1698175906
transform -1 0 61936 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._127__CLK
timestamp 1698175906
transform 1 0 63840 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._128__CLK
timestamp 1698175906
transform 1 0 43680 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._129__CLK
timestamp 1698175906
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._130__CLK
timestamp 1698175906
transform 1 0 33152 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._131__CLK
timestamp 1698175906
transform 1 0 26320 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._132__CLK
timestamp 1698175906
transform 1 0 39872 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._132__RN
timestamp 1698175906
transform -1 0 40544 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._133__CLK
timestamp 1698175906
transform 1 0 45472 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_CTRL._133__RN
timestamp 1698175906
transform -1 0 46144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout93_I
timestamp 1698175906
transform -1 0 7392 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout94_I
timestamp 1698175906
transform 1 0 5712 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout95_I
timestamp 1698175906
transform 1 0 17472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout96_I
timestamp 1698175906
transform 1 0 7280 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout97_I
timestamp 1698175906
transform 1 0 7168 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout98_I
timestamp 1698175906
transform 1 0 18368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout99_I
timestamp 1698175906
transform 1 0 7056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout100_I
timestamp 1698175906
transform -1 0 4368 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout101_I
timestamp 1698175906
transform 1 0 29680 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout102_I
timestamp 1698175906
transform -1 0 29008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout103_I
timestamp 1698175906
transform 1 0 29568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout104_I
timestamp 1698175906
transform 1 0 42560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout105_I
timestamp 1698175906
transform 1 0 64288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout106_I
timestamp 1698175906
transform 1 0 53424 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout107_I
timestamp 1698175906
transform -1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout108_I
timestamp 1698175906
transform 1 0 66864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout109_I
timestamp 1698175906
transform 1 0 75488 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout110_I
timestamp 1698175906
transform 1 0 76832 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout111_I
timestamp 1698175906
transform 1 0 87136 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout112_I
timestamp 1698175906
transform 1 0 73696 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout113_I
timestamp 1698175906
transform 1 0 6832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout115_I
timestamp 1698175906
transform 1 0 50400 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout116_I
timestamp 1698175906
transform 1 0 84672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698175906
transform -1 0 93968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698175906
transform -1 0 86016 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698175906
transform 1 0 78848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698175906
transform 1 0 63168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698175906
transform -1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698175906
transform -1 0 37184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698175906
transform -1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698175906
transform -1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698175906
transform 1 0 2464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698175906
transform 1 0 2464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698175906
transform 1 0 2464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698175906
transform 1 0 3136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698175906
transform -1 0 2240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698175906
transform 1 0 2464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698175906
transform 1 0 2464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698175906
transform 1 0 1792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698175906
transform 1 0 2464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698175906
transform 1 0 2464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698175906
transform 1 0 1792 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698175906
transform 1 0 2464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698175906
transform -1 0 2240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698175906
transform 1 0 3136 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698175906
transform 1 0 1792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698175906
transform 1 0 2464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698175906
transform 1 0 3248 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698175906
transform 1 0 1792 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698175906
transform 1 0 2912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698175906
transform 1 0 2464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698175906
transform 1 0 2464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698175906
transform 1 0 2464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698175906
transform 1 0 2912 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698175906
transform 1 0 2464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698175906
transform 1 0 2464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698175906
transform 1 0 2464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698175906
transform 1 0 3136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698175906
transform 1 0 2464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698175906
transform 1 0 3584 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698175906
transform 1 0 3136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698175906
transform 1 0 2464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698175906
transform 1 0 2912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698175906
transform 1 0 2464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698175906
transform 1 0 2464 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698175906
transform 1 0 2464 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698175906
transform 1 0 2464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698175906
transform 1 0 3136 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698175906
transform 1 0 2464 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698175906
transform 1 0 1792 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698175906
transform 1 0 2464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698175906
transform 1 0 1792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698175906
transform -1 0 6160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_net299_2_I
timestamp 1698175906
transform 1 0 78960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output52_I
timestamp 1698175906
transform 1 0 96544 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output53_I
timestamp 1698175906
transform 1 0 98112 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output57_I
timestamp 1698175906
transform 1 0 96544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output58_I
timestamp 1698175906
transform -1 0 96768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output59_I
timestamp 1698175906
transform -1 0 96768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output60_I
timestamp 1698175906
transform 1 0 96544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output61_I
timestamp 1698175906
transform 1 0 96544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output63_I
timestamp 1698175906
transform 1 0 96544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output65_I
timestamp 1698175906
transform 1 0 96544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output66_I
timestamp 1698175906
transform -1 0 96768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output67_I
timestamp 1698175906
transform -1 0 96768 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output68_I
timestamp 1698175906
transform -1 0 96768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output70_I
timestamp 1698175906
transform 1 0 96544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output71_I
timestamp 1698175906
transform -1 0 96768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output72_I
timestamp 1698175906
transform -1 0 96768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output73_I
timestamp 1698175906
transform -1 0 96768 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output74_I
timestamp 1698175906
transform 1 0 96544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output76_I
timestamp 1698175906
transform 1 0 96320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output77_I
timestamp 1698175906
transform -1 0 96768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output92_I
timestamp 1698175906
transform -1 0 8848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._287__I
timestamp 1698175906
transform 1 0 43008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._288__A2
timestamp 1698175906
transform 1 0 42672 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._289__A1
timestamp 1698175906
transform 1 0 34496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._289__A2
timestamp 1698175906
transform 1 0 34048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._291__A1
timestamp 1698175906
transform 1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._291__A2
timestamp 1698175906
transform 1 0 41216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._291__A3
timestamp 1698175906
transform 1 0 36176 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._291__A4
timestamp 1698175906
transform 1 0 35280 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._293__I
timestamp 1698175906
transform 1 0 39760 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._294__A1
timestamp 1698175906
transform -1 0 38192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._295__I
timestamp 1698175906
transform -1 0 12096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._296__A2
timestamp 1698175906
transform -1 0 57680 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._298__I
timestamp 1698175906
transform -1 0 74256 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._299__I
timestamp 1698175906
transform 1 0 83440 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._300__A1
timestamp 1698175906
transform -1 0 54656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._301__A1
timestamp 1698175906
transform -1 0 57680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._302__I
timestamp 1698175906
transform 1 0 46816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._303__A1
timestamp 1698175906
transform 1 0 38864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._303__A2
timestamp 1698175906
transform -1 0 39536 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._307__I
timestamp 1698175906
transform -1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._308__I
timestamp 1698175906
transform 1 0 45472 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._311__A1
timestamp 1698175906
transform 1 0 46928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._316__I
timestamp 1698175906
transform 1 0 40992 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._317__A1
timestamp 1698175906
transform 1 0 41440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._317__B
timestamp 1698175906
transform 1 0 38192 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._317__C
timestamp 1698175906
transform 1 0 38640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._318__A1
timestamp 1698175906
transform 1 0 38416 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._318__A2
timestamp 1698175906
transform 1 0 38864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._318__A3
timestamp 1698175906
transform 1 0 42672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._318__A4
timestamp 1698175906
transform 1 0 42896 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._319__A2
timestamp 1698175906
transform 1 0 49728 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._321__I1
timestamp 1698175906
transform 1 0 56336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._321__S
timestamp 1698175906
transform 1 0 55328 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._323__I1
timestamp 1698175906
transform 1 0 76720 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._323__S
timestamp 1698175906
transform -1 0 76720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._325__I1
timestamp 1698175906
transform 1 0 71232 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._325__S
timestamp 1698175906
transform 1 0 71680 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._327__I1
timestamp 1698175906
transform 1 0 72912 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._327__S
timestamp 1698175906
transform 1 0 72464 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._329__I1
timestamp 1698175906
transform -1 0 63168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._329__S
timestamp 1698175906
transform -1 0 63616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._331__I1
timestamp 1698175906
transform 1 0 44464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._331__S
timestamp 1698175906
transform -1 0 46816 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._333__I1
timestamp 1698175906
transform -1 0 64960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._333__S
timestamp 1698175906
transform 1 0 63840 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._335__I1
timestamp 1698175906
transform 1 0 44464 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._335__S
timestamp 1698175906
transform 1 0 46592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._339__I1
timestamp 1698175906
transform 1 0 61040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._339__S
timestamp 1698175906
transform -1 0 61712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._341__I1
timestamp 1698175906
transform 1 0 77616 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._341__S
timestamp 1698175906
transform 1 0 77392 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._343__I1
timestamp 1698175906
transform 1 0 72128 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._343__S
timestamp 1698175906
transform -1 0 71904 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._345__I1
timestamp 1698175906
transform 1 0 76384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._345__S
timestamp 1698175906
transform 1 0 76832 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._347__I1
timestamp 1698175906
transform 1 0 63616 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._347__S
timestamp 1698175906
transform -1 0 64288 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._349__I1
timestamp 1698175906
transform 1 0 44240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._349__S
timestamp 1698175906
transform 1 0 46368 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._351__I1
timestamp 1698175906
transform -1 0 67536 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._351__S
timestamp 1698175906
transform 1 0 67760 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._353__I1
timestamp 1698175906
transform 1 0 44352 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._353__S
timestamp 1698175906
transform 1 0 46480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._357__I1
timestamp 1698175906
transform 1 0 55328 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._357__S
timestamp 1698175906
transform 1 0 53872 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._359__I1
timestamp 1698175906
transform 1 0 75712 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._359__S
timestamp 1698175906
transform 1 0 76160 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._361__I1
timestamp 1698175906
transform 1 0 71232 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._361__S
timestamp 1698175906
transform 1 0 71680 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._363__I1
timestamp 1698175906
transform 1 0 72688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._363__S
timestamp 1698175906
transform 1 0 71680 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._365__I1
timestamp 1698175906
transform 1 0 61264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._365__S
timestamp 1698175906
transform 1 0 60592 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._367__I1
timestamp 1698175906
transform 1 0 38528 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._367__S
timestamp 1698175906
transform 1 0 40992 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._369__I1
timestamp 1698175906
transform 1 0 60144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._369__S
timestamp 1698175906
transform 1 0 59920 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._371__I1
timestamp 1698175906
transform 1 0 40320 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._371__S
timestamp 1698175906
transform 1 0 42672 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._373__A1
timestamp 1698175906
transform 1 0 38416 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._373__A2
timestamp 1698175906
transform 1 0 38864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._373__A3
timestamp 1698175906
transform 1 0 41440 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._373__A4
timestamp 1698175906
transform 1 0 40992 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._375__I0
timestamp 1698175906
transform -1 0 55328 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._375__S
timestamp 1698175906
transform -1 0 53200 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._377__I0
timestamp 1698175906
transform 1 0 58352 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._377__S
timestamp 1698175906
transform -1 0 56448 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._379__I0
timestamp 1698175906
transform 1 0 58464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._379__S
timestamp 1698175906
transform 1 0 55888 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._381__I0
timestamp 1698175906
transform 1 0 55552 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._381__S
timestamp 1698175906
transform 1 0 56000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._383__I0
timestamp 1698175906
transform 1 0 35728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._383__S
timestamp 1698175906
transform 1 0 35280 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._385__I0
timestamp 1698175906
transform 1 0 35952 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._385__S
timestamp 1698175906
transform 1 0 35504 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._387__I0
timestamp 1698175906
transform 1 0 33264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._387__S
timestamp 1698175906
transform 1 0 35840 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._389__I0
timestamp 1698175906
transform 1 0 32928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._389__S
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._391__A1
timestamp 1698175906
transform -1 0 44688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._393__I0
timestamp 1698175906
transform -1 0 61264 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._393__S
timestamp 1698175906
transform 1 0 60816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._395__I0
timestamp 1698175906
transform 1 0 77952 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._395__S
timestamp 1698175906
transform 1 0 76272 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._397__I0
timestamp 1698175906
transform 1 0 69664 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._397__S
timestamp 1698175906
transform 1 0 69440 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._399__I0
timestamp 1698175906
transform -1 0 77280 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._399__S
timestamp 1698175906
transform 1 0 76832 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._401__I0
timestamp 1698175906
transform 1 0 61264 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._401__S
timestamp 1698175906
transform 1 0 61712 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._403__I0
timestamp 1698175906
transform 1 0 40656 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._403__S
timestamp 1698175906
transform 1 0 42672 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._405__I0
timestamp 1698175906
transform 1 0 66080 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._405__S
timestamp 1698175906
transform 1 0 65968 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._407__I0
timestamp 1698175906
transform -1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._407__S
timestamp 1698175906
transform 1 0 42672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._410__I0
timestamp 1698175906
transform -1 0 55776 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._410__S
timestamp 1698175906
transform 1 0 56000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._412__I0
timestamp 1698175906
transform 1 0 53536 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._412__S
timestamp 1698175906
transform 1 0 51408 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._414__I0
timestamp 1698175906
transform 1 0 55552 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._414__S
timestamp 1698175906
transform 1 0 54096 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._416__I0
timestamp 1698175906
transform 1 0 55328 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._416__S
timestamp 1698175906
transform 1 0 53200 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._418__I0
timestamp 1698175906
transform 1 0 31584 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._418__S
timestamp 1698175906
transform 1 0 31136 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._420__I0
timestamp 1698175906
transform 1 0 31024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._420__S
timestamp 1698175906
transform 1 0 31248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._422__I0
timestamp 1698175906
transform 1 0 31360 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._422__S
timestamp 1698175906
transform 1 0 30912 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._424__I0
timestamp 1698175906
transform 1 0 28784 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._424__S
timestamp 1698175906
transform 1 0 30016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._426__A2
timestamp 1698175906
transform 1 0 91280 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._427__I
timestamp 1698175906
transform 1 0 45472 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._428__A1
timestamp 1698175906
transform 1 0 45024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._428__A2
timestamp 1698175906
transform 1 0 45920 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._429__A2
timestamp 1698175906
transform 1 0 45248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._431__I
timestamp 1698175906
transform 1 0 46368 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._432__A2
timestamp 1698175906
transform 1 0 46368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._432__A3
timestamp 1698175906
transform 1 0 45920 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._433__I
timestamp 1698175906
transform 1 0 51184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._434__A1
timestamp 1698175906
transform 1 0 45920 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._434__A2
timestamp 1698175906
transform -1 0 51744 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._434__A3
timestamp 1698175906
transform 1 0 44912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._435__A2
timestamp 1698175906
transform -1 0 59920 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._435__B1
timestamp 1698175906
transform -1 0 60368 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._435__C2
timestamp 1698175906
transform -1 0 60816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._436__A1
timestamp 1698175906
transform 1 0 50400 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._436__A2
timestamp 1698175906
transform -1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._436__A3
timestamp 1698175906
transform -1 0 47936 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._437__A1
timestamp 1698175906
transform 1 0 52080 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._438__I
timestamp 1698175906
transform -1 0 49056 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._440__A1
timestamp 1698175906
transform 1 0 52416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._440__A2
timestamp 1698175906
transform 1 0 51968 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._440__A4
timestamp 1698175906
transform 1 0 51520 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._441__A1
timestamp 1698175906
transform 1 0 56000 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._441__A2
timestamp 1698175906
transform 1 0 56784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._441__A4
timestamp 1698175906
transform 1 0 56672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._442__A1
timestamp 1698175906
transform 1 0 38640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._444__I
timestamp 1698175906
transform 1 0 73808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._445__B
timestamp 1698175906
transform 1 0 65408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._446__A2
timestamp 1698175906
transform -1 0 89152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._448__A1
timestamp 1698175906
transform 1 0 75376 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._448__A2
timestamp 1698175906
transform 1 0 75376 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._448__A4
timestamp 1698175906
transform 1 0 74928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._449__A2
timestamp 1698175906
transform -1 0 77168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._450__A1
timestamp 1698175906
transform 1 0 50960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._451__A1
timestamp 1698175906
transform 1 0 55552 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._451__A2
timestamp 1698175906
transform 1 0 54208 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._451__B1
timestamp 1698175906
transform 1 0 56000 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._451__C2
timestamp 1698175906
transform -1 0 55328 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._452__A1
timestamp 1698175906
transform 1 0 50848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._452__A2
timestamp 1698175906
transform 1 0 48944 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._452__A3
timestamp 1698175906
transform 1 0 49392 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._453__A2
timestamp 1698175906
transform 1 0 75936 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._453__B1
timestamp 1698175906
transform 1 0 76384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._454__A3
timestamp 1698175906
transform -1 0 76720 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._455__S
timestamp 1698175906
transform -1 0 84784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._457__A1
timestamp 1698175906
transform -1 0 73696 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._457__A2
timestamp 1698175906
transform -1 0 73696 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._457__A4
timestamp 1698175906
transform 1 0 73024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._458__A2
timestamp 1698175906
transform -1 0 72800 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._459__A1
timestamp 1698175906
transform -1 0 54208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._459__A2
timestamp 1698175906
transform 1 0 54656 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._459__B1
timestamp 1698175906
transform 1 0 54432 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._459__C2
timestamp 1698175906
transform 1 0 54432 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._460__A2
timestamp 1698175906
transform -1 0 74032 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._460__B1
timestamp 1698175906
transform -1 0 73584 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._461__A3
timestamp 1698175906
transform 1 0 73360 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._462__I0
timestamp 1698175906
transform 1 0 91616 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._462__S
timestamp 1698175906
transform 1 0 91168 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._464__A1
timestamp 1698175906
transform 1 0 74928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._464__A2
timestamp 1698175906
transform 1 0 76384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._464__A4
timestamp 1698175906
transform 1 0 75376 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._465__A2
timestamp 1698175906
transform 1 0 77840 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._466__A1
timestamp 1698175906
transform 1 0 53312 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._466__A2
timestamp 1698175906
transform 1 0 54656 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._466__B1
timestamp 1698175906
transform 1 0 53760 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._466__C2
timestamp 1698175906
transform 1 0 54208 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._467__A2
timestamp 1698175906
transform 1 0 75936 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._467__B1
timestamp 1698175906
transform 1 0 75600 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._468__A3
timestamp 1698175906
transform -1 0 76384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._469__S
timestamp 1698175906
transform 1 0 87584 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._471__A1
timestamp 1698175906
transform 1 0 65408 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._471__A2
timestamp 1698175906
transform 1 0 64512 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._471__A4
timestamp 1698175906
transform 1 0 64960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._472__A2
timestamp 1698175906
transform -1 0 65408 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._473__A1
timestamp 1698175906
transform 1 0 33264 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._473__B1
timestamp 1698175906
transform 1 0 38976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._473__C2
timestamp 1698175906
transform 1 0 39424 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._474__A2
timestamp 1698175906
transform 1 0 63840 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._474__B1
timestamp 1698175906
transform 1 0 64512 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._475__A3
timestamp 1698175906
transform -1 0 65072 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._476__I0
timestamp 1698175906
transform 1 0 85456 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._476__S
timestamp 1698175906
transform 1 0 85008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._478__A1
timestamp 1698175906
transform -1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._478__A2
timestamp 1698175906
transform -1 0 51744 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._478__A4
timestamp 1698175906
transform 1 0 47712 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._479__A2
timestamp 1698175906
transform 1 0 48048 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._480__A1
timestamp 1698175906
transform 1 0 32480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._480__B1
timestamp 1698175906
transform 1 0 39200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._480__C2
timestamp 1698175906
transform 1 0 39648 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._481__A2
timestamp 1698175906
transform 1 0 49168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._481__B1
timestamp 1698175906
transform 1 0 48720 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._483__I0
timestamp 1698175906
transform -1 0 91280 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._483__S
timestamp 1698175906
transform 1 0 90608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._485__A1
timestamp 1698175906
transform 1 0 67200 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._485__A2
timestamp 1698175906
transform 1 0 67648 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._485__A4
timestamp 1698175906
transform 1 0 66640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._486__A2
timestamp 1698175906
transform 1 0 68992 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._487__A1
timestamp 1698175906
transform 1 0 33712 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._487__B1
timestamp 1698175906
transform 1 0 39424 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._487__C2
timestamp 1698175906
transform 1 0 39872 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._488__A2
timestamp 1698175906
transform 1 0 68208 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._488__B1
timestamp 1698175906
transform 1 0 67760 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._489__A3
timestamp 1698175906
transform -1 0 68656 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._490__I0
timestamp 1698175906
transform -1 0 91504 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._490__S
timestamp 1698175906
transform 1 0 90832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._492__A1
timestamp 1698175906
transform 1 0 52864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._492__A2
timestamp 1698175906
transform 1 0 52416 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._492__A4
timestamp 1698175906
transform -1 0 47824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._493__A2
timestamp 1698175906
transform 1 0 48384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._494__A1
timestamp 1698175906
transform 1 0 33376 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._494__B1
timestamp 1698175906
transform 1 0 39088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._494__C2
timestamp 1698175906
transform 1 0 38864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._495__A2
timestamp 1698175906
transform 1 0 48832 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._495__B1
timestamp 1698175906
transform 1 0 50288 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._497__I0
timestamp 1698175906
transform 1 0 90160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._497__S
timestamp 1698175906
transform 1 0 89712 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._499__A1
timestamp 1698175906
transform 1 0 35840 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._500__I
timestamp 1698175906
transform 1 0 73136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._501__A2
timestamp 1698175906
transform 1 0 83664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._502__A1
timestamp 1698175906
transform 1 0 83440 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._502__A2
timestamp 1698175906
transform 1 0 82096 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._503__A1
timestamp 1698175906
transform 1 0 37632 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._504__A2
timestamp 1698175906
transform 1 0 85680 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._505__A1
timestamp 1698175906
transform -1 0 84672 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._505__A2
timestamp 1698175906
transform -1 0 84448 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._507__A2
timestamp 1698175906
transform 1 0 85904 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._508__A1
timestamp 1698175906
transform 1 0 85232 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._508__A2
timestamp 1698175906
transform 1 0 83440 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._509__A1
timestamp 1698175906
transform 1 0 37632 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._510__A2
timestamp 1698175906
transform 1 0 80752 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._511__A1
timestamp 1698175906
transform 1 0 78960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._511__A2
timestamp 1698175906
transform -1 0 78064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._512__A1
timestamp 1698175906
transform 1 0 37296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._513__A2
timestamp 1698175906
transform 1 0 85344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._514__A1
timestamp 1698175906
transform 1 0 86016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._514__A2
timestamp 1698175906
transform 1 0 84224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._516__I
timestamp 1698175906
transform 1 0 74704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._517__A2
timestamp 1698175906
transform 1 0 75040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._518__A1
timestamp 1698175906
transform 1 0 73696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._518__A2
timestamp 1698175906
transform -1 0 72576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._520__A2
timestamp 1698175906
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._521__A1
timestamp 1698175906
transform 1 0 70672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._521__A2
timestamp 1698175906
transform -1 0 69552 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._522__A1
timestamp 1698175906
transform 1 0 35840 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._523__A2
timestamp 1698175906
transform 1 0 67200 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._524__A1
timestamp 1698175906
transform 1 0 66528 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._524__A2
timestamp 1698175906
transform -1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._526__A2
timestamp 1698175906
transform 1 0 71232 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._527__A1
timestamp 1698175906
transform -1 0 69776 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._527__A2
timestamp 1698175906
transform -1 0 68432 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._528__I
timestamp 1698175906
transform 1 0 75824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._529__I
timestamp 1698175906
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._530__A1
timestamp 1698175906
transform 1 0 60704 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._531__A2
timestamp 1698175906
transform 1 0 66192 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._532__A1
timestamp 1698175906
transform 1 0 64400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._533__A1
timestamp 1698175906
transform 1 0 62272 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._534__A2
timestamp 1698175906
transform 1 0 78064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._535__A1
timestamp 1698175906
transform 1 0 77056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._536__A1
timestamp 1698175906
transform 1 0 59920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._537__A2
timestamp 1698175906
transform -1 0 75152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._538__A1
timestamp 1698175906
transform 1 0 73472 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._539__A1
timestamp 1698175906
transform 1 0 62272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._540__A2
timestamp 1698175906
transform 1 0 65744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._541__A1
timestamp 1698175906
transform 1 0 63280 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._542__A1
timestamp 1698175906
transform -1 0 60928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._543__A2
timestamp 1698175906
transform 1 0 69328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._544__A1
timestamp 1698175906
transform 1 0 68096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._545__A1
timestamp 1698175906
transform 1 0 59584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._546__A2
timestamp 1698175906
transform -1 0 77840 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._547__A1
timestamp 1698175906
transform 1 0 76944 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._547__A2
timestamp 1698175906
transform 1 0 76720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._548__A1
timestamp 1698175906
transform 1 0 60144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._549__A2
timestamp 1698175906
transform 1 0 65072 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._550__A1
timestamp 1698175906
transform 1 0 63280 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._551__A1
timestamp 1698175906
transform -1 0 60368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._552__A2
timestamp 1698175906
transform 1 0 80976 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._553__A1
timestamp 1698175906
transform 1 0 77392 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._554__A1
timestamp 1698175906
transform 1 0 59360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._555__A2
timestamp 1698175906
transform 1 0 70336 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._556__A1
timestamp 1698175906
transform 1 0 69888 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._557__A1
timestamp 1698175906
transform -1 0 60928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._558__A2
timestamp 1698175906
transform 1 0 75712 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._559__A1
timestamp 1698175906
transform 1 0 74480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._560__A1
timestamp 1698175906
transform 1 0 45136 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._560__A2
timestamp 1698175906
transform 1 0 45584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._561__A2
timestamp 1698175906
transform 1 0 84336 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._562__A1
timestamp 1698175906
transform 1 0 80976 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._562__A2
timestamp 1698175906
transform 1 0 81424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._563__A2
timestamp 1698175906
transform 1 0 43344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._564__A2
timestamp 1698175906
transform -1 0 85344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._565__A1
timestamp 1698175906
transform -1 0 84784 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._565__A2
timestamp 1698175906
transform 1 0 84336 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._566__A2
timestamp 1698175906
transform 1 0 43456 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._567__A2
timestamp 1698175906
transform -1 0 78848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._568__A1
timestamp 1698175906
transform -1 0 77504 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._568__A2
timestamp 1698175906
transform 1 0 76272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._569__A1
timestamp 1698175906
transform 1 0 55440 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._569__A2
timestamp 1698175906
transform 1 0 56672 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._570__A2
timestamp 1698175906
transform -1 0 73136 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._571__A1
timestamp 1698175906
transform 1 0 73024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._572__A2
timestamp 1698175906
transform -1 0 39984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._573__A2
timestamp 1698175906
transform -1 0 82992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._574__A1
timestamp 1698175906
transform 1 0 80640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._574__A2
timestamp 1698175906
transform 1 0 80416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._575__RN
timestamp 1698175906
transform 1 0 52864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._576__RN
timestamp 1698175906
transform 1 0 54208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._577__RN
timestamp 1698175906
transform 1 0 39872 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._578__RN
timestamp 1698175906
transform -1 0 38640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._579__RN
timestamp 1698175906
transform -1 0 54768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._580__RN
timestamp 1698175906
transform 1 0 80528 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._581__RN
timestamp 1698175906
transform 1 0 69328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._582__RN
timestamp 1698175906
transform 1 0 76160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._583__RN
timestamp 1698175906
transform 1 0 61824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._584__RN
timestamp 1698175906
transform 1 0 43232 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._585__RN
timestamp 1698175906
transform 1 0 67088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._586__RN
timestamp 1698175906
transform -1 0 43456 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._587__RN
timestamp 1698175906
transform 1 0 66976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._588__RN
timestamp 1698175906
transform 1 0 79744 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._589__RN
timestamp 1698175906
transform 1 0 74928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._590__RN
timestamp 1698175906
transform 1 0 77616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._591__RN
timestamp 1698175906
transform 1 0 69216 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._592__RN
timestamp 1698175906
transform 1 0 43008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._593__RN
timestamp 1698175906
transform -1 0 67984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._594__RN
timestamp 1698175906
transform 1 0 44464 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._595__RN
timestamp 1698175906
transform 1 0 56672 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._596__RN
timestamp 1698175906
transform -1 0 76720 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._597__RN
timestamp 1698175906
transform 1 0 74256 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._598__RN
timestamp 1698175906
transform 1 0 75040 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._599__RN
timestamp 1698175906
transform -1 0 64624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._600__RN
timestamp 1698175906
transform 1 0 40992 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._601__RN
timestamp 1698175906
transform -1 0 58016 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._602__RN
timestamp 1698175906
transform 1 0 42336 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._603__RN
timestamp 1698175906
transform 1 0 53200 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._604__RN
timestamp 1698175906
transform 1 0 54432 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._605__RN
timestamp 1698175906
transform 1 0 56000 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._606__RN
timestamp 1698175906
transform 1 0 57792 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._607__RN
timestamp 1698175906
transform 1 0 30576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._608__RN
timestamp 1698175906
transform 1 0 31136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._609__RN
timestamp 1698175906
transform 1 0 30912 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._610__RN
timestamp 1698175906
transform 1 0 31136 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._611__RN
timestamp 1698175906
transform 1 0 64400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._612__RN
timestamp 1698175906
transform -1 0 79184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._613__RN
timestamp 1698175906
transform 1 0 67760 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._614__RN
timestamp 1698175906
transform 1 0 78512 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._615__RN
timestamp 1698175906
transform 1 0 64512 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._616__RN
timestamp 1698175906
transform 1 0 41776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._617__RN
timestamp 1698175906
transform 1 0 67760 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._618__RN
timestamp 1698175906
transform 1 0 42112 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._619__RN
timestamp 1698175906
transform 1 0 54992 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._620__RN
timestamp 1698175906
transform 1 0 53200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._621__RN
timestamp 1698175906
transform 1 0 53872 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._622__RN
timestamp 1698175906
transform 1 0 53648 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._623__RN
timestamp 1698175906
transform 1 0 29232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._624__RN
timestamp 1698175906
transform 1 0 29344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._625__RN
timestamp 1698175906
transform 1 0 29232 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._626__RN
timestamp 1698175906
transform 1 0 29792 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._627__RN
timestamp 1698175906
transform 1 0 56000 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._628__RN
timestamp 1698175906
transform 1 0 58016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._629__RN
timestamp 1698175906
transform 1 0 34832 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._630__D
timestamp 1698175906
transform -1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._630__RN
timestamp 1698175906
transform 1 0 8512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._631__D
timestamp 1698175906
transform -1 0 32256 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._631__RN
timestamp 1698175906
transform 1 0 32480 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._632__D
timestamp 1698175906
transform -1 0 25872 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._632__RN
timestamp 1698175906
transform 1 0 30128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._633__D
timestamp 1698175906
transform -1 0 27104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._633__RN
timestamp 1698175906
transform 1 0 31360 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._634__RN
timestamp 1698175906
transform 1 0 9520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._635__RN
timestamp 1698175906
transform 1 0 6048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._636__RN
timestamp 1698175906
transform -1 0 6608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._637__RN
timestamp 1698175906
transform -1 0 6160 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._638__RN
timestamp 1698175906
transform 1 0 11312 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._639__RN
timestamp 1698175906
transform 1 0 5600 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._640__D
timestamp 1698175906
transform -1 0 16240 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._640__RN
timestamp 1698175906
transform -1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._641__RN
timestamp 1698175906
transform 1 0 10080 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._646__RN
timestamp 1698175906
transform 1 0 9184 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._647__RN
timestamp 1698175906
transform 1 0 6608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._648__RN
timestamp 1698175906
transform 1 0 5712 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._649__RN
timestamp 1698175906
transform 1 0 5936 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._650__RN
timestamp 1698175906
transform 1 0 9296 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._651__RN
timestamp 1698175906
transform -1 0 6720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._652__RN
timestamp 1698175906
transform 1 0 5600 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._658__D
timestamp 1698175906
transform 1 0 20384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._658__RN
timestamp 1698175906
transform 1 0 19936 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._660__D
timestamp 1698175906
transform 1 0 17696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._660__RN
timestamp 1698175906
transform 1 0 22400 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._663__RN
timestamp 1698175906
transform 1 0 9520 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._664__RN
timestamp 1698175906
transform 1 0 5600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._665__RN
timestamp 1698175906
transform 1 0 19600 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._666__D
timestamp 1698175906
transform 1 0 26320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._666__RN
timestamp 1698175906
transform 1 0 30576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._667__D
timestamp 1698175906
transform 1 0 26992 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._667__RN
timestamp 1698175906
transform -1 0 28560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._668__RN
timestamp 1698175906
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._669__D
timestamp 1698175906
transform 1 0 18480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._669__RN
timestamp 1698175906
transform -1 0 18256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._670__D
timestamp 1698175906
transform 1 0 43792 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._670__RN
timestamp 1698175906
transform 1 0 44240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._671__RN
timestamp 1698175906
transform 1 0 53648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._672__RN
timestamp 1698175906
transform -1 0 90048 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._673__RN
timestamp 1698175906
transform 1 0 90496 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._674__RN
timestamp 1698175906
transform -1 0 92512 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._675__RN
timestamp 1698175906
transform 1 0 90384 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._676__RN
timestamp 1698175906
transform 1 0 89936 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._677__RN
timestamp 1698175906
transform 1 0 91280 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._678__RN
timestamp 1698175906
transform 1 0 90944 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._679__RN
timestamp 1698175906
transform 1 0 90720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._680__RN
timestamp 1698175906
transform 1 0 86240 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._681__RN
timestamp 1698175906
transform 1 0 90608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._682__RN
timestamp 1698175906
transform 1 0 88032 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._683__RN
timestamp 1698175906
transform 1 0 77616 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._684__RN
timestamp 1698175906
transform -1 0 84448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._685__RN
timestamp 1698175906
transform -1 0 76496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._686__RN
timestamp 1698175906
transform 1 0 68544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._687__RN
timestamp 1698175906
transform 1 0 68880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._688__RN
timestamp 1698175906
transform 1 0 67312 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._689__RN
timestamp 1698175906
transform 1 0 62272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._690__RN
timestamp 1698175906
transform 1 0 75712 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._691__RN
timestamp 1698175906
transform 1 0 76272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._692__RN
timestamp 1698175906
transform 1 0 65520 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._693__RN
timestamp 1698175906
transform 1 0 66304 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._694__RN
timestamp 1698175906
transform 1 0 77952 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._695__RN
timestamp 1698175906
transform 1 0 65520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._696__RN
timestamp 1698175906
transform 1 0 77728 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._697__RN
timestamp 1698175906
transform 1 0 65968 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._698__RN
timestamp 1698175906
transform 1 0 76272 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._699__RN
timestamp 1698175906
transform 1 0 82544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._700__RN
timestamp 1698175906
transform 1 0 85120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._701__RN
timestamp 1698175906
transform 1 0 75600 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._702__RN
timestamp 1698175906
transform 1 0 74704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg._703__RN
timestamp 1698175906
transform -1 0 79744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._069__I1
timestamp 1698175906
transform 1 0 21840 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._069__S
timestamp 1698175906
transform 1 0 18928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._071__I1
timestamp 1698175906
transform 1 0 11760 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._071__S
timestamp 1698175906
transform 1 0 11312 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._073__I1
timestamp 1698175906
transform -1 0 22176 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._073__S
timestamp 1698175906
transform 1 0 19824 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._075__I1
timestamp 1698175906
transform 1 0 11536 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._075__S
timestamp 1698175906
transform 1 0 11088 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._077__I1
timestamp 1698175906
transform -1 0 16576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._077__S
timestamp 1698175906
transform 1 0 13552 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._079__I1
timestamp 1698175906
transform -1 0 17696 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._079__S
timestamp 1698175906
transform 1 0 14896 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._081__I1
timestamp 1698175906
transform 1 0 23072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._081__S
timestamp 1698175906
transform 1 0 20720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._083__I1
timestamp 1698175906
transform 1 0 15232 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._083__S
timestamp 1698175906
transform 1 0 12208 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._086__I1
timestamp 1698175906
transform -1 0 13664 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._086__S
timestamp 1698175906
transform 1 0 11200 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._088__I1
timestamp 1698175906
transform -1 0 19152 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._088__S
timestamp 1698175906
transform 1 0 16800 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._090__I0
timestamp 1698175906
transform -1 0 20272 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._090__S
timestamp 1698175906
transform 1 0 19600 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._092__I1
timestamp 1698175906
transform -1 0 11984 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._092__S
timestamp 1698175906
transform 1 0 11312 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._094__I1
timestamp 1698175906
transform 1 0 17472 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._094__S
timestamp 1698175906
transform 1 0 14896 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._096__S
timestamp 1698175906
transform 1 0 19712 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._098__S
timestamp 1698175906
transform 1 0 19040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._100__I1
timestamp 1698175906
transform 1 0 16688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._100__S
timestamp 1698175906
transform 1 0 14560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._103__I0
timestamp 1698175906
transform 1 0 26656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._103__S
timestamp 1698175906
transform 1 0 26208 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._105__I1
timestamp 1698175906
transform 1 0 16800 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._105__S
timestamp 1698175906
transform 1 0 14672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._107__I0
timestamp 1698175906
transform -1 0 30688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._107__I1
timestamp 1698175906
transform 1 0 33152 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._107__S
timestamp 1698175906
transform 1 0 30240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._109__I0
timestamp 1698175906
transform 1 0 29904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._109__I1
timestamp 1698175906
transform 1 0 32032 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._109__S
timestamp 1698175906
transform 1 0 29456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._111__I1
timestamp 1698175906
transform 1 0 26768 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._111__S
timestamp 1698175906
transform 1 0 24192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._113__I1
timestamp 1698175906
transform -1 0 13888 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._113__S
timestamp 1698175906
transform 1 0 11760 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._115__I1
timestamp 1698175906
transform 1 0 23072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._115__S
timestamp 1698175906
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._117__I0
timestamp 1698175906
transform 1 0 25648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._117__I1
timestamp 1698175906
transform 1 0 28224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._117__S
timestamp 1698175906
transform 1 0 25200 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._120__I0
timestamp 1698175906
transform -1 0 38192 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._120__I1
timestamp 1698175906
transform -1 0 40320 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._120__S
timestamp 1698175906
transform 1 0 37520 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._122__I0
timestamp 1698175906
transform 1 0 32592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._122__I1
timestamp 1698175906
transform 1 0 34720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._122__S
timestamp 1698175906
transform 1 0 32144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._124__I1
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._124__S
timestamp 1698175906
transform -1 0 12432 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._126__I1
timestamp 1698175906
transform 1 0 23072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._126__S
timestamp 1698175906
transform 1 0 20272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._128__S
timestamp 1698175906
transform 1 0 38080 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._130__S
timestamp 1698175906
transform 1 0 32592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._132__I1
timestamp 1698175906
transform -1 0 16912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._132__S
timestamp 1698175906
transform 1 0 14560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._134__S
timestamp 1698175906
transform 1 0 22960 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._136__RN
timestamp 1698175906
transform 1 0 19712 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._138__RN
timestamp 1698175906
transform 1 0 20944 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._140__RN
timestamp 1698175906
transform 1 0 18144 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._141__RN
timestamp 1698175906
transform 1 0 14000 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._142__RN
timestamp 1698175906
transform 1 0 19600 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._143__RN
timestamp 1698175906
transform 1 0 17472 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._144__RN
timestamp 1698175906
transform 1 0 17472 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._145__RN
timestamp 1698175906
transform 1 0 22960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._146__RN
timestamp 1698175906
transform 1 0 21056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._147__RN
timestamp 1698175906
transform 1 0 8400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._148__RN
timestamp 1698175906
transform 1 0 18592 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._149__RN
timestamp 1698175906
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._150__RN
timestamp 1698175906
transform 1 0 20272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._151__RN
timestamp 1698175906
transform 1 0 18368 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._152__RN
timestamp 1698175906
transform 1 0 30016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._153__RN
timestamp 1698175906
transform 1 0 12992 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._154__RN
timestamp 1698175906
transform 1 0 32704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._155__RN
timestamp 1698175906
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._156__RN
timestamp 1698175906
transform 1 0 29232 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._157__RN
timestamp 1698175906
transform 1 0 17696 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._158__RN
timestamp 1698175906
transform 1 0 19152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._159__RN
timestamp 1698175906
transform 1 0 30464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._160__RN
timestamp 1698175906
transform 1 0 38416 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._161__RN
timestamp 1698175906
transform 1 0 32032 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._162__RN
timestamp 1698175906
transform 1 0 12432 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._163__RN
timestamp 1698175906
transform 1 0 20272 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._164__RN
timestamp 1698175906
transform 1 0 38976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._165__RN
timestamp 1698175906
transform 1 0 33040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._166__RN
timestamp 1698175906
transform 1 0 18704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_u_adc_reg.u_reg_0._167__RN
timestamp 1698175906
transform -1 0 29456 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_wire26_I
timestamp 1698175906
transform 1 0 20720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_wire114_I
timestamp 1698175906
transform 1 0 26544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_20  clkbuf_0_clk open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 52528 0 1 29792
box -86 -86 7030 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_0.net1 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 87808 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_0.net2
timestamp 1698175906
transform 1 0 83888 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_0.net3
timestamp 1698175906
transform 1 0 83888 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_0.net4
timestamp 1698175906
transform 1 0 79968 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_0.Q
timestamp 1698175906
transform -1 0 77728 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_1.net1
timestamp 1698175906
transform 1 0 76048 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_1.net2
timestamp 1698175906
transform 1 0 79968 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_1.net3
timestamp 1698175906
transform 1 0 79968 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_1.net4
timestamp 1698175906
transform 1 0 72128 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_1.Q
timestamp 1698175906
transform -1 0 73808 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_2.net1
timestamp 1698175906
transform 1 0 64288 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_2.net2
timestamp 1698175906
transform 1 0 60368 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_2.net3
timestamp 1698175906
transform 1 0 58464 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_2.net4
timestamp 1698175906
transform 1 0 68208 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_2.Q
timestamp 1698175906
transform -1 0 62048 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_3.net1
timestamp 1698175906
transform 1 0 50624 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_3.net2
timestamp 1698175906
transform 1 0 46704 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_3.net3
timestamp 1698175906
transform 1 0 50400 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_3.net4
timestamp 1698175906
transform 1 0 46704 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_3.Q
timestamp 1698175906
transform 1 0 50624 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_4.net1
timestamp 1698175906
transform -1 0 40544 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_4.net2
timestamp 1698175906
transform 1 0 42224 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_4.net3
timestamp 1698175906
transform -1 0 44464 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_4.net4
timestamp 1698175906
transform -1 0 40544 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_4.Q
timestamp 1698175906
transform -1 0 44464 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_5.net1
timestamp 1698175906
transform 1 0 27104 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_5.net2
timestamp 1698175906
transform 1 0 34496 0 -1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_5.net3
timestamp 1698175906
transform -1 0 36624 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_5.net4
timestamp 1698175906
transform -1 0 32704 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_COMP_5.Q
timestamp 1698175906
transform 1 0 38864 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_CTRL.cmp
timestamp 1698175906
transform -1 0 47712 0 -1 53312
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_0.net1
timestamp 1698175906
transform -1 0 82880 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_0.net2
timestamp 1698175906
transform -1 0 81648 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_16  clkbuf_1_0__f_COMP_0.net3 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 82096 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_16  clkbuf_1_0__f_COMP_0.net4
timestamp 1698175906
transform 1 0 87808 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_16  clkbuf_1_0__f_COMP_0.Q
timestamp 1698175906
transform -1 0 69888 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_1.net1
timestamp 1698175906
transform -1 0 73808 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_1.net2
timestamp 1698175906
transform -1 0 74032 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_1.net3
timestamp 1698175906
transform -1 0 77728 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_1.net4
timestamp 1698175906
transform -1 0 77728 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_1.Q
timestamp 1698175906
transform -1 0 65968 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_2.net1
timestamp 1698175906
transform -1 0 69888 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_2.net2
timestamp 1698175906
transform -1 0 64064 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_2.net3
timestamp 1698175906
transform -1 0 63280 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_2.net4
timestamp 1698175906
transform -1 0 66304 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_2.Q
timestamp 1698175906
transform -1 0 58128 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_3.net1
timestamp 1698175906
transform -1 0 48384 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_3.net2
timestamp 1698175906
transform 1 0 52528 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_3.net3
timestamp 1698175906
transform -1 0 48384 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_3.net4
timestamp 1698175906
transform -1 0 54208 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_3.Q
timestamp 1698175906
transform -1 0 52304 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_4.net1
timestamp 1698175906
transform 1 0 42112 0 -1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_4.net2
timestamp 1698175906
transform -1 0 32704 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_4.net3
timestamp 1698175906
transform -1 0 36624 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_4.net4
timestamp 1698175906
transform -1 0 36624 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_4.Q
timestamp 1698175906
transform -1 0 40544 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_5.net1
timestamp 1698175906
transform 1 0 31024 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_5.net2
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_5.net3
timestamp 1698175906
transform -1 0 28784 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_5.net4
timestamp 1698175906
transform -1 0 32704 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_COMP_5.Q
timestamp 1698175906
transform -1 0 40544 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_16  clkbuf_1_0__f_CTRL.cmp
timestamp 1698175906
transform -1 0 44016 0 1 51744
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_0.net1
timestamp 1698175906
transform -1 0 89488 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_0.net2
timestamp 1698175906
transform 1 0 87808 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_0.net3
timestamp 1698175906
transform -1 0 85568 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_0.net4
timestamp 1698175906
transform -1 0 89488 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_0.Q
timestamp 1698175906
transform 1 0 76048 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_1.net1
timestamp 1698175906
transform -1 0 77728 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_1.net2
timestamp 1698175906
transform -1 0 81648 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_1.net3
timestamp 1698175906
transform -1 0 85568 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_1.net4
timestamp 1698175906
transform -1 0 75264 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_1.Q
timestamp 1698175906
transform 1 0 68208 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_2.net1
timestamp 1698175906
transform -1 0 69888 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_2.net2
timestamp 1698175906
transform -1 0 65968 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_2.net3
timestamp 1698175906
transform 1 0 72128 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_2.net4
timestamp 1698175906
transform 1 0 60368 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_2.Q
timestamp 1698175906
transform 1 0 64288 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_3.net1
timestamp 1698175906
transform 1 0 52528 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_3.net2
timestamp 1698175906
transform 1 0 50624 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_3.net3
timestamp 1698175906
transform 1 0 52752 0 1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_3.net4
timestamp 1698175906
transform 1 0 56448 0 -1 6272
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_3.Q
timestamp 1698175906
transform 1 0 56448 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_4.net1
timestamp 1698175906
transform 1 0 42784 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_4.net2
timestamp 1698175906
transform -1 0 48384 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_4.net3
timestamp 1698175906
transform 1 0 42784 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_4.net4
timestamp 1698175906
transform 1 0 44912 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_4.Q
timestamp 1698175906
transform 1 0 46480 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_5.net1
timestamp 1698175906
transform 1 0 38864 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_5.net2
timestamp 1698175906
transform -1 0 36624 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_5.net3
timestamp 1698175906
transform 1 0 34944 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_5.net4
timestamp 1698175906
transform 1 0 34944 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_COMP_5.Q
timestamp 1698175906
transform 1 0 38864 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_16  clkbuf_1_1__f_CTRL.cmp
timestamp 1698175906
transform 1 0 45920 0 1 53312
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1698175906
transform 1 0 38416 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1698175906
transform -1 0 43456 0 1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_16  clkbuf_2_2__f_clk
timestamp 1698175906
transform 1 0 62384 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1698175906
transform 1 0 61824 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  clone1 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 66304 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_8  COMP_0.x2_21 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 77728 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_0.x3_15 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 81648 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  COMP_0.x6 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 79968 0 -1 12544
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  COMP_0.x6_118 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 78288 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  COMP_0.x7 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 78176 0 1 14112
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  COMP_0.x7_291 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 79744 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  COMP_0.x8
timestamp 1698175906
transform 1 0 79968 0 -1 14112
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  COMP_0.x8_292
timestamp 1698175906
transform 1 0 77728 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  COMP_0.x9
timestamp 1698175906
transform -1 0 79072 0 -1 14112
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  COMP_0.x9_119
timestamp 1698175906
transform 1 0 77840 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  COMP_0.x10 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 84448 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  COMP_0.x11
timestamp 1698175906
transform -1 0 77504 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  COMP_0.x15_1 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 77728 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_1.x2_16
timestamp 1698175906
transform -1 0 74256 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_1.x3_13
timestamp 1698175906
transform 1 0 70112 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  COMP_1.x6_120
timestamp 1698175906
transform -1 0 75152 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  COMP_1.x6 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 71904 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  COMP_1.x7
timestamp 1698175906
transform 1 0 67424 0 -1 12544
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  COMP_1.x7_293
timestamp 1698175906
transform -1 0 75152 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  COMP_1.x8
timestamp 1698175906
transform 1 0 69888 0 1 14112
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  COMP_1.x8_294
timestamp 1698175906
transform 1 0 67536 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  COMP_1.x9_121
timestamp 1698175906
transform -1 0 75600 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  COMP_1.x9
timestamp 1698175906
transform -1 0 71904 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  COMP_1.x10
timestamp 1698175906
transform -1 0 73024 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  COMP_1.x11 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 70784 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  COMP_1.x15_3
timestamp 1698175906
transform 1 0 69888 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_1.x15_4
timestamp 1698175906
transform -1 0 69888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_2.x2_22
timestamp 1698175906
transform -1 0 60032 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_2.x3_17
timestamp 1698175906
transform -1 0 64064 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  COMP_2.x6_122
timestamp 1698175906
transform -1 0 63840 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  COMP_2.x6
timestamp 1698175906
transform -1 0 61040 0 1 3136
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  COMP_2.x7
timestamp 1698175906
transform 1 0 58352 0 -1 14112
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  COMP_2.x7_295
timestamp 1698175906
transform -1 0 62496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  COMP_2.x8
timestamp 1698175906
transform 1 0 55664 0 1 10976
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  COMP_2.x8_296
timestamp 1698175906
transform -1 0 58576 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  COMP_2.x9_123
timestamp 1698175906
transform -1 0 62496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  COMP_2.x9
timestamp 1698175906
transform -1 0 60144 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  COMP_2.x10 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 62048 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  COMP_2.x11
timestamp 1698175906
transform 1 0 58576 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  COMP_2.x15_5
timestamp 1698175906
transform -1 0 59584 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_2.x15_6
timestamp 1698175906
transform 1 0 58016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_3.x2_18
timestamp 1698175906
transform -1 0 50176 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_3.x3_14
timestamp 1698175906
transform -1 0 50400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  COMP_3.x6
timestamp 1698175906
transform 1 0 49168 0 1 3136
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  COMP_3.x6_124
timestamp 1698175906
transform 1 0 46144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  COMP_3.x7
timestamp 1698175906
transform 1 0 48608 0 -1 12544
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  COMP_3.x7_297
timestamp 1698175906
transform 1 0 45696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  COMP_3.x8
timestamp 1698175906
transform -1 0 50624 0 1 12544
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  COMP_3.x8_298
timestamp 1698175906
transform 1 0 49504 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  COMP_3.x9_125
timestamp 1698175906
transform -1 0 49504 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  COMP_3.x9
timestamp 1698175906
transform 1 0 48944 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  COMP_3.x10
timestamp 1698175906
transform -1 0 46704 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  COMP_3.x11
timestamp 1698175906
transform -1 0 49728 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  COMP_3.x15_7
timestamp 1698175906
transform -1 0 48160 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_3.x15_8
timestamp 1698175906
transform 1 0 46592 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_4.x2_23
timestamp 1698175906
transform 1 0 40768 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_4.x3_19
timestamp 1698175906
transform 1 0 42784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  COMP_4.x6_126
timestamp 1698175906
transform 1 0 38416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  COMP_4.x6
timestamp 1698175906
transform 1 0 40768 0 1 3136
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  COMP_4.x7
timestamp 1698175906
transform 1 0 41216 0 -1 15680
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  COMP_4.x7_299
timestamp 1698175906
transform 1 0 40768 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  COMP_4.x8_300
timestamp 1698175906
transform 1 0 41440 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  COMP_4.x8 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 43456 0 1 3136
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  COMP_4.x9_127
timestamp 1698175906
transform 1 0 40992 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  COMP_4.x9
timestamp 1698175906
transform 1 0 41216 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  COMP_4.x10
timestamp 1698175906
transform -1 0 45584 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  COMP_4.x11
timestamp 1698175906
transform -1 0 42784 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_4.x15_9
timestamp 1698175906
transform 1 0 42336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_4.x15_10
timestamp 1698175906
transform 1 0 38976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_5.x2_24
timestamp 1698175906
transform 1 0 34496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_5.x3_20
timestamp 1698175906
transform -1 0 38192 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  COMP_5.x6_128
timestamp 1698175906
transform 1 0 33264 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  COMP_5.x6
timestamp 1698175906
transform -1 0 34496 0 1 3136
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  COMP_5.x7
timestamp 1698175906
transform -1 0 28784 0 1 6272
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  COMP_5.x7_301
timestamp 1698175906
transform -1 0 31024 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  COMP_5.x8
timestamp 1698175906
transform 1 0 33712 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  COMP_5.x8_302
timestamp 1698175906
transform 1 0 33152 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  COMP_5.x9_129
timestamp 1698175906
transform 1 0 33264 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  COMP_5.x9
timestamp 1698175906
transform 1 0 33600 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  COMP_5.x10
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  COMP_5.x11
timestamp 1698175906
transform -1 0 37744 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_5.x15_11
timestamp 1698175906
transform -1 0 34496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  COMP_5.x15_12
timestamp 1698175906
transform -1 0 34944 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  CTRL._052_
timestamp 1698175906
transform 1 0 49840 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  CTRL._053_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 42896 0 -1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  CTRL._054_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 44016 0 -1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  CTRL._055_
timestamp 1698175906
transform 1 0 38864 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  CTRL._056_
timestamp 1698175906
transform 1 0 49728 0 -1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__inv_4  CTRL._057_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 46928 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  CTRL._058_
timestamp 1698175906
transform -1 0 54544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  CTRL._059_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 59472 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  CTRL._060_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 39088 0 1 53312
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  CTRL._061_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 48272 0 -1 54880
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  CTRL._062_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 36848 0 -1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  CTRL._063_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40768 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  CTRL._064_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 41328 0 -1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  CTRL._065_
timestamp 1698175906
transform 1 0 45808 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  CTRL._066_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 46032 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  CTRL._067_
timestamp 1698175906
transform -1 0 47600 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  CTRL._068_
timestamp 1698175906
transform -1 0 62384 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  CTRL._069_
timestamp 1698175906
transform -1 0 67424 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  CTRL._070_
timestamp 1698175906
transform -1 0 66304 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  CTRL._071_
timestamp 1698175906
transform 1 0 55552 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  CTRL._072_
timestamp 1698175906
transform -1 0 43008 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  CTRL._073_
timestamp 1698175906
transform 1 0 32144 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  CTRL._074_
timestamp 1698175906
transform -1 0 29680 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  CTRL._075_
timestamp 1698175906
transform -1 0 28224 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  CTRL._077_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 50624 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  CTRL._078_
timestamp 1698175906
transform -1 0 49952 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  CTRL._079_
timestamp 1698175906
transform -1 0 49280 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  CTRL._080_
timestamp 1698175906
transform 1 0 49392 0 -1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  CTRL._081_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 57904 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  CTRL._082_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 56784 0 1 53312
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  CTRL._083_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 66976 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  CTRL._084_
timestamp 1698175906
transform 1 0 57568 0 1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  CTRL._085_
timestamp 1698175906
transform -1 0 58688 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  CTRL._086_
timestamp 1698175906
transform 1 0 56784 0 -1 53312
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  CTRL._087_
timestamp 1698175906
transform 1 0 64736 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  CTRL._088_
timestamp 1698175906
transform -1 0 45248 0 -1 54880
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  CTRL._089_
timestamp 1698175906
transform -1 0 58800 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  CTRL._090_
timestamp 1698175906
transform 1 0 54208 0 1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  CTRL._091_
timestamp 1698175906
transform 1 0 56224 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  CTRL._092_
timestamp 1698175906
transform -1 0 39872 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  CTRL._093_
timestamp 1698175906
transform 1 0 40096 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  CTRL._094_
timestamp 1698175906
transform -1 0 43568 0 1 53312
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  CTRL._095_
timestamp 1698175906
transform 1 0 40768 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  CTRL._096_
timestamp 1698175906
transform -1 0 36064 0 1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  CTRL._097_
timestamp 1698175906
transform -1 0 36512 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  CTRL._098_
timestamp 1698175906
transform 1 0 33488 0 -1 53312
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  CTRL._099_
timestamp 1698175906
transform -1 0 33936 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  CTRL._100_
timestamp 1698175906
transform -1 0 36288 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  CTRL._101_
timestamp 1698175906
transform -1 0 31024 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  CTRL._102_
timestamp 1698175906
transform -1 0 31472 0 1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  CTRL._103_
timestamp 1698175906
transform 1 0 29456 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  CTRL._104_
timestamp 1698175906
transform -1 0 28784 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  CTRL._105_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28784 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  CTRL._106_
timestamp 1698175906
transform -1 0 29344 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  CTRL._107_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26768 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  CTRL._108_
timestamp 1698175906
transform 1 0 48608 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  CTRL._109_
timestamp 1698175906
transform 1 0 52528 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  CTRL._110_
timestamp 1698175906
transform 1 0 57344 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  CTRL._111_
timestamp 1698175906
transform -1 0 57680 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  CTRL._112_
timestamp 1698175906
transform -1 0 41664 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  CTRL._113_
timestamp 1698175906
transform 1 0 34272 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  CTRL._114_
timestamp 1698175906
transform -1 0 30352 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  CTRL._115_
timestamp 1698175906
transform -1 0 28336 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  CTRL._116_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 50624 0 -1 50176
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  CTRL._117_
timestamp 1698175906
transform 1 0 69776 0 1 53312
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  CTRL._118_
timestamp 1698175906
transform 1 0 65072 0 -1 53312
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  CTRL._119_
timestamp 1698175906
transform -1 0 58352 0 1 50176
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  CTRL._120_
timestamp 1698175906
transform -1 0 38640 0 -1 50176
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  CTRL._121_
timestamp 1698175906
transform 1 0 32032 0 1 48608
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  CTRL._122_
timestamp 1698175906
transform 1 0 28784 0 -1 50176
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  CTRL._123_
timestamp 1698175906
transform 1 0 25312 0 -1 50176
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  CTRL._124_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 45024 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  CTRL._125_
timestamp 1698175906
transform 1 0 50848 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  CTRL._126_
timestamp 1698175906
transform -1 0 61488 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  CTRL._127_
timestamp 1698175906
transform -1 0 63616 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  CTRL._128_
timestamp 1698175906
transform 1 0 39536 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  CTRL._129_
timestamp 1698175906
transform 1 0 33376 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  CTRL._130_
timestamp 1698175906
transform 1 0 29008 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  CTRL._131_
timestamp 1698175906
transform -1 0 26096 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  CTRL._132_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40544 0 1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  CTRL._133_
timestamp 1698175906
transform 1 0 46144 0 1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout93
timestamp 1698175906
transform 1 0 5376 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  fanout94
timestamp 1698175906
transform 1 0 5936 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout95
timestamp 1698175906
transform 1 0 17696 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout96
timestamp 1698175906
transform -1 0 7056 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout97 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 6944 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout98
timestamp 1698175906
transform -1 0 20160 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout99
timestamp 1698175906
transform -1 0 6832 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout100
timestamp 1698175906
transform 1 0 4368 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout101
timestamp 1698175906
transform -1 0 28784 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout102
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout103
timestamp 1698175906
transform 1 0 29792 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  fanout104
timestamp 1698175906
transform 1 0 42112 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout105
timestamp 1698175906
transform 1 0 64512 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout106
timestamp 1698175906
transform 1 0 53648 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout107
timestamp 1698175906
transform 1 0 52528 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout108
timestamp 1698175906
transform 1 0 67088 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout109
timestamp 1698175906
transform -1 0 75264 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout110
timestamp 1698175906
transform 1 0 74592 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout111
timestamp 1698175906
transform 1 0 87360 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  fanout112 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 73920 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout113
timestamp 1698175906
transform -1 0 6608 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout115
timestamp 1698175906
transform -1 0 50624 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  fanout116
timestamp 1698175906
transform -1 0 81312 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  fanout117
timestamp 1698175906
transform -1 0 83440 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_36 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_40 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5824 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_49 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6832 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_65 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698175906
transform 1 0 8848 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_120 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14784 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_128
timestamp 1698175906
transform 1 0 15680 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_132
timestamp 1698175906
transform 1 0 16128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_140
timestamp 1698175906
transform 1 0 17024 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_149
timestamp 1698175906
transform 1 0 18032 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165
timestamp 1698175906
transform 1 0 19824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_206
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_222
timestamp 1698175906
transform 1 0 26208 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_230
timestamp 1698175906
transform 1 0 27104 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_234
timestamp 1698175906
transform 1 0 27552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_248
timestamp 1698175906
transform 1 0 29120 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_264
timestamp 1698175906
transform 1 0 30912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_268
timestamp 1698175906
transform 1 0 31360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_280
timestamp 1698175906
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_300
timestamp 1698175906
transform 1 0 34944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_304
timestamp 1698175906
transform 1 0 35392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_312
timestamp 1698175906
transform 1 0 36288 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_316
timestamp 1698175906
transform 1 0 36736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_320
timestamp 1698175906
transform 1 0 37184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_324
timestamp 1698175906
transform 1 0 37632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_328
timestamp 1698175906
transform 1 0 38080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_332
timestamp 1698175906
transform 1 0 38528 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_350
timestamp 1698175906
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_364
timestamp 1698175906
transform 1 0 42112 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_395
timestamp 1698175906
transform 1 0 45584 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_410
timestamp 1698175906
transform 1 0 47264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_418
timestamp 1698175906
transform 1 0 48160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_422
timestamp 1698175906
transform 1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_426
timestamp 1698175906
transform 1 0 49056 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_439
timestamp 1698175906
transform 1 0 50512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_441
timestamp 1698175906
transform 1 0 50736 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_444
timestamp 1698175906
transform 1 0 51072 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_448
timestamp 1698175906
transform 1 0 51520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_452
timestamp 1698175906
transform 1 0 51968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_456
timestamp 1698175906
transform 1 0 52416 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_460
timestamp 1698175906
transform 1 0 52864 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_468
timestamp 1698175906
transform 1 0 53760 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_472
timestamp 1698175906
transform 1 0 54208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_486
timestamp 1698175906
transform 1 0 55776 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_494
timestamp 1698175906
transform 1 0 56672 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_498
timestamp 1698175906
transform 1 0 57120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_502
timestamp 1698175906
transform 1 0 57568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_512
timestamp 1698175906
transform 1 0 58688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_520
timestamp 1698175906
transform 1 0 59584 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_541
timestamp 1698175906
transform 1 0 61936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_543
timestamp 1698175906
transform 1 0 62160 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_546
timestamp 1698175906
transform 1 0 62496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_550
timestamp 1698175906
transform 1 0 62944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_554
timestamp 1698175906
transform 1 0 63392 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_570
timestamp 1698175906
transform 1 0 65184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_574
timestamp 1698175906
transform 1 0 65632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_606
timestamp 1698175906
transform 1 0 69216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_640
timestamp 1698175906
transform 1 0 73024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_644
timestamp 1698175906
transform 1 0 73472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_648
timestamp 1698175906
transform 1 0 73920 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_652
timestamp 1698175906
transform 1 0 74368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_742
timestamp 1698175906
transform 1 0 84448 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_746
timestamp 1698175906
transform 1 0 84896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_760
timestamp 1698175906
transform 1 0 86464 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_776
timestamp 1698175906
transform 1 0 88256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_780
timestamp 1698175906
transform 1 0 88704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_784
timestamp 1698175906
transform 1 0 89152 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_818
timestamp 1698175906
transform 1 0 92960 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_822
timestamp 1698175906
transform 1 0 93408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_824
timestamp 1698175906
transform 1 0 93632 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_833
timestamp 1698175906
transform 1 0 94640 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_841
timestamp 1698175906
transform 1 0 95536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_845
timestamp 1698175906
transform 1 0 95984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_847
timestamp 1698175906
transform 1 0 96208 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_862
timestamp 1698175906
transform 1 0 97888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_228
timestamp 1698175906
transform 1 0 26880 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_368
timestamp 1698175906
transform 1 0 42560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_422
timestamp 1698175906
transform 1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_424
timestamp 1698175906
transform 1 0 48832 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_437
timestamp 1698175906
transform 1 0 50288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_439
timestamp 1698175906
transform 1 0 50512 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_546
timestamp 1698175906
transform 1 0 62496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_550
timestamp 1698175906
transform 1 0 62944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_558
timestamp 1698175906
transform 1 0 63840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_690
timestamp 1698175906
transform 1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_694
timestamp 1698175906
transform 1 0 79072 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_752
timestamp 1698175906
transform 1 0 85568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_756
timestamp 1698175906
transform 1 0 86016 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_764
timestamp 1698175906
transform 1 0 86912 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_768
timestamp 1698175906
transform 1 0 87360 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_822
timestamp 1698175906
transform 1 0 93408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_838
timestamp 1698175906
transform 1 0 95200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_842
timestamp 1698175906
transform 1 0 95648 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_862
timestamp 1698175906
transform 1 0 97888 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_6
timestamp 1698175906
transform 1 0 2016 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_22
timestamp 1698175906
transform 1 0 3808 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_30
timestamp 1698175906
transform 1 0 4704 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_193
timestamp 1698175906
transform 1 0 22960 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_255
timestamp 1698175906
transform 1 0 29904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_259
timestamp 1698175906
transform 1 0 30352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_329
timestamp 1698175906
transform 1 0 38192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_387
timestamp 1698175906
transform 1 0 44688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_511
timestamp 1698175906
transform 1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_577
timestamp 1698175906
transform 1 0 65968 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_585
timestamp 1698175906
transform 1 0 66864 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_663
timestamp 1698175906
transform 1 0 75600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_717
timestamp 1698175906
transform 1 0 81648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_733
timestamp 1698175906
transform 1 0 83440 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_787
timestamp 1698175906
transform 1 0 89488 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_803
timestamp 1698175906
transform 1 0 91280 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_807
timestamp 1698175906
transform 1 0 91728 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_839
timestamp 1698175906
transform 1 0 95312 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_847
timestamp 1698175906
transform 1 0 96208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_849
timestamp 1698175906
transform 1 0 96432 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_862
timestamp 1698175906
transform 1 0 97888 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_10
timestamp 1698175906
transform 1 0 2464 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_42
timestamp 1698175906
transform 1 0 6048 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_58
timestamp 1698175906
transform 1 0 7840 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_228
timestamp 1698175906
transform 1 0 26880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_284
timestamp 1698175906
transform 1 0 33152 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_356
timestamp 1698175906
transform 1 0 41216 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_362
timestamp 1698175906
transform 1 0 41888 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_366
timestamp 1698175906
transform 1 0 42336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_422
timestamp 1698175906
transform 1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_436
timestamp 1698175906
transform 1 0 50176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_612
timestamp 1698175906
transform 1 0 69888 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_682
timestamp 1698175906
transform 1 0 77728 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_691
timestamp 1698175906
transform 1 0 78736 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_695
timestamp 1698175906
transform 1 0 79184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_699
timestamp 1698175906
transform 1 0 79632 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_752
timestamp 1698175906
transform 1 0 85568 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_768
timestamp 1698175906
transform 1 0 87360 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_822
timestamp 1698175906
transform 1 0 93408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_838
timestamp 1698175906
transform 1 0 95200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_842
timestamp 1698175906
transform 1 0 95648 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_858
timestamp 1698175906
transform 1 0 97440 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_10
timestamp 1698175906
transform 1 0 2464 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_26
timestamp 1698175906
transform 1 0 4256 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_193
timestamp 1698175906
transform 1 0 22960 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_201
timestamp 1698175906
transform 1 0 23856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_251
timestamp 1698175906
transform 1 0 29456 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_259
timestamp 1698175906
transform 1 0 30352 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_263
timestamp 1698175906
transform 1 0 30800 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_325
timestamp 1698175906
transform 1 0 37744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_329
timestamp 1698175906
transform 1 0 38192 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_333
timestamp 1698175906
transform 1 0 38640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_387
timestamp 1698175906
transform 1 0 44688 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_391
timestamp 1698175906
transform 1 0 45136 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_404
timestamp 1698175906
transform 1 0 46592 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_457
timestamp 1698175906
transform 1 0 52528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_509
timestamp 1698175906
transform 1 0 58352 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_517
timestamp 1698175906
transform 1 0 59248 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_524
timestamp 1698175906
transform 1 0 60032 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_577
timestamp 1698175906
transform 1 0 65968 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_593
timestamp 1698175906
transform 1 0 67760 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_651
timestamp 1698175906
transform 1 0 74256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_659
timestamp 1698175906
transform 1 0 75152 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_663
timestamp 1698175906
transform 1 0 75600 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_721
timestamp 1698175906
transform 1 0 82096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_725
timestamp 1698175906
transform 1 0 82544 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_733
timestamp 1698175906
transform 1 0 83440 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_787
timestamp 1698175906
transform 1 0 89488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_803
timestamp 1698175906
transform 1 0 91280 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_807
timestamp 1698175906
transform 1 0 91728 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_839
timestamp 1698175906
transform 1 0 95312 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_847
timestamp 1698175906
transform 1 0 96208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_849
timestamp 1698175906
transform 1 0 96432 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_6
timestamp 1698175906
transform 1 0 2016 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_228
timestamp 1698175906
transform 1 0 26880 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_284
timestamp 1698175906
transform 1 0 33152 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_289
timestamp 1698175906
transform 1 0 33712 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_291
timestamp 1698175906
transform 1 0 33936 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_352
timestamp 1698175906
transform 1 0 40768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_422
timestamp 1698175906
transform 1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_546
timestamp 1698175906
transform 1 0 62496 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_554
timestamp 1698175906
transform 1 0 63392 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_558
timestamp 1698175906
transform 1 0 63840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_612
timestamp 1698175906
transform 1 0 69888 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_618
timestamp 1698175906
transform 1 0 70560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_628
timestamp 1698175906
transform 1 0 71680 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_752
timestamp 1698175906
transform 1 0 85568 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_768
timestamp 1698175906
transform 1 0 87360 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_822
timestamp 1698175906
transform 1 0 93408 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_838
timestamp 1698175906
transform 1 0 95200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_842
timestamp 1698175906
transform 1 0 95648 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_858
timestamp 1698175906
transform 1 0 97440 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_263
timestamp 1698175906
transform 1 0 30800 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_333
timestamp 1698175906
transform 1 0 38640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_507
timestamp 1698175906
transform 1 0 58128 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_519
timestamp 1698175906
transform 1 0 59472 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_523
timestamp 1698175906
transform 1 0 59920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_577
timestamp 1698175906
transform 1 0 65968 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_581
timestamp 1698175906
transform 1 0 66416 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_589
timestamp 1698175906
transform 1 0 67312 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_593
timestamp 1698175906
transform 1 0 67760 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_647
timestamp 1698175906
transform 1 0 73808 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_663
timestamp 1698175906
transform 1 0 75600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_717
timestamp 1698175906
transform 1 0 81648 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_721
timestamp 1698175906
transform 1 0 82096 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_729
timestamp 1698175906
transform 1 0 82992 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_733
timestamp 1698175906
transform 1 0 83440 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_787
timestamp 1698175906
transform 1 0 89488 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_803
timestamp 1698175906
transform 1 0 91280 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_807
timestamp 1698175906
transform 1 0 91728 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_839
timestamp 1698175906
transform 1 0 95312 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_855
timestamp 1698175906
transform 1 0 97104 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_863
timestamp 1698175906
transform 1 0 98000 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_865
timestamp 1698175906
transform 1 0 98224 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_228
timestamp 1698175906
transform 1 0 26880 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_290
timestamp 1698175906
transform 1 0 33824 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_294
timestamp 1698175906
transform 1 0 34272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_298
timestamp 1698175906
transform 1 0 34720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_352
timestamp 1698175906
transform 1 0 40768 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_488
timestamp 1698175906
transform 1 0 56000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_492
timestamp 1698175906
transform 1 0 56448 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_500
timestamp 1698175906
transform 1 0 57344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_502
timestamp 1698175906
transform 1 0 57568 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_553
timestamp 1698175906
transform 1 0 63280 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_557
timestamp 1698175906
transform 1 0 63728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_559
timestamp 1698175906
transform 1 0 63952 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_612
timestamp 1698175906
transform 1 0 69888 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_628
timestamp 1698175906
transform 1 0 71680 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_682
timestamp 1698175906
transform 1 0 77728 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_698
timestamp 1698175906
transform 1 0 79520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_752
timestamp 1698175906
transform 1 0 85568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_768
timestamp 1698175906
transform 1 0 87360 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_772
timestamp 1698175906
transform 1 0 87808 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_836
timestamp 1698175906
transform 1 0 94976 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_842
timestamp 1698175906
transform 1 0 95648 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_862
timestamp 1698175906
transform 1 0 97888 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_8
timestamp 1698175906
transform 1 0 2240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_12
timestamp 1698175906
transform 1 0 2688 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_28
timestamp 1698175906
transform 1 0 4480 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698175906
transform 1 0 4928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_263
timestamp 1698175906
transform 1 0 30800 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_333
timestamp 1698175906
transform 1 0 38640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_387
timestamp 1698175906
transform 1 0 44688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_393
timestamp 1698175906
transform 1 0 45360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_401
timestamp 1698175906
transform 1 0 46256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_453
timestamp 1698175906
transform 1 0 52080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_507
timestamp 1698175906
transform 1 0 58128 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_523
timestamp 1698175906
transform 1 0 59920 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_577
timestamp 1698175906
transform 1 0 65968 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_593
timestamp 1698175906
transform 1 0 67760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_597
timestamp 1698175906
transform 1 0 68208 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_605
timestamp 1698175906
transform 1 0 69104 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_609
timestamp 1698175906
transform 1 0 69552 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_660
timestamp 1698175906
transform 1 0 75264 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_664
timestamp 1698175906
transform 1 0 75712 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_717
timestamp 1698175906
transform 1 0 81648 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_733
timestamp 1698175906
transform 1 0 83440 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_787
timestamp 1698175906
transform 1 0 89488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_803
timestamp 1698175906
transform 1 0 91280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_807
timestamp 1698175906
transform 1 0 91728 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_839
timestamp 1698175906
transform 1 0 95312 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_855
timestamp 1698175906
transform 1 0 97104 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_863
timestamp 1698175906
transform 1 0 98000 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_865
timestamp 1698175906
transform 1 0 98224 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_298
timestamp 1698175906
transform 1 0 34720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_352
timestamp 1698175906
transform 1 0 40768 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_368
timestamp 1698175906
transform 1 0 42560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_472
timestamp 1698175906
transform 1 0 54208 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_488
timestamp 1698175906
transform 1 0 56000 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_492
timestamp 1698175906
transform 1 0 56448 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_508
timestamp 1698175906
transform 1 0 58240 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_612
timestamp 1698175906
transform 1 0 69888 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_628
timestamp 1698175906
transform 1 0 71680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_688
timestamp 1698175906
transform 1 0 78400 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_696
timestamp 1698175906
transform 1 0 79296 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_752
timestamp 1698175906
transform 1 0 85568 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_768
timestamp 1698175906
transform 1 0 87360 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_772
timestamp 1698175906
transform 1 0 87808 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_836
timestamp 1698175906
transform 1 0 94976 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_842
timestamp 1698175906
transform 1 0 95648 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_8
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_12
timestamp 1698175906
transform 1 0 2688 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_28
timestamp 1698175906
transform 1 0 4480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1698175906
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_263
timestamp 1698175906
transform 1 0 30800 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_333
timestamp 1698175906
transform 1 0 38640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_387
timestamp 1698175906
transform 1 0 44688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_439
timestamp 1698175906
transform 1 0 50512 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_457
timestamp 1698175906
transform 1 0 52528 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_473
timestamp 1698175906
transform 1 0 54320 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_481
timestamp 1698175906
transform 1 0 55216 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_527
timestamp 1698175906
transform 1 0 60368 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_531
timestamp 1698175906
transform 1 0 60816 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_535
timestamp 1698175906
transform 1 0 61264 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_647
timestamp 1698175906
transform 1 0 73808 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_663
timestamp 1698175906
transform 1 0 75600 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_667
timestamp 1698175906
transform 1 0 76048 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_721
timestamp 1698175906
transform 1 0 82096 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_729
timestamp 1698175906
transform 1 0 82992 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_733
timestamp 1698175906
transform 1 0 83440 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_737
timestamp 1698175906
transform 1 0 83888 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_801
timestamp 1698175906
transform 1 0 91056 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_807
timestamp 1698175906
transform 1 0 91728 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_839
timestamp 1698175906
transform 1 0 95312 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_855
timestamp 1698175906
transform 1 0 97104 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_863
timestamp 1698175906
transform 1 0 98000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_865
timestamp 1698175906
transform 1 0 98224 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_8
timestamp 1698175906
transform 1 0 2240 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_12
timestamp 1698175906
transform 1 0 2688 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_44
timestamp 1698175906
transform 1 0 6272 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_60
timestamp 1698175906
transform 1 0 8064 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_68
timestamp 1698175906
transform 1 0 8960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_298
timestamp 1698175906
transform 1 0 34720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_352
timestamp 1698175906
transform 1 0 40768 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_360
timestamp 1698175906
transform 1 0 41664 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_364
timestamp 1698175906
transform 1 0 42112 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_415
timestamp 1698175906
transform 1 0 47824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_417
timestamp 1698175906
transform 1 0 48048 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_462
timestamp 1698175906
transform 1 0 53088 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_478
timestamp 1698175906
transform 1 0 54880 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698175906
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698175906
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_508
timestamp 1698175906
transform 1 0 58240 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_562
timestamp 1698175906
transform 1 0 64288 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_578
timestamp 1698175906
transform 1 0 66080 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_586
timestamp 1698175906
transform 1 0 66976 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_682
timestamp 1698175906
transform 1 0 77728 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_690
timestamp 1698175906
transform 1 0 78624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_694
timestamp 1698175906
transform 1 0 79072 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_698
timestamp 1698175906
transform 1 0 79520 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_745
timestamp 1698175906
transform 1 0 84784 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_761
timestamp 1698175906
transform 1 0 86576 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_769
timestamp 1698175906
transform 1 0 87472 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_772
timestamp 1698175906
transform 1 0 87808 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_836
timestamp 1698175906
transform 1 0 94976 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_842
timestamp 1698175906
transform 1 0 95648 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_367
timestamp 1698175906
transform 1 0 42448 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_383
timestamp 1698175906
transform 1 0 44240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_387
timestamp 1698175906
transform 1 0 44688 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_391
timestamp 1698175906
transform 1 0 45136 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_395
timestamp 1698175906
transform 1 0 45584 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_399
timestamp 1698175906
transform 1 0 46032 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_440
timestamp 1698175906
transform 1 0 50624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_444
timestamp 1698175906
transform 1 0 51072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_448
timestamp 1698175906
transform 1 0 51520 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_452
timestamp 1698175906
transform 1 0 51968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_454
timestamp 1698175906
transform 1 0 52192 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_457
timestamp 1698175906
transform 1 0 52528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_521
timestamp 1698175906
transform 1 0 59696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_527
timestamp 1698175906
transform 1 0 60368 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_529
timestamp 1698175906
transform 1 0 60592 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_580
timestamp 1698175906
transform 1 0 66304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_584
timestamp 1698175906
transform 1 0 66752 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_592
timestamp 1698175906
transform 1 0 67648 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_594
timestamp 1698175906
transform 1 0 67872 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_597
timestamp 1698175906
transform 1 0 68208 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_649
timestamp 1698175906
transform 1 0 74032 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_653
timestamp 1698175906
transform 1 0 74480 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_661
timestamp 1698175906
transform 1 0 75376 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_667
timestamp 1698175906
transform 1 0 76048 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_675
timestamp 1698175906
transform 1 0 76944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_677
timestamp 1698175906
transform 1 0 77168 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_728
timestamp 1698175906
transform 1 0 82880 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_732
timestamp 1698175906
transform 1 0 83328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_734
timestamp 1698175906
transform 1 0 83552 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_737
timestamp 1698175906
transform 1 0 83888 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_801
timestamp 1698175906
transform 1 0 91056 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_807
timestamp 1698175906
transform 1 0 91728 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_839
timestamp 1698175906
transform 1 0 95312 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_855
timestamp 1698175906
transform 1 0 97104 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_863
timestamp 1698175906
transform 1 0 98000 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_865
timestamp 1698175906
transform 1 0 98224 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_8
timestamp 1698175906
transform 1 0 2240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_12
timestamp 1698175906
transform 1 0 2688 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_44
timestamp 1698175906
transform 1 0 6272 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_60
timestamp 1698175906
transform 1 0 8064 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_68
timestamp 1698175906
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_290
timestamp 1698175906
transform 1 0 33824 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_294
timestamp 1698175906
transform 1 0 34272 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_352
timestamp 1698175906
transform 1 0 40768 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_360
timestamp 1698175906
transform 1 0 41664 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_414
timestamp 1698175906
transform 1 0 47712 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_418
timestamp 1698175906
transform 1 0 48160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_422
timestamp 1698175906
transform 1 0 48608 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_438
timestamp 1698175906
transform 1 0 50400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_442
timestamp 1698175906
transform 1 0 50848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_478
timestamp 1698175906
transform 1 0 54880 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_482
timestamp 1698175906
transform 1 0 55328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_486
timestamp 1698175906
transform 1 0 55776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_492
timestamp 1698175906
transform 1 0 56448 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1698175906
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_549
timestamp 1698175906
transform 1 0 62832 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_557
timestamp 1698175906
transform 1 0 63728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_559
timestamp 1698175906
transform 1 0 63952 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_562
timestamp 1698175906
transform 1 0 64288 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_626
timestamp 1698175906
transform 1 0 71456 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_638
timestamp 1698175906
transform 1 0 72800 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_646
timestamp 1698175906
transform 1 0 73696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_648
timestamp 1698175906
transform 1 0 73920 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_694
timestamp 1698175906
transform 1 0 79072 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_698
timestamp 1698175906
transform 1 0 79520 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_742
timestamp 1698175906
transform 1 0 84448 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_758
timestamp 1698175906
transform 1 0 86240 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_766
timestamp 1698175906
transform 1 0 87136 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_772
timestamp 1698175906
transform 1 0 87808 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_836
timestamp 1698175906
transform 1 0 94976 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_842
timestamp 1698175906
transform 1 0 95648 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_858
timestamp 1698175906
transform 1 0 97440 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_171
timestamp 1698175906
transform 1 0 20496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698175906
transform 1 0 28112 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_381
timestamp 1698175906
transform 1 0 44016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_387
timestamp 1698175906
transform 1 0 44688 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_423
timestamp 1698175906
transform 1 0 48720 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_457
timestamp 1698175906
transform 1 0 52528 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_521
timestamp 1698175906
transform 1 0 59696 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_527
timestamp 1698175906
transform 1 0 60368 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_591
timestamp 1698175906
transform 1 0 67536 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_597
timestamp 1698175906
transform 1 0 68208 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_605
timestamp 1698175906
transform 1 0 69104 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_609
timestamp 1698175906
transform 1 0 69552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_611
timestamp 1698175906
transform 1 0 69776 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_652
timestamp 1698175906
transform 1 0 74368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_656
timestamp 1698175906
transform 1 0 74816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_660
timestamp 1698175906
transform 1 0 75264 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_664
timestamp 1698175906
transform 1 0 75712 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_667
timestamp 1698175906
transform 1 0 76048 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_683
timestamp 1698175906
transform 1 0 77840 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_685
timestamp 1698175906
transform 1 0 78064 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_732
timestamp 1698175906
transform 1 0 83328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_734
timestamp 1698175906
transform 1 0 83552 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_737
timestamp 1698175906
transform 1 0 83888 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_801
timestamp 1698175906
transform 1 0 91056 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_807
timestamp 1698175906
transform 1 0 91728 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_839
timestamp 1698175906
transform 1 0 95312 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_847
timestamp 1698175906
transform 1 0 96208 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_851
timestamp 1698175906
transform 1 0 96656 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698175906
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_352
timestamp 1698175906
transform 1 0 40768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_396
timestamp 1698175906
transform 1 0 45696 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_412
timestamp 1698175906
transform 1 0 47488 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_422
timestamp 1698175906
transform 1 0 48608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698175906
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_492
timestamp 1698175906
transform 1 0 56448 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_556
timestamp 1698175906
transform 1 0 63616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_562
timestamp 1698175906
transform 1 0 64288 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_626
timestamp 1698175906
transform 1 0 71456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_632
timestamp 1698175906
transform 1 0 72128 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_696
timestamp 1698175906
transform 1 0 79296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_702
timestamp 1698175906
transform 1 0 79968 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_706
timestamp 1698175906
transform 1 0 80416 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_722
timestamp 1698175906
transform 1 0 82208 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_728
timestamp 1698175906
transform 1 0 82880 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_760
timestamp 1698175906
transform 1 0 86464 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_768
timestamp 1698175906
transform 1 0 87360 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_772
timestamp 1698175906
transform 1 0 87808 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_836
timestamp 1698175906
transform 1 0 94976 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_842
timestamp 1698175906
transform 1 0 95648 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_858
timestamp 1698175906
transform 1 0 97440 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698175906
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_387
timestamp 1698175906
transform 1 0 44688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1698175906
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_457
timestamp 1698175906
transform 1 0 52528 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_521
timestamp 1698175906
transform 1 0 59696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_527
timestamp 1698175906
transform 1 0 60368 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_591
timestamp 1698175906
transform 1 0 67536 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_597
timestamp 1698175906
transform 1 0 68208 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_661
timestamp 1698175906
transform 1 0 75376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_667
timestamp 1698175906
transform 1 0 76048 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_731
timestamp 1698175906
transform 1 0 83216 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_737
timestamp 1698175906
transform 1 0 83888 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_801
timestamp 1698175906
transform 1 0 91056 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_807
timestamp 1698175906
transform 1 0 91728 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_839
timestamp 1698175906
transform 1 0 95312 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_847
timestamp 1698175906
transform 1 0 96208 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_849
timestamp 1698175906
transform 1 0 96432 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_8
timestamp 1698175906
transform 1 0 2240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_12
timestamp 1698175906
transform 1 0 2688 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_44
timestamp 1698175906
transform 1 0 6272 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698175906
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698175906
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_352
timestamp 1698175906
transform 1 0 40768 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698175906
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_422
timestamp 1698175906
transform 1 0 48608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_486
timestamp 1698175906
transform 1 0 55776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_492
timestamp 1698175906
transform 1 0 56448 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_556
timestamp 1698175906
transform 1 0 63616 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_562
timestamp 1698175906
transform 1 0 64288 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_626
timestamp 1698175906
transform 1 0 71456 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_632
timestamp 1698175906
transform 1 0 72128 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_696
timestamp 1698175906
transform 1 0 79296 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_702
timestamp 1698175906
transform 1 0 79968 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_766
timestamp 1698175906
transform 1 0 87136 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_772
timestamp 1698175906
transform 1 0 87808 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_836
timestamp 1698175906
transform 1 0 94976 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_842
timestamp 1698175906
transform 1 0 95648 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_858
timestamp 1698175906
transform 1 0 97440 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_8
timestamp 1698175906
transform 1 0 2240 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_12
timestamp 1698175906
transform 1 0 2688 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698175906
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_381
timestamp 1698175906
transform 1 0 44016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_387
timestamp 1698175906
transform 1 0 44688 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698175906
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_457
timestamp 1698175906
transform 1 0 52528 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_521
timestamp 1698175906
transform 1 0 59696 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_527
timestamp 1698175906
transform 1 0 60368 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_591
timestamp 1698175906
transform 1 0 67536 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_597
timestamp 1698175906
transform 1 0 68208 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_661
timestamp 1698175906
transform 1 0 75376 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_667
timestamp 1698175906
transform 1 0 76048 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_731
timestamp 1698175906
transform 1 0 83216 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_737
timestamp 1698175906
transform 1 0 83888 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_745
timestamp 1698175906
transform 1 0 84784 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_749
timestamp 1698175906
transform 1 0 85232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_751
timestamp 1698175906
transform 1 0 85456 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_758
timestamp 1698175906
transform 1 0 86240 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_790
timestamp 1698175906
transform 1 0 89824 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_798
timestamp 1698175906
transform 1 0 90720 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_802
timestamp 1698175906
transform 1 0 91168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_804
timestamp 1698175906
transform 1 0 91392 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_807
timestamp 1698175906
transform 1 0 91728 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_839
timestamp 1698175906
transform 1 0 95312 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_847
timestamp 1698175906
transform 1 0 96208 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_849
timestamp 1698175906
transform 1 0 96432 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_8
timestamp 1698175906
transform 1 0 2240 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_40
timestamp 1698175906
transform 1 0 5824 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_56
timestamp 1698175906
transform 1 0 7616 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_64
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_352
timestamp 1698175906
transform 1 0 40768 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698175906
transform 1 0 47936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_422
timestamp 1698175906
transform 1 0 48608 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_486
timestamp 1698175906
transform 1 0 55776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_492
timestamp 1698175906
transform 1 0 56448 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_556
timestamp 1698175906
transform 1 0 63616 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_562
timestamp 1698175906
transform 1 0 64288 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_626
timestamp 1698175906
transform 1 0 71456 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_632
timestamp 1698175906
transform 1 0 72128 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_648
timestamp 1698175906
transform 1 0 73920 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_656
timestamp 1698175906
transform 1 0 74816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_664
timestamp 1698175906
transform 1 0 75712 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_696
timestamp 1698175906
transform 1 0 79296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_702
timestamp 1698175906
transform 1 0 79968 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_709
timestamp 1698175906
transform 1 0 80752 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_741
timestamp 1698175906
transform 1 0 84336 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_757
timestamp 1698175906
transform 1 0 86128 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_765
timestamp 1698175906
transform 1 0 87024 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_769
timestamp 1698175906
transform 1 0 87472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_772
timestamp 1698175906
transform 1 0 87808 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_788
timestamp 1698175906
transform 1 0 89600 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_796
timestamp 1698175906
transform 1 0 90496 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_828
timestamp 1698175906
transform 1 0 94080 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_836
timestamp 1698175906
transform 1 0 94976 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_842
timestamp 1698175906
transform 1 0 95648 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_858
timestamp 1698175906
transform 1 0 97440 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_14
timestamp 1698175906
transform 1 0 2912 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_18
timestamp 1698175906
transform 1 0 3360 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_43
timestamp 1698175906
transform 1 0 6160 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_47
timestamp 1698175906
transform 1 0 6608 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_79
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_95
timestamp 1698175906
transform 1 0 11984 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_103
timestamp 1698175906
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698175906
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698175906
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_325
timestamp 1698175906
transform 1 0 37744 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_329
timestamp 1698175906
transform 1 0 38192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_381
timestamp 1698175906
transform 1 0 44016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_387
timestamp 1698175906
transform 1 0 44688 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_451
timestamp 1698175906
transform 1 0 51856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_457
timestamp 1698175906
transform 1 0 52528 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_521
timestamp 1698175906
transform 1 0 59696 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_527
timestamp 1698175906
transform 1 0 60368 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_591
timestamp 1698175906
transform 1 0 67536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_597
timestamp 1698175906
transform 1 0 68208 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_613
timestamp 1698175906
transform 1 0 70000 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_617
timestamp 1698175906
transform 1 0 70448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_653
timestamp 1698175906
transform 1 0 74480 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_657
timestamp 1698175906
transform 1 0 74928 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_661
timestamp 1698175906
transform 1 0 75376 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_737
timestamp 1698175906
transform 1 0 83888 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_745
timestamp 1698175906
transform 1 0 84784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_747
timestamp 1698175906
transform 1 0 85008 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_784
timestamp 1698175906
transform 1 0 89152 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_800
timestamp 1698175906
transform 1 0 90944 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_804
timestamp 1698175906
transform 1 0 91392 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_807
timestamp 1698175906
transform 1 0 91728 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_839
timestamp 1698175906
transform 1 0 95312 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_847
timestamp 1698175906
transform 1 0 96208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_849
timestamp 1698175906
transform 1 0 96432 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_50
timestamp 1698175906
transform 1 0 6944 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_54
timestamp 1698175906
transform 1 0 7392 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698175906
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_146
timestamp 1698175906
transform 1 0 17696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_148
timestamp 1698175906
transform 1 0 17920 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_151
timestamp 1698175906
transform 1 0 18256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_189
timestamp 1698175906
transform 1 0 22512 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_205
timestamp 1698175906
transform 1 0 24304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_218
timestamp 1698175906
transform 1 0 25760 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_234
timestamp 1698175906
transform 1 0 27552 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_238
timestamp 1698175906
transform 1 0 28000 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_240
timestamp 1698175906
transform 1 0 28224 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_243
timestamp 1698175906
transform 1 0 28560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_247
timestamp 1698175906
transform 1 0 29008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_251
timestamp 1698175906
transform 1 0 29456 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_267
timestamp 1698175906
transform 1 0 31248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_275
timestamp 1698175906
transform 1 0 32144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698175906
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_330
timestamp 1698175906
transform 1 0 38304 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_338
timestamp 1698175906
transform 1 0 39200 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_342
timestamp 1698175906
transform 1 0 39648 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_352
timestamp 1698175906
transform 1 0 40768 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_416
timestamp 1698175906
transform 1 0 47936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_422
timestamp 1698175906
transform 1 0 48608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698175906
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_492
timestamp 1698175906
transform 1 0 56448 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_556
timestamp 1698175906
transform 1 0 63616 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_562
timestamp 1698175906
transform 1 0 64288 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_570
timestamp 1698175906
transform 1 0 65184 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_574
timestamp 1698175906
transform 1 0 65632 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_581
timestamp 1698175906
transform 1 0 66416 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_613
timestamp 1698175906
transform 1 0 70000 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_625
timestamp 1698175906
transform 1 0 71344 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_629
timestamp 1698175906
transform 1 0 71792 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_632
timestamp 1698175906
transform 1 0 72128 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_636
timestamp 1698175906
transform 1 0 72576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_638
timestamp 1698175906
transform 1 0 72800 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_660
timestamp 1698175906
transform 1 0 75264 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_676
timestamp 1698175906
transform 1 0 77056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_680
timestamp 1698175906
transform 1 0 77504 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_682
timestamp 1698175906
transform 1 0 77728 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_688
timestamp 1698175906
transform 1 0 78400 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_692
timestamp 1698175906
transform 1 0 78848 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_702
timestamp 1698175906
transform 1 0 79968 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_708
timestamp 1698175906
transform 1 0 80640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_722
timestamp 1698175906
transform 1 0 82208 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_726
timestamp 1698175906
transform 1 0 82656 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_734
timestamp 1698175906
transform 1 0 83552 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_742
timestamp 1698175906
transform 1 0 84448 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_745
timestamp 1698175906
transform 1 0 84784 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_747
timestamp 1698175906
transform 1 0 85008 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_759
timestamp 1698175906
transform 1 0 86352 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_767
timestamp 1698175906
transform 1 0 87248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_769
timestamp 1698175906
transform 1 0 87472 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_772
timestamp 1698175906
transform 1 0 87808 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_836
timestamp 1698175906
transform 1 0 94976 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_842
timestamp 1698175906
transform 1 0 95648 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_858
timestamp 1698175906
transform 1 0 97440 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_8
timestamp 1698175906
transform 1 0 2240 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_24
timestamp 1698175906
transform 1 0 4032 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_77
timestamp 1698175906
transform 1 0 9968 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_93
timestamp 1698175906
transform 1 0 11760 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_115
timestamp 1698175906
transform 1 0 14224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_153
timestamp 1698175906
transform 1 0 18480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_161
timestamp 1698175906
transform 1 0 19376 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_169
timestamp 1698175906
transform 1 0 20272 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698175906
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_261
timestamp 1698175906
transform 1 0 30576 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_277
timestamp 1698175906
transform 1 0 32368 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_281
timestamp 1698175906
transform 1 0 32816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_285
timestamp 1698175906
transform 1 0 33264 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_301
timestamp 1698175906
transform 1 0 35056 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_309
timestamp 1698175906
transform 1 0 35952 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_313
timestamp 1698175906
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_333
timestamp 1698175906
transform 1 0 38640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_335
timestamp 1698175906
transform 1 0 38864 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_372
timestamp 1698175906
transform 1 0 43008 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_383
timestamp 1698175906
transform 1 0 44240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_387
timestamp 1698175906
transform 1 0 44688 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_451
timestamp 1698175906
transform 1 0 51856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_457
timestamp 1698175906
transform 1 0 52528 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_473
timestamp 1698175906
transform 1 0 54320 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_481
timestamp 1698175906
transform 1 0 55216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_485
timestamp 1698175906
transform 1 0 55664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_492
timestamp 1698175906
transform 1 0 56448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_496
timestamp 1698175906
transform 1 0 56896 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_512
timestamp 1698175906
transform 1 0 58688 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_520
timestamp 1698175906
transform 1 0 59584 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_524
timestamp 1698175906
transform 1 0 60032 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_527
timestamp 1698175906
transform 1 0 60368 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_535
timestamp 1698175906
transform 1 0 61264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_571
timestamp 1698175906
transform 1 0 65296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_575
timestamp 1698175906
transform 1 0 65744 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_591
timestamp 1698175906
transform 1 0 67536 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_597
timestamp 1698175906
transform 1 0 68208 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_629
timestamp 1698175906
transform 1 0 71792 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_638
timestamp 1698175906
transform 1 0 72800 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_642
timestamp 1698175906
transform 1 0 73248 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_658
timestamp 1698175906
transform 1 0 75040 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_662
timestamp 1698175906
transform 1 0 75488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_664
timestamp 1698175906
transform 1 0 75712 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_667
timestamp 1698175906
transform 1 0 76048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_671
timestamp 1698175906
transform 1 0 76496 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_703
timestamp 1698175906
transform 1 0 80080 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_707
timestamp 1698175906
transform 1 0 80528 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_710
timestamp 1698175906
transform 1 0 80864 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_726
timestamp 1698175906
transform 1 0 82656 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_734
timestamp 1698175906
transform 1 0 83552 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_737
timestamp 1698175906
transform 1 0 83888 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_743
timestamp 1698175906
transform 1 0 84560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_753
timestamp 1698175906
transform 1 0 85680 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_785
timestamp 1698175906
transform 1 0 89264 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_801
timestamp 1698175906
transform 1 0 91056 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_807
timestamp 1698175906
transform 1 0 91728 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_839
timestamp 1698175906
transform 1 0 95312 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_855
timestamp 1698175906
transform 1 0 97104 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_863
timestamp 1698175906
transform 1 0 98000 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_865
timestamp 1698175906
transform 1 0 98224 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_8
timestamp 1698175906
transform 1 0 2240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_12
timestamp 1698175906
transform 1 0 2688 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_28
timestamp 1698175906
transform 1 0 4480 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_32
timestamp 1698175906
transform 1 0 4928 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_47
timestamp 1698175906
transform 1 0 6608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_51
timestamp 1698175906
transform 1 0 7056 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_67
timestamp 1698175906
transform 1 0 8848 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_112
timestamp 1698175906
transform 1 0 13888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_135
timestamp 1698175906
transform 1 0 16464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_160
timestamp 1698175906
transform 1 0 19264 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_192
timestamp 1698175906
transform 1 0 22848 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_216
timestamp 1698175906
transform 1 0 25536 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_224
timestamp 1698175906
transform 1 0 26432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_227
timestamp 1698175906
transform 1 0 26768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_284
timestamp 1698175906
transform 1 0 33152 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_319
timestamp 1698175906
transform 1 0 37072 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_341
timestamp 1698175906
transform 1 0 39536 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698175906
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_352
timestamp 1698175906
transform 1 0 40768 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_368
timestamp 1698175906
transform 1 0 42560 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_372
timestamp 1698175906
transform 1 0 43008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_374
timestamp 1698175906
transform 1 0 43232 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_382
timestamp 1698175906
transform 1 0 44128 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_414
timestamp 1698175906
transform 1 0 47712 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_418
timestamp 1698175906
transform 1 0 48160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_422
timestamp 1698175906
transform 1 0 48608 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1698175906
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_492
timestamp 1698175906
transform 1 0 56448 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_556
timestamp 1698175906
transform 1 0 63616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_567
timestamp 1698175906
transform 1 0 64848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_571
timestamp 1698175906
transform 1 0 65296 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_603
timestamp 1698175906
transform 1 0 68880 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_619
timestamp 1698175906
transform 1 0 70672 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_627
timestamp 1698175906
transform 1 0 71568 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_629
timestamp 1698175906
transform 1 0 71792 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_632
timestamp 1698175906
transform 1 0 72128 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_648
timestamp 1698175906
transform 1 0 73920 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_656
timestamp 1698175906
transform 1 0 74816 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_662
timestamp 1698175906
transform 1 0 75488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_666
timestamp 1698175906
transform 1 0 75936 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_698
timestamp 1698175906
transform 1 0 79520 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_702
timestamp 1698175906
transform 1 0 79968 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_709
timestamp 1698175906
transform 1 0 80752 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_713
timestamp 1698175906
transform 1 0 81200 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_745
timestamp 1698175906
transform 1 0 84784 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_761
timestamp 1698175906
transform 1 0 86576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_763
timestamp 1698175906
transform 1 0 86800 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_772
timestamp 1698175906
transform 1 0 87808 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_836
timestamp 1698175906
transform 1 0 94976 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_842
timestamp 1698175906
transform 1 0 95648 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_12
timestamp 1698175906
transform 1 0 2688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_16
timestamp 1698175906
transform 1 0 3136 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_71
timestamp 1698175906
transform 1 0 9296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_75
timestamp 1698175906
transform 1 0 9744 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_79
timestamp 1698175906
transform 1 0 10192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_97
timestamp 1698175906
transform 1 0 12208 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_115
timestamp 1698175906
transform 1 0 14224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_117
timestamp 1698175906
transform 1 0 14448 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_124
timestamp 1698175906
transform 1 0 15232 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_156
timestamp 1698175906
transform 1 0 18816 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698175906
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_183
timestamp 1698175906
transform 1 0 21840 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_215
timestamp 1698175906
transform 1 0 25424 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_251
timestamp 1698175906
transform 1 0 29456 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_255
timestamp 1698175906
transform 1 0 29904 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_271
timestamp 1698175906
transform 1 0 31696 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_279
timestamp 1698175906
transform 1 0 32592 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_283
timestamp 1698175906
transform 1 0 33040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_285
timestamp 1698175906
transform 1 0 33264 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_296
timestamp 1698175906
transform 1 0 34496 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698175906
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698175906
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_325
timestamp 1698175906
transform 1 0 37744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_327
timestamp 1698175906
transform 1 0 37968 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_349
timestamp 1698175906
transform 1 0 40432 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_381
timestamp 1698175906
transform 1 0 44016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_387
timestamp 1698175906
transform 1 0 44688 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_451
timestamp 1698175906
transform 1 0 51856 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_457
timestamp 1698175906
transform 1 0 52528 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_521
timestamp 1698175906
transform 1 0 59696 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_527
timestamp 1698175906
transform 1 0 60368 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_535
timestamp 1698175906
transform 1 0 61264 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_543
timestamp 1698175906
transform 1 0 62160 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_559
timestamp 1698175906
transform 1 0 63952 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_561
timestamp 1698175906
transform 1 0 64176 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_578
timestamp 1698175906
transform 1 0 66080 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_590
timestamp 1698175906
transform 1 0 67424 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_594
timestamp 1698175906
transform 1 0 67872 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_610
timestamp 1698175906
transform 1 0 69664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_614
timestamp 1698175906
transform 1 0 70112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_618
timestamp 1698175906
transform 1 0 70560 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_626
timestamp 1698175906
transform 1 0 71456 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_630
timestamp 1698175906
transform 1 0 71904 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_667
timestamp 1698175906
transform 1 0 76048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_671
timestamp 1698175906
transform 1 0 76496 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_679
timestamp 1698175906
transform 1 0 77392 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_681
timestamp 1698175906
transform 1 0 77616 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_718
timestamp 1698175906
transform 1 0 81760 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_722
timestamp 1698175906
transform 1 0 82208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_724
timestamp 1698175906
transform 1 0 82432 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_727
timestamp 1698175906
transform 1 0 82768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_733
timestamp 1698175906
transform 1 0 83440 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_737
timestamp 1698175906
transform 1 0 83888 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_748
timestamp 1698175906
transform 1 0 85120 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_780
timestamp 1698175906
transform 1 0 88704 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_796
timestamp 1698175906
transform 1 0 90496 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_804
timestamp 1698175906
transform 1 0 91392 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_807
timestamp 1698175906
transform 1 0 91728 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_839
timestamp 1698175906
transform 1 0 95312 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_855
timestamp 1698175906
transform 1 0 97104 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_863
timestamp 1698175906
transform 1 0 98000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_865
timestamp 1698175906
transform 1 0 98224 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_40
timestamp 1698175906
transform 1 0 5824 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_44
timestamp 1698175906
transform 1 0 6272 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_90
timestamp 1698175906
transform 1 0 11424 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_122
timestamp 1698175906
transform 1 0 15008 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698175906
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_158
timestamp 1698175906
transform 1 0 19040 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_166
timestamp 1698175906
transform 1 0 19936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_168
timestamp 1698175906
transform 1 0 20160 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_205
timestamp 1698175906
transform 1 0 24304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_220
timestamp 1698175906
transform 1 0 25984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_222
timestamp 1698175906
transform 1 0 26208 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_259
timestamp 1698175906
transform 1 0 30352 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_263
timestamp 1698175906
transform 1 0 30800 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_352
timestamp 1698175906
transform 1 0 40768 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_384
timestamp 1698175906
transform 1 0 44352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_388
timestamp 1698175906
transform 1 0 44800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_390
timestamp 1698175906
transform 1 0 45024 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_393
timestamp 1698175906
transform 1 0 45360 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_402
timestamp 1698175906
transform 1 0 46368 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_418
timestamp 1698175906
transform 1 0 48160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_422
timestamp 1698175906
transform 1 0 48608 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_486
timestamp 1698175906
transform 1 0 55776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_492
timestamp 1698175906
transform 1 0 56448 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_524
timestamp 1698175906
transform 1 0 60032 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_527
timestamp 1698175906
transform 1 0 60368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_529
timestamp 1698175906
transform 1 0 60592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_532
timestamp 1698175906
transform 1 0 60928 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_540
timestamp 1698175906
transform 1 0 61824 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_542
timestamp 1698175906
transform 1 0 62048 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_551
timestamp 1698175906
transform 1 0 63056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_555
timestamp 1698175906
transform 1 0 63504 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_559
timestamp 1698175906
transform 1 0 63952 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_562
timestamp 1698175906
transform 1 0 64288 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_570
timestamp 1698175906
transform 1 0 65184 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_574
timestamp 1698175906
transform 1 0 65632 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_576
timestamp 1698175906
transform 1 0 65856 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_619
timestamp 1698175906
transform 1 0 70672 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_627
timestamp 1698175906
transform 1 0 71568 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_629
timestamp 1698175906
transform 1 0 71792 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_632
timestamp 1698175906
transform 1 0 72128 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_636
timestamp 1698175906
transform 1 0 72576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_642
timestamp 1698175906
transform 1 0 73248 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_651
timestamp 1698175906
transform 1 0 74256 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_655
timestamp 1698175906
transform 1 0 74704 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_671
timestamp 1698175906
transform 1 0 76496 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_693
timestamp 1698175906
transform 1 0 78960 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_697
timestamp 1698175906
transform 1 0 79408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_699
timestamp 1698175906
transform 1 0 79632 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_702
timestamp 1698175906
transform 1 0 79968 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_710
timestamp 1698175906
transform 1 0 80864 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_713
timestamp 1698175906
transform 1 0 81200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_717
timestamp 1698175906
transform 1 0 81648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_761
timestamp 1698175906
transform 1 0 86576 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_769
timestamp 1698175906
transform 1 0 87472 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_772
timestamp 1698175906
transform 1 0 87808 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_836
timestamp 1698175906
transform 1 0 94976 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_842
timestamp 1698175906
transform 1 0 95648 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_14
timestamp 1698175906
transform 1 0 2912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_18
timestamp 1698175906
transform 1 0 3360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_22
timestamp 1698175906
transform 1 0 3808 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_30
timestamp 1698175906
transform 1 0 4704 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_69
timestamp 1698175906
transform 1 0 9072 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_77
timestamp 1698175906
transform 1 0 9968 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_94
timestamp 1698175906
transform 1 0 11872 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_98
timestamp 1698175906
transform 1 0 12320 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_123
timestamp 1698175906
transform 1 0 15120 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_161
timestamp 1698175906
transform 1 0 19376 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_165
timestamp 1698175906
transform 1 0 19824 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_192
timestamp 1698175906
transform 1 0 22848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_196
timestamp 1698175906
transform 1 0 23296 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_212
timestamp 1698175906
transform 1 0 25088 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_220
timestamp 1698175906
transform 1 0 25984 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_224
timestamp 1698175906
transform 1 0 26432 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_226
timestamp 1698175906
transform 1 0 26656 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_231
timestamp 1698175906
transform 1 0 27216 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_239
timestamp 1698175906
transform 1 0 28112 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_263
timestamp 1698175906
transform 1 0 30800 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_271
timestamp 1698175906
transform 1 0 31696 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_277
timestamp 1698175906
transform 1 0 32368 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_296
timestamp 1698175906
transform 1 0 34496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_300
timestamp 1698175906
transform 1 0 34944 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_308
timestamp 1698175906
transform 1 0 35840 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698175906
transform 1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698175906
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_325
timestamp 1698175906
transform 1 0 37744 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_329
timestamp 1698175906
transform 1 0 38192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_367
timestamp 1698175906
transform 1 0 42448 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_383
timestamp 1698175906
transform 1 0 44240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_387
timestamp 1698175906
transform 1 0 44688 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_451
timestamp 1698175906
transform 1 0 51856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_457
timestamp 1698175906
transform 1 0 52528 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_489
timestamp 1698175906
transform 1 0 56112 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_505
timestamp 1698175906
transform 1 0 57904 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_513
timestamp 1698175906
transform 1 0 58800 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_517
timestamp 1698175906
transform 1 0 59248 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_571
timestamp 1698175906
transform 1 0 65296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_575
timestamp 1698175906
transform 1 0 65744 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_591
timestamp 1698175906
transform 1 0 67536 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_597
timestamp 1698175906
transform 1 0 68208 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_613
timestamp 1698175906
transform 1 0 70000 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_621
timestamp 1698175906
transform 1 0 70896 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_628
timestamp 1698175906
transform 1 0 71680 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_660
timestamp 1698175906
transform 1 0 75264 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_664
timestamp 1698175906
transform 1 0 75712 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_667
timestamp 1698175906
transform 1 0 76048 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_674
timestamp 1698175906
transform 1 0 76832 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_706
timestamp 1698175906
transform 1 0 80416 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_722
timestamp 1698175906
transform 1 0 82208 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_730
timestamp 1698175906
transform 1 0 83104 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_734
timestamp 1698175906
transform 1 0 83552 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_737
timestamp 1698175906
transform 1 0 83888 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_801
timestamp 1698175906
transform 1 0 91056 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_807
timestamp 1698175906
transform 1 0 91728 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_839
timestamp 1698175906
transform 1 0 95312 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_855
timestamp 1698175906
transform 1 0 97104 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_863
timestamp 1698175906
transform 1 0 98000 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_865
timestamp 1698175906
transform 1 0 98224 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_36
timestamp 1698175906
transform 1 0 5376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_40
timestamp 1698175906
transform 1 0 5824 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_56
timestamp 1698175906
transform 1 0 7616 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_64
timestamp 1698175906
transform 1 0 8512 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_96
timestamp 1698175906
transform 1 0 12096 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698175906
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_220
timestamp 1698175906
transform 1 0 25984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_258
timestamp 1698175906
transform 1 0 30240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_262
timestamp 1698175906
transform 1 0 30688 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_270
timestamp 1698175906
transform 1 0 31584 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_316
timestamp 1698175906
transform 1 0 36736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_320
timestamp 1698175906
transform 1 0 37184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 37408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_325
timestamp 1698175906
transform 1 0 37744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_344
timestamp 1698175906
transform 1 0 39872 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_352
timestamp 1698175906
transform 1 0 40768 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_368
timestamp 1698175906
transform 1 0 42560 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_378
timestamp 1698175906
transform 1 0 43680 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_382
timestamp 1698175906
transform 1 0 44128 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_385
timestamp 1698175906
transform 1 0 44464 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_417
timestamp 1698175906
transform 1 0 48048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_419
timestamp 1698175906
transform 1 0 48272 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_422
timestamp 1698175906
transform 1 0 48608 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_486
timestamp 1698175906
transform 1 0 55776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_492
timestamp 1698175906
transform 1 0 56448 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_524
timestamp 1698175906
transform 1 0 60032 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_532
timestamp 1698175906
transform 1 0 60928 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_548
timestamp 1698175906
transform 1 0 62720 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_556
timestamp 1698175906
transform 1 0 63616 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_562
timestamp 1698175906
transform 1 0 64288 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_578
timestamp 1698175906
transform 1 0 66080 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_616
timestamp 1698175906
transform 1 0 70336 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_624
timestamp 1698175906
transform 1 0 71232 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_628
timestamp 1698175906
transform 1 0 71680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_632
timestamp 1698175906
transform 1 0 72128 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_648
timestamp 1698175906
transform 1 0 73920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_655
timestamp 1698175906
transform 1 0 74704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_659
timestamp 1698175906
transform 1 0 75152 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_677
timestamp 1698175906
transform 1 0 77168 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_692
timestamp 1698175906
transform 1 0 78848 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_702
timestamp 1698175906
transform 1 0 79968 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_718
timestamp 1698175906
transform 1 0 81760 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_726
timestamp 1698175906
transform 1 0 82656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_728
timestamp 1698175906
transform 1 0 82880 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_735
timestamp 1698175906
transform 1 0 83664 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_767
timestamp 1698175906
transform 1 0 87248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_769
timestamp 1698175906
transform 1 0 87472 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_772
timestamp 1698175906
transform 1 0 87808 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_836
timestamp 1698175906
transform 1 0 94976 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_842
timestamp 1698175906
transform 1 0 95648 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_850
timestamp 1698175906
transform 1 0 96544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_8
timestamp 1698175906
transform 1 0 2240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_12
timestamp 1698175906
transform 1 0 2688 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_71
timestamp 1698175906
transform 1 0 9296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_75
timestamp 1698175906
transform 1 0 9744 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_79
timestamp 1698175906
transform 1 0 10192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_95
timestamp 1698175906
transform 1 0 11984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_99
timestamp 1698175906
transform 1 0 12432 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_103
timestamp 1698175906
transform 1 0 12880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_139
timestamp 1698175906
transform 1 0 16912 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_155
timestamp 1698175906
transform 1 0 18704 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_163
timestamp 1698175906
transform 1 0 19600 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_167
timestamp 1698175906
transform 1 0 20048 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_209
timestamp 1698175906
transform 1 0 24752 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_215
timestamp 1698175906
transform 1 0 25424 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_238
timestamp 1698175906
transform 1 0 28000 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_279
timestamp 1698175906
transform 1 0 32592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_281
timestamp 1698175906
transform 1 0 32816 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_288
timestamp 1698175906
transform 1 0 33600 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_294
timestamp 1698175906
transform 1 0 34272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_306
timestamp 1698175906
transform 1 0 35616 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698175906
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_343
timestamp 1698175906
transform 1 0 39760 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_359
timestamp 1698175906
transform 1 0 41552 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_367
timestamp 1698175906
transform 1 0 42448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_377
timestamp 1698175906
transform 1 0 43568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_421
timestamp 1698175906
transform 1 0 48496 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_453
timestamp 1698175906
transform 1 0 52080 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_457
timestamp 1698175906
transform 1 0 52528 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_467
timestamp 1698175906
transform 1 0 53648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_469
timestamp 1698175906
transform 1 0 53872 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_504
timestamp 1698175906
transform 1 0 57792 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_508
timestamp 1698175906
transform 1 0 58240 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_524
timestamp 1698175906
transform 1 0 60032 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_527
timestamp 1698175906
transform 1 0 60368 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_535
timestamp 1698175906
transform 1 0 61264 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_551
timestamp 1698175906
transform 1 0 63056 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_555
timestamp 1698175906
transform 1 0 63504 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_563
timestamp 1698175906
transform 1 0 64400 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_567
timestamp 1698175906
transform 1 0 64848 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_573
timestamp 1698175906
transform 1 0 65520 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_577
timestamp 1698175906
transform 1 0 65968 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_593
timestamp 1698175906
transform 1 0 67760 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_597
timestamp 1698175906
transform 1 0 68208 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_599
timestamp 1698175906
transform 1 0 68432 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_605
timestamp 1698175906
transform 1 0 69104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_609
timestamp 1698175906
transform 1 0 69552 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_625
timestamp 1698175906
transform 1 0 71344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_667
timestamp 1698175906
transform 1 0 76048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_671
timestamp 1698175906
transform 1 0 76496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_675
timestamp 1698175906
transform 1 0 76944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_685
timestamp 1698175906
transform 1 0 78064 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_720
timestamp 1698175906
transform 1 0 81984 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_728
timestamp 1698175906
transform 1 0 82880 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_732
timestamp 1698175906
transform 1 0 83328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_734
timestamp 1698175906
transform 1 0 83552 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_737
timestamp 1698175906
transform 1 0 83888 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_801
timestamp 1698175906
transform 1 0 91056 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_807
timestamp 1698175906
transform 1 0 91728 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_839
timestamp 1698175906
transform 1 0 95312 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_855
timestamp 1698175906
transform 1 0 97104 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_863
timestamp 1698175906
transform 1 0 98000 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_865
timestamp 1698175906
transform 1 0 98224 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_8
timestamp 1698175906
transform 1 0 2240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_12
timestamp 1698175906
transform 1 0 2688 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_28
timestamp 1698175906
transform 1 0 4480 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_32
timestamp 1698175906
transform 1 0 4928 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_37
timestamp 1698175906
transform 1 0 5488 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_69
timestamp 1698175906
transform 1 0 9072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_80
timestamp 1698175906
transform 1 0 10304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_92
timestamp 1698175906
transform 1 0 11648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_96
timestamp 1698175906
transform 1 0 12096 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_128
timestamp 1698175906
transform 1 0 15680 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698175906
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_158
timestamp 1698175906
transform 1 0 19040 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_195
timestamp 1698175906
transform 1 0 23184 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_203
timestamp 1698175906
transform 1 0 24080 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698175906
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_220
timestamp 1698175906
transform 1 0 25984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_228
timestamp 1698175906
transform 1 0 26880 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_260
timestamp 1698175906
transform 1 0 30464 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_352
timestamp 1698175906
transform 1 0 40768 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_416
timestamp 1698175906
transform 1 0 47936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_422
timestamp 1698175906
transform 1 0 48608 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_426
timestamp 1698175906
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_428
timestamp 1698175906
transform 1 0 49280 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_481
timestamp 1698175906
transform 1 0 55216 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_489
timestamp 1698175906
transform 1 0 56112 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_492
timestamp 1698175906
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_496
timestamp 1698175906
transform 1 0 56896 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_499
timestamp 1698175906
transform 1 0 57232 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_503
timestamp 1698175906
transform 1 0 57680 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_512
timestamp 1698175906
transform 1 0 58688 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_527
timestamp 1698175906
transform 1 0 60368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_529
timestamp 1698175906
transform 1 0 60592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_532
timestamp 1698175906
transform 1 0 60928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_540
timestamp 1698175906
transform 1 0 61824 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_546
timestamp 1698175906
transform 1 0 62496 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_554
timestamp 1698175906
transform 1 0 63392 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_558
timestamp 1698175906
transform 1 0 63840 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_562
timestamp 1698175906
transform 1 0 64288 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_578
timestamp 1698175906
transform 1 0 66080 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_594
timestamp 1698175906
transform 1 0 67872 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_598
timestamp 1698175906
transform 1 0 68320 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_632
timestamp 1698175906
transform 1 0 72128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_642
timestamp 1698175906
transform 1 0 73248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_646
timestamp 1698175906
transform 1 0 73696 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_654
timestamp 1698175906
transform 1 0 74592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_671
timestamp 1698175906
transform 1 0 76496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_675
timestamp 1698175906
transform 1 0 76944 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_678
timestamp 1698175906
transform 1 0 77280 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_682
timestamp 1698175906
transform 1 0 77728 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_686
timestamp 1698175906
transform 1 0 78176 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_694
timestamp 1698175906
transform 1 0 79072 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_698
timestamp 1698175906
transform 1 0 79520 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_702
timestamp 1698175906
transform 1 0 79968 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_734
timestamp 1698175906
transform 1 0 83552 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_742
timestamp 1698175906
transform 1 0 84448 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_758
timestamp 1698175906
transform 1 0 86240 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_766
timestamp 1698175906
transform 1 0 87136 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_772
timestamp 1698175906
transform 1 0 87808 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_836
timestamp 1698175906
transform 1 0 94976 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_842
timestamp 1698175906
transform 1 0 95648 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_858
timestamp 1698175906
transform 1 0 97440 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_14
timestamp 1698175906
transform 1 0 2912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_18
timestamp 1698175906
transform 1 0 3360 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_41
timestamp 1698175906
transform 1 0 5936 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_49
timestamp 1698175906
transform 1 0 6832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_85
timestamp 1698175906
transform 1 0 10864 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_109
timestamp 1698175906
transform 1 0 13552 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_144
timestamp 1698175906
transform 1 0 17472 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_148
timestamp 1698175906
transform 1 0 17920 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_156
timestamp 1698175906
transform 1 0 18816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_160
timestamp 1698175906
transform 1 0 19264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_162
timestamp 1698175906
transform 1 0 19488 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_167
timestamp 1698175906
transform 1 0 20048 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_171
timestamp 1698175906
transform 1 0 20496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_192
timestamp 1698175906
transform 1 0 22848 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_196
timestamp 1698175906
transform 1 0 23296 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_228
timestamp 1698175906
transform 1 0 26880 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_253
timestamp 1698175906
transform 1 0 29680 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_272
timestamp 1698175906
transform 1 0 31808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_276
timestamp 1698175906
transform 1 0 32256 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_292
timestamp 1698175906
transform 1 0 34048 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_300
timestamp 1698175906
transform 1 0 34944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_308
timestamp 1698175906
transform 1 0 35840 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1698175906
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698175906
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_325
timestamp 1698175906
transform 1 0 37744 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_329
timestamp 1698175906
transform 1 0 38192 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_361
timestamp 1698175906
transform 1 0 41776 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_377
timestamp 1698175906
transform 1 0 43568 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_387
timestamp 1698175906
transform 1 0 44688 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698175906
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_457
timestamp 1698175906
transform 1 0 52528 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_465
timestamp 1698175906
transform 1 0 53424 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_469
timestamp 1698175906
transform 1 0 53872 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_475
timestamp 1698175906
transform 1 0 54544 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_491
timestamp 1698175906
transform 1 0 56336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_501
timestamp 1698175906
transform 1 0 57456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_512
timestamp 1698175906
transform 1 0 58688 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_520
timestamp 1698175906
transform 1 0 59584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_522
timestamp 1698175906
transform 1 0 59808 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_542
timestamp 1698175906
transform 1 0 62048 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_580
timestamp 1698175906
transform 1 0 66304 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_584
timestamp 1698175906
transform 1 0 66752 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_586
timestamp 1698175906
transform 1 0 66976 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_593
timestamp 1698175906
transform 1 0 67760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_597
timestamp 1698175906
transform 1 0 68208 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_629
timestamp 1698175906
transform 1 0 71792 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_645
timestamp 1698175906
transform 1 0 73584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_663
timestamp 1698175906
transform 1 0 75600 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_667
timestamp 1698175906
transform 1 0 76048 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_676
timestamp 1698175906
transform 1 0 77056 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_683
timestamp 1698175906
transform 1 0 77840 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_687
timestamp 1698175906
transform 1 0 78288 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_719
timestamp 1698175906
transform 1 0 81872 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_737
timestamp 1698175906
transform 1 0 83888 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_801
timestamp 1698175906
transform 1 0 91056 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_807
timestamp 1698175906
transform 1 0 91728 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_839
timestamp 1698175906
transform 1 0 95312 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_847
timestamp 1698175906
transform 1 0 96208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_849
timestamp 1698175906
transform 1 0 96432 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_862
timestamp 1698175906
transform 1 0 97888 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_55
timestamp 1698175906
transform 1 0 7504 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_63
timestamp 1698175906
transform 1 0 8400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_67
timestamp 1698175906
transform 1 0 8848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_69
timestamp 1698175906
transform 1 0 9072 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_88
timestamp 1698175906
transform 1 0 11200 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_92
timestamp 1698175906
transform 1 0 11648 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_120
timestamp 1698175906
transform 1 0 14784 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_174
timestamp 1698175906
transform 1 0 20832 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_190
timestamp 1698175906
transform 1 0 22624 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_198
timestamp 1698175906
transform 1 0 23520 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_202
timestamp 1698175906
transform 1 0 23968 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_286
timestamp 1698175906
transform 1 0 33376 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_294
timestamp 1698175906
transform 1 0 34272 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_298
timestamp 1698175906
transform 1 0 34720 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_335
timestamp 1698175906
transform 1 0 38864 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_343
timestamp 1698175906
transform 1 0 39760 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_388
timestamp 1698175906
transform 1 0 44800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_404
timestamp 1698175906
transform 1 0 46592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_408
timestamp 1698175906
transform 1 0 47040 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_416
timestamp 1698175906
transform 1 0 47936 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_458
timestamp 1698175906
transform 1 0 52640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_462
timestamp 1698175906
transform 1 0 53088 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_478
timestamp 1698175906
transform 1 0 54880 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_481
timestamp 1698175906
transform 1 0 55216 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_485
timestamp 1698175906
transform 1 0 55664 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_487
timestamp 1698175906
transform 1 0 55888 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_526
timestamp 1698175906
transform 1 0 60256 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_558
timestamp 1698175906
transform 1 0 63840 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_562
timestamp 1698175906
transform 1 0 64288 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_570
timestamp 1698175906
transform 1 0 65184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_577
timestamp 1698175906
transform 1 0 65968 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_581
timestamp 1698175906
transform 1 0 66416 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_613
timestamp 1698175906
transform 1 0 70000 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_622
timestamp 1698175906
transform 1 0 71008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_626
timestamp 1698175906
transform 1 0 71456 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_632
timestamp 1698175906
transform 1 0 72128 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_640
timestamp 1698175906
transform 1 0 73024 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_657
timestamp 1698175906
transform 1 0 74928 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_661
timestamp 1698175906
transform 1 0 75376 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_663
timestamp 1698175906
transform 1 0 75600 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_702
timestamp 1698175906
transform 1 0 79968 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_766
timestamp 1698175906
transform 1 0 87136 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_772
timestamp 1698175906
transform 1 0 87808 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_836
timestamp 1698175906
transform 1 0 94976 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_842
timestamp 1698175906
transform 1 0 95648 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_858
timestamp 1698175906
transform 1 0 97440 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_8
timestamp 1698175906
transform 1 0 2240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_12
timestamp 1698175906
transform 1 0 2688 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_28
timestamp 1698175906
transform 1 0 4480 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_32
timestamp 1698175906
transform 1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_57
timestamp 1698175906
transform 1 0 7728 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_89
timestamp 1698175906
transform 1 0 11312 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_109
timestamp 1698175906
transform 1 0 13552 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_112
timestamp 1698175906
transform 1 0 13888 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_144
timestamp 1698175906
transform 1 0 17472 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_160
timestamp 1698175906
transform 1 0 19264 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_168
timestamp 1698175906
transform 1 0 20160 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698175906
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_193
timestamp 1698175906
transform 1 0 22960 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_201
timestamp 1698175906
transform 1 0 23856 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_203
timestamp 1698175906
transform 1 0 24080 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_225
timestamp 1698175906
transform 1 0 26544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_229
timestamp 1698175906
transform 1 0 26992 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_251
timestamp 1698175906
transform 1 0 29456 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_255
timestamp 1698175906
transform 1 0 29904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_267
timestamp 1698175906
transform 1 0 31248 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_299
timestamp 1698175906
transform 1 0 34832 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_307
timestamp 1698175906
transform 1 0 35728 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_349
timestamp 1698175906
transform 1 0 40432 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_353
timestamp 1698175906
transform 1 0 40880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_355
timestamp 1698175906
transform 1 0 41104 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_362
timestamp 1698175906
transform 1 0 41888 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_378
timestamp 1698175906
transform 1 0 43680 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_382
timestamp 1698175906
transform 1 0 44128 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_423
timestamp 1698175906
transform 1 0 48720 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_457
timestamp 1698175906
transform 1 0 52528 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_473
timestamp 1698175906
transform 1 0 54320 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_515
timestamp 1698175906
transform 1 0 59024 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_523
timestamp 1698175906
transform 1 0 59920 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_527
timestamp 1698175906
transform 1 0 60368 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_529
timestamp 1698175906
transform 1 0 60592 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_542
timestamp 1698175906
transform 1 0 62048 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_546
timestamp 1698175906
transform 1 0 62496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_548
timestamp 1698175906
transform 1 0 62720 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_561
timestamp 1698175906
transform 1 0 64176 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_565
timestamp 1698175906
transform 1 0 64624 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_581
timestamp 1698175906
transform 1 0 66416 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_631
timestamp 1698175906
transform 1 0 72016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_639
timestamp 1698175906
transform 1 0 72912 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_647
timestamp 1698175906
transform 1 0 73808 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_685
timestamp 1698175906
transform 1 0 78064 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_717
timestamp 1698175906
transform 1 0 81648 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_733
timestamp 1698175906
transform 1 0 83440 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_737
timestamp 1698175906
transform 1 0 83888 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_801
timestamp 1698175906
transform 1 0 91056 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_807
timestamp 1698175906
transform 1 0 91728 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_839
timestamp 1698175906
transform 1 0 95312 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_847
timestamp 1698175906
transform 1 0 96208 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_849
timestamp 1698175906
transform 1 0 96432 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_862
timestamp 1698175906
transform 1 0 97888 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_41
timestamp 1698175906
transform 1 0 5936 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_57
timestamp 1698175906
transform 1 0 7728 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_65
timestamp 1698175906
transform 1 0 8624 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_69
timestamp 1698175906
transform 1 0 9072 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_186
timestamp 1698175906
transform 1 0 22176 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_190
timestamp 1698175906
transform 1 0 22624 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_314
timestamp 1698175906
transform 1 0 36512 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_330
timestamp 1698175906
transform 1 0 38304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_332
timestamp 1698175906
transform 1 0 38528 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_341
timestamp 1698175906
transform 1 0 39536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_345
timestamp 1698175906
transform 1 0 39984 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_349
timestamp 1698175906
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_352
timestamp 1698175906
transform 1 0 40768 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_360
timestamp 1698175906
transform 1 0 41664 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_377
timestamp 1698175906
transform 1 0 43568 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_392
timestamp 1698175906
transform 1 0 45248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_405
timestamp 1698175906
transform 1 0 46704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_409
timestamp 1698175906
transform 1 0 47152 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_417
timestamp 1698175906
transform 1 0 48048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_419
timestamp 1698175906
transform 1 0 48272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_422
timestamp 1698175906
transform 1 0 48608 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_430
timestamp 1698175906
transform 1 0 49504 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_470
timestamp 1698175906
transform 1 0 53984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_474
timestamp 1698175906
transform 1 0 54432 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_482
timestamp 1698175906
transform 1 0 55328 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_492
timestamp 1698175906
transform 1 0 56448 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_499
timestamp 1698175906
transform 1 0 57232 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_503
timestamp 1698175906
transform 1 0 57680 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_535
timestamp 1698175906
transform 1 0 61264 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_551
timestamp 1698175906
transform 1 0 63056 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_559
timestamp 1698175906
transform 1 0 63952 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_562
timestamp 1698175906
transform 1 0 64288 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_594
timestamp 1698175906
transform 1 0 67872 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_596
timestamp 1698175906
transform 1 0 68096 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_607
timestamp 1698175906
transform 1 0 69328 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_611
timestamp 1698175906
transform 1 0 69776 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_627
timestamp 1698175906
transform 1 0 71568 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_629
timestamp 1698175906
transform 1 0 71792 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_632
timestamp 1698175906
transform 1 0 72128 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_664
timestamp 1698175906
transform 1 0 75712 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_667
timestamp 1698175906
transform 1 0 76048 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_699
timestamp 1698175906
transform 1 0 79632 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_702
timestamp 1698175906
transform 1 0 79968 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_766
timestamp 1698175906
transform 1 0 87136 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_772
timestamp 1698175906
transform 1 0 87808 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_836
timestamp 1698175906
transform 1 0 94976 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_842
timestamp 1698175906
transform 1 0 95648 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_858
timestamp 1698175906
transform 1 0 97440 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_8
timestamp 1698175906
transform 1 0 2240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_12
timestamp 1698175906
transform 1 0 2688 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_28
timestamp 1698175906
transform 1 0 4480 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_32
timestamp 1698175906
transform 1 0 4928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_53
timestamp 1698175906
transform 1 0 7280 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_61
timestamp 1698175906
transform 1 0 8176 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_136
timestamp 1698175906
transform 1 0 16576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_140
timestamp 1698175906
transform 1 0 17024 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_172
timestamp 1698175906
transform 1 0 20608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698175906
transform 1 0 20832 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_209
timestamp 1698175906
transform 1 0 24752 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_217
timestamp 1698175906
transform 1 0 25648 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_221
timestamp 1698175906
transform 1 0 26096 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_224
timestamp 1698175906
transform 1 0 26432 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_243
timestamp 1698175906
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_255
timestamp 1698175906
transform 1 0 29904 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_257
timestamp 1698175906
transform 1 0 30128 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_260
timestamp 1698175906
transform 1 0 30464 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_268
timestamp 1698175906
transform 1 0 31360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_276
timestamp 1698175906
transform 1 0 32256 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_282
timestamp 1698175906
transform 1 0 32928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_286
timestamp 1698175906
transform 1 0 33376 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_302
timestamp 1698175906
transform 1 0 35168 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_310
timestamp 1698175906
transform 1 0 36064 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698175906
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_322
timestamp 1698175906
transform 1 0 37408 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_338
timestamp 1698175906
transform 1 0 39200 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_346
timestamp 1698175906
transform 1 0 40096 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_387
timestamp 1698175906
transform 1 0 44688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_430
timestamp 1698175906
transform 1 0 49504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_434
timestamp 1698175906
transform 1 0 49952 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_439
timestamp 1698175906
transform 1 0 50512 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_447
timestamp 1698175906
transform 1 0 51408 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_451
timestamp 1698175906
transform 1 0 51856 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_519
timestamp 1698175906
transform 1 0 59472 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_523
timestamp 1698175906
transform 1 0 59920 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_527
timestamp 1698175906
transform 1 0 60368 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_559
timestamp 1698175906
transform 1 0 63952 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_575
timestamp 1698175906
transform 1 0 65744 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_579
timestamp 1698175906
transform 1 0 66192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_586
timestamp 1698175906
transform 1 0 66976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_590
timestamp 1698175906
transform 1 0 67424 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_594
timestamp 1698175906
transform 1 0 67872 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_597
timestamp 1698175906
transform 1 0 68208 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_629
timestamp 1698175906
transform 1 0 71792 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_633
timestamp 1698175906
transform 1 0 72240 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_640
timestamp 1698175906
transform 1 0 73024 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_656
timestamp 1698175906
transform 1 0 74816 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_664
timestamp 1698175906
transform 1 0 75712 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_667
timestamp 1698175906
transform 1 0 76048 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_731
timestamp 1698175906
transform 1 0 83216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_737
timestamp 1698175906
transform 1 0 83888 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_753
timestamp 1698175906
transform 1 0 85680 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_785
timestamp 1698175906
transform 1 0 89264 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_801
timestamp 1698175906
transform 1 0 91056 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_807
timestamp 1698175906
transform 1 0 91728 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_839
timestamp 1698175906
transform 1 0 95312 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_847
timestamp 1698175906
transform 1 0 96208 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_849
timestamp 1698175906
transform 1 0 96432 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_36
timestamp 1698175906
transform 1 0 5376 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_68
timestamp 1698175906
transform 1 0 8960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_104
timestamp 1698175906
transform 1 0 12992 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_112
timestamp 1698175906
transform 1 0 13888 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_116
timestamp 1698175906
transform 1 0 14336 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_118
timestamp 1698175906
transform 1 0 14560 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_121
timestamp 1698175906
transform 1 0 14896 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_137
timestamp 1698175906
transform 1 0 16688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698175906
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_158
timestamp 1698175906
transform 1 0 19040 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_168
timestamp 1698175906
transform 1 0 20160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_220
timestamp 1698175906
transform 1 0 25984 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_256
timestamp 1698175906
transform 1 0 30016 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_277
timestamp 1698175906
transform 1 0 32368 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_279
timestamp 1698175906
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_316
timestamp 1698175906
transform 1 0 36736 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_332
timestamp 1698175906
transform 1 0 38528 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_334
timestamp 1698175906
transform 1 0 38752 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_337
timestamp 1698175906
transform 1 0 39088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_352
timestamp 1698175906
transform 1 0 40768 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_368
timestamp 1698175906
transform 1 0 42560 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_371
timestamp 1698175906
transform 1 0 42896 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_411
timestamp 1698175906
transform 1 0 47376 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_419
timestamp 1698175906
transform 1 0 48272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_422
timestamp 1698175906
transform 1 0 48608 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_486
timestamp 1698175906
transform 1 0 55776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_492
timestamp 1698175906
transform 1 0 56448 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_524
timestamp 1698175906
transform 1 0 60032 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_532
timestamp 1698175906
transform 1 0 60928 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_539
timestamp 1698175906
transform 1 0 61712 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_555
timestamp 1698175906
transform 1 0 63504 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_559
timestamp 1698175906
transform 1 0 63952 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_562
timestamp 1698175906
transform 1 0 64288 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_566
timestamp 1698175906
transform 1 0 64736 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_601
timestamp 1698175906
transform 1 0 68656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_605
timestamp 1698175906
transform 1 0 69104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_617
timestamp 1698175906
transform 1 0 70448 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_621
timestamp 1698175906
transform 1 0 70896 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_629
timestamp 1698175906
transform 1 0 71792 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_637
timestamp 1698175906
transform 1 0 72688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_641
timestamp 1698175906
transform 1 0 73136 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_673
timestamp 1698175906
transform 1 0 76720 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_689
timestamp 1698175906
transform 1 0 78512 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_697
timestamp 1698175906
transform 1 0 79408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_699
timestamp 1698175906
transform 1 0 79632 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_702
timestamp 1698175906
transform 1 0 79968 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_766
timestamp 1698175906
transform 1 0 87136 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_772
timestamp 1698175906
transform 1 0 87808 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_836
timestamp 1698175906
transform 1 0 94976 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_842
timestamp 1698175906
transform 1 0 95648 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_858
timestamp 1698175906
transform 1 0 97440 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_12
timestamp 1698175906
transform 1 0 2688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_16
timestamp 1698175906
transform 1 0 3136 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_24
timestamp 1698175906
transform 1 0 4032 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_28
timestamp 1698175906
transform 1 0 4480 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_30
timestamp 1698175906
transform 1 0 4704 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_71
timestamp 1698175906
transform 1 0 9296 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_103
timestamp 1698175906
transform 1 0 12880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_115
timestamp 1698175906
transform 1 0 14224 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_150
timestamp 1698175906
transform 1 0 18144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_154
timestamp 1698175906
transform 1 0 18592 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_170
timestamp 1698175906
transform 1 0 20384 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_174
timestamp 1698175906
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_209
timestamp 1698175906
transform 1 0 24752 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_225
timestamp 1698175906
transform 1 0 26544 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_236
timestamp 1698175906
transform 1 0 27776 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_244
timestamp 1698175906
transform 1 0 28672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_255
timestamp 1698175906
transform 1 0 29904 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_258
timestamp 1698175906
transform 1 0 30240 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_274
timestamp 1698175906
transform 1 0 32032 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_282
timestamp 1698175906
transform 1 0 32928 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_298
timestamp 1698175906
transform 1 0 34720 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_306
timestamp 1698175906
transform 1 0 35616 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_325
timestamp 1698175906
transform 1 0 37744 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_329
timestamp 1698175906
transform 1 0 38192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_333
timestamp 1698175906
transform 1 0 38640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_369
timestamp 1698175906
transform 1 0 42672 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_383
timestamp 1698175906
transform 1 0 44240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_413
timestamp 1698175906
transform 1 0 47600 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_429
timestamp 1698175906
transform 1 0 49392 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_437
timestamp 1698175906
transform 1 0 50288 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_447
timestamp 1698175906
transform 1 0 51408 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_457
timestamp 1698175906
transform 1 0 52528 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_463
timestamp 1698175906
transform 1 0 53200 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_479
timestamp 1698175906
transform 1 0 54992 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_483
timestamp 1698175906
transform 1 0 55440 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_495
timestamp 1698175906
transform 1 0 56784 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_511
timestamp 1698175906
transform 1 0 58576 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_519
timestamp 1698175906
transform 1 0 59472 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_561
timestamp 1698175906
transform 1 0 64176 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_565
timestamp 1698175906
transform 1 0 64624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_567
timestamp 1698175906
transform 1 0 64848 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_580
timestamp 1698175906
transform 1 0 66304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_584
timestamp 1698175906
transform 1 0 66752 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_592
timestamp 1698175906
transform 1 0 67648 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_594
timestamp 1698175906
transform 1 0 67872 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_597
timestamp 1698175906
transform 1 0 68208 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_599
timestamp 1698175906
transform 1 0 68432 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_640
timestamp 1698175906
transform 1 0 73024 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_654
timestamp 1698175906
transform 1 0 74592 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_662
timestamp 1698175906
transform 1 0 75488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_664
timestamp 1698175906
transform 1 0 75712 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_667
timestamp 1698175906
transform 1 0 76048 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_731
timestamp 1698175906
transform 1 0 83216 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_737
timestamp 1698175906
transform 1 0 83888 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_801
timestamp 1698175906
transform 1 0 91056 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_807
timestamp 1698175906
transform 1 0 91728 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_839
timestamp 1698175906
transform 1 0 95312 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_847
timestamp 1698175906
transform 1 0 96208 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_849
timestamp 1698175906
transform 1 0 96432 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_8
timestamp 1698175906
transform 1 0 2240 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_12
timestamp 1698175906
transform 1 0 2688 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_44
timestamp 1698175906
transform 1 0 6272 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_60
timestamp 1698175906
transform 1 0 8064 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_108
timestamp 1698175906
transform 1 0 13440 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_116
timestamp 1698175906
transform 1 0 14336 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_118
timestamp 1698175906
transform 1 0 14560 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_129
timestamp 1698175906
transform 1 0 15792 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_137
timestamp 1698175906
transform 1 0 16688 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_139
timestamp 1698175906
transform 1 0 16912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_158
timestamp 1698175906
transform 1 0 19040 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_166
timestamp 1698175906
transform 1 0 19936 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_168
timestamp 1698175906
transform 1 0 20160 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_205
timestamp 1698175906
transform 1 0 24304 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_209
timestamp 1698175906
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_216
timestamp 1698175906
transform 1 0 25536 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_255
timestamp 1698175906
transform 1 0 29904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_259
timestamp 1698175906
transform 1 0 30352 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_275
timestamp 1698175906
transform 1 0 32144 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698175906
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_298
timestamp 1698175906
transform 1 0 34720 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_306
timestamp 1698175906
transform 1 0 35616 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_312
timestamp 1698175906
transform 1 0 36288 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_328
timestamp 1698175906
transform 1 0 38080 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_330
timestamp 1698175906
transform 1 0 38304 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_333
timestamp 1698175906
transform 1 0 38640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_352
timestamp 1698175906
transform 1 0 40768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_356
timestamp 1698175906
transform 1 0 41216 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_360
timestamp 1698175906
transform 1 0 41664 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_368
timestamp 1698175906
transform 1 0 42560 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_372
timestamp 1698175906
transform 1 0 43008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_405
timestamp 1698175906
transform 1 0 46704 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_413
timestamp 1698175906
transform 1 0 47600 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_416
timestamp 1698175906
transform 1 0 47936 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_422
timestamp 1698175906
transform 1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_424
timestamp 1698175906
transform 1 0 48832 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_478
timestamp 1698175906
transform 1 0 54880 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_482
timestamp 1698175906
transform 1 0 55328 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_486
timestamp 1698175906
transform 1 0 55776 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_507
timestamp 1698175906
transform 1 0 58128 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_515
timestamp 1698175906
transform 1 0 59024 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_519
timestamp 1698175906
transform 1 0 59472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_523
timestamp 1698175906
transform 1 0 59920 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_527
timestamp 1698175906
transform 1 0 60368 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_531
timestamp 1698175906
transform 1 0 60816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_562
timestamp 1698175906
transform 1 0 64288 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_568
timestamp 1698175906
transform 1 0 64960 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_600
timestamp 1698175906
transform 1 0 68544 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_616
timestamp 1698175906
transform 1 0 70336 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_624
timestamp 1698175906
transform 1 0 71232 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_628
timestamp 1698175906
transform 1 0 71680 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_632
timestamp 1698175906
transform 1 0 72128 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_696
timestamp 1698175906
transform 1 0 79296 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_702
timestamp 1698175906
transform 1 0 79968 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_766
timestamp 1698175906
transform 1 0 87136 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_772
timestamp 1698175906
transform 1 0 87808 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_836
timestamp 1698175906
transform 1 0 94976 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_842
timestamp 1698175906
transform 1 0 95648 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_858
timestamp 1698175906
transform 1 0 97440 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_8
timestamp 1698175906
transform 1 0 2240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_12
timestamp 1698175906
transform 1 0 2688 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_28
timestamp 1698175906
transform 1 0 4480 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_32
timestamp 1698175906
transform 1 0 4928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_53
timestamp 1698175906
transform 1 0 7280 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_61
timestamp 1698175906
transform 1 0 8176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_69
timestamp 1698175906
transform 1 0 9072 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_115
timestamp 1698175906
transform 1 0 14224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_117
timestamp 1698175906
transform 1 0 14448 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_135
timestamp 1698175906
transform 1 0 16464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_139
timestamp 1698175906
transform 1 0 16912 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_155
timestamp 1698175906
transform 1 0 18704 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_157
timestamp 1698175906
transform 1 0 18928 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_183
timestamp 1698175906
transform 1 0 21840 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_215
timestamp 1698175906
transform 1 0 25424 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_231
timestamp 1698175906
transform 1 0 27216 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_239
timestamp 1698175906
transform 1 0 28112 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_243
timestamp 1698175906
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_263
timestamp 1698175906
transform 1 0 30800 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_271
timestamp 1698175906
transform 1 0 31696 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_275
timestamp 1698175906
transform 1 0 32144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_277
timestamp 1698175906
transform 1 0 32368 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_280
timestamp 1698175906
transform 1 0 32704 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_312
timestamp 1698175906
transform 1 0 36288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698175906
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_325
timestamp 1698175906
transform 1 0 37744 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_329
timestamp 1698175906
transform 1 0 38192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_367
timestamp 1698175906
transform 1 0 42448 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_375
timestamp 1698175906
transform 1 0 43344 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_387
timestamp 1698175906
transform 1 0 44688 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_396
timestamp 1698175906
transform 1 0 45696 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_400
timestamp 1698175906
transform 1 0 46144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_441
timestamp 1698175906
transform 1 0 50736 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_449
timestamp 1698175906
transform 1 0 51632 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_453
timestamp 1698175906
transform 1 0 52080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_457
timestamp 1698175906
transform 1 0 52528 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_461
timestamp 1698175906
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_465
timestamp 1698175906
transform 1 0 53424 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_481
timestamp 1698175906
transform 1 0 55216 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_489
timestamp 1698175906
transform 1 0 56112 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_493
timestamp 1698175906
transform 1 0 56560 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_527
timestamp 1698175906
transform 1 0 60368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_533
timestamp 1698175906
transform 1 0 61040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_584
timestamp 1698175906
transform 1 0 66752 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_588
timestamp 1698175906
transform 1 0 67200 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_592
timestamp 1698175906
transform 1 0 67648 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_594
timestamp 1698175906
transform 1 0 67872 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_597
timestamp 1698175906
transform 1 0 68208 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_661
timestamp 1698175906
transform 1 0 75376 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_667
timestamp 1698175906
transform 1 0 76048 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_731
timestamp 1698175906
transform 1 0 83216 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_737
timestamp 1698175906
transform 1 0 83888 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_801
timestamp 1698175906
transform 1 0 91056 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_807
timestamp 1698175906
transform 1 0 91728 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_839
timestamp 1698175906
transform 1 0 95312 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_855
timestamp 1698175906
transform 1 0 97104 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_863
timestamp 1698175906
transform 1 0 98000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_865
timestamp 1698175906
transform 1 0 98224 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_36
timestamp 1698175906
transform 1 0 5376 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_40
timestamp 1698175906
transform 1 0 5824 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_56
timestamp 1698175906
transform 1 0 7616 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_64
timestamp 1698175906
transform 1 0 8512 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_68
timestamp 1698175906
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_80
timestamp 1698175906
transform 1 0 10304 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_84
timestamp 1698175906
transform 1 0 10752 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_86
timestamp 1698175906
transform 1 0 10976 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_121
timestamp 1698175906
transform 1 0 14896 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_137
timestamp 1698175906
transform 1 0 16688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698175906
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_158
timestamp 1698175906
transform 1 0 19040 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_166
timestamp 1698175906
transform 1 0 19936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_170
timestamp 1698175906
transform 1 0 20384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_172
timestamp 1698175906
transform 1 0 20608 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_177
timestamp 1698175906
transform 1 0 21168 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_209
timestamp 1698175906
transform 1 0 24752 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_266
timestamp 1698175906
transform 1 0 31136 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_270
timestamp 1698175906
transform 1 0 31584 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_322
timestamp 1698175906
transform 1 0 37408 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_326
timestamp 1698175906
transform 1 0 37856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_328
timestamp 1698175906
transform 1 0 38080 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_331
timestamp 1698175906
transform 1 0 38416 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_349
timestamp 1698175906
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_352
timestamp 1698175906
transform 1 0 40768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_356
timestamp 1698175906
transform 1 0 41216 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_360
timestamp 1698175906
transform 1 0 41664 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_376
timestamp 1698175906
transform 1 0 43456 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_384
timestamp 1698175906
transform 1 0 44352 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_387
timestamp 1698175906
transform 1 0 44688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_391
timestamp 1698175906
transform 1 0 45136 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_418
timestamp 1698175906
transform 1 0 48160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_436
timestamp 1698175906
transform 1 0 50176 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_440
timestamp 1698175906
transform 1 0 50624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_442
timestamp 1698175906
transform 1 0 50848 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_462
timestamp 1698175906
transform 1 0 53088 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_478
timestamp 1698175906
transform 1 0 54880 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_492
timestamp 1698175906
transform 1 0 56448 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_508
timestamp 1698175906
transform 1 0 58240 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_524
timestamp 1698175906
transform 1 0 60032 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_532
timestamp 1698175906
transform 1 0 60928 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_535
timestamp 1698175906
transform 1 0 61264 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_539
timestamp 1698175906
transform 1 0 61712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_570
timestamp 1698175906
transform 1 0 65184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_574
timestamp 1698175906
transform 1 0 65632 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_606
timestamp 1698175906
transform 1 0 69216 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_622
timestamp 1698175906
transform 1 0 71008 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_632
timestamp 1698175906
transform 1 0 72128 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_644
timestamp 1698175906
transform 1 0 73472 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_648
timestamp 1698175906
transform 1 0 73920 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_650
timestamp 1698175906
transform 1 0 74144 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_656
timestamp 1698175906
transform 1 0 74816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_660
timestamp 1698175906
transform 1 0 75264 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_664
timestamp 1698175906
transform 1 0 75712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_666
timestamp 1698175906
transform 1 0 75936 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_673
timestamp 1698175906
transform 1 0 76720 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_689
timestamp 1698175906
transform 1 0 78512 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_697
timestamp 1698175906
transform 1 0 79408 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_699
timestamp 1698175906
transform 1 0 79632 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_702
timestamp 1698175906
transform 1 0 79968 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_734
timestamp 1698175906
transform 1 0 83552 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_757
timestamp 1698175906
transform 1 0 86128 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_765
timestamp 1698175906
transform 1 0 87024 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_769
timestamp 1698175906
transform 1 0 87472 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_772
timestamp 1698175906
transform 1 0 87808 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_836
timestamp 1698175906
transform 1 0 94976 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_842
timestamp 1698175906
transform 1 0 95648 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_862
timestamp 1698175906
transform 1 0 97888 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_12
timestamp 1698175906
transform 1 0 2688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_16
timestamp 1698175906
transform 1 0 3136 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_24
timestamp 1698175906
transform 1 0 4032 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_28
timestamp 1698175906
transform 1 0 4480 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_30
timestamp 1698175906
transform 1 0 4704 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_71
timestamp 1698175906
transform 1 0 9296 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_87
timestamp 1698175906
transform 1 0 11088 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_92
timestamp 1698175906
transform 1 0 11648 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_100
timestamp 1698175906
transform 1 0 12544 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698175906
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_211
timestamp 1698175906
transform 1 0 24976 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_219
timestamp 1698175906
transform 1 0 25872 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_225
timestamp 1698175906
transform 1 0 26544 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_229
timestamp 1698175906
transform 1 0 26992 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_231
timestamp 1698175906
transform 1 0 27216 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_236
timestamp 1698175906
transform 1 0 27776 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698175906
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_279
timestamp 1698175906
transform 1 0 32592 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_295
timestamp 1698175906
transform 1 0 34384 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_310
timestamp 1698175906
transform 1 0 36064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_312
timestamp 1698175906
transform 1 0 36288 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_354
timestamp 1698175906
transform 1 0 40992 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_358
timestamp 1698175906
transform 1 0 41440 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_366
timestamp 1698175906
transform 1 0 42336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_370
timestamp 1698175906
transform 1 0 42784 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_387
timestamp 1698175906
transform 1 0 44688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_446
timestamp 1698175906
transform 1 0 51296 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_450
timestamp 1698175906
transform 1 0 51744 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_452
timestamp 1698175906
transform 1 0 51968 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_464
timestamp 1698175906
transform 1 0 53312 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_472
timestamp 1698175906
transform 1 0 54208 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_474
timestamp 1698175906
transform 1 0 54432 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_515
timestamp 1698175906
transform 1 0 59024 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_523
timestamp 1698175906
transform 1 0 59920 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_527
timestamp 1698175906
transform 1 0 60368 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_535
timestamp 1698175906
transform 1 0 61264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_537
timestamp 1698175906
transform 1 0 61488 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_590
timestamp 1698175906
transform 1 0 67424 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_592
timestamp 1698175906
transform 1 0 67648 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_667
timestamp 1698175906
transform 1 0 76048 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_671
timestamp 1698175906
transform 1 0 76496 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_679
timestamp 1698175906
transform 1 0 77392 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_717
timestamp 1698175906
transform 1 0 81648 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_733
timestamp 1698175906
transform 1 0 83440 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_737
timestamp 1698175906
transform 1 0 83888 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_739
timestamp 1698175906
transform 1 0 84112 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_776
timestamp 1698175906
transform 1 0 88256 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_784
timestamp 1698175906
transform 1 0 89152 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_788
timestamp 1698175906
transform 1 0 89600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_792
timestamp 1698175906
transform 1 0 90048 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_800
timestamp 1698175906
transform 1 0 90944 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_804
timestamp 1698175906
transform 1 0 91392 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_807
timestamp 1698175906
transform 1 0 91728 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_839
timestamp 1698175906
transform 1 0 95312 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_843
timestamp 1698175906
transform 1 0 95760 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_845
timestamp 1698175906
transform 1 0 95984 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_852
timestamp 1698175906
transform 1 0 96768 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_860
timestamp 1698175906
transform 1 0 97664 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_864
timestamp 1698175906
transform 1 0 98112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_8
timestamp 1698175906
transform 1 0 2240 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_44
timestamp 1698175906
transform 1 0 6272 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_48
timestamp 1698175906
transform 1 0 6720 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_64
timestamp 1698175906
transform 1 0 8512 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_68
timestamp 1698175906
transform 1 0 8960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_104
timestamp 1698175906
transform 1 0 12992 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_120
timestamp 1698175906
transform 1 0 14784 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_138
timestamp 1698175906
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_146
timestamp 1698175906
transform 1 0 17696 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_156
timestamp 1698175906
transform 1 0 18816 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_187
timestamp 1698175906
transform 1 0 22288 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_203
timestamp 1698175906
transform 1 0 24080 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_207
timestamp 1698175906
transform 1 0 24528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_209
timestamp 1698175906
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_298
timestamp 1698175906
transform 1 0 34720 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_306
timestamp 1698175906
transform 1 0 35616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_310
timestamp 1698175906
transform 1 0 36064 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_313
timestamp 1698175906
transform 1 0 36400 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_319
timestamp 1698175906
transform 1 0 37072 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_323
timestamp 1698175906
transform 1 0 37520 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_331
timestamp 1698175906
transform 1 0 38416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_344
timestamp 1698175906
transform 1 0 39872 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_352
timestamp 1698175906
transform 1 0 40768 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_384
timestamp 1698175906
transform 1 0 44352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_388
timestamp 1698175906
transform 1 0 44800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_392
timestamp 1698175906
transform 1 0 45248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_396
timestamp 1698175906
transform 1 0 45696 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_422
timestamp 1698175906
transform 1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_438
timestamp 1698175906
transform 1 0 50400 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_454
timestamp 1698175906
transform 1 0 52192 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_458
timestamp 1698175906
transform 1 0 52640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_460
timestamp 1698175906
transform 1 0 52864 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_472
timestamp 1698175906
transform 1 0 54208 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_492
timestamp 1698175906
transform 1 0 56448 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_496
timestamp 1698175906
transform 1 0 56896 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_506
timestamp 1698175906
transform 1 0 58016 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_538
timestamp 1698175906
transform 1 0 61600 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_552
timestamp 1698175906
transform 1 0 63168 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_562
timestamp 1698175906
transform 1 0 64288 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_604
timestamp 1698175906
transform 1 0 68992 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_620
timestamp 1698175906
transform 1 0 70784 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_628
timestamp 1698175906
transform 1 0 71680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_632
timestamp 1698175906
transform 1 0 72128 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_637
timestamp 1698175906
transform 1 0 72688 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_669
timestamp 1698175906
transform 1 0 76272 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_677
timestamp 1698175906
transform 1 0 77168 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_681
timestamp 1698175906
transform 1 0 77616 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_697
timestamp 1698175906
transform 1 0 79408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_699
timestamp 1698175906
transform 1 0 79632 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_707
timestamp 1698175906
transform 1 0 80528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_711
timestamp 1698175906
transform 1 0 80976 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_727
timestamp 1698175906
transform 1 0 82768 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_735
timestamp 1698175906
transform 1 0 83664 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_739
timestamp 1698175906
transform 1 0 84112 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_754
timestamp 1698175906
transform 1 0 85792 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_758
timestamp 1698175906
transform 1 0 86240 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_766
timestamp 1698175906
transform 1 0 87136 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_772
timestamp 1698175906
transform 1 0 87808 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_780
timestamp 1698175906
transform 1 0 88704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_826
timestamp 1698175906
transform 1 0 93856 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_834
timestamp 1698175906
transform 1 0 94752 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_838
timestamp 1698175906
transform 1 0 95200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_842
timestamp 1698175906
transform 1 0 95648 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_850
timestamp 1698175906
transform 1 0 96544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_862
timestamp 1698175906
transform 1 0 97888 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_8
timestamp 1698175906
transform 1 0 2240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_10
timestamp 1698175906
transform 1 0 2464 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_15
timestamp 1698175906
transform 1 0 3024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_19
timestamp 1698175906
transform 1 0 3472 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_51
timestamp 1698175906
transform 1 0 7056 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_55
timestamp 1698175906
transform 1 0 7504 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_99
timestamp 1698175906
transform 1 0 12432 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_103
timestamp 1698175906
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_115
timestamp 1698175906
transform 1 0 14224 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_168
timestamp 1698175906
transform 1 0 20160 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_172
timestamp 1698175906
transform 1 0 20608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698175906
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_181
timestamp 1698175906
transform 1 0 21616 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_213
timestamp 1698175906
transform 1 0 25200 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_235
timestamp 1698175906
transform 1 0 27664 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1698175906
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_251
timestamp 1698175906
transform 1 0 29456 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_253
timestamp 1698175906
transform 1 0 29680 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_256
timestamp 1698175906
transform 1 0 30016 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_264
timestamp 1698175906
transform 1 0 30912 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_302
timestamp 1698175906
transform 1 0 35168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_310
timestamp 1698175906
transform 1 0 36064 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_314
timestamp 1698175906
transform 1 0 36512 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_322
timestamp 1698175906
transform 1 0 37408 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_326
timestamp 1698175906
transform 1 0 37856 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_334
timestamp 1698175906
transform 1 0 38752 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_337
timestamp 1698175906
transform 1 0 39088 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_369
timestamp 1698175906
transform 1 0 42672 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_387
timestamp 1698175906
transform 1 0 44688 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_395
timestamp 1698175906
transform 1 0 45584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_397
timestamp 1698175906
transform 1 0 45808 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_400
timestamp 1698175906
transform 1 0 46144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_410
timestamp 1698175906
transform 1 0 47264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_422
timestamp 1698175906
transform 1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_426
timestamp 1698175906
transform 1 0 49056 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_444
timestamp 1698175906
transform 1 0 51072 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_450
timestamp 1698175906
transform 1 0 51744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_454
timestamp 1698175906
transform 1 0 52192 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_457
timestamp 1698175906
transform 1 0 52528 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_467
timestamp 1698175906
transform 1 0 53648 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_471
timestamp 1698175906
transform 1 0 54096 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_487
timestamp 1698175906
transform 1 0 55888 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_497
timestamp 1698175906
transform 1 0 57008 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_513
timestamp 1698175906
transform 1 0 58800 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_521
timestamp 1698175906
transform 1 0 59696 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_527
timestamp 1698175906
transform 1 0 60368 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_559
timestamp 1698175906
transform 1 0 63952 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_563
timestamp 1698175906
transform 1 0 64400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_565
timestamp 1698175906
transform 1 0 64624 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_568
timestamp 1698175906
transform 1 0 64960 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_584
timestamp 1698175906
transform 1 0 66752 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_588
timestamp 1698175906
transform 1 0 67200 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_591
timestamp 1698175906
transform 1 0 67536 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_612
timestamp 1698175906
transform 1 0 69888 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_644
timestamp 1698175906
transform 1 0 73472 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_660
timestamp 1698175906
transform 1 0 75264 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_664
timestamp 1698175906
transform 1 0 75712 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_667
timestamp 1698175906
transform 1 0 76048 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_675
timestamp 1698175906
transform 1 0 76944 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_678
timestamp 1698175906
transform 1 0 77280 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_686
timestamp 1698175906
transform 1 0 78176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_690
timestamp 1698175906
transform 1 0 78624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_692
timestamp 1698175906
transform 1 0 78848 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_695
timestamp 1698175906
transform 1 0 79184 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_727
timestamp 1698175906
transform 1 0 82768 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_737
timestamp 1698175906
transform 1 0 83888 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_769
timestamp 1698175906
transform 1 0 87472 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_785
timestamp 1698175906
transform 1 0 89264 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_793
timestamp 1698175906
transform 1 0 90160 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_801
timestamp 1698175906
transform 1 0 91056 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_815
timestamp 1698175906
transform 1 0 92624 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_831
timestamp 1698175906
transform 1 0 94416 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_839
timestamp 1698175906
transform 1 0 95312 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_843
timestamp 1698175906
transform 1 0 95760 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_845
timestamp 1698175906
transform 1 0 95984 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_852
timestamp 1698175906
transform 1 0 96768 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_860
timestamp 1698175906
transform 1 0 97664 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_864
timestamp 1698175906
transform 1 0 98112 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_6
timestamp 1698175906
transform 1 0 2016 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_49
timestamp 1698175906
transform 1 0 6832 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_53
timestamp 1698175906
transform 1 0 7280 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_57
timestamp 1698175906
transform 1 0 7728 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_59
timestamp 1698175906
transform 1 0 7952 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_87
timestamp 1698175906
transform 1 0 11088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_91
timestamp 1698175906
transform 1 0 11536 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_95
timestamp 1698175906
transform 1 0 11984 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_111
timestamp 1698175906
transform 1 0 13776 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_119
timestamp 1698175906
transform 1 0 14672 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_129
timestamp 1698175906
transform 1 0 15792 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_137
timestamp 1698175906
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698175906
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_150
timestamp 1698175906
transform 1 0 18144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_154
timestamp 1698175906
transform 1 0 18592 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_162
timestamp 1698175906
transform 1 0 19488 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_165
timestamp 1698175906
transform 1 0 19824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_184
timestamp 1698175906
transform 1 0 21952 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_200
timestamp 1698175906
transform 1 0 23744 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698175906
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_268
timestamp 1698175906
transform 1 0 31360 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_274
timestamp 1698175906
transform 1 0 32032 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_335
timestamp 1698175906
transform 1 0 38864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_345
timestamp 1698175906
transform 1 0 39984 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_347
timestamp 1698175906
transform 1 0 40208 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_367
timestamp 1698175906
transform 1 0 42448 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_371
timestamp 1698175906
transform 1 0 42896 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_373
timestamp 1698175906
transform 1 0 43120 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_410
timestamp 1698175906
transform 1 0 47264 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_418
timestamp 1698175906
transform 1 0 48160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_422
timestamp 1698175906
transform 1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_424
timestamp 1698175906
transform 1 0 48832 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_427
timestamp 1698175906
transform 1 0 49168 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_442
timestamp 1698175906
transform 1 0 50848 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_444
timestamp 1698175906
transform 1 0 51072 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_480
timestamp 1698175906
transform 1 0 55104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_484
timestamp 1698175906
transform 1 0 55552 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_488
timestamp 1698175906
transform 1 0 56000 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_492
timestamp 1698175906
transform 1 0 56448 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_500
timestamp 1698175906
transform 1 0 57344 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_540
timestamp 1698175906
transform 1 0 61824 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_556
timestamp 1698175906
transform 1 0 63616 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_583
timestamp 1698175906
transform 1 0 66640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_587
timestamp 1698175906
transform 1 0 67088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_591
timestamp 1698175906
transform 1 0 67536 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_595
timestamp 1698175906
transform 1 0 67984 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_599
timestamp 1698175906
transform 1 0 68432 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_615
timestamp 1698175906
transform 1 0 70224 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_623
timestamp 1698175906
transform 1 0 71120 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_627
timestamp 1698175906
transform 1 0 71568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_629
timestamp 1698175906
transform 1 0 71792 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_666
timestamp 1698175906
transform 1 0 75936 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_670
timestamp 1698175906
transform 1 0 76384 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_676
timestamp 1698175906
transform 1 0 77056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_693
timestamp 1698175906
transform 1 0 78960 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_697
timestamp 1698175906
transform 1 0 79408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_699
timestamp 1698175906
transform 1 0 79632 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_702
timestamp 1698175906
transform 1 0 79968 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_734
timestamp 1698175906
transform 1 0 83552 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_772
timestamp 1698175906
transform 1 0 87808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_776
timestamp 1698175906
transform 1 0 88256 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_792
timestamp 1698175906
transform 1 0 90048 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_798
timestamp 1698175906
transform 1 0 90720 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_830
timestamp 1698175906
transform 1 0 94304 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_838
timestamp 1698175906
transform 1 0 95200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_842
timestamp 1698175906
transform 1 0 95648 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_844
timestamp 1698175906
transform 1 0 95872 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_851
timestamp 1698175906
transform 1 0 96656 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_8
timestamp 1698175906
transform 1 0 2240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_12
timestamp 1698175906
transform 1 0 2688 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_28
timestamp 1698175906
transform 1 0 4480 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_32
timestamp 1698175906
transform 1 0 4928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_37
timestamp 1698175906
transform 1 0 5488 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_43
timestamp 1698175906
transform 1 0 6160 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_75
timestamp 1698175906
transform 1 0 9744 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_91
timestamp 1698175906
transform 1 0 11536 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_99
timestamp 1698175906
transform 1 0 12432 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_103
timestamp 1698175906
transform 1 0 12880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_107
timestamp 1698175906
transform 1 0 13328 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_139
timestamp 1698175906
transform 1 0 16912 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_155
timestamp 1698175906
transform 1 0 18704 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_163
timestamp 1698175906
transform 1 0 19600 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_167
timestamp 1698175906
transform 1 0 20048 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_177
timestamp 1698175906
transform 1 0 21168 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_212
timestamp 1698175906
transform 1 0 25088 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_220
timestamp 1698175906
transform 1 0 25984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_226
timestamp 1698175906
transform 1 0 26656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_247
timestamp 1698175906
transform 1 0 29008 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_251
timestamp 1698175906
transform 1 0 29456 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_254
timestamp 1698175906
transform 1 0 29792 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_258
timestamp 1698175906
transform 1 0 30240 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_284
timestamp 1698175906
transform 1 0 33152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_288
timestamp 1698175906
transform 1 0 33600 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_304
timestamp 1698175906
transform 1 0 35392 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_312
timestamp 1698175906
transform 1 0 36288 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_314
timestamp 1698175906
transform 1 0 36512 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_322
timestamp 1698175906
transform 1 0 37408 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_378
timestamp 1698175906
transform 1 0 43680 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_402
timestamp 1698175906
transform 1 0 46368 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_406
timestamp 1698175906
transform 1 0 46816 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_414
timestamp 1698175906
transform 1 0 47712 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_416
timestamp 1698175906
transform 1 0 47936 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_449
timestamp 1698175906
transform 1 0 51632 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_453
timestamp 1698175906
transform 1 0 52080 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_457
timestamp 1698175906
transform 1 0 52528 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_492
timestamp 1698175906
transform 1 0 56448 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_496
timestamp 1698175906
transform 1 0 56896 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_512
timestamp 1698175906
transform 1 0 58688 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_519
timestamp 1698175906
transform 1 0 59472 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_542
timestamp 1698175906
transform 1 0 62048 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_546
timestamp 1698175906
transform 1 0 62496 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_548
timestamp 1698175906
transform 1 0 62720 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_606
timestamp 1698175906
transform 1 0 69216 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_622
timestamp 1698175906
transform 1 0 71008 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_626
timestamp 1698175906
transform 1 0 71456 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_632
timestamp 1698175906
transform 1 0 72128 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_654
timestamp 1698175906
transform 1 0 74592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_656
timestamp 1698175906
transform 1 0 74816 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_659
timestamp 1698175906
transform 1 0 75152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_663
timestamp 1698175906
transform 1 0 75600 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_683
timestamp 1698175906
transform 1 0 77840 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_725
timestamp 1698175906
transform 1 0 82544 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_737
timestamp 1698175906
transform 1 0 83888 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_747
timestamp 1698175906
transform 1 0 85008 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_753
timestamp 1698175906
transform 1 0 85680 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_757
timestamp 1698175906
transform 1 0 86128 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_765
timestamp 1698175906
transform 1 0 87024 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_782
timestamp 1698175906
transform 1 0 88928 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_798
timestamp 1698175906
transform 1 0 90720 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_802
timestamp 1698175906
transform 1 0 91168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_804
timestamp 1698175906
transform 1 0 91392 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_807
timestamp 1698175906
transform 1 0 91728 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_839
timestamp 1698175906
transform 1 0 95312 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_843
timestamp 1698175906
transform 1 0 95760 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_845
timestamp 1698175906
transform 1 0 95984 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_852
timestamp 1698175906
transform 1 0 96768 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_860
timestamp 1698175906
transform 1 0 97664 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_864
timestamp 1698175906
transform 1 0 98112 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_2
timestamp 1698175906
transform 1 0 1568 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_6
timestamp 1698175906
transform 1 0 2016 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_12
timestamp 1698175906
transform 1 0 2688 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_44
timestamp 1698175906
transform 1 0 6272 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_60
timestamp 1698175906
transform 1 0 8064 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_68
timestamp 1698175906
transform 1 0 8960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_72
timestamp 1698175906
transform 1 0 9408 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_104
timestamp 1698175906
transform 1 0 12992 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_139
timestamp 1698175906
transform 1 0 16912 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_142
timestamp 1698175906
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_146
timestamp 1698175906
transform 1 0 17696 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_162
timestamp 1698175906
transform 1 0 19488 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_170
timestamp 1698175906
transform 1 0 20384 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_174
timestamp 1698175906
transform 1 0 20832 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_178
timestamp 1698175906
transform 1 0 21280 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_184
timestamp 1698175906
transform 1 0 21952 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_200
timestamp 1698175906
transform 1 0 23744 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_208
timestamp 1698175906
transform 1 0 24640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_212
timestamp 1698175906
transform 1 0 25088 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_244
timestamp 1698175906
transform 1 0 28672 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_247
timestamp 1698175906
transform 1 0 29008 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_279
timestamp 1698175906
transform 1 0 32592 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_282
timestamp 1698175906
transform 1 0 32928 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_314
timestamp 1698175906
transform 1 0 36512 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_330
timestamp 1698175906
transform 1 0 38304 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_335
timestamp 1698175906
transform 1 0 38864 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_343
timestamp 1698175906
transform 1 0 39760 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_347
timestamp 1698175906
transform 1 0 40208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_349
timestamp 1698175906
transform 1 0 40432 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_352
timestamp 1698175906
transform 1 0 40768 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_360
timestamp 1698175906
transform 1 0 41664 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_366
timestamp 1698175906
transform 1 0 42336 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_370
timestamp 1698175906
transform 1 0 42784 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_382
timestamp 1698175906
transform 1 0 44128 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_384
timestamp 1698175906
transform 1 0 44352 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_387
timestamp 1698175906
transform 1 0 44688 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_403
timestamp 1698175906
transform 1 0 46480 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_411
timestamp 1698175906
transform 1 0 47376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_454
timestamp 1698175906
transform 1 0 52192 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_458
timestamp 1698175906
transform 1 0 52640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_472
timestamp 1698175906
transform 1 0 54208 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_488
timestamp 1698175906
transform 1 0 56000 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_492
timestamp 1698175906
transform 1 0 56448 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_512
timestamp 1698175906
transform 1 0 58688 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_520
timestamp 1698175906
transform 1 0 59584 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_524
timestamp 1698175906
transform 1 0 60032 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_527
timestamp 1698175906
transform 1 0 60368 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_559
timestamp 1698175906
transform 1 0 63952 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_562
timestamp 1698175906
transform 1 0 64288 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_578
timestamp 1698175906
transform 1 0 66080 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_582
timestamp 1698175906
transform 1 0 66528 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_585
timestamp 1698175906
transform 1 0 66864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_589
timestamp 1698175906
transform 1 0 67312 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_591
timestamp 1698175906
transform 1 0 67536 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_608
timestamp 1698175906
transform 1 0 69440 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_624
timestamp 1698175906
transform 1 0 71232 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_628
timestamp 1698175906
transform 1 0 71680 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_632
timestamp 1698175906
transform 1 0 72128 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_634
timestamp 1698175906
transform 1 0 72352 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_637
timestamp 1698175906
transform 1 0 72688 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_641
timestamp 1698175906
transform 1 0 73136 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_649
timestamp 1698175906
transform 1 0 74032 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_653
timestamp 1698175906
transform 1 0 74480 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_668
timestamp 1698175906
transform 1 0 76160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_672
timestamp 1698175906
transform 1 0 76608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_681
timestamp 1698175906
transform 1 0 77616 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_685
timestamp 1698175906
transform 1 0 78064 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_691
timestamp 1698175906
transform 1 0 78736 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_696
timestamp 1698175906
transform 1 0 79296 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_702
timestamp 1698175906
transform 1 0 79968 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_734
timestamp 1698175906
transform 1 0 83552 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_737
timestamp 1698175906
transform 1 0 83888 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_739
timestamp 1698175906
transform 1 0 84112 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_742
timestamp 1698175906
transform 1 0 84448 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_747
timestamp 1698175906
transform 1 0 85008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_751
timestamp 1698175906
transform 1 0 85456 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_755
timestamp 1698175906
transform 1 0 85904 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_763
timestamp 1698175906
transform 1 0 86800 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_767
timestamp 1698175906
transform 1 0 87248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_769
timestamp 1698175906
transform 1 0 87472 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_772
timestamp 1698175906
transform 1 0 87808 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_788
timestamp 1698175906
transform 1 0 89600 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_791
timestamp 1698175906
transform 1 0 89936 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_795
timestamp 1698175906
transform 1 0 90384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_812
timestamp 1698175906
transform 1 0 92288 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_828
timestamp 1698175906
transform 1 0 94080 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_836
timestamp 1698175906
transform 1 0 94976 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_842
timestamp 1698175906
transform 1 0 95648 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_858
timestamp 1698175906
transform 1 0 97440 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_12
timestamp 1698175906
transform 1 0 2688 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_28
timestamp 1698175906
transform 1 0 4480 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_32
timestamp 1698175906
transform 1 0 4928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698175906
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_41
timestamp 1698175906
transform 1 0 5936 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_57
timestamp 1698175906
transform 1 0 7728 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_65
timestamp 1698175906
transform 1 0 8624 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_69
timestamp 1698175906
transform 1 0 9072 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_72
timestamp 1698175906
transform 1 0 9408 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_117
timestamp 1698175906
transform 1 0 14448 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_149
timestamp 1698175906
transform 1 0 18032 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_156
timestamp 1698175906
transform 1 0 18816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_158
timestamp 1698175906
transform 1 0 19040 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_163
timestamp 1698175906
transform 1 0 19600 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698175906
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_177
timestamp 1698175906
transform 1 0 21168 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_209
timestamp 1698175906
transform 1 0 24752 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_217
timestamp 1698175906
transform 1 0 25648 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_221
timestamp 1698175906
transform 1 0 26096 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_223
timestamp 1698175906
transform 1 0 26320 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_230
timestamp 1698175906
transform 1 0 27104 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_238
timestamp 1698175906
transform 1 0 28000 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_242
timestamp 1698175906
transform 1 0 28448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698175906
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_247
timestamp 1698175906
transform 1 0 29008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_251
timestamp 1698175906
transform 1 0 29456 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_259
timestamp 1698175906
transform 1 0 30352 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_263
timestamp 1698175906
transform 1 0 30800 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_300
timestamp 1698175906
transform 1 0 34944 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_322
timestamp 1698175906
transform 1 0 37408 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_326
timestamp 1698175906
transform 1 0 37856 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_358
timestamp 1698175906
transform 1 0 41440 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_374
timestamp 1698175906
transform 1 0 43232 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_382
timestamp 1698175906
transform 1 0 44128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698175906
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_387
timestamp 1698175906
transform 1 0 44688 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_419
timestamp 1698175906
transform 1 0 48272 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_422
timestamp 1698175906
transform 1 0 48608 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_454
timestamp 1698175906
transform 1 0 52192 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_457
timestamp 1698175906
transform 1 0 52528 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_461
timestamp 1698175906
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_465
timestamp 1698175906
transform 1 0 53424 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_469
timestamp 1698175906
transform 1 0 53872 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_501
timestamp 1698175906
transform 1 0 57456 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_517
timestamp 1698175906
transform 1 0 59248 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_527
timestamp 1698175906
transform 1 0 60368 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_559
timestamp 1698175906
transform 1 0 63952 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_575
timestamp 1698175906
transform 1 0 65744 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_577
timestamp 1698175906
transform 1 0 65968 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_580
timestamp 1698175906
transform 1 0 66304 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_590
timestamp 1698175906
transform 1 0 67424 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_594
timestamp 1698175906
transform 1 0 67872 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_602
timestamp 1698175906
transform 1 0 68768 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_606
timestamp 1698175906
transform 1 0 69216 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_622
timestamp 1698175906
transform 1 0 71008 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_630
timestamp 1698175906
transform 1 0 71904 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_634
timestamp 1698175906
transform 1 0 72352 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_636
timestamp 1698175906
transform 1 0 72576 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_639
timestamp 1698175906
transform 1 0 72912 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_655
timestamp 1698175906
transform 1 0 74704 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_663
timestamp 1698175906
transform 1 0 75600 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_667
timestamp 1698175906
transform 1 0 76048 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_699
timestamp 1698175906
transform 1 0 79632 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_715
timestamp 1698175906
transform 1 0 81424 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_719
timestamp 1698175906
transform 1 0 81872 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_731
timestamp 1698175906
transform 1 0 83216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_742
timestamp 1698175906
transform 1 0 84448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_795
timestamp 1698175906
transform 1 0 90384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_799
timestamp 1698175906
transform 1 0 90832 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_803
timestamp 1698175906
transform 1 0 91280 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_807
timestamp 1698175906
transform 1 0 91728 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_813
timestamp 1698175906
transform 1 0 92400 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_845
timestamp 1698175906
transform 1 0 95984 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_849
timestamp 1698175906
transform 1 0 96432 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_851
timestamp 1698175906
transform 1 0 96656 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_106
timestamp 1698175906
transform 1 0 13216 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_110
timestamp 1698175906
transform 1 0 13664 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_126
timestamp 1698175906
transform 1 0 15456 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_134
timestamp 1698175906
transform 1 0 16352 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_191
timestamp 1698175906
transform 1 0 22736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_195
timestamp 1698175906
transform 1 0 23184 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_203
timestamp 1698175906
transform 1 0 24080 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_207
timestamp 1698175906
transform 1 0 24528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698175906
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_212
timestamp 1698175906
transform 1 0 25088 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_262
timestamp 1698175906
transform 1 0 30688 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_266
timestamp 1698175906
transform 1 0 31136 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_270
timestamp 1698175906
transform 1 0 31584 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_278
timestamp 1698175906
transform 1 0 32480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_288
timestamp 1698175906
transform 1 0 33600 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_290
timestamp 1698175906
transform 1 0 33824 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_338
timestamp 1698175906
transform 1 0 39200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_342
timestamp 1698175906
transform 1 0 39648 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_346
timestamp 1698175906
transform 1 0 40096 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_367
timestamp 1698175906
transform 1 0 42448 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_371
timestamp 1698175906
transform 1 0 42896 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_379
timestamp 1698175906
transform 1 0 43792 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_383
timestamp 1698175906
transform 1 0 44240 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_401
timestamp 1698175906
transform 1 0 46256 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_405
timestamp 1698175906
transform 1 0 46704 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_413
timestamp 1698175906
transform 1 0 47600 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_417
timestamp 1698175906
transform 1 0 48048 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_419
timestamp 1698175906
transform 1 0 48272 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_422
timestamp 1698175906
transform 1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_426
timestamp 1698175906
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_428
timestamp 1698175906
transform 1 0 49280 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_463
timestamp 1698175906
transform 1 0 53200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_480
timestamp 1698175906
transform 1 0 55104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_484
timestamp 1698175906
transform 1 0 55552 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_488
timestamp 1698175906
transform 1 0 56000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_492
timestamp 1698175906
transform 1 0 56448 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_502
timestamp 1698175906
transform 1 0 57568 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_540
timestamp 1698175906
transform 1 0 61824 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_556
timestamp 1698175906
transform 1 0 63616 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_562
timestamp 1698175906
transform 1 0 64288 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_566
timestamp 1698175906
transform 1 0 64736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_568
timestamp 1698175906
transform 1 0 64960 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_575
timestamp 1698175906
transform 1 0 65744 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_579
timestamp 1698175906
transform 1 0 66192 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_611
timestamp 1698175906
transform 1 0 69776 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_627
timestamp 1698175906
transform 1 0 71568 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_638
timestamp 1698175906
transform 1 0 72800 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_654
timestamp 1698175906
transform 1 0 74592 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_662
timestamp 1698175906
transform 1 0 75488 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_666
timestamp 1698175906
transform 1 0 75936 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_686
timestamp 1698175906
transform 1 0 78176 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_694
timestamp 1698175906
transform 1 0 79072 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_698
timestamp 1698175906
transform 1 0 79520 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_702
timestamp 1698175906
transform 1 0 79968 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_718
timestamp 1698175906
transform 1 0 81760 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_756
timestamp 1698175906
transform 1 0 86016 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_760
timestamp 1698175906
transform 1 0 86464 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_768
timestamp 1698175906
transform 1 0 87360 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_772
timestamp 1698175906
transform 1 0 87808 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_788
timestamp 1698175906
transform 1 0 89600 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_796
timestamp 1698175906
transform 1 0 90496 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_842
timestamp 1698175906
transform 1 0 95648 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_852
timestamp 1698175906
transform 1 0 96768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_860
timestamp 1698175906
transform 1 0 97664 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_864
timestamp 1698175906
transform 1 0 98112 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_14
timestamp 1698175906
transform 1 0 2912 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_18
timestamp 1698175906
transform 1 0 3360 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698175906
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_37
timestamp 1698175906
transform 1 0 5488 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_41
timestamp 1698175906
transform 1 0 5936 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_57
timestamp 1698175906
transform 1 0 7728 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_69
timestamp 1698175906
transform 1 0 9072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_73
timestamp 1698175906
transform 1 0 9520 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_107
timestamp 1698175906
transform 1 0 13328 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_139
timestamp 1698175906
transform 1 0 16912 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_155
timestamp 1698175906
transform 1 0 18704 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_159
timestamp 1698175906
transform 1 0 19152 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_177
timestamp 1698175906
transform 1 0 21168 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_209
timestamp 1698175906
transform 1 0 24752 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_213
timestamp 1698175906
transform 1 0 25200 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_218
timestamp 1698175906
transform 1 0 25760 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_234
timestamp 1698175906
transform 1 0 27552 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_242
timestamp 1698175906
transform 1 0 28448 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_244
timestamp 1698175906
transform 1 0 28672 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_247
timestamp 1698175906
transform 1 0 29008 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_263
timestamp 1698175906
transform 1 0 30800 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_267
timestamp 1698175906
transform 1 0 31248 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_272
timestamp 1698175906
transform 1 0 31808 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_280
timestamp 1698175906
transform 1 0 32704 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_284
timestamp 1698175906
transform 1 0 33152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_287
timestamp 1698175906
transform 1 0 33488 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_306
timestamp 1698175906
transform 1 0 35616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_310
timestamp 1698175906
transform 1 0 36064 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698175906
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_317
timestamp 1698175906
transform 1 0 36848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_325
timestamp 1698175906
transform 1 0 37744 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_329
timestamp 1698175906
transform 1 0 38192 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_364
timestamp 1698175906
transform 1 0 42112 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_368
timestamp 1698175906
transform 1 0 42560 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_376
timestamp 1698175906
transform 1 0 43456 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_378
timestamp 1698175906
transform 1 0 43680 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_437
timestamp 1698175906
transform 1 0 50288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_445
timestamp 1698175906
transform 1 0 51184 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_471
timestamp 1698175906
transform 1 0 54096 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_519
timestamp 1698175906
transform 1 0 59472 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_523
timestamp 1698175906
transform 1 0 59920 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_527
timestamp 1698175906
transform 1 0 60368 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_543
timestamp 1698175906
transform 1 0 62160 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_551
timestamp 1698175906
transform 1 0 63056 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_593
timestamp 1698175906
transform 1 0 67760 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_597
timestamp 1698175906
transform 1 0 68208 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_601
timestamp 1698175906
transform 1 0 68656 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_617
timestamp 1698175906
transform 1 0 70448 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_656
timestamp 1698175906
transform 1 0 74816 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_660
timestamp 1698175906
transform 1 0 75264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_662
timestamp 1698175906
transform 1 0 75488 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_667
timestamp 1698175906
transform 1 0 76048 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_677
timestamp 1698175906
transform 1 0 77168 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_717
timestamp 1698175906
transform 1 0 81648 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_721
timestamp 1698175906
transform 1 0 82096 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_723
timestamp 1698175906
transform 1 0 82320 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_728
timestamp 1698175906
transform 1 0 82880 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_732
timestamp 1698175906
transform 1 0 83328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_734
timestamp 1698175906
transform 1 0 83552 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_737
timestamp 1698175906
transform 1 0 83888 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_741
timestamp 1698175906
transform 1 0 84336 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_744
timestamp 1698175906
transform 1 0 84672 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_760
timestamp 1698175906
transform 1 0 86464 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_768
timestamp 1698175906
transform 1 0 87360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_772
timestamp 1698175906
transform 1 0 87808 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_804
timestamp 1698175906
transform 1 0 91392 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_807
timestamp 1698175906
transform 1 0 91728 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_839
timestamp 1698175906
transform 1 0 95312 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_843
timestamp 1698175906
transform 1 0 95760 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_845
timestamp 1698175906
transform 1 0 95984 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_2
timestamp 1698175906
transform 1 0 1568 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_8
timestamp 1698175906
transform 1 0 2240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_10
timestamp 1698175906
transform 1 0 2464 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_45
timestamp 1698175906
transform 1 0 6384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_49
timestamp 1698175906
transform 1 0 6832 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_65
timestamp 1698175906
transform 1 0 8624 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_69
timestamp 1698175906
transform 1 0 9072 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_72
timestamp 1698175906
transform 1 0 9408 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_104
timestamp 1698175906
transform 1 0 12992 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_142
timestamp 1698175906
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_146
timestamp 1698175906
transform 1 0 17696 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_162
timestamp 1698175906
transform 1 0 19488 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_208
timestamp 1698175906
transform 1 0 24640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_212
timestamp 1698175906
transform 1 0 25088 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_276
timestamp 1698175906
transform 1 0 32256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_282
timestamp 1698175906
transform 1 0 32928 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_314
timestamp 1698175906
transform 1 0 36512 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_330
timestamp 1698175906
transform 1 0 38304 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_335
timestamp 1698175906
transform 1 0 38864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_343
timestamp 1698175906
transform 1 0 39760 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_347
timestamp 1698175906
transform 1 0 40208 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_349
timestamp 1698175906
transform 1 0 40432 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_352
timestamp 1698175906
transform 1 0 40768 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_368
timestamp 1698175906
transform 1 0 42560 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_376
timestamp 1698175906
transform 1 0 43456 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_378
timestamp 1698175906
transform 1 0 43680 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_383
timestamp 1698175906
transform 1 0 44240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_387
timestamp 1698175906
transform 1 0 44688 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_419
timestamp 1698175906
transform 1 0 48272 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_422
timestamp 1698175906
transform 1 0 48608 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_434
timestamp 1698175906
transform 1 0 49952 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_436
timestamp 1698175906
transform 1 0 50176 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_439
timestamp 1698175906
transform 1 0 50512 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_455
timestamp 1698175906
transform 1 0 52304 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_463
timestamp 1698175906
transform 1 0 53200 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_466
timestamp 1698175906
transform 1 0 53536 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_470
timestamp 1698175906
transform 1 0 53984 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_474
timestamp 1698175906
transform 1 0 54432 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_478
timestamp 1698175906
transform 1 0 54880 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_482
timestamp 1698175906
transform 1 0 55328 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_486
timestamp 1698175906
transform 1 0 55776 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_507
timestamp 1698175906
transform 1 0 58128 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_512
timestamp 1698175906
transform 1 0 58688 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_544
timestamp 1698175906
transform 1 0 62272 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_562
timestamp 1698175906
transform 1 0 64288 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_578
timestamp 1698175906
transform 1 0 66080 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_586
timestamp 1698175906
transform 1 0 66976 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_590
timestamp 1698175906
transform 1 0 67424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_592
timestamp 1698175906
transform 1 0 67648 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_595
timestamp 1698175906
transform 1 0 67984 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_627
timestamp 1698175906
transform 1 0 71568 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_629
timestamp 1698175906
transform 1 0 71792 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_632
timestamp 1698175906
transform 1 0 72128 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_664
timestamp 1698175906
transform 1 0 75712 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_668
timestamp 1698175906
transform 1 0 76160 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_672
timestamp 1698175906
transform 1 0 76608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_676
timestamp 1698175906
transform 1 0 77056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_697
timestamp 1698175906
transform 1 0 79408 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_699
timestamp 1698175906
transform 1 0 79632 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_702
timestamp 1698175906
transform 1 0 79968 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_734
timestamp 1698175906
transform 1 0 83552 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_750
timestamp 1698175906
transform 1 0 85344 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_758
timestamp 1698175906
transform 1 0 86240 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_768
timestamp 1698175906
transform 1 0 87360 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_787
timestamp 1698175906
transform 1 0 89488 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_803
timestamp 1698175906
transform 1 0 91280 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_807
timestamp 1698175906
transform 1 0 91728 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_814
timestamp 1698175906
transform 1 0 92512 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_830
timestamp 1698175906
transform 1 0 94304 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_838
timestamp 1698175906
transform 1 0 95200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_842
timestamp 1698175906
transform 1 0 95648 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_858
timestamp 1698175906
transform 1 0 97440 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_8
timestamp 1698175906
transform 1 0 2240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_12
timestamp 1698175906
transform 1 0 2688 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_17
timestamp 1698175906
transform 1 0 3248 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_33
timestamp 1698175906
transform 1 0 5040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_37
timestamp 1698175906
transform 1 0 5488 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_69
timestamp 1698175906
transform 1 0 9072 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_85
timestamp 1698175906
transform 1 0 10864 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_93
timestamp 1698175906
transform 1 0 11760 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_122
timestamp 1698175906
transform 1 0 15008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_126
timestamp 1698175906
transform 1 0 15456 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_142
timestamp 1698175906
transform 1 0 17248 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_150
timestamp 1698175906
transform 1 0 18144 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_154
timestamp 1698175906
transform 1 0 18592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_156
timestamp 1698175906
transform 1 0 18816 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698175906
transform 1 0 20832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_181
timestamp 1698175906
transform 1 0 21616 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_185
timestamp 1698175906
transform 1 0 22064 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_217
timestamp 1698175906
transform 1 0 25648 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_225
timestamp 1698175906
transform 1 0 26544 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_233
timestamp 1698175906
transform 1 0 27440 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_241
timestamp 1698175906
transform 1 0 28336 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_247
timestamp 1698175906
transform 1 0 29008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_249
timestamp 1698175906
transform 1 0 29232 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_252
timestamp 1698175906
transform 1 0 29568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_260
timestamp 1698175906
transform 1 0 30464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_264
timestamp 1698175906
transform 1 0 30912 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_302
timestamp 1698175906
transform 1 0 35168 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_310
timestamp 1698175906
transform 1 0 36064 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_314
timestamp 1698175906
transform 1 0 36512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_317
timestamp 1698175906
transform 1 0 36848 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698175906
transform 1 0 44016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_387
timestamp 1698175906
transform 1 0 44688 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_451
timestamp 1698175906
transform 1 0 51856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_457
timestamp 1698175906
transform 1 0 52528 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_521
timestamp 1698175906
transform 1 0 59696 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_527
timestamp 1698175906
transform 1 0 60368 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_535
timestamp 1698175906
transform 1 0 61264 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_539
timestamp 1698175906
transform 1 0 61712 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_576
timestamp 1698175906
transform 1 0 65856 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_592
timestamp 1698175906
transform 1 0 67648 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_594
timestamp 1698175906
transform 1 0 67872 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_597
timestamp 1698175906
transform 1 0 68208 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_605
timestamp 1698175906
transform 1 0 69104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_643
timestamp 1698175906
transform 1 0 73360 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_659
timestamp 1698175906
transform 1 0 75152 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_663
timestamp 1698175906
transform 1 0 75600 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_667
timestamp 1698175906
transform 1 0 76048 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_675
timestamp 1698175906
transform 1 0 76944 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_679
timestamp 1698175906
transform 1 0 77392 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_687
timestamp 1698175906
transform 1 0 78288 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_719
timestamp 1698175906
transform 1 0 81872 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_737
timestamp 1698175906
transform 1 0 83888 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_753
timestamp 1698175906
transform 1 0 85680 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_757
timestamp 1698175906
transform 1 0 86128 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_793
timestamp 1698175906
transform 1 0 90160 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_797
timestamp 1698175906
transform 1 0 90608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_801
timestamp 1698175906
transform 1 0 91056 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_822
timestamp 1698175906
transform 1 0 93408 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_838
timestamp 1698175906
transform 1 0 95200 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_50
timestamp 1698175906
transform 1 0 6944 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_54
timestamp 1698175906
transform 1 0 7392 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_108
timestamp 1698175906
transform 1 0 13440 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_110
timestamp 1698175906
transform 1 0 13664 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_115
timestamp 1698175906
transform 1 0 14224 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_131
timestamp 1698175906
transform 1 0 16016 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_139
timestamp 1698175906
transform 1 0 16912 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_142
timestamp 1698175906
transform 1 0 17248 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_206
timestamp 1698175906
transform 1 0 24416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_265
timestamp 1698175906
transform 1 0 31024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_269
timestamp 1698175906
transform 1 0 31472 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_274
timestamp 1698175906
transform 1 0 32032 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_288
timestamp 1698175906
transform 1 0 33600 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_336
timestamp 1698175906
transform 1 0 38976 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_340
timestamp 1698175906
transform 1 0 39424 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_344
timestamp 1698175906
transform 1 0 39872 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_348
timestamp 1698175906
transform 1 0 40320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_352
timestamp 1698175906
transform 1 0 40768 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_368
timestamp 1698175906
transform 1 0 42560 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_372
timestamp 1698175906
transform 1 0 43008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_410
timestamp 1698175906
transform 1 0 47264 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_418
timestamp 1698175906
transform 1 0 48160 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_422
timestamp 1698175906
transform 1 0 48608 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_430
timestamp 1698175906
transform 1 0 49504 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_432
timestamp 1698175906
transform 1 0 49728 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_467
timestamp 1698175906
transform 1 0 53648 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_471
timestamp 1698175906
transform 1 0 54096 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_479
timestamp 1698175906
transform 1 0 54992 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_483
timestamp 1698175906
transform 1 0 55440 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_486
timestamp 1698175906
transform 1 0 55776 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_526
timestamp 1698175906
transform 1 0 60256 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_542
timestamp 1698175906
transform 1 0 62048 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_548
timestamp 1698175906
transform 1 0 62720 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_556
timestamp 1698175906
transform 1 0 63616 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_562
timestamp 1698175906
transform 1 0 64288 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_566
timestamp 1698175906
transform 1 0 64736 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_570
timestamp 1698175906
transform 1 0 65184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_590
timestamp 1698175906
transform 1 0 67424 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_606
timestamp 1698175906
transform 1 0 69216 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_610
timestamp 1698175906
transform 1 0 69664 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_621
timestamp 1698175906
transform 1 0 70896 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_623
timestamp 1698175906
transform 1 0 71120 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_626
timestamp 1698175906
transform 1 0 71456 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_647
timestamp 1698175906
transform 1 0 73808 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_655
timestamp 1698175906
transform 1 0 74704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_659
timestamp 1698175906
transform 1 0 75152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_679
timestamp 1698175906
transform 1 0 77392 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_695
timestamp 1698175906
transform 1 0 79184 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_699
timestamp 1698175906
transform 1 0 79632 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_702
timestamp 1698175906
transform 1 0 79968 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_706
timestamp 1698175906
transform 1 0 80416 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_743
timestamp 1698175906
transform 1 0 84560 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_759
timestamp 1698175906
transform 1 0 86352 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_764
timestamp 1698175906
transform 1 0 86912 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_768
timestamp 1698175906
transform 1 0 87360 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_772
timestamp 1698175906
transform 1 0 87808 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_788
timestamp 1698175906
transform 1 0 89600 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_796
timestamp 1698175906
transform 1 0 90496 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_842
timestamp 1698175906
transform 1 0 95648 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_858
timestamp 1698175906
transform 1 0 97440 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_2
timestamp 1698175906
transform 1 0 1568 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_6
timestamp 1698175906
transform 1 0 2016 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_14
timestamp 1698175906
transform 1 0 2912 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_30
timestamp 1698175906
transform 1 0 4704 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698175906
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_37
timestamp 1698175906
transform 1 0 5488 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_53
timestamp 1698175906
transform 1 0 7280 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_57
timestamp 1698175906
transform 1 0 7728 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_59
timestamp 1698175906
transform 1 0 7952 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_85
timestamp 1698175906
transform 1 0 10864 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_89
timestamp 1698175906
transform 1 0 11312 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_93
timestamp 1698175906
transform 1 0 11760 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_101
timestamp 1698175906
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_107
timestamp 1698175906
transform 1 0 13328 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_111
timestamp 1698175906
transform 1 0 13776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_149
timestamp 1698175906
transform 1 0 18032 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_165
timestamp 1698175906
transform 1 0 19824 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_192
timestamp 1698175906
transform 1 0 22848 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_196
timestamp 1698175906
transform 1 0 23296 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_228
timestamp 1698175906
transform 1 0 26880 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_244
timestamp 1698175906
transform 1 0 28672 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_247
timestamp 1698175906
transform 1 0 29008 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_263
timestamp 1698175906
transform 1 0 30800 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_267
timestamp 1698175906
transform 1 0 31248 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_283
timestamp 1698175906
transform 1 0 33040 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_287
timestamp 1698175906
transform 1 0 33488 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_303
timestamp 1698175906
transform 1 0 35280 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_307
timestamp 1698175906
transform 1 0 35728 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_311
timestamp 1698175906
transform 1 0 36176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_317
timestamp 1698175906
transform 1 0 36848 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_359
timestamp 1698175906
transform 1 0 41552 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_363
timestamp 1698175906
transform 1 0 42000 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_402
timestamp 1698175906
transform 1 0 46368 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_406
timestamp 1698175906
transform 1 0 46816 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_454
timestamp 1698175906
transform 1 0 52192 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_457
timestamp 1698175906
transform 1 0 52528 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_461
timestamp 1698175906
transform 1 0 52976 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_469
timestamp 1698175906
transform 1 0 53872 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_488
timestamp 1698175906
transform 1 0 56000 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_508
timestamp 1698175906
transform 1 0 58240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_512
timestamp 1698175906
transform 1 0 58688 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_520
timestamp 1698175906
transform 1 0 59584 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_524
timestamp 1698175906
transform 1 0 60032 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_527
timestamp 1698175906
transform 1 0 60368 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_543
timestamp 1698175906
transform 1 0 62160 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_547
timestamp 1698175906
transform 1 0 62608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_549
timestamp 1698175906
transform 1 0 62832 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_552
timestamp 1698175906
transform 1 0 63168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_556
timestamp 1698175906
transform 1 0 63616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_573
timestamp 1698175906
transform 1 0 65520 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_589
timestamp 1698175906
transform 1 0 67312 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_593
timestamp 1698175906
transform 1 0 67760 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_597
timestamp 1698175906
transform 1 0 68208 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_605
timestamp 1698175906
transform 1 0 69104 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_609
timestamp 1698175906
transform 1 0 69552 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_612
timestamp 1698175906
transform 1 0 69888 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_628
timestamp 1698175906
transform 1 0 71680 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_636
timestamp 1698175906
transform 1 0 72576 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_642
timestamp 1698175906
transform 1 0 73248 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_662
timestamp 1698175906
transform 1 0 75488 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_664
timestamp 1698175906
transform 1 0 75712 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_667
timestamp 1698175906
transform 1 0 76048 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_673
timestamp 1698175906
transform 1 0 76720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_690
timestamp 1698175906
transform 1 0 78624 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_698
timestamp 1698175906
transform 1 0 79520 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_705
timestamp 1698175906
transform 1 0 80304 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_709
timestamp 1698175906
transform 1 0 80752 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_715
timestamp 1698175906
transform 1 0 81424 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_731
timestamp 1698175906
transform 1 0 83216 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_737
timestamp 1698175906
transform 1 0 83888 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_801
timestamp 1698175906
transform 1 0 91056 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_807
timestamp 1698175906
transform 1 0 91728 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_839
timestamp 1698175906
transform 1 0 95312 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_8
timestamp 1698175906
transform 1 0 2240 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_12
timestamp 1698175906
transform 1 0 2688 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_47
timestamp 1698175906
transform 1 0 6608 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_63
timestamp 1698175906
transform 1 0 8400 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_67
timestamp 1698175906
transform 1 0 8848 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_69
timestamp 1698175906
transform 1 0 9072 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_72
timestamp 1698175906
transform 1 0 9408 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_104
timestamp 1698175906
transform 1 0 12992 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_112
timestamp 1698175906
transform 1 0 13888 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_138
timestamp 1698175906
transform 1 0 16800 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_142
timestamp 1698175906
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_146
timestamp 1698175906
transform 1 0 17696 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_162
timestamp 1698175906
transform 1 0 19488 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_205
timestamp 1698175906
transform 1 0 24304 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_209
timestamp 1698175906
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_212
timestamp 1698175906
transform 1 0 25088 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_276
timestamp 1698175906
transform 1 0 32256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_282
timestamp 1698175906
transform 1 0 32928 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_314
timestamp 1698175906
transform 1 0 36512 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_318
timestamp 1698175906
transform 1 0 36960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_367
timestamp 1698175906
transform 1 0 42448 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_371
timestamp 1698175906
transform 1 0 42896 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_375
timestamp 1698175906
transform 1 0 43344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_377
timestamp 1698175906
transform 1 0 43568 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_382
timestamp 1698175906
transform 1 0 44128 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_384
timestamp 1698175906
transform 1 0 44352 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_387
timestamp 1698175906
transform 1 0 44688 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_403
timestamp 1698175906
transform 1 0 46480 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_407
timestamp 1698175906
transform 1 0 46928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_409
timestamp 1698175906
transform 1 0 47152 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_415
timestamp 1698175906
transform 1 0 47824 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_419
timestamp 1698175906
transform 1 0 48272 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_422
timestamp 1698175906
transform 1 0 48608 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_430
timestamp 1698175906
transform 1 0 49504 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_434
timestamp 1698175906
transform 1 0 49952 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_439
timestamp 1698175906
transform 1 0 50512 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_447
timestamp 1698175906
transform 1 0 51408 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_450
timestamp 1698175906
transform 1 0 51744 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_466
timestamp 1698175906
transform 1 0 53536 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_476
timestamp 1698175906
transform 1 0 54656 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_484
timestamp 1698175906
transform 1 0 55552 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_486
timestamp 1698175906
transform 1 0 55776 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_489
timestamp 1698175906
transform 1 0 56112 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_498
timestamp 1698175906
transform 1 0 57120 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_530
timestamp 1698175906
transform 1 0 60704 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_534
timestamp 1698175906
transform 1 0 61152 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_537
timestamp 1698175906
transform 1 0 61488 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_541
timestamp 1698175906
transform 1 0 61936 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_558
timestamp 1698175906
transform 1 0 63840 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_562
timestamp 1698175906
transform 1 0 64288 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_566
timestamp 1698175906
transform 1 0 64736 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_598
timestamp 1698175906
transform 1 0 68320 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_605
timestamp 1698175906
transform 1 0 69104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_607
timestamp 1698175906
transform 1 0 69328 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_610
timestamp 1698175906
transform 1 0 69664 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_627
timestamp 1698175906
transform 1 0 71568 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_629
timestamp 1698175906
transform 1 0 71792 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_632
timestamp 1698175906
transform 1 0 72128 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_640
timestamp 1698175906
transform 1 0 73024 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_646
timestamp 1698175906
transform 1 0 73696 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_662
timestamp 1698175906
transform 1 0 75488 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_666
timestamp 1698175906
transform 1 0 75936 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_668
timestamp 1698175906
transform 1 0 76160 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_671
timestamp 1698175906
transform 1 0 76496 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_675
timestamp 1698175906
transform 1 0 76944 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_677
timestamp 1698175906
transform 1 0 77168 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_693
timestamp 1698175906
transform 1 0 78960 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_697
timestamp 1698175906
transform 1 0 79408 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_699
timestamp 1698175906
transform 1 0 79632 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_702
timestamp 1698175906
transform 1 0 79968 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_714
timestamp 1698175906
transform 1 0 81312 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_746
timestamp 1698175906
transform 1 0 84896 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_762
timestamp 1698175906
transform 1 0 86688 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_772
timestamp 1698175906
transform 1 0 87808 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_788
timestamp 1698175906
transform 1 0 89600 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_796
timestamp 1698175906
transform 1 0 90496 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_799
timestamp 1698175906
transform 1 0 90832 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_803
timestamp 1698175906
transform 1 0 91280 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_820
timestamp 1698175906
transform 1 0 93184 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_836
timestamp 1698175906
transform 1 0 94976 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_842
timestamp 1698175906
transform 1 0 95648 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_858
timestamp 1698175906
transform 1 0 97440 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_8
timestamp 1698175906
transform 1 0 2240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_12
timestamp 1698175906
transform 1 0 2688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_14
timestamp 1698175906
transform 1 0 2912 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_19
timestamp 1698175906
transform 1 0 3472 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_37
timestamp 1698175906
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_101
timestamp 1698175906
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_107
timestamp 1698175906
transform 1 0 13328 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_115
timestamp 1698175906
transform 1 0 14224 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_119
timestamp 1698175906
transform 1 0 14672 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_123
timestamp 1698175906
transform 1 0 15120 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_155
timestamp 1698175906
transform 1 0 18704 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_171
timestamp 1698175906
transform 1 0 20496 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_181
timestamp 1698175906
transform 1 0 21616 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_213
timestamp 1698175906
transform 1 0 25200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_215
timestamp 1698175906
transform 1 0 25424 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_220
timestamp 1698175906
transform 1 0 25984 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_224
timestamp 1698175906
transform 1 0 26432 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_226
timestamp 1698175906
transform 1 0 26656 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_233
timestamp 1698175906
transform 1 0 27440 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_241
timestamp 1698175906
transform 1 0 28336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_247
timestamp 1698175906
transform 1 0 29008 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_251
timestamp 1698175906
transform 1 0 29456 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_259
timestamp 1698175906
transform 1 0 30352 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_297
timestamp 1698175906
transform 1 0 34608 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_313
timestamp 1698175906
transform 1 0 36400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_317
timestamp 1698175906
transform 1 0 36848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_325
timestamp 1698175906
transform 1 0 37744 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_329
timestamp 1698175906
transform 1 0 38192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_331
timestamp 1698175906
transform 1 0 38416 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_334
timestamp 1698175906
transform 1 0 38752 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_338
timestamp 1698175906
transform 1 0 39200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_342
timestamp 1698175906
transform 1 0 39648 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_349
timestamp 1698175906
transform 1 0 40432 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_353
timestamp 1698175906
transform 1 0 40880 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_387
timestamp 1698175906
transform 1 0 44688 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_403
timestamp 1698175906
transform 1 0 46480 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_443
timestamp 1698175906
transform 1 0 50960 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_451
timestamp 1698175906
transform 1 0 51856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_457
timestamp 1698175906
transform 1 0 52528 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_465
timestamp 1698175906
transform 1 0 53424 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_469
timestamp 1698175906
transform 1 0 53872 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_472
timestamp 1698175906
transform 1 0 54208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_476
timestamp 1698175906
transform 1 0 54656 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_561
timestamp 1698175906
transform 1 0 64176 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_568
timestamp 1698175906
transform 1 0 64960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_572
timestamp 1698175906
transform 1 0 65408 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_588
timestamp 1698175906
transform 1 0 67200 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_592
timestamp 1698175906
transform 1 0 67648 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_631
timestamp 1698175906
transform 1 0 72016 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_635
timestamp 1698175906
transform 1 0 72464 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_643
timestamp 1698175906
transform 1 0 73360 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_659
timestamp 1698175906
transform 1 0 75152 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_663
timestamp 1698175906
transform 1 0 75600 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_667
timestamp 1698175906
transform 1 0 76048 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_682
timestamp 1698175906
transform 1 0 77728 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_686
timestamp 1698175906
transform 1 0 78176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_690
timestamp 1698175906
transform 1 0 78624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_692
timestamp 1698175906
transform 1 0 78848 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_737
timestamp 1698175906
transform 1 0 83888 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_753
timestamp 1698175906
transform 1 0 85680 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_789
timestamp 1698175906
transform 1 0 89712 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_793
timestamp 1698175906
transform 1 0 90160 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_801
timestamp 1698175906
transform 1 0 91056 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_807
timestamp 1698175906
transform 1 0 91728 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_843
timestamp 1698175906
transform 1 0 95760 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_859
timestamp 1698175906
transform 1 0 97552 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_863
timestamp 1698175906
transform 1 0 98000 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_865
timestamp 1698175906
transform 1 0 98224 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_2
timestamp 1698175906
transform 1 0 1568 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_6
timestamp 1698175906
transform 1 0 2016 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_42
timestamp 1698175906
transform 1 0 6048 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_58
timestamp 1698175906
transform 1 0 7840 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_62
timestamp 1698175906
transform 1 0 8288 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_108
timestamp 1698175906
transform 1 0 13440 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_142
timestamp 1698175906
transform 1 0 17248 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_174
timestamp 1698175906
transform 1 0 20832 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_177
timestamp 1698175906
transform 1 0 21168 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_209
timestamp 1698175906
transform 1 0 24752 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_212
timestamp 1698175906
transform 1 0 25088 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_214
timestamp 1698175906
transform 1 0 25312 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_264
timestamp 1698175906
transform 1 0 30912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_268
timestamp 1698175906
transform 1 0 31360 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_272
timestamp 1698175906
transform 1 0 31808 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_282
timestamp 1698175906
transform 1 0 32928 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_284
timestamp 1698175906
transform 1 0 33152 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_334
timestamp 1698175906
transform 1 0 38752 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_352
timestamp 1698175906
transform 1 0 40768 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_356
timestamp 1698175906
transform 1 0 41216 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_408
timestamp 1698175906
transform 1 0 47040 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_416
timestamp 1698175906
transform 1 0 47936 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_422
timestamp 1698175906
transform 1 0 48608 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_438
timestamp 1698175906
transform 1 0 50400 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_446
timestamp 1698175906
transform 1 0 51296 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_464
timestamp 1698175906
transform 1 0 53312 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_468
timestamp 1698175906
transform 1 0 53760 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_474
timestamp 1698175906
transform 1 0 54432 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_478
timestamp 1698175906
transform 1 0 54880 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_482
timestamp 1698175906
transform 1 0 55328 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_486
timestamp 1698175906
transform 1 0 55776 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_545
timestamp 1698175906
transform 1 0 62384 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_553
timestamp 1698175906
transform 1 0 63280 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_557
timestamp 1698175906
transform 1 0 63728 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_559
timestamp 1698175906
transform 1 0 63952 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_562
timestamp 1698175906
transform 1 0 64288 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_566
timestamp 1698175906
transform 1 0 64736 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_585
timestamp 1698175906
transform 1 0 66864 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_593
timestamp 1698175906
transform 1 0 67760 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_625
timestamp 1698175906
transform 1 0 71344 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_629
timestamp 1698175906
transform 1 0 71792 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_632
timestamp 1698175906
transform 1 0 72128 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_640
timestamp 1698175906
transform 1 0 73024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_642
timestamp 1698175906
transform 1 0 73248 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_661
timestamp 1698175906
transform 1 0 75376 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_669
timestamp 1698175906
transform 1 0 76272 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_689
timestamp 1698175906
transform 1 0 78512 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_697
timestamp 1698175906
transform 1 0 79408 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_699
timestamp 1698175906
transform 1 0 79632 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_702
timestamp 1698175906
transform 1 0 79968 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_734
timestamp 1698175906
transform 1 0 83552 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_742
timestamp 1698175906
transform 1 0 84448 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_746
timestamp 1698175906
transform 1 0 84896 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_749
timestamp 1698175906
transform 1 0 85232 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_753
timestamp 1698175906
transform 1 0 85680 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_772
timestamp 1698175906
transform 1 0 87808 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_804
timestamp 1698175906
transform 1 0 91392 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_806
timestamp 1698175906
transform 1 0 91616 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_817
timestamp 1698175906
transform 1 0 92848 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_833
timestamp 1698175906
transform 1 0 94640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_837
timestamp 1698175906
transform 1 0 95088 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_839
timestamp 1698175906
transform 1 0 95312 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_842
timestamp 1698175906
transform 1 0 95648 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_8
timestamp 1698175906
transform 1 0 2240 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_14
timestamp 1698175906
transform 1 0 2912 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_30
timestamp 1698175906
transform 1 0 4704 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698175906
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_37
timestamp 1698175906
transform 1 0 5488 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_53
timestamp 1698175906
transform 1 0 7280 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_61
timestamp 1698175906
transform 1 0 8176 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_65
timestamp 1698175906
transform 1 0 8624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_71
timestamp 1698175906
transform 1 0 9296 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_87
timestamp 1698175906
transform 1 0 11088 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_91
timestamp 1698175906
transform 1 0 11536 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_95
timestamp 1698175906
transform 1 0 11984 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_103
timestamp 1698175906
transform 1 0 12880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_107
timestamp 1698175906
transform 1 0 13328 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_111
timestamp 1698175906
transform 1 0 13776 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_113
timestamp 1698175906
transform 1 0 14000 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_148
timestamp 1698175906
transform 1 0 17920 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_152
timestamp 1698175906
transform 1 0 18368 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_168
timestamp 1698175906
transform 1 0 20160 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_211
timestamp 1698175906
transform 1 0 24976 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_243
timestamp 1698175906
transform 1 0 28560 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_247
timestamp 1698175906
transform 1 0 29008 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_263
timestamp 1698175906
transform 1 0 30800 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_269
timestamp 1698175906
transform 1 0 31472 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_285
timestamp 1698175906
transform 1 0 33264 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_301
timestamp 1698175906
transform 1 0 35056 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_305
timestamp 1698175906
transform 1 0 35504 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_309
timestamp 1698175906
transform 1 0 35952 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_317
timestamp 1698175906
transform 1 0 36848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_319
timestamp 1698175906
transform 1 0 37072 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_376
timestamp 1698175906
transform 1 0 43456 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_380
timestamp 1698175906
transform 1 0 43904 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_382
timestamp 1698175906
transform 1 0 44128 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_402
timestamp 1698175906
transform 1 0 46368 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_404
timestamp 1698175906
transform 1 0 46592 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_421
timestamp 1698175906
transform 1 0 48496 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_425
timestamp 1698175906
transform 1 0 48944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_429
timestamp 1698175906
transform 1 0 49392 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_437
timestamp 1698175906
transform 1 0 50288 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_444
timestamp 1698175906
transform 1 0 51072 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_452
timestamp 1698175906
transform 1 0 51968 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_454
timestamp 1698175906
transform 1 0 52192 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_457
timestamp 1698175906
transform 1 0 52528 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_473
timestamp 1698175906
transform 1 0 54320 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_510
timestamp 1698175906
transform 1 0 58464 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_518
timestamp 1698175906
transform 1 0 59360 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_522
timestamp 1698175906
transform 1 0 59808 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_524
timestamp 1698175906
transform 1 0 60032 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_527
timestamp 1698175906
transform 1 0 60368 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_533
timestamp 1698175906
transform 1 0 61040 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_565
timestamp 1698175906
transform 1 0 64624 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_581
timestamp 1698175906
transform 1 0 66416 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_589
timestamp 1698175906
transform 1 0 67312 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_593
timestamp 1698175906
transform 1 0 67760 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_597
timestamp 1698175906
transform 1 0 68208 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_613
timestamp 1698175906
transform 1 0 70000 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_655
timestamp 1698175906
transform 1 0 74704 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_659
timestamp 1698175906
transform 1 0 75152 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_663
timestamp 1698175906
transform 1 0 75600 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_667
timestamp 1698175906
transform 1 0 76048 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_675
timestamp 1698175906
transform 1 0 76944 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_681
timestamp 1698175906
transform 1 0 77616 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_689
timestamp 1698175906
transform 1 0 78512 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_693
timestamp 1698175906
transform 1 0 78960 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_700
timestamp 1698175906
transform 1 0 79744 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_732
timestamp 1698175906
transform 1 0 83328 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_734
timestamp 1698175906
transform 1 0 83552 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_737
timestamp 1698175906
transform 1 0 83888 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_753
timestamp 1698175906
transform 1 0 85680 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_757
timestamp 1698175906
transform 1 0 86128 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_768
timestamp 1698175906
transform 1 0 87360 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_800
timestamp 1698175906
transform 1 0 90944 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_804
timestamp 1698175906
transform 1 0 91392 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_807
timestamp 1698175906
transform 1 0 91728 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_811
timestamp 1698175906
transform 1 0 92176 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_819
timestamp 1698175906
transform 1 0 93072 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_851
timestamp 1698175906
transform 1 0 96656 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_859
timestamp 1698175906
transform 1 0 97552 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_863
timestamp 1698175906
transform 1 0 98000 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_865
timestamp 1698175906
transform 1 0 98224 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_36
timestamp 1698175906
transform 1 0 5376 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_40
timestamp 1698175906
transform 1 0 5824 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_56
timestamp 1698175906
transform 1 0 7616 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_64
timestamp 1698175906
transform 1 0 8512 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_68
timestamp 1698175906
transform 1 0 8960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_72
timestamp 1698175906
transform 1 0 9408 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_104
timestamp 1698175906
transform 1 0 12992 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_108
timestamp 1698175906
transform 1 0 13440 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_132
timestamp 1698175906
transform 1 0 16128 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_136
timestamp 1698175906
transform 1 0 16576 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_142
timestamp 1698175906
transform 1 0 17248 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_158
timestamp 1698175906
transform 1 0 19040 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_162
timestamp 1698175906
transform 1 0 19488 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_164
timestamp 1698175906
transform 1 0 19712 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_182
timestamp 1698175906
transform 1 0 21728 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_186
timestamp 1698175906
transform 1 0 22176 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_202
timestamp 1698175906
transform 1 0 23968 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_212
timestamp 1698175906
transform 1 0 25088 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_276
timestamp 1698175906
transform 1 0 32256 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_282
timestamp 1698175906
transform 1 0 32928 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_314
timestamp 1698175906
transform 1 0 36512 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_352
timestamp 1698175906
transform 1 0 40768 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_356
timestamp 1698175906
transform 1 0 41216 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_372
timestamp 1698175906
transform 1 0 43008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_374
timestamp 1698175906
transform 1 0 43232 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_385
timestamp 1698175906
transform 1 0 44464 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_401
timestamp 1698175906
transform 1 0 46256 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_404
timestamp 1698175906
transform 1 0 46592 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_422
timestamp 1698175906
transform 1 0 48608 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_461
timestamp 1698175906
transform 1 0 52976 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_465
timestamp 1698175906
transform 1 0 53424 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_481
timestamp 1698175906
transform 1 0 55216 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_483
timestamp 1698175906
transform 1 0 55440 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_507
timestamp 1698175906
transform 1 0 58128 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_511
timestamp 1698175906
transform 1 0 58576 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_543
timestamp 1698175906
transform 1 0 62160 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_551
timestamp 1698175906
transform 1 0 63056 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_555
timestamp 1698175906
transform 1 0 63504 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_557
timestamp 1698175906
transform 1 0 63728 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_562
timestamp 1698175906
transform 1 0 64288 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_575
timestamp 1698175906
transform 1 0 65744 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_607
timestamp 1698175906
transform 1 0 69328 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_615
timestamp 1698175906
transform 1 0 70224 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_619
timestamp 1698175906
transform 1 0 70672 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_656
timestamp 1698175906
transform 1 0 74816 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_664
timestamp 1698175906
transform 1 0 75712 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_668
timestamp 1698175906
transform 1 0 76160 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_672
timestamp 1698175906
transform 1 0 76608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_698
timestamp 1698175906
transform 1 0 79520 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_736
timestamp 1698175906
transform 1 0 83776 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_768
timestamp 1698175906
transform 1 0 87360 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_772
timestamp 1698175906
transform 1 0 87808 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_788
timestamp 1698175906
transform 1 0 89600 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_796
timestamp 1698175906
transform 1 0 90496 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_800
timestamp 1698175906
transform 1 0 90944 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_804
timestamp 1698175906
transform 1 0 91392 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_808
timestamp 1698175906
transform 1 0 91840 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_825
timestamp 1698175906
transform 1 0 93744 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_833
timestamp 1698175906
transform 1 0 94640 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_837
timestamp 1698175906
transform 1 0 95088 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_839
timestamp 1698175906
transform 1 0 95312 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_842
timestamp 1698175906
transform 1 0 95648 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_14
timestamp 1698175906
transform 1 0 2912 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_18
timestamp 1698175906
transform 1 0 3360 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698175906
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_37
timestamp 1698175906
transform 1 0 5488 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_53
timestamp 1698175906
transform 1 0 7280 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_61
timestamp 1698175906
transform 1 0 8176 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_65
timestamp 1698175906
transform 1 0 8624 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_100
timestamp 1698175906
transform 1 0 12544 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_104
timestamp 1698175906
transform 1 0 12992 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_107
timestamp 1698175906
transform 1 0 13328 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_115
timestamp 1698175906
transform 1 0 14224 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_120
timestamp 1698175906
transform 1 0 14784 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_152
timestamp 1698175906
transform 1 0 18368 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_168
timestamp 1698175906
transform 1 0 20160 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_170
timestamp 1698175906
transform 1 0 20384 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_177
timestamp 1698175906
transform 1 0 21168 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_241
timestamp 1698175906
transform 1 0 28336 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_247
timestamp 1698175906
transform 1 0 29008 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_251
timestamp 1698175906
transform 1 0 29456 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_267
timestamp 1698175906
transform 1 0 31248 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_271
timestamp 1698175906
transform 1 0 31696 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_273
timestamp 1698175906
transform 1 0 31920 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_305
timestamp 1698175906
transform 1 0 35504 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_309
timestamp 1698175906
transform 1 0 35952 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_313
timestamp 1698175906
transform 1 0 36400 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_317
timestamp 1698175906
transform 1 0 36848 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_381
timestamp 1698175906
transform 1 0 44016 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_387
timestamp 1698175906
transform 1 0 44688 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_451
timestamp 1698175906
transform 1 0 51856 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_457
timestamp 1698175906
transform 1 0 52528 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_473
timestamp 1698175906
transform 1 0 54320 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_477
timestamp 1698175906
transform 1 0 54768 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_482
timestamp 1698175906
transform 1 0 55328 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_492
timestamp 1698175906
transform 1 0 56448 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_524
timestamp 1698175906
transform 1 0 60032 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_527
timestamp 1698175906
transform 1 0 60368 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_537
timestamp 1698175906
transform 1 0 61488 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_553
timestamp 1698175906
transform 1 0 63280 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_555
timestamp 1698175906
transform 1 0 63504 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_558
timestamp 1698175906
transform 1 0 63840 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_562
timestamp 1698175906
transform 1 0 64288 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_579
timestamp 1698175906
transform 1 0 66192 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_597
timestamp 1698175906
transform 1 0 68208 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_613
timestamp 1698175906
transform 1 0 70000 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_621
timestamp 1698175906
transform 1 0 70896 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_625
timestamp 1698175906
transform 1 0 71344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_627
timestamp 1698175906
transform 1 0 71568 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_630
timestamp 1698175906
transform 1 0 71904 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_634
timestamp 1698175906
transform 1 0 72352 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_642
timestamp 1698175906
transform 1 0 73248 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_645
timestamp 1698175906
transform 1 0 73584 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_649
timestamp 1698175906
transform 1 0 74032 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_667
timestamp 1698175906
transform 1 0 76048 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_675
timestamp 1698175906
transform 1 0 76944 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_679
timestamp 1698175906
transform 1 0 77392 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_683
timestamp 1698175906
transform 1 0 77840 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_699
timestamp 1698175906
transform 1 0 79632 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_702
timestamp 1698175906
transform 1 0 79968 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_707
timestamp 1698175906
transform 1 0 80528 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_723
timestamp 1698175906
transform 1 0 82320 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_731
timestamp 1698175906
transform 1 0 83216 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_737
timestamp 1698175906
transform 1 0 83888 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_741
timestamp 1698175906
transform 1 0 84336 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_794
timestamp 1698175906
transform 1 0 90272 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_798
timestamp 1698175906
transform 1 0 90720 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_802
timestamp 1698175906
transform 1 0 91168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_804
timestamp 1698175906
transform 1 0 91392 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_807
timestamp 1698175906
transform 1 0 91728 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_809
timestamp 1698175906
transform 1 0 91952 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_848
timestamp 1698175906
transform 1 0 96320 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_864
timestamp 1698175906
transform 1 0 98112 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_2
timestamp 1698175906
transform 1 0 1568 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_8
timestamp 1698175906
transform 1 0 2240 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_12
timestamp 1698175906
transform 1 0 2688 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_28
timestamp 1698175906
transform 1 0 4480 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_32
timestamp 1698175906
transform 1 0 4928 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_34
timestamp 1698175906
transform 1 0 5152 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_69
timestamp 1698175906
transform 1 0 9072 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_76
timestamp 1698175906
transform 1 0 9856 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_80
timestamp 1698175906
transform 1 0 10304 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_88
timestamp 1698175906
transform 1 0 11200 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_125
timestamp 1698175906
transform 1 0 15344 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_133
timestamp 1698175906
transform 1 0 16240 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_137
timestamp 1698175906
transform 1 0 16688 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_139
timestamp 1698175906
transform 1 0 16912 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_142
timestamp 1698175906
transform 1 0 17248 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_206
timestamp 1698175906
transform 1 0 24416 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_212
timestamp 1698175906
transform 1 0 25088 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_276
timestamp 1698175906
transform 1 0 32256 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_282
timestamp 1698175906
transform 1 0 32928 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_298
timestamp 1698175906
transform 1 0 34720 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_333
timestamp 1698175906
transform 1 0 38640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_337
timestamp 1698175906
transform 1 0 39088 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_345
timestamp 1698175906
transform 1 0 39984 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_349
timestamp 1698175906
transform 1 0 40432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_352
timestamp 1698175906
transform 1 0 40768 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_360
timestamp 1698175906
transform 1 0 41664 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_364
timestamp 1698175906
transform 1 0 42112 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_368
timestamp 1698175906
transform 1 0 42560 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_400
timestamp 1698175906
transform 1 0 46144 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_416
timestamp 1698175906
transform 1 0 47936 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_422
timestamp 1698175906
transform 1 0 48608 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_471
timestamp 1698175906
transform 1 0 54096 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_487
timestamp 1698175906
transform 1 0 55888 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_489
timestamp 1698175906
transform 1 0 56112 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_492
timestamp 1698175906
transform 1 0 56448 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_524
timestamp 1698175906
transform 1 0 60032 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_528
timestamp 1698175906
transform 1 0 60480 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_552
timestamp 1698175906
transform 1 0 63168 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_562
timestamp 1698175906
transform 1 0 64288 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_604
timestamp 1698175906
transform 1 0 68992 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_608
timestamp 1698175906
transform 1 0 69440 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_626
timestamp 1698175906
transform 1 0 71456 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_647
timestamp 1698175906
transform 1 0 73808 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_663
timestamp 1698175906
transform 1 0 75600 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_666
timestamp 1698175906
transform 1 0 75936 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_670
timestamp 1698175906
transform 1 0 76384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_687
timestamp 1698175906
transform 1 0 78288 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_695
timestamp 1698175906
transform 1 0 79184 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_699
timestamp 1698175906
transform 1 0 79632 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_702
timestamp 1698175906
transform 1 0 79968 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_734
timestamp 1698175906
transform 1 0 83552 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_750
timestamp 1698175906
transform 1 0 85344 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_760
timestamp 1698175906
transform 1 0 86464 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_768
timestamp 1698175906
transform 1 0 87360 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_772
timestamp 1698175906
transform 1 0 87808 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_804
timestamp 1698175906
transform 1 0 91392 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_814
timestamp 1698175906
transform 1 0 92512 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_830
timestamp 1698175906
transform 1 0 94304 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_838
timestamp 1698175906
transform 1 0 95200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_842
timestamp 1698175906
transform 1 0 95648 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_850
timestamp 1698175906
transform 1 0 96544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_8
timestamp 1698175906
transform 1 0 2240 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_12
timestamp 1698175906
transform 1 0 2688 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_28
timestamp 1698175906
transform 1 0 4480 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_32
timestamp 1698175906
transform 1 0 4928 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698175906
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_41
timestamp 1698175906
transform 1 0 5936 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_107
timestamp 1698175906
transform 1 0 13328 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_123
timestamp 1698175906
transform 1 0 15120 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_171
timestamp 1698175906
transform 1 0 20496 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_177
timestamp 1698175906
transform 1 0 21168 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_209
timestamp 1698175906
transform 1 0 24752 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_225
timestamp 1698175906
transform 1 0 26544 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_233
timestamp 1698175906
transform 1 0 27440 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_235
timestamp 1698175906
transform 1 0 27664 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_240
timestamp 1698175906
transform 1 0 28224 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_244
timestamp 1698175906
transform 1 0 28672 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_247
timestamp 1698175906
transform 1 0 29008 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_253
timestamp 1698175906
transform 1 0 29680 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_257
timestamp 1698175906
transform 1 0 30128 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_273
timestamp 1698175906
transform 1 0 31920 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_279
timestamp 1698175906
transform 1 0 32592 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_283
timestamp 1698175906
transform 1 0 33040 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_317
timestamp 1698175906
transform 1 0 36848 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_325
timestamp 1698175906
transform 1 0 37744 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_329
timestamp 1698175906
transform 1 0 38192 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_331
timestamp 1698175906
transform 1 0 38416 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_334
timestamp 1698175906
transform 1 0 38752 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_338
timestamp 1698175906
transform 1 0 39200 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_342
timestamp 1698175906
transform 1 0 39648 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_346
timestamp 1698175906
transform 1 0 40096 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_384
timestamp 1698175906
transform 1 0 44352 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_387
timestamp 1698175906
transform 1 0 44688 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_391
timestamp 1698175906
transform 1 0 45136 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_393
timestamp 1698175906
transform 1 0 45360 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_396
timestamp 1698175906
transform 1 0 45696 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_434
timestamp 1698175906
transform 1 0 49952 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_450
timestamp 1698175906
transform 1 0 51744 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_454
timestamp 1698175906
transform 1 0 52192 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_457
timestamp 1698175906
transform 1 0 52528 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_473
timestamp 1698175906
transform 1 0 54320 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_477
timestamp 1698175906
transform 1 0 54768 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_509
timestamp 1698175906
transform 1 0 58352 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_513
timestamp 1698175906
transform 1 0 58800 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_561
timestamp 1698175906
transform 1 0 64176 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_565
timestamp 1698175906
transform 1 0 64624 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_569
timestamp 1698175906
transform 1 0 65072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_571
timestamp 1698175906
transform 1 0 65296 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_576
timestamp 1698175906
transform 1 0 65856 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_592
timestamp 1698175906
transform 1 0 67648 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_594
timestamp 1698175906
transform 1 0 67872 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_597
timestamp 1698175906
transform 1 0 68208 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_613
timestamp 1698175906
transform 1 0 70000 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_649
timestamp 1698175906
transform 1 0 74032 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_653
timestamp 1698175906
transform 1 0 74480 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_661
timestamp 1698175906
transform 1 0 75376 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_707
timestamp 1698175906
transform 1 0 80528 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_723
timestamp 1698175906
transform 1 0 82320 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_731
timestamp 1698175906
transform 1 0 83216 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_737
timestamp 1698175906
transform 1 0 83888 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_753
timestamp 1698175906
transform 1 0 85680 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_761
timestamp 1698175906
transform 1 0 86576 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_766
timestamp 1698175906
transform 1 0 87136 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_798
timestamp 1698175906
transform 1 0 90720 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_802
timestamp 1698175906
transform 1 0 91168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_804
timestamp 1698175906
transform 1 0 91392 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_807
timestamp 1698175906
transform 1 0 91728 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_839
timestamp 1698175906
transform 1 0 95312 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_843
timestamp 1698175906
transform 1 0 95760 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_845
timestamp 1698175906
transform 1 0 95984 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_852
timestamp 1698175906
transform 1 0 96768 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_860
timestamp 1698175906
transform 1 0 97664 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_864
timestamp 1698175906
transform 1 0 98112 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_8
timestamp 1698175906
transform 1 0 2240 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_12
timestamp 1698175906
transform 1 0 2688 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_44
timestamp 1698175906
transform 1 0 6272 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_60
timestamp 1698175906
transform 1 0 8064 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_68
timestamp 1698175906
transform 1 0 8960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_72
timestamp 1698175906
transform 1 0 9408 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_88
timestamp 1698175906
transform 1 0 11200 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_92
timestamp 1698175906
transform 1 0 11648 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_97
timestamp 1698175906
transform 1 0 12208 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_129
timestamp 1698175906
transform 1 0 15792 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_137
timestamp 1698175906
transform 1 0 16688 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_139
timestamp 1698175906
transform 1 0 16912 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_142
timestamp 1698175906
transform 1 0 17248 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_206
timestamp 1698175906
transform 1 0 24416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_212
timestamp 1698175906
transform 1 0 25088 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_244
timestamp 1698175906
transform 1 0 28672 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_247
timestamp 1698175906
transform 1 0 29008 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_279
timestamp 1698175906
transform 1 0 32592 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_282
timestamp 1698175906
transform 1 0 32928 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_314
timestamp 1698175906
transform 1 0 36512 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_316
timestamp 1698175906
transform 1 0 36736 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_345
timestamp 1698175906
transform 1 0 39984 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_347
timestamp 1698175906
transform 1 0 40208 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_372
timestamp 1698175906
transform 1 0 43008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_376
timestamp 1698175906
transform 1 0 43456 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_380
timestamp 1698175906
transform 1 0 43904 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_395
timestamp 1698175906
transform 1 0 45584 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_413
timestamp 1698175906
transform 1 0 47600 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_417
timestamp 1698175906
transform 1 0 48048 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_419
timestamp 1698175906
transform 1 0 48272 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_422
timestamp 1698175906
transform 1 0 48608 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_430
timestamp 1698175906
transform 1 0 49504 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_446
timestamp 1698175906
transform 1 0 51296 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_478
timestamp 1698175906
transform 1 0 54880 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_488
timestamp 1698175906
transform 1 0 56000 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_492
timestamp 1698175906
transform 1 0 56448 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_496
timestamp 1698175906
transform 1 0 56896 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_500
timestamp 1698175906
transform 1 0 57344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_504
timestamp 1698175906
transform 1 0 57792 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_536
timestamp 1698175906
transform 1 0 61376 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_538
timestamp 1698175906
transform 1 0 61600 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_545
timestamp 1698175906
transform 1 0 62384 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_553
timestamp 1698175906
transform 1 0 63280 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_557
timestamp 1698175906
transform 1 0 63728 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_559
timestamp 1698175906
transform 1 0 63952 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_562
timestamp 1698175906
transform 1 0 64288 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_594
timestamp 1698175906
transform 1 0 67872 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_610
timestamp 1698175906
transform 1 0 69664 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_614
timestamp 1698175906
transform 1 0 70112 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_616
timestamp 1698175906
transform 1 0 70336 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_627
timestamp 1698175906
transform 1 0 71568 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_629
timestamp 1698175906
transform 1 0 71792 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_632
timestamp 1698175906
transform 1 0 72128 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_664
timestamp 1698175906
transform 1 0 75712 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_668
timestamp 1698175906
transform 1 0 76160 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_670
timestamp 1698175906
transform 1 0 76384 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_673
timestamp 1698175906
transform 1 0 76720 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_679
timestamp 1698175906
transform 1 0 77392 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_695
timestamp 1698175906
transform 1 0 79184 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_699
timestamp 1698175906
transform 1 0 79632 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_702
timestamp 1698175906
transform 1 0 79968 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_766
timestamp 1698175906
transform 1 0 87136 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_772
timestamp 1698175906
transform 1 0 87808 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_788
timestamp 1698175906
transform 1 0 89600 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_802
timestamp 1698175906
transform 1 0 91168 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_834
timestamp 1698175906
transform 1 0 94752 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_838
timestamp 1698175906
transform 1 0 95200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_842
timestamp 1698175906
transform 1 0 95648 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_858
timestamp 1698175906
transform 1 0 97440 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698175906
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698175906
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_37
timestamp 1698175906
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_101
timestamp 1698175906
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_107
timestamp 1698175906
transform 1 0 13328 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_171
timestamp 1698175906
transform 1 0 20496 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_177
timestamp 1698175906
transform 1 0 21168 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_185
timestamp 1698175906
transform 1 0 22064 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_189
timestamp 1698175906
transform 1 0 22512 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_191
timestamp 1698175906
transform 1 0 22736 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_221
timestamp 1698175906
transform 1 0 26096 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_225
timestamp 1698175906
transform 1 0 26544 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_247
timestamp 1698175906
transform 1 0 29008 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_269
timestamp 1698175906
transform 1 0 31472 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_273
timestamp 1698175906
transform 1 0 31920 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_277
timestamp 1698175906
transform 1 0 32368 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_291
timestamp 1698175906
transform 1 0 33936 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_295
timestamp 1698175906
transform 1 0 34384 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_303
timestamp 1698175906
transform 1 0 35280 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_309
timestamp 1698175906
transform 1 0 35952 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_313
timestamp 1698175906
transform 1 0 36400 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_317
timestamp 1698175906
transform 1 0 36848 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_325
timestamp 1698175906
transform 1 0 37744 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_329
timestamp 1698175906
transform 1 0 38192 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_381
timestamp 1698175906
transform 1 0 44016 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_387
timestamp 1698175906
transform 1 0 44688 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_417
timestamp 1698175906
transform 1 0 48048 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_421
timestamp 1698175906
transform 1 0 48496 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_425
timestamp 1698175906
transform 1 0 48944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_429
timestamp 1698175906
transform 1 0 49392 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_439
timestamp 1698175906
transform 1 0 50512 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_443
timestamp 1698175906
transform 1 0 50960 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_447
timestamp 1698175906
transform 1 0 51408 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_457
timestamp 1698175906
transform 1 0 52528 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_461
timestamp 1698175906
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_463
timestamp 1698175906
transform 1 0 53200 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_466
timestamp 1698175906
transform 1 0 53536 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_470
timestamp 1698175906
transform 1 0 53984 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_500
timestamp 1698175906
transform 1 0 57344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_513
timestamp 1698175906
transform 1 0 58800 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_521
timestamp 1698175906
transform 1 0 59696 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_556
timestamp 1698175906
transform 1 0 63616 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_560
timestamp 1698175906
transform 1 0 64064 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_580
timestamp 1698175906
transform 1 0 66304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_584
timestamp 1698175906
transform 1 0 66752 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_592
timestamp 1698175906
transform 1 0 67648 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_594
timestamp 1698175906
transform 1 0 67872 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_597
timestamp 1698175906
transform 1 0 68208 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_661
timestamp 1698175906
transform 1 0 75376 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_667
timestamp 1698175906
transform 1 0 76048 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_731
timestamp 1698175906
transform 1 0 83216 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_737
timestamp 1698175906
transform 1 0 83888 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_801
timestamp 1698175906
transform 1 0 91056 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_807
timestamp 1698175906
transform 1 0 91728 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_839
timestamp 1698175906
transform 1 0 95312 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_847
timestamp 1698175906
transform 1 0 96208 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_851
timestamp 1698175906
transform 1 0 96656 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_862
timestamp 1698175906
transform 1 0 97888 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_8
timestamp 1698175906
transform 1 0 2240 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_12
timestamp 1698175906
transform 1 0 2688 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_44
timestamp 1698175906
transform 1 0 6272 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_60
timestamp 1698175906
transform 1 0 8064 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_68
timestamp 1698175906
transform 1 0 8960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_72
timestamp 1698175906
transform 1 0 9408 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_136
timestamp 1698175906
transform 1 0 16576 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_142
timestamp 1698175906
transform 1 0 17248 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_206
timestamp 1698175906
transform 1 0 24416 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_212
timestamp 1698175906
transform 1 0 25088 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_228
timestamp 1698175906
transform 1 0 26880 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_232
timestamp 1698175906
transform 1 0 27328 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_250
timestamp 1698175906
transform 1 0 29344 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_261
timestamp 1698175906
transform 1 0 30576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_265
timestamp 1698175906
transform 1 0 31024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_269
timestamp 1698175906
transform 1 0 31472 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_277
timestamp 1698175906
transform 1 0 32368 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_279
timestamp 1698175906
transform 1 0 32592 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_282
timestamp 1698175906
transform 1 0 32928 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_286
timestamp 1698175906
transform 1 0 33376 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_312
timestamp 1698175906
transform 1 0 36288 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_316
timestamp 1698175906
transform 1 0 36736 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_320
timestamp 1698175906
transform 1 0 37184 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_328
timestamp 1698175906
transform 1 0 38080 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_330
timestamp 1698175906
transform 1 0 38304 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_333
timestamp 1698175906
transform 1 0 38640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_344
timestamp 1698175906
transform 1 0 39872 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_348
timestamp 1698175906
transform 1 0 40320 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_362
timestamp 1698175906
transform 1 0 41888 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_414
timestamp 1698175906
transform 1 0 47712 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_428
timestamp 1698175906
transform 1 0 49280 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_447
timestamp 1698175906
transform 1 0 51408 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_451
timestamp 1698175906
transform 1 0 51856 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_455
timestamp 1698175906
transform 1 0 52304 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_458
timestamp 1698175906
transform 1 0 52640 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_474
timestamp 1698175906
transform 1 0 54432 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_478
timestamp 1698175906
transform 1 0 54880 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_482
timestamp 1698175906
transform 1 0 55328 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_486
timestamp 1698175906
transform 1 0 55776 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_492
timestamp 1698175906
transform 1 0 56448 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_494
timestamp 1698175906
transform 1 0 56672 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_532
timestamp 1698175906
transform 1 0 60928 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_548
timestamp 1698175906
transform 1 0 62720 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_556
timestamp 1698175906
transform 1 0 63616 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_562
timestamp 1698175906
transform 1 0 64288 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_566
timestamp 1698175906
transform 1 0 64736 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_568
timestamp 1698175906
transform 1 0 64960 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_600
timestamp 1698175906
transform 1 0 68544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_604
timestamp 1698175906
transform 1 0 68992 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_620
timestamp 1698175906
transform 1 0 70784 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_628
timestamp 1698175906
transform 1 0 71680 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_632
timestamp 1698175906
transform 1 0 72128 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_696
timestamp 1698175906
transform 1 0 79296 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_702
timestamp 1698175906
transform 1 0 79968 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_766
timestamp 1698175906
transform 1 0 87136 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_772
timestamp 1698175906
transform 1 0 87808 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_836
timestamp 1698175906
transform 1 0 94976 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_842
timestamp 1698175906
transform 1 0 95648 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_858
timestamp 1698175906
transform 1 0 97440 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_8
timestamp 1698175906
transform 1 0 2240 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_12
timestamp 1698175906
transform 1 0 2688 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_28
timestamp 1698175906
transform 1 0 4480 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_32
timestamp 1698175906
transform 1 0 4928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698175906
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1698175906
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698175906
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_107
timestamp 1698175906
transform 1 0 13328 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_171
timestamp 1698175906
transform 1 0 20496 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_177
timestamp 1698175906
transform 1 0 21168 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_243
timestamp 1698175906
transform 1 0 28560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_247
timestamp 1698175906
transform 1 0 29008 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_259
timestamp 1698175906
transform 1 0 30352 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_265
timestamp 1698175906
transform 1 0 31024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_269
timestamp 1698175906
transform 1 0 31472 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_285
timestamp 1698175906
transform 1 0 33264 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_293
timestamp 1698175906
transform 1 0 34160 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_302
timestamp 1698175906
transform 1 0 35168 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_314
timestamp 1698175906
transform 1 0 36512 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_317
timestamp 1698175906
transform 1 0 36848 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_337
timestamp 1698175906
transform 1 0 39088 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_339
timestamp 1698175906
transform 1 0 39312 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_377
timestamp 1698175906
transform 1 0 43568 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_381
timestamp 1698175906
transform 1 0 44016 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_387
timestamp 1698175906
transform 1 0 44688 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_391
timestamp 1698175906
transform 1 0 45136 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_395
timestamp 1698175906
transform 1 0 45584 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_397
timestamp 1698175906
transform 1 0 45808 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_448
timestamp 1698175906
transform 1 0 51520 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_452
timestamp 1698175906
transform 1 0 51968 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_457
timestamp 1698175906
transform 1 0 52528 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_503
timestamp 1698175906
transform 1 0 57680 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_507
timestamp 1698175906
transform 1 0 58128 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_511
timestamp 1698175906
transform 1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_519
timestamp 1698175906
transform 1 0 59472 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_523
timestamp 1698175906
transform 1 0 59920 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_527
timestamp 1698175906
transform 1 0 60368 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_559
timestamp 1698175906
transform 1 0 63952 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_563
timestamp 1698175906
transform 1 0 64400 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_590
timestamp 1698175906
transform 1 0 67424 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_594
timestamp 1698175906
transform 1 0 67872 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_597
timestamp 1698175906
transform 1 0 68208 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_605
timestamp 1698175906
transform 1 0 69104 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_642
timestamp 1698175906
transform 1 0 73248 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_658
timestamp 1698175906
transform 1 0 75040 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_662
timestamp 1698175906
transform 1 0 75488 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_664
timestamp 1698175906
transform 1 0 75712 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_667
timestamp 1698175906
transform 1 0 76048 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_731
timestamp 1698175906
transform 1 0 83216 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_737
timestamp 1698175906
transform 1 0 83888 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_801
timestamp 1698175906
transform 1 0 91056 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_807
timestamp 1698175906
transform 1 0 91728 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_839
timestamp 1698175906
transform 1 0 95312 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_847
timestamp 1698175906
transform 1 0 96208 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_851
timestamp 1698175906
transform 1 0 96656 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_2
timestamp 1698175906
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_66
timestamp 1698175906
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_72
timestamp 1698175906
transform 1 0 9408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_136
timestamp 1698175906
transform 1 0 16576 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_142
timestamp 1698175906
transform 1 0 17248 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_206
timestamp 1698175906
transform 1 0 24416 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_212
timestamp 1698175906
transform 1 0 25088 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_276
timestamp 1698175906
transform 1 0 32256 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_282
timestamp 1698175906
transform 1 0 32928 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_298
timestamp 1698175906
transform 1 0 34720 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_304
timestamp 1698175906
transform 1 0 35392 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_314
timestamp 1698175906
transform 1 0 36512 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_318
timestamp 1698175906
transform 1 0 36960 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_334
timestamp 1698175906
transform 1 0 38752 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_342
timestamp 1698175906
transform 1 0 39648 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_360
timestamp 1698175906
transform 1 0 41664 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_364
timestamp 1698175906
transform 1 0 42112 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_368
timestamp 1698175906
transform 1 0 42560 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_370
timestamp 1698175906
transform 1 0 42784 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_392
timestamp 1698175906
transform 1 0 45248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_396
timestamp 1698175906
transform 1 0 45696 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_400
timestamp 1698175906
transform 1 0 46144 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_419
timestamp 1698175906
transform 1 0 48272 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_434
timestamp 1698175906
transform 1 0 49952 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_438
timestamp 1698175906
transform 1 0 50400 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_475
timestamp 1698175906
transform 1 0 54544 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_483
timestamp 1698175906
transform 1 0 55440 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_486
timestamp 1698175906
transform 1 0 55776 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_505
timestamp 1698175906
transform 1 0 57904 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_507
timestamp 1698175906
transform 1 0 58128 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_537
timestamp 1698175906
transform 1 0 61488 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_541
timestamp 1698175906
transform 1 0 61936 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_557
timestamp 1698175906
transform 1 0 63728 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_559
timestamp 1698175906
transform 1 0 63952 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_562
timestamp 1698175906
transform 1 0 64288 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_570
timestamp 1698175906
transform 1 0 65184 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_576
timestamp 1698175906
transform 1 0 65856 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_608
timestamp 1698175906
transform 1 0 69440 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_624
timestamp 1698175906
transform 1 0 71232 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_628
timestamp 1698175906
transform 1 0 71680 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_632
timestamp 1698175906
transform 1 0 72128 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_696
timestamp 1698175906
transform 1 0 79296 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_702
timestamp 1698175906
transform 1 0 79968 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_710
timestamp 1698175906
transform 1 0 80864 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_714
timestamp 1698175906
transform 1 0 81312 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_723
timestamp 1698175906
transform 1 0 82320 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_755
timestamp 1698175906
transform 1 0 85904 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_763
timestamp 1698175906
transform 1 0 86800 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_767
timestamp 1698175906
transform 1 0 87248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_769
timestamp 1698175906
transform 1 0 87472 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_772
timestamp 1698175906
transform 1 0 87808 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_836
timestamp 1698175906
transform 1 0 94976 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_842
timestamp 1698175906
transform 1 0 95648 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_858
timestamp 1698175906
transform 1 0 97440 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_8
timestamp 1698175906
transform 1 0 2240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_12
timestamp 1698175906
transform 1 0 2688 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_28
timestamp 1698175906
transform 1 0 4480 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_32
timestamp 1698175906
transform 1 0 4928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698175906
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_37
timestamp 1698175906
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_101
timestamp 1698175906
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_107
timestamp 1698175906
transform 1 0 13328 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_171
timestamp 1698175906
transform 1 0 20496 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_177
timestamp 1698175906
transform 1 0 21168 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_209
timestamp 1698175906
transform 1 0 24752 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_213
timestamp 1698175906
transform 1 0 25200 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_226
timestamp 1698175906
transform 1 0 26656 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_242
timestamp 1698175906
transform 1 0 28448 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_244
timestamp 1698175906
transform 1 0 28672 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_282
timestamp 1698175906
transform 1 0 32928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_317
timestamp 1698175906
transform 1 0 36848 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_321
timestamp 1698175906
transform 1 0 37296 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_337
timestamp 1698175906
transform 1 0 39088 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_376
timestamp 1698175906
transform 1 0 43456 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_380
timestamp 1698175906
transform 1 0 43904 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_382
timestamp 1698175906
transform 1 0 44128 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_387
timestamp 1698175906
transform 1 0 44688 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_389
timestamp 1698175906
transform 1 0 44912 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_419
timestamp 1698175906
transform 1 0 48272 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_423
timestamp 1698175906
transform 1 0 48720 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_439
timestamp 1698175906
transform 1 0 50512 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_447
timestamp 1698175906
transform 1 0 51408 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_451
timestamp 1698175906
transform 1 0 51856 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_465
timestamp 1698175906
transform 1 0 53424 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_481
timestamp 1698175906
transform 1 0 55216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_483
timestamp 1698175906
transform 1 0 55440 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_490
timestamp 1698175906
transform 1 0 56224 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_512
timestamp 1698175906
transform 1 0 58688 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_520
timestamp 1698175906
transform 1 0 59584 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_524
timestamp 1698175906
transform 1 0 60032 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_527
timestamp 1698175906
transform 1 0 60368 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_559
timestamp 1698175906
transform 1 0 63952 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_575
timestamp 1698175906
transform 1 0 65744 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_589
timestamp 1698175906
transform 1 0 67312 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_593
timestamp 1698175906
transform 1 0 67760 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_603
timestamp 1698175906
transform 1 0 68880 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_635
timestamp 1698175906
transform 1 0 72464 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_651
timestamp 1698175906
transform 1 0 74256 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_659
timestamp 1698175906
transform 1 0 75152 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_663
timestamp 1698175906
transform 1 0 75600 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_667
timestamp 1698175906
transform 1 0 76048 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_731
timestamp 1698175906
transform 1 0 83216 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_737
timestamp 1698175906
transform 1 0 83888 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_801
timestamp 1698175906
transform 1 0 91056 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_807
timestamp 1698175906
transform 1 0 91728 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_839
timestamp 1698175906
transform 1 0 95312 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_847
timestamp 1698175906
transform 1 0 96208 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_849
timestamp 1698175906
transform 1 0 96432 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_8
timestamp 1698175906
transform 1 0 2240 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_12
timestamp 1698175906
transform 1 0 2688 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_28
timestamp 1698175906
transform 1 0 4480 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_32
timestamp 1698175906
transform 1 0 4928 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_36
timestamp 1698175906
transform 1 0 5376 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_44
timestamp 1698175906
transform 1 0 6272 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_48
timestamp 1698175906
transform 1 0 6720 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_63
timestamp 1698175906
transform 1 0 8400 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_67
timestamp 1698175906
transform 1 0 8848 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_70
timestamp 1698175906
transform 1 0 9184 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_104
timestamp 1698175906
transform 1 0 12992 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_138
timestamp 1698175906
transform 1 0 16800 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_154
timestamp 1698175906
transform 1 0 18592 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_172
timestamp 1698175906
transform 1 0 20608 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_206
timestamp 1698175906
transform 1 0 24416 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_240
timestamp 1698175906
transform 1 0 28224 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_284
timestamp 1698175906
transform 1 0 33152 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_300
timestamp 1698175906
transform 1 0 34944 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_304
timestamp 1698175906
transform 1 0 35392 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_308
timestamp 1698175906
transform 1 0 35840 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_342
timestamp 1698175906
transform 1 0 39648 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_376
timestamp 1698175906
transform 1 0 43456 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_378
timestamp 1698175906
transform 1 0 43680 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_389
timestamp 1698175906
transform 1 0 44912 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_405
timestamp 1698175906
transform 1 0 46704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_407
timestamp 1698175906
transform 1 0 46928 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_410
timestamp 1698175906
transform 1 0 47264 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_444
timestamp 1698175906
transform 1 0 51072 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_478
timestamp 1698175906
transform 1 0 54880 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_486
timestamp 1698175906
transform 1 0 55776 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_488
timestamp 1698175906
transform 1 0 56000 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_499
timestamp 1698175906
transform 1 0 57232 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_507
timestamp 1698175906
transform 1 0 58128 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_509
timestamp 1698175906
transform 1 0 58352 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_512
timestamp 1698175906
transform 1 0 58688 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_546
timestamp 1698175906
transform 1 0 62496 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_580
timestamp 1698175906
transform 1 0 66304 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_596
timestamp 1698175906
transform 1 0 68096 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_608
timestamp 1698175906
transform 1 0 69440 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_614
timestamp 1698175906
transform 1 0 70112 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_648
timestamp 1698175906
transform 1 0 73920 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_682
timestamp 1698175906
transform 1 0 77728 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_726
timestamp 1698175906
transform 1 0 82656 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_742
timestamp 1698175906
transform 1 0 84448 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_746
timestamp 1698175906
transform 1 0 84896 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_750
timestamp 1698175906
transform 1 0 85344 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_784
timestamp 1698175906
transform 1 0 89152 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_818
timestamp 1698175906
transform 1 0 92960 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_829
timestamp 1698175906
transform 1 0 94192 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_837
timestamp 1698175906
transform 1 0 95088 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_839
timestamp 1698175906
transform 1 0 95312 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_862
timestamp 1698175906
transform 1 0 97888 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698175906
transform -1 0 94640 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  input2
timestamp 1698175906
transform -1 0 86464 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input3
timestamp 1698175906
transform -1 0 74704 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input4
timestamp 1698175906
transform 1 0 61040 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input5
timestamp 1698175906
transform 1 0 54880 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input6
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input7
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input8
timestamp 1698175906
transform 1 0 17136 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input10 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input12
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698175906
transform -1 0 2912 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input17 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698175906
transform 1 0 1568 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698175906
transform 1 0 1568 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698175906
transform 1 0 1568 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698175906
transform 1 0 1568 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698175906
transform 1 0 2240 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698175906
transform 1 0 1568 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698175906
transform 1 0 1568 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698175906
transform 1 0 1568 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698175906
transform -1 0 2912 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698175906
transform 1 0 2240 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698175906
transform 1 0 1568 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698175906
transform 1 0 1568 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698175906
transform 1 0 1568 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1698175906
transform 1 0 1568 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698175906
transform 1 0 2240 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698175906
transform 1 0 1568 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698175906
transform 1 0 1568 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1698175906
transform 1 0 1568 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input50
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1698175906
transform 1 0 6160 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  net299_2
timestamp 1698175906
transform 1 0 78176 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output52
timestamp 1698175906
transform 1 0 96768 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output53
timestamp 1698175906
transform -1 0 96544 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output54
timestamp 1698175906
transform 1 0 96768 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output55
timestamp 1698175906
transform 1 0 96768 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output56
timestamp 1698175906
transform 1 0 96768 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output57
timestamp 1698175906
transform 1 0 96768 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output58
timestamp 1698175906
transform 1 0 96768 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output59
timestamp 1698175906
transform 1 0 96768 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output60
timestamp 1698175906
transform 1 0 96768 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output61
timestamp 1698175906
transform 1 0 96768 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output62
timestamp 1698175906
transform 1 0 96768 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output63
timestamp 1698175906
transform 1 0 96768 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output64
timestamp 1698175906
transform 1 0 96768 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output65
timestamp 1698175906
transform 1 0 96768 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output66
timestamp 1698175906
transform 1 0 96768 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output67
timestamp 1698175906
transform 1 0 96768 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output68
timestamp 1698175906
transform 1 0 96768 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output69
timestamp 1698175906
transform 1 0 96768 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output70
timestamp 1698175906
transform 1 0 96768 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output71
timestamp 1698175906
transform 1 0 96768 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output72
timestamp 1698175906
transform 1 0 96768 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output73
timestamp 1698175906
transform 1 0 96768 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output74
timestamp 1698175906
transform 1 0 96768 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output75
timestamp 1698175906
transform 1 0 96768 0 1 53312
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output76
timestamp 1698175906
transform 1 0 96768 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output77
timestamp 1698175906
transform 1 0 96768 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output78
timestamp 1698175906
transform 1 0 96768 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output79
timestamp 1698175906
transform 1 0 96768 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output80
timestamp 1698175906
transform 1 0 96768 0 -1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output81
timestamp 1698175906
transform 1 0 96768 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output82
timestamp 1698175906
transform 1 0 96768 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output83
timestamp 1698175906
transform 1 0 96768 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output84
timestamp 1698175906
transform 1 0 96768 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output85
timestamp 1698175906
transform 1 0 93072 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output86
timestamp 1698175906
transform 1 0 81536 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output87
timestamp 1698175906
transform 1 0 68320 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output88
timestamp 1698175906
transform 1 0 56112 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output89
timestamp 1698175906
transform 1 0 43792 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output90
timestamp 1698175906
transform -1 0 33152 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output91 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 20384 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output92
timestamp 1698175906
transform -1 0 8400 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 98560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 98560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 98560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 98560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 98560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 98560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 98560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 98560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 98560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 98560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 98560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 98560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 98560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 98560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 98560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 98560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 98560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 98560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 98560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 98560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 98560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 98560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 98560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 98560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 98560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 98560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 98560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 98560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 98560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 98560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 98560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 98560 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 98560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 98560 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 98560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 98560 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 98560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 98560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 98560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 98560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 98560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 98560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 98560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 98560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 98560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698175906
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698175906
transform -1 0 98560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698175906
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698175906
transform -1 0 98560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698175906
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698175906
transform -1 0 98560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698175906
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698175906
transform -1 0 98560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698175906
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698175906
transform -1 0 98560 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698175906
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698175906
transform -1 0 98560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698175906
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698175906
transform -1 0 98560 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698175906
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698175906
transform -1 0 98560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698175906
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698175906
transform -1 0 98560 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698175906
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698175906
transform -1 0 98560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698175906
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698175906
transform -1 0 98560 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698175906
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698175906
transform -1 0 98560 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698175906
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698175906
transform -1 0 98560 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698175906
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698175906
transform -1 0 98560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698175906
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698175906
transform -1 0 98560 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698175906
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698175906
transform -1 0 98560 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698175906
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698175906
transform -1 0 98560 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698175906
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698175906
transform -1 0 98560 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698175906
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698175906
transform -1 0 98560 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698175906
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698175906
transform -1 0 98560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698175906
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698175906
transform -1 0 98560 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698175906
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698175906
transform -1 0 98560 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698175906
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698175906
transform -1 0 98560 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698175906
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698175906
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698175906
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698175906
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_150
timestamp 1698175906
transform 1 0 58464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_151
timestamp 1698175906
transform 1 0 62272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_152
timestamp 1698175906
transform 1 0 66080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_153
timestamp 1698175906
transform 1 0 69888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_154
timestamp 1698175906
transform 1 0 73696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_155
timestamp 1698175906
transform 1 0 77504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_156
timestamp 1698175906
transform 1 0 81312 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_157
timestamp 1698175906
transform 1 0 85120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_158
timestamp 1698175906
transform 1 0 88928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_159
timestamp 1698175906
transform 1 0 92736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_160
timestamp 1698175906
transform 1 0 96544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_161
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_162
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_163
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_164
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_165
timestamp 1698175906
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_166
timestamp 1698175906
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_167
timestamp 1698175906
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_168
timestamp 1698175906
transform 1 0 64064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_169
timestamp 1698175906
transform 1 0 71904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_170
timestamp 1698175906
transform 1 0 79744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_171
timestamp 1698175906
transform 1 0 87584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_172
timestamp 1698175906
transform 1 0 95424 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_173
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_174
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_175
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_176
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_177
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_178
timestamp 1698175906
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_179
timestamp 1698175906
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_180
timestamp 1698175906
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_181
timestamp 1698175906
transform 1 0 67984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_182
timestamp 1698175906
transform 1 0 75824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_183
timestamp 1698175906
transform 1 0 83664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_184
timestamp 1698175906
transform 1 0 91504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_185
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_186
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_187
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_188
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_189
timestamp 1698175906
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_190
timestamp 1698175906
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_191
timestamp 1698175906
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_192
timestamp 1698175906
transform 1 0 64064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_193
timestamp 1698175906
transform 1 0 71904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_194
timestamp 1698175906
transform 1 0 79744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_195
timestamp 1698175906
transform 1 0 87584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_196
timestamp 1698175906
transform 1 0 95424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_197
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_198
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_199
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_200
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_201
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_202
timestamp 1698175906
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_203
timestamp 1698175906
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_204
timestamp 1698175906
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_205
timestamp 1698175906
transform 1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_206
timestamp 1698175906
transform 1 0 75824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_207
timestamp 1698175906
transform 1 0 83664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_208
timestamp 1698175906
transform 1 0 91504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_209
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_210
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_211
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_212
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_213
timestamp 1698175906
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_214
timestamp 1698175906
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_215
timestamp 1698175906
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_216
timestamp 1698175906
transform 1 0 64064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_217
timestamp 1698175906
transform 1 0 71904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_218
timestamp 1698175906
transform 1 0 79744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_219
timestamp 1698175906
transform 1 0 87584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_220
timestamp 1698175906
transform 1 0 95424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_221
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_222
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_223
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_224
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_225
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_226
timestamp 1698175906
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_227
timestamp 1698175906
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_228
timestamp 1698175906
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_229
timestamp 1698175906
transform 1 0 67984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_230
timestamp 1698175906
transform 1 0 75824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_231
timestamp 1698175906
transform 1 0 83664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_232
timestamp 1698175906
transform 1 0 91504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_233
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_234
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_235
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_236
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_237
timestamp 1698175906
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_238
timestamp 1698175906
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_239
timestamp 1698175906
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_240
timestamp 1698175906
transform 1 0 64064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_241
timestamp 1698175906
transform 1 0 71904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_242
timestamp 1698175906
transform 1 0 79744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_243
timestamp 1698175906
transform 1 0 87584 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_244
timestamp 1698175906
transform 1 0 95424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_245
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_246
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_247
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_248
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_249
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_250
timestamp 1698175906
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_251
timestamp 1698175906
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_252
timestamp 1698175906
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_253
timestamp 1698175906
transform 1 0 67984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_254
timestamp 1698175906
transform 1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_255
timestamp 1698175906
transform 1 0 83664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_256
timestamp 1698175906
transform 1 0 91504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_257
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_258
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_259
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_260
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_261
timestamp 1698175906
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_262
timestamp 1698175906
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_263
timestamp 1698175906
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_264
timestamp 1698175906
transform 1 0 64064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_265
timestamp 1698175906
transform 1 0 71904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_266
timestamp 1698175906
transform 1 0 79744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_267
timestamp 1698175906
transform 1 0 87584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_268
timestamp 1698175906
transform 1 0 95424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_269
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_270
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_271
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_272
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_273
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_274
timestamp 1698175906
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_275
timestamp 1698175906
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_276
timestamp 1698175906
transform 1 0 60144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_277
timestamp 1698175906
transform 1 0 67984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_278
timestamp 1698175906
transform 1 0 75824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_279
timestamp 1698175906
transform 1 0 83664 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_280
timestamp 1698175906
transform 1 0 91504 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_281
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_282
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_283
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_284
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_285
timestamp 1698175906
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_286
timestamp 1698175906
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_287
timestamp 1698175906
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_288
timestamp 1698175906
transform 1 0 64064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_289
timestamp 1698175906
transform 1 0 71904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_290
timestamp 1698175906
transform 1 0 79744 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_291
timestamp 1698175906
transform 1 0 87584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_292
timestamp 1698175906
transform 1 0 95424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_293
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_294
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_295
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_296
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_297
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_298
timestamp 1698175906
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_299
timestamp 1698175906
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_300
timestamp 1698175906
transform 1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_301
timestamp 1698175906
transform 1 0 67984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_302
timestamp 1698175906
transform 1 0 75824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_303
timestamp 1698175906
transform 1 0 83664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_304
timestamp 1698175906
transform 1 0 91504 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_305
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_306
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_307
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_308
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_309
timestamp 1698175906
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_310
timestamp 1698175906
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_311
timestamp 1698175906
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_312
timestamp 1698175906
transform 1 0 64064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_313
timestamp 1698175906
transform 1 0 71904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_314
timestamp 1698175906
transform 1 0 79744 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_315
timestamp 1698175906
transform 1 0 87584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_316
timestamp 1698175906
transform 1 0 95424 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_317
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_318
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_319
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_320
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_321
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_322
timestamp 1698175906
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_323
timestamp 1698175906
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_324
timestamp 1698175906
transform 1 0 60144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_325
timestamp 1698175906
transform 1 0 67984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_326
timestamp 1698175906
transform 1 0 75824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_327
timestamp 1698175906
transform 1 0 83664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_328
timestamp 1698175906
transform 1 0 91504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_329
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_330
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_331
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_332
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_333
timestamp 1698175906
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_334
timestamp 1698175906
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_335
timestamp 1698175906
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_336
timestamp 1698175906
transform 1 0 64064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_337
timestamp 1698175906
transform 1 0 71904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_338
timestamp 1698175906
transform 1 0 79744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_339
timestamp 1698175906
transform 1 0 87584 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_340
timestamp 1698175906
transform 1 0 95424 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_341
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_342
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_343
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_344
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_345
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_346
timestamp 1698175906
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_347
timestamp 1698175906
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_348
timestamp 1698175906
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_349
timestamp 1698175906
transform 1 0 67984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_350
timestamp 1698175906
transform 1 0 75824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_351
timestamp 1698175906
transform 1 0 83664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_352
timestamp 1698175906
transform 1 0 91504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_353
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_354
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_355
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_356
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_357
timestamp 1698175906
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_358
timestamp 1698175906
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_359
timestamp 1698175906
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_360
timestamp 1698175906
transform 1 0 64064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_361
timestamp 1698175906
transform 1 0 71904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_362
timestamp 1698175906
transform 1 0 79744 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_363
timestamp 1698175906
transform 1 0 87584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_364
timestamp 1698175906
transform 1 0 95424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_365
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_366
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_367
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_368
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_369
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_370
timestamp 1698175906
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_371
timestamp 1698175906
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_372
timestamp 1698175906
transform 1 0 60144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_373
timestamp 1698175906
transform 1 0 67984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_374
timestamp 1698175906
transform 1 0 75824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_375
timestamp 1698175906
transform 1 0 83664 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_376
timestamp 1698175906
transform 1 0 91504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_377
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_378
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_379
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_380
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_381
timestamp 1698175906
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_382
timestamp 1698175906
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_383
timestamp 1698175906
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_384
timestamp 1698175906
transform 1 0 64064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_385
timestamp 1698175906
transform 1 0 71904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_386
timestamp 1698175906
transform 1 0 79744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_387
timestamp 1698175906
transform 1 0 87584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_388
timestamp 1698175906
transform 1 0 95424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_389
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_390
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_391
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_392
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_393
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_394
timestamp 1698175906
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_395
timestamp 1698175906
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_396
timestamp 1698175906
transform 1 0 60144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_397
timestamp 1698175906
transform 1 0 67984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_398
timestamp 1698175906
transform 1 0 75824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_399
timestamp 1698175906
transform 1 0 83664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_400
timestamp 1698175906
transform 1 0 91504 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_401
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_402
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_403
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_404
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_405
timestamp 1698175906
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_406
timestamp 1698175906
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_407
timestamp 1698175906
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_408
timestamp 1698175906
transform 1 0 64064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_409
timestamp 1698175906
transform 1 0 71904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_410
timestamp 1698175906
transform 1 0 79744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_411
timestamp 1698175906
transform 1 0 87584 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_412
timestamp 1698175906
transform 1 0 95424 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_413
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_414
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_415
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_416
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_417
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_418
timestamp 1698175906
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_419
timestamp 1698175906
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_420
timestamp 1698175906
transform 1 0 60144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_421
timestamp 1698175906
transform 1 0 67984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_422
timestamp 1698175906
transform 1 0 75824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_423
timestamp 1698175906
transform 1 0 83664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_424
timestamp 1698175906
transform 1 0 91504 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_425
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_426
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_427
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_428
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_429
timestamp 1698175906
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_430
timestamp 1698175906
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_431
timestamp 1698175906
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_432
timestamp 1698175906
transform 1 0 64064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_433
timestamp 1698175906
transform 1 0 71904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_434
timestamp 1698175906
transform 1 0 79744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_435
timestamp 1698175906
transform 1 0 87584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_436
timestamp 1698175906
transform 1 0 95424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_437
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_438
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_439
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_440
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_441
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_442
timestamp 1698175906
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_443
timestamp 1698175906
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_444
timestamp 1698175906
transform 1 0 60144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_445
timestamp 1698175906
transform 1 0 67984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_446
timestamp 1698175906
transform 1 0 75824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_447
timestamp 1698175906
transform 1 0 83664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_448
timestamp 1698175906
transform 1 0 91504 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_449
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_450
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_451
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_452
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_453
timestamp 1698175906
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_454
timestamp 1698175906
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_455
timestamp 1698175906
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_456
timestamp 1698175906
transform 1 0 64064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_457
timestamp 1698175906
transform 1 0 71904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_458
timestamp 1698175906
transform 1 0 79744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_459
timestamp 1698175906
transform 1 0 87584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_460
timestamp 1698175906
transform 1 0 95424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_461
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_462
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_463
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_464
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_465
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_466
timestamp 1698175906
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_467
timestamp 1698175906
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_468
timestamp 1698175906
transform 1 0 60144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_469
timestamp 1698175906
transform 1 0 67984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_470
timestamp 1698175906
transform 1 0 75824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_471
timestamp 1698175906
transform 1 0 83664 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_472
timestamp 1698175906
transform 1 0 91504 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_473
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_474
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_475
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_476
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_477
timestamp 1698175906
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_478
timestamp 1698175906
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_479
timestamp 1698175906
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_480
timestamp 1698175906
transform 1 0 64064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_481
timestamp 1698175906
transform 1 0 71904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_482
timestamp 1698175906
transform 1 0 79744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_483
timestamp 1698175906
transform 1 0 87584 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_484
timestamp 1698175906
transform 1 0 95424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_485
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_486
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_487
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_488
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_489
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_490
timestamp 1698175906
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_491
timestamp 1698175906
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_492
timestamp 1698175906
transform 1 0 60144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_493
timestamp 1698175906
transform 1 0 67984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_494
timestamp 1698175906
transform 1 0 75824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_495
timestamp 1698175906
transform 1 0 83664 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_496
timestamp 1698175906
transform 1 0 91504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_497
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_498
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_499
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_500
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_501
timestamp 1698175906
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_502
timestamp 1698175906
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_503
timestamp 1698175906
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_504
timestamp 1698175906
transform 1 0 64064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_505
timestamp 1698175906
transform 1 0 71904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_506
timestamp 1698175906
transform 1 0 79744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_507
timestamp 1698175906
transform 1 0 87584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_508
timestamp 1698175906
transform 1 0 95424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_509
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_510
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_511
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_512
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_513
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_514
timestamp 1698175906
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_515
timestamp 1698175906
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_516
timestamp 1698175906
transform 1 0 60144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_517
timestamp 1698175906
transform 1 0 67984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_518
timestamp 1698175906
transform 1 0 75824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_519
timestamp 1698175906
transform 1 0 83664 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_520
timestamp 1698175906
transform 1 0 91504 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_521
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_522
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_523
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_524
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_525
timestamp 1698175906
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_526
timestamp 1698175906
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_527
timestamp 1698175906
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_528
timestamp 1698175906
transform 1 0 64064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_529
timestamp 1698175906
transform 1 0 71904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_530
timestamp 1698175906
transform 1 0 79744 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_531
timestamp 1698175906
transform 1 0 87584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_532
timestamp 1698175906
transform 1 0 95424 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_533
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_534
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_535
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_536
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_537
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_538
timestamp 1698175906
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_539
timestamp 1698175906
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_540
timestamp 1698175906
transform 1 0 60144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_541
timestamp 1698175906
transform 1 0 67984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_542
timestamp 1698175906
transform 1 0 75824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_543
timestamp 1698175906
transform 1 0 83664 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_544
timestamp 1698175906
transform 1 0 91504 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_545
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_546
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_547
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_548
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_549
timestamp 1698175906
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_550
timestamp 1698175906
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_551
timestamp 1698175906
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_552
timestamp 1698175906
transform 1 0 64064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_553
timestamp 1698175906
transform 1 0 71904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_554
timestamp 1698175906
transform 1 0 79744 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_555
timestamp 1698175906
transform 1 0 87584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_556
timestamp 1698175906
transform 1 0 95424 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_557
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_558
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_559
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_560
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_561
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_562
timestamp 1698175906
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_563
timestamp 1698175906
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_564
timestamp 1698175906
transform 1 0 60144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_565
timestamp 1698175906
transform 1 0 67984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_566
timestamp 1698175906
transform 1 0 75824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_567
timestamp 1698175906
transform 1 0 83664 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_568
timestamp 1698175906
transform 1 0 91504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_569
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_570
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_571
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_572
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_573
timestamp 1698175906
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_574
timestamp 1698175906
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_575
timestamp 1698175906
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_576
timestamp 1698175906
transform 1 0 64064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_577
timestamp 1698175906
transform 1 0 71904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_578
timestamp 1698175906
transform 1 0 79744 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_579
timestamp 1698175906
transform 1 0 87584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_580
timestamp 1698175906
transform 1 0 95424 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_581
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_582
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_583
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_584
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_585
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_586
timestamp 1698175906
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_587
timestamp 1698175906
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_588
timestamp 1698175906
transform 1 0 60144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_589
timestamp 1698175906
transform 1 0 67984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_590
timestamp 1698175906
transform 1 0 75824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_591
timestamp 1698175906
transform 1 0 83664 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_592
timestamp 1698175906
transform 1 0 91504 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_593
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_594
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_595
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_596
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_597
timestamp 1698175906
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_598
timestamp 1698175906
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_599
timestamp 1698175906
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_600
timestamp 1698175906
transform 1 0 64064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_601
timestamp 1698175906
transform 1 0 71904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_602
timestamp 1698175906
transform 1 0 79744 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_603
timestamp 1698175906
transform 1 0 87584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_604
timestamp 1698175906
transform 1 0 95424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_605
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_606
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_607
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_608
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_609
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_610
timestamp 1698175906
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_611
timestamp 1698175906
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_612
timestamp 1698175906
transform 1 0 60144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_613
timestamp 1698175906
transform 1 0 67984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_614
timestamp 1698175906
transform 1 0 75824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_615
timestamp 1698175906
transform 1 0 83664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_616
timestamp 1698175906
transform 1 0 91504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_617
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_618
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_619
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_620
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_621
timestamp 1698175906
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_622
timestamp 1698175906
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_623
timestamp 1698175906
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_624
timestamp 1698175906
transform 1 0 64064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_625
timestamp 1698175906
transform 1 0 71904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_626
timestamp 1698175906
transform 1 0 79744 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_627
timestamp 1698175906
transform 1 0 87584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_628
timestamp 1698175906
transform 1 0 95424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_629
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_630
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_631
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_632
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_633
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_634
timestamp 1698175906
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_635
timestamp 1698175906
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_636
timestamp 1698175906
transform 1 0 60144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_637
timestamp 1698175906
transform 1 0 67984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_638
timestamp 1698175906
transform 1 0 75824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_639
timestamp 1698175906
transform 1 0 83664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_640
timestamp 1698175906
transform 1 0 91504 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_641
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_642
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_643
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_644
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_645
timestamp 1698175906
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_646
timestamp 1698175906
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_647
timestamp 1698175906
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_648
timestamp 1698175906
transform 1 0 64064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_649
timestamp 1698175906
transform 1 0 71904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_650
timestamp 1698175906
transform 1 0 79744 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_651
timestamp 1698175906
transform 1 0 87584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_652
timestamp 1698175906
transform 1 0 95424 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_653
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_654
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_655
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_656
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_657
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_658
timestamp 1698175906
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_659
timestamp 1698175906
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_660
timestamp 1698175906
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_661
timestamp 1698175906
transform 1 0 67984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_662
timestamp 1698175906
transform 1 0 75824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_663
timestamp 1698175906
transform 1 0 83664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_664
timestamp 1698175906
transform 1 0 91504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_665
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_666
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_667
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_668
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_669
timestamp 1698175906
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_670
timestamp 1698175906
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_671
timestamp 1698175906
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_672
timestamp 1698175906
transform 1 0 64064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_673
timestamp 1698175906
transform 1 0 71904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_674
timestamp 1698175906
transform 1 0 79744 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_675
timestamp 1698175906
transform 1 0 87584 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_676
timestamp 1698175906
transform 1 0 95424 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_677
timestamp 1698175906
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_678
timestamp 1698175906
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_679
timestamp 1698175906
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_680
timestamp 1698175906
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_681
timestamp 1698175906
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_682
timestamp 1698175906
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_683
timestamp 1698175906
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_684
timestamp 1698175906
transform 1 0 60144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_685
timestamp 1698175906
transform 1 0 67984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_686
timestamp 1698175906
transform 1 0 75824 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_687
timestamp 1698175906
transform 1 0 83664 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_688
timestamp 1698175906
transform 1 0 91504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_689
timestamp 1698175906
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_690
timestamp 1698175906
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_691
timestamp 1698175906
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_692
timestamp 1698175906
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_693
timestamp 1698175906
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_694
timestamp 1698175906
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_695
timestamp 1698175906
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_696
timestamp 1698175906
transform 1 0 64064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_697
timestamp 1698175906
transform 1 0 71904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_698
timestamp 1698175906
transform 1 0 79744 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_699
timestamp 1698175906
transform 1 0 87584 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_700
timestamp 1698175906
transform 1 0 95424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_701
timestamp 1698175906
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_702
timestamp 1698175906
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_703
timestamp 1698175906
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_704
timestamp 1698175906
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_705
timestamp 1698175906
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_706
timestamp 1698175906
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_707
timestamp 1698175906
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_708
timestamp 1698175906
transform 1 0 60144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_709
timestamp 1698175906
transform 1 0 67984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_710
timestamp 1698175906
transform 1 0 75824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_711
timestamp 1698175906
transform 1 0 83664 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_712
timestamp 1698175906
transform 1 0 91504 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_713
timestamp 1698175906
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_714
timestamp 1698175906
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_715
timestamp 1698175906
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_716
timestamp 1698175906
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_717
timestamp 1698175906
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_718
timestamp 1698175906
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_719
timestamp 1698175906
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_720
timestamp 1698175906
transform 1 0 64064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_721
timestamp 1698175906
transform 1 0 71904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_722
timestamp 1698175906
transform 1 0 79744 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_723
timestamp 1698175906
transform 1 0 87584 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_724
timestamp 1698175906
transform 1 0 95424 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_725
timestamp 1698175906
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_726
timestamp 1698175906
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_727
timestamp 1698175906
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_728
timestamp 1698175906
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_729
timestamp 1698175906
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_730
timestamp 1698175906
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_731
timestamp 1698175906
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_732
timestamp 1698175906
transform 1 0 60144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_733
timestamp 1698175906
transform 1 0 67984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_734
timestamp 1698175906
transform 1 0 75824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_735
timestamp 1698175906
transform 1 0 83664 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_736
timestamp 1698175906
transform 1 0 91504 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_737
timestamp 1698175906
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_738
timestamp 1698175906
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_739
timestamp 1698175906
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_740
timestamp 1698175906
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_741
timestamp 1698175906
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_742
timestamp 1698175906
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_743
timestamp 1698175906
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_744
timestamp 1698175906
transform 1 0 64064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_745
timestamp 1698175906
transform 1 0 71904 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_746
timestamp 1698175906
transform 1 0 79744 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_747
timestamp 1698175906
transform 1 0 87584 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_748
timestamp 1698175906
transform 1 0 95424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_749
timestamp 1698175906
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_750
timestamp 1698175906
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_751
timestamp 1698175906
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_752
timestamp 1698175906
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_753
timestamp 1698175906
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_754
timestamp 1698175906
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_755
timestamp 1698175906
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_756
timestamp 1698175906
transform 1 0 60144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_757
timestamp 1698175906
transform 1 0 67984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_758
timestamp 1698175906
transform 1 0 75824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_759
timestamp 1698175906
transform 1 0 83664 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_760
timestamp 1698175906
transform 1 0 91504 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_761
timestamp 1698175906
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_762
timestamp 1698175906
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_763
timestamp 1698175906
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_764
timestamp 1698175906
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_765
timestamp 1698175906
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_766
timestamp 1698175906
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_767
timestamp 1698175906
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_768
timestamp 1698175906
transform 1 0 64064 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_769
timestamp 1698175906
transform 1 0 71904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_770
timestamp 1698175906
transform 1 0 79744 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_771
timestamp 1698175906
transform 1 0 87584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_772
timestamp 1698175906
transform 1 0 95424 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_773
timestamp 1698175906
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_774
timestamp 1698175906
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_775
timestamp 1698175906
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_776
timestamp 1698175906
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_777
timestamp 1698175906
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_778
timestamp 1698175906
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_779
timestamp 1698175906
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_780
timestamp 1698175906
transform 1 0 60144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_781
timestamp 1698175906
transform 1 0 67984 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_782
timestamp 1698175906
transform 1 0 75824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_783
timestamp 1698175906
transform 1 0 83664 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_784
timestamp 1698175906
transform 1 0 91504 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_785
timestamp 1698175906
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_786
timestamp 1698175906
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_787
timestamp 1698175906
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_788
timestamp 1698175906
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_789
timestamp 1698175906
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_790
timestamp 1698175906
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_791
timestamp 1698175906
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_792
timestamp 1698175906
transform 1 0 64064 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_793
timestamp 1698175906
transform 1 0 71904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_794
timestamp 1698175906
transform 1 0 79744 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_795
timestamp 1698175906
transform 1 0 87584 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_796
timestamp 1698175906
transform 1 0 95424 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_797
timestamp 1698175906
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_798
timestamp 1698175906
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_799
timestamp 1698175906
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_800
timestamp 1698175906
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_801
timestamp 1698175906
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_802
timestamp 1698175906
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_803
timestamp 1698175906
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_804
timestamp 1698175906
transform 1 0 60144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_805
timestamp 1698175906
transform 1 0 67984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_806
timestamp 1698175906
transform 1 0 75824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_807
timestamp 1698175906
transform 1 0 83664 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_808
timestamp 1698175906
transform 1 0 91504 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_809
timestamp 1698175906
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_810
timestamp 1698175906
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_811
timestamp 1698175906
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_812
timestamp 1698175906
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_813
timestamp 1698175906
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_814
timestamp 1698175906
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_815
timestamp 1698175906
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_816
timestamp 1698175906
transform 1 0 64064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_817
timestamp 1698175906
transform 1 0 71904 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_818
timestamp 1698175906
transform 1 0 79744 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_819
timestamp 1698175906
transform 1 0 87584 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_820
timestamp 1698175906
transform 1 0 95424 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_821
timestamp 1698175906
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_822
timestamp 1698175906
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_823
timestamp 1698175906
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_824
timestamp 1698175906
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_825
timestamp 1698175906
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_826
timestamp 1698175906
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_827
timestamp 1698175906
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_828
timestamp 1698175906
transform 1 0 60144 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_829
timestamp 1698175906
transform 1 0 67984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_830
timestamp 1698175906
transform 1 0 75824 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_831
timestamp 1698175906
transform 1 0 83664 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_832
timestamp 1698175906
transform 1 0 91504 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_833
timestamp 1698175906
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_834
timestamp 1698175906
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_835
timestamp 1698175906
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_836
timestamp 1698175906
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_837
timestamp 1698175906
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_838
timestamp 1698175906
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_839
timestamp 1698175906
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_840
timestamp 1698175906
transform 1 0 64064 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_841
timestamp 1698175906
transform 1 0 71904 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_842
timestamp 1698175906
transform 1 0 79744 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_843
timestamp 1698175906
transform 1 0 87584 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_844
timestamp 1698175906
transform 1 0 95424 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_845
timestamp 1698175906
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_846
timestamp 1698175906
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_847
timestamp 1698175906
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_848
timestamp 1698175906
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_849
timestamp 1698175906
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_850
timestamp 1698175906
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_851
timestamp 1698175906
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_852
timestamp 1698175906
transform 1 0 60144 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_853
timestamp 1698175906
transform 1 0 67984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_854
timestamp 1698175906
transform 1 0 75824 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_855
timestamp 1698175906
transform 1 0 83664 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_856
timestamp 1698175906
transform 1 0 91504 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_857
timestamp 1698175906
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_858
timestamp 1698175906
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_859
timestamp 1698175906
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_860
timestamp 1698175906
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_861
timestamp 1698175906
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_862
timestamp 1698175906
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_863
timestamp 1698175906
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_864
timestamp 1698175906
transform 1 0 64064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_865
timestamp 1698175906
transform 1 0 71904 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_866
timestamp 1698175906
transform 1 0 79744 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_867
timestamp 1698175906
transform 1 0 87584 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_868
timestamp 1698175906
transform 1 0 95424 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_869
timestamp 1698175906
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_870
timestamp 1698175906
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_871
timestamp 1698175906
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_872
timestamp 1698175906
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_873
timestamp 1698175906
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_874
timestamp 1698175906
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_875
timestamp 1698175906
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_876
timestamp 1698175906
transform 1 0 60144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_877
timestamp 1698175906
transform 1 0 67984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_878
timestamp 1698175906
transform 1 0 75824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_879
timestamp 1698175906
transform 1 0 83664 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_880
timestamp 1698175906
transform 1 0 91504 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_881
timestamp 1698175906
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_882
timestamp 1698175906
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_883
timestamp 1698175906
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_884
timestamp 1698175906
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_885
timestamp 1698175906
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_886
timestamp 1698175906
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_887
timestamp 1698175906
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_888
timestamp 1698175906
transform 1 0 64064 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_889
timestamp 1698175906
transform 1 0 71904 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_890
timestamp 1698175906
transform 1 0 79744 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_891
timestamp 1698175906
transform 1 0 87584 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_892
timestamp 1698175906
transform 1 0 95424 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_893
timestamp 1698175906
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_894
timestamp 1698175906
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_895
timestamp 1698175906
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_896
timestamp 1698175906
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_897
timestamp 1698175906
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_898
timestamp 1698175906
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_899
timestamp 1698175906
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_900
timestamp 1698175906
transform 1 0 60144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_901
timestamp 1698175906
transform 1 0 67984 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_902
timestamp 1698175906
transform 1 0 75824 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_903
timestamp 1698175906
transform 1 0 83664 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_904
timestamp 1698175906
transform 1 0 91504 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_905
timestamp 1698175906
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_906
timestamp 1698175906
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_907
timestamp 1698175906
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_908
timestamp 1698175906
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_909
timestamp 1698175906
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_910
timestamp 1698175906
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_911
timestamp 1698175906
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_912
timestamp 1698175906
transform 1 0 64064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_913
timestamp 1698175906
transform 1 0 71904 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_914
timestamp 1698175906
transform 1 0 79744 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_915
timestamp 1698175906
transform 1 0 87584 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_916
timestamp 1698175906
transform 1 0 95424 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_917
timestamp 1698175906
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_918
timestamp 1698175906
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_919
timestamp 1698175906
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_920
timestamp 1698175906
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_921
timestamp 1698175906
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_922
timestamp 1698175906
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_923
timestamp 1698175906
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_924
timestamp 1698175906
transform 1 0 60144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_925
timestamp 1698175906
transform 1 0 67984 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_926
timestamp 1698175906
transform 1 0 75824 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_927
timestamp 1698175906
transform 1 0 83664 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_928
timestamp 1698175906
transform 1 0 91504 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_929
timestamp 1698175906
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_930
timestamp 1698175906
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_931
timestamp 1698175906
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_932
timestamp 1698175906
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_933
timestamp 1698175906
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_934
timestamp 1698175906
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_935
timestamp 1698175906
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_936
timestamp 1698175906
transform 1 0 64064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_937
timestamp 1698175906
transform 1 0 71904 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_938
timestamp 1698175906
transform 1 0 79744 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_939
timestamp 1698175906
transform 1 0 87584 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_940
timestamp 1698175906
transform 1 0 95424 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_941
timestamp 1698175906
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_942
timestamp 1698175906
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_943
timestamp 1698175906
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_944
timestamp 1698175906
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_945
timestamp 1698175906
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_946
timestamp 1698175906
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_947
timestamp 1698175906
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_948
timestamp 1698175906
transform 1 0 60144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_949
timestamp 1698175906
transform 1 0 67984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_950
timestamp 1698175906
transform 1 0 75824 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_951
timestamp 1698175906
transform 1 0 83664 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_952
timestamp 1698175906
transform 1 0 91504 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_953
timestamp 1698175906
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_954
timestamp 1698175906
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_955
timestamp 1698175906
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_956
timestamp 1698175906
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_957
timestamp 1698175906
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_958
timestamp 1698175906
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_959
timestamp 1698175906
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_960
timestamp 1698175906
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_961
timestamp 1698175906
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_962
timestamp 1698175906
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_963
timestamp 1698175906
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_964
timestamp 1698175906
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_965
timestamp 1698175906
transform 1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_966
timestamp 1698175906
transform 1 0 54656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_967
timestamp 1698175906
transform 1 0 58464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_968
timestamp 1698175906
transform 1 0 62272 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_969
timestamp 1698175906
transform 1 0 66080 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_970
timestamp 1698175906
transform 1 0 69888 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_971
timestamp 1698175906
transform 1 0 73696 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_972
timestamp 1698175906
transform 1 0 77504 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_973
timestamp 1698175906
transform 1 0 81312 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_974
timestamp 1698175906
transform 1 0 85120 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_975
timestamp 1698175906
transform 1 0 88928 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_976
timestamp 1698175906
transform 1 0 92736 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_977
timestamp 1698175906
transform 1 0 96544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_adc_reg._287_
timestamp 1698175906
transform -1 0 43680 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_adc_reg._288_
timestamp 1698175906
transform 1 0 42896 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_adc_reg._289_
timestamp 1698175906
transform 1 0 34720 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._290_
timestamp 1698175906
transform 1 0 35168 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  u_adc_reg._291_
timestamp 1698175906
transform -1 0 40992 0 1 34496
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  u_adc_reg._292_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37632 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  u_adc_reg._293_
timestamp 1698175906
transform -1 0 39536 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_adc_reg._294_
timestamp 1698175906
transform -1 0 37744 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  u_adc_reg._295_
timestamp 1698175906
transform -1 0 11648 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_adc_reg._296_
timestamp 1698175906
transform -1 0 57456 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  u_adc_reg._297_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 57680 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  u_adc_reg._298_
timestamp 1698175906
transform 1 0 74256 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  u_adc_reg._299_
timestamp 1698175906
transform 1 0 84112 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._300_
timestamp 1698175906
transform -1 0 55216 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._301_
timestamp 1698175906
transform 1 0 56672 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  u_adc_reg._302_
timestamp 1698175906
transform -1 0 46592 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._303_
timestamp 1698175906
transform 1 0 39536 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  u_adc_reg._304_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 46256 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._305_
timestamp 1698175906
transform 1 0 47600 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._306_
timestamp 1698175906
transform -1 0 44352 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  u_adc_reg._307_
timestamp 1698175906
transform -1 0 46256 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  u_adc_reg._308_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 45248 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._309_
timestamp 1698175906
transform -1 0 46704 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_adc_reg._310_
timestamp 1698175906
transform 1 0 46704 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_adc_reg._311_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 46704 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_adc_reg._312_
timestamp 1698175906
transform 1 0 49056 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  u_adc_reg._313_
timestamp 1698175906
transform -1 0 44240 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._314_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 41888 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._315_
timestamp 1698175906
transform -1 0 41888 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  u_adc_reg._316_
timestamp 1698175906
transform -1 0 40432 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  u_adc_reg._317_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 39984 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  u_adc_reg._318_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 42672 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  u_adc_reg._319_
timestamp 1698175906
transform 1 0 44912 0 1 29792
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  u_adc_reg._320_
timestamp 1698175906
transform -1 0 47040 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._321_
timestamp 1698175906
transform 1 0 56560 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._322_
timestamp 1698175906
transform -1 0 56224 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._323_
timestamp 1698175906
transform -1 0 78624 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._324_
timestamp 1698175906
transform 1 0 79632 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._325_
timestamp 1698175906
transform 1 0 72128 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._326_
timestamp 1698175906
transform -1 0 70896 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._327_
timestamp 1698175906
transform 1 0 72912 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._328_
timestamp 1698175906
transform 1 0 72240 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._329_
timestamp 1698175906
transform 1 0 63840 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._330_
timestamp 1698175906
transform -1 0 63616 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._331_
timestamp 1698175906
transform 1 0 44688 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._332_
timestamp 1698175906
transform -1 0 44464 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._333_
timestamp 1698175906
transform 1 0 64960 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._334_
timestamp 1698175906
transform -1 0 64960 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._335_
timestamp 1698175906
transform 1 0 44688 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._336_
timestamp 1698175906
transform -1 0 44464 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  u_adc_reg._337_
timestamp 1698175906
transform 1 0 44800 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  u_adc_reg._338_
timestamp 1698175906
transform 1 0 45136 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._339_
timestamp 1698175906
transform 1 0 61936 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._340_
timestamp 1698175906
transform 1 0 62496 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._341_
timestamp 1698175906
transform -1 0 79520 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._342_
timestamp 1698175906
transform 1 0 79072 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._343_
timestamp 1698175906
transform 1 0 72128 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._344_
timestamp 1698175906
transform -1 0 71904 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._345_
timestamp 1698175906
transform 1 0 77280 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._346_
timestamp 1698175906
transform 1 0 77616 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._347_
timestamp 1698175906
transform 1 0 64512 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._348_
timestamp 1698175906
transform 1 0 64512 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._349_
timestamp 1698175906
transform 1 0 44688 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._350_
timestamp 1698175906
transform -1 0 44464 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._351_
timestamp 1698175906
transform 1 0 68208 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._352_
timestamp 1698175906
transform 1 0 67872 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._353_
timestamp 1698175906
transform 1 0 44576 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._354_
timestamp 1698175906
transform 1 0 43792 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  u_adc_reg._355_
timestamp 1698175906
transform 1 0 40320 0 1 29792
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  u_adc_reg._356_
timestamp 1698175906
transform 1 0 42896 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._357_
timestamp 1698175906
transform 1 0 53424 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._358_
timestamp 1698175906
transform -1 0 53760 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._359_
timestamp 1698175906
transform 1 0 76608 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._360_
timestamp 1698175906
transform 1 0 76048 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._361_
timestamp 1698175906
transform 1 0 72128 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._362_
timestamp 1698175906
transform -1 0 71568 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._363_
timestamp 1698175906
transform 1 0 72912 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._364_
timestamp 1698175906
transform -1 0 72800 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._365_
timestamp 1698175906
transform 1 0 61488 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._366_
timestamp 1698175906
transform -1 0 61488 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._367_
timestamp 1698175906
transform 1 0 38864 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._368_
timestamp 1698175906
transform -1 0 37856 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._369_
timestamp 1698175906
transform 1 0 60368 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._370_
timestamp 1698175906
transform -1 0 59472 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._371_
timestamp 1698175906
transform 1 0 40768 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._372_
timestamp 1698175906
transform -1 0 39760 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  u_adc_reg._373_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 39088 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  u_adc_reg._374_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 44688 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._375_
timestamp 1698175906
transform 1 0 53200 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._376_
timestamp 1698175906
transform -1 0 51408 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._377_
timestamp 1698175906
transform 1 0 56448 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._378_
timestamp 1698175906
transform -1 0 56224 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._379_
timestamp 1698175906
transform 1 0 56112 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._380_
timestamp 1698175906
transform 1 0 56448 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._381_
timestamp 1698175906
transform 1 0 56448 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._382_
timestamp 1698175906
transform 1 0 56896 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._383_
timestamp 1698175906
transform 1 0 33376 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._384_
timestamp 1698175906
transform -1 0 32704 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._385_
timestamp 1698175906
transform 1 0 33600 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._386_
timestamp 1698175906
transform -1 0 33600 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._387_
timestamp 1698175906
transform 1 0 33936 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._388_
timestamp 1698175906
transform -1 0 33600 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._389_
timestamp 1698175906
transform 1 0 33712 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._390_
timestamp 1698175906
transform -1 0 33600 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_adc_reg._391_
timestamp 1698175906
transform 1 0 43792 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  u_adc_reg._392_
timestamp 1698175906
transform 1 0 43232 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._393_
timestamp 1698175906
transform 1 0 61264 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._394_
timestamp 1698175906
transform -1 0 61712 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._395_
timestamp 1698175906
transform -1 0 78960 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._396_
timestamp 1698175906
transform 1 0 79184 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._397_
timestamp 1698175906
transform 1 0 69888 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._398_
timestamp 1698175906
transform -1 0 69104 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._399_
timestamp 1698175906
transform -1 0 78960 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._400_
timestamp 1698175906
transform 1 0 78064 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._401_
timestamp 1698175906
transform 1 0 62160 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._402_
timestamp 1698175906
transform -1 0 62384 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._403_
timestamp 1698175906
transform 1 0 40768 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._404_
timestamp 1698175906
transform -1 0 40432 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._405_
timestamp 1698175906
transform 1 0 66304 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._406_
timestamp 1698175906
transform -1 0 65744 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._407_
timestamp 1698175906
transform 1 0 40768 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._408_
timestamp 1698175906
transform -1 0 39984 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  u_adc_reg._409_
timestamp 1698175906
transform 1 0 43120 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._410_
timestamp 1698175906
transform 1 0 56448 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._411_
timestamp 1698175906
transform -1 0 56336 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._412_
timestamp 1698175906
transform 1 0 51632 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._413_
timestamp 1698175906
transform -1 0 51072 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._414_
timestamp 1698175906
transform 1 0 54320 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._415_
timestamp 1698175906
transform -1 0 52192 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._416_
timestamp 1698175906
transform 1 0 53424 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._417_
timestamp 1698175906
transform -1 0 51184 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._418_
timestamp 1698175906
transform 1 0 29232 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._419_
timestamp 1698175906
transform -1 0 27440 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._420_
timestamp 1698175906
transform 1 0 29344 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._421_
timestamp 1698175906
transform -1 0 27440 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._422_
timestamp 1698175906
transform 1 0 29008 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._423_
timestamp 1698175906
transform -1 0 27104 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._424_
timestamp 1698175906
transform 1 0 27104 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._425_
timestamp 1698175906
transform -1 0 27664 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  u_adc_reg._426_
timestamp 1698175906
transform -1 0 92624 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  u_adc_reg._427_
timestamp 1698175906
transform 1 0 46704 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  u_adc_reg._428_
timestamp 1698175906
transform 1 0 46144 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  u_adc_reg._429_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 47040 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  u_adc_reg._430_
timestamp 1698175906
transform 1 0 47488 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  u_adc_reg._431_
timestamp 1698175906
transform 1 0 46592 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  u_adc_reg._432_
timestamp 1698175906
transform -1 0 50736 0 1 32928
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_8  u_adc_reg._433_
timestamp 1698175906
transform 1 0 51408 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  u_adc_reg._434_
timestamp 1698175906
transform 1 0 47152 0 1 34496
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  u_adc_reg._435_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 61264 0 -1 32928
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  u_adc_reg._436_
timestamp 1698175906
transform -1 0 50176 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  u_adc_reg._437_
timestamp 1698175906
transform 1 0 52528 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  u_adc_reg._438_
timestamp 1698175906
transform 1 0 48832 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  u_adc_reg._439_
timestamp 1698175906
transform 1 0 46816 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  u_adc_reg._440_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 53648 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  u_adc_reg._441_
timestamp 1698175906
transform -1 0 58016 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._442_
timestamp 1698175906
transform 1 0 38864 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  u_adc_reg._443_
timestamp 1698175906
transform 1 0 52976 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  u_adc_reg._444_
timestamp 1698175906
transform 1 0 74032 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  u_adc_reg._445_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 64288 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  u_adc_reg._446_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 89152 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._447_
timestamp 1698175906
transform 1 0 90384 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_adc_reg._448_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 75600 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._449_
timestamp 1698175906
transform 1 0 77168 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  u_adc_reg._450_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 53088 0 -1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  u_adc_reg._451_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 61712 0 -1 47040
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  u_adc_reg._452_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 50848 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_adc_reg._453_
timestamp 1698175906
transform -1 0 77840 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_adc_reg._454_
timestamp 1698175906
transform 1 0 76720 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._455_
timestamp 1698175906
transform -1 0 86464 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._456_
timestamp 1698175906
transform 1 0 85792 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_adc_reg._457_
timestamp 1698175906
transform -1 0 75488 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._458_
timestamp 1698175906
transform 1 0 72800 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  u_adc_reg._459_
timestamp 1698175906
transform -1 0 60144 0 1 45472
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_adc_reg._460_
timestamp 1698175906
transform 1 0 73808 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_adc_reg._461_
timestamp 1698175906
transform 1 0 73584 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._462_
timestamp 1698175906
transform -1 0 93744 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._463_
timestamp 1698175906
transform 1 0 92400 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_adc_reg._464_
timestamp 1698175906
transform 1 0 76048 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._465_
timestamp 1698175906
transform 1 0 77056 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  u_adc_reg._466_
timestamp 1698175906
transform 1 0 54208 0 1 40768
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_adc_reg._467_
timestamp 1698175906
transform 1 0 76160 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_adc_reg._468_
timestamp 1698175906
transform 1 0 76384 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._469_
timestamp 1698175906
transform -1 0 89488 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._470_
timestamp 1698175906
transform -1 0 87360 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_adc_reg._471_
timestamp 1698175906
transform -1 0 67424 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._472_
timestamp 1698175906
transform 1 0 64400 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  u_adc_reg._473_
timestamp 1698175906
transform 1 0 33488 0 -1 47040
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_adc_reg._474_
timestamp 1698175906
transform 1 0 64736 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_adc_reg._475_
timestamp 1698175906
transform -1 0 66864 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._476_
timestamp 1698175906
transform -1 0 87584 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._477_
timestamp 1698175906
transform -1 0 86912 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  u_adc_reg._478_
timestamp 1698175906
transform 1 0 47936 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._479_
timestamp 1698175906
transform -1 0 47824 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  u_adc_reg._480_
timestamp 1698175906
transform 1 0 33712 0 -1 43904
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  u_adc_reg._481_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 48496 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  u_adc_reg._482_
timestamp 1698175906
transform 1 0 47376 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._483_
timestamp 1698175906
transform -1 0 93184 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._484_
timestamp 1698175906
transform 1 0 91728 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_adc_reg._485_
timestamp 1698175906
transform -1 0 69440 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._486_
timestamp 1698175906
transform 1 0 68208 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  u_adc_reg._487_
timestamp 1698175906
transform 1 0 33936 0 -1 40768
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  u_adc_reg._488_
timestamp 1698175906
transform 1 0 68208 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  u_adc_reg._489_
timestamp 1698175906
transform 1 0 67984 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._490_
timestamp 1698175906
transform -1 0 93408 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._491_
timestamp 1698175906
transform -1 0 92512 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  u_adc_reg._492_
timestamp 1698175906
transform 1 0 48608 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._493_
timestamp 1698175906
transform 1 0 47824 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  u_adc_reg._494_
timestamp 1698175906
transform 1 0 33600 0 -1 37632
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  u_adc_reg._495_
timestamp 1698175906
transform -1 0 50288 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  u_adc_reg._496_
timestamp 1698175906
transform 1 0 48048 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg._497_
timestamp 1698175906
transform -1 0 92288 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg._498_
timestamp 1698175906
transform 1 0 90944 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._499_
timestamp 1698175906
transform 1 0 36064 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  u_adc_reg._500_
timestamp 1698175906
transform 1 0 73360 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._501_
timestamp 1698175906
transform -1 0 84448 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._502_
timestamp 1698175906
transform 1 0 82320 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._503_
timestamp 1698175906
transform 1 0 36848 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._504_
timestamp 1698175906
transform -1 0 86128 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._505_
timestamp 1698175906
transform 1 0 84672 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._506_
timestamp 1698175906
transform 1 0 36848 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._507_
timestamp 1698175906
transform -1 0 85680 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._508_
timestamp 1698175906
transform 1 0 84112 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._509_
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._510_
timestamp 1698175906
transform -1 0 80528 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._511_
timestamp 1698175906
transform 1 0 78064 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._512_
timestamp 1698175906
transform 1 0 36512 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._513_
timestamp 1698175906
transform -1 0 86128 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._514_
timestamp 1698175906
transform 1 0 84448 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._515_
timestamp 1698175906
transform -1 0 36064 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  u_adc_reg._516_
timestamp 1698175906
transform 1 0 74928 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._517_
timestamp 1698175906
transform -1 0 74816 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._518_
timestamp 1698175906
transform 1 0 72576 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._519_
timestamp 1698175906
transform 1 0 35728 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._520_
timestamp 1698175906
transform -1 0 72688 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._521_
timestamp 1698175906
transform 1 0 69552 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._522_
timestamp 1698175906
transform 1 0 36064 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._523_
timestamp 1698175906
transform -1 0 66976 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._524_
timestamp 1698175906
transform 1 0 64960 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._525_
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._526_
timestamp 1698175906
transform -1 0 71008 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._527_
timestamp 1698175906
transform 1 0 68432 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  u_adc_reg._528_
timestamp 1698175906
transform -1 0 77616 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  u_adc_reg._529_
timestamp 1698175906
transform 1 0 57792 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._530_
timestamp 1698175906
transform 1 0 60928 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._531_
timestamp 1698175906
transform -1 0 65968 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._532_
timestamp 1698175906
transform 1 0 62832 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._533_
timestamp 1698175906
transform 1 0 61488 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._534_
timestamp 1698175906
transform -1 0 77840 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._535_
timestamp 1698175906
transform 1 0 76160 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._536_
timestamp 1698175906
transform 1 0 60368 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._537_
timestamp 1698175906
transform -1 0 74704 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._538_
timestamp 1698175906
transform 1 0 72352 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._539_
timestamp 1698175906
transform 1 0 61488 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._540_
timestamp 1698175906
transform -1 0 65520 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._541_
timestamp 1698175906
transform 1 0 62160 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._542_
timestamp 1698175906
transform 1 0 60928 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._543_
timestamp 1698175906
transform -1 0 69104 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._544_
timestamp 1698175906
transform 1 0 66976 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._545_
timestamp 1698175906
transform 1 0 59808 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._546_
timestamp 1698175906
transform -1 0 78400 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._547_
timestamp 1698175906
transform 1 0 77168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._548_
timestamp 1698175906
transform 1 0 60368 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._549_
timestamp 1698175906
transform -1 0 64848 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._550_
timestamp 1698175906
transform 1 0 62160 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._551_
timestamp 1698175906
transform 1 0 60368 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._552_
timestamp 1698175906
transform -1 0 80752 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._553_
timestamp 1698175906
transform 1 0 77616 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._554_
timestamp 1698175906
transform 1 0 59584 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._555_
timestamp 1698175906
transform -1 0 69664 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._556_
timestamp 1698175906
transform 1 0 68208 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._557_
timestamp 1698175906
transform 1 0 60928 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._558_
timestamp 1698175906
transform -1 0 75488 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._559_
timestamp 1698175906
transform 1 0 73360 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._560_
timestamp 1698175906
transform 1 0 45808 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._561_
timestamp 1698175906
transform -1 0 85120 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._562_
timestamp 1698175906
transform 1 0 81872 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._563_
timestamp 1698175906
transform 1 0 43568 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._564_
timestamp 1698175906
transform 1 0 85344 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._565_
timestamp 1698175906
transform 1 0 84784 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._566_
timestamp 1698175906
transform 1 0 43680 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._567_
timestamp 1698175906
transform -1 0 78400 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._568_
timestamp 1698175906
transform 1 0 76160 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._569_
timestamp 1698175906
transform 1 0 55888 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._570_
timestamp 1698175906
transform -1 0 73696 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._571_
timestamp 1698175906
transform 1 0 71904 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._572_
timestamp 1698175906
transform 1 0 39984 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  u_adc_reg._573_
timestamp 1698175906
transform -1 0 83552 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  u_adc_reg._574_
timestamp 1698175906
transform 1 0 80864 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._575__130
timestamp 1698175906
transform 1 0 48272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_adc_reg._575_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 48608 0 -1 28224
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_adc_reg._576_
timestamp 1698175906
transform 1 0 49952 0 -1 29792
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._576__131
timestamp 1698175906
transform -1 0 50512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._577__132
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_adc_reg._577_
timestamp 1698175906
transform 1 0 40768 0 -1 28224
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._578__133
timestamp 1698175906
transform -1 0 39872 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._578_
timestamp 1698175906
transform 1 0 38640 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._579__134
timestamp 1698175906
transform 1 0 54768 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._579_
timestamp 1698175906
transform 1 0 55216 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._580__135
timestamp 1698175906
transform -1 0 81424 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._580_
timestamp 1698175906
transform 1 0 80752 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._581__136
timestamp 1698175906
transform -1 0 70224 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._581_
timestamp 1698175906
transform 1 0 69552 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._582__137
timestamp 1698175906
transform 1 0 71680 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._582_
timestamp 1698175906
transform 1 0 72128 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._583__138
timestamp 1698175906
transform -1 0 62720 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._583_
timestamp 1698175906
transform 1 0 62048 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._584__139
timestamp 1698175906
transform -1 0 44128 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._584_
timestamp 1698175906
transform 1 0 43456 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._585_
timestamp 1698175906
transform 1 0 63280 0 1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._585__140
timestamp 1698175906
transform 1 0 62832 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._586__141
timestamp 1698175906
transform -1 0 44128 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._586_
timestamp 1698175906
transform 1 0 43456 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._587_
timestamp 1698175906
transform 1 0 62944 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._587__142
timestamp 1698175906
transform -1 0 64064 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._588__143
timestamp 1698175906
transform -1 0 80528 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._588_
timestamp 1698175906
transform 1 0 79968 0 -1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._589__144
timestamp 1698175906
transform 1 0 70784 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._589_
timestamp 1698175906
transform 1 0 70896 0 1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._590__145
timestamp 1698175906
transform -1 0 79408 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._590_
timestamp 1698175906
transform 1 0 77840 0 1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._591__146
timestamp 1698175906
transform -1 0 65856 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._591_
timestamp 1698175906
transform 1 0 65184 0 -1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._592__147
timestamp 1698175906
transform -1 0 43792 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._592_
timestamp 1698175906
transform 1 0 43232 0 -1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._593__148
timestamp 1698175906
transform -1 0 68992 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._593_
timestamp 1698175906
transform 1 0 68208 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._594__149
timestamp 1698175906
transform 1 0 43792 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._594_
timestamp 1698175906
transform 1 0 44688 0 1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._595__150
timestamp 1698175906
transform -1 0 54208 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._595_
timestamp 1698175906
transform 1 0 52640 0 1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._596_
timestamp 1698175906
transform 1 0 76720 0 1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._596__151
timestamp 1698175906
transform -1 0 77392 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._597_
timestamp 1698175906
transform 1 0 70224 0 1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._597__152
timestamp 1698175906
transform -1 0 70896 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._598__153
timestamp 1698175906
transform 1 0 70560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._598_
timestamp 1698175906
transform 1 0 71008 0 1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._599_
timestamp 1698175906
transform 1 0 60368 0 1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._599__154
timestamp 1698175906
transform 1 0 59696 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._600_
timestamp 1698175906
transform 1 0 36736 0 -1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._600__155
timestamp 1698175906
transform 1 0 36176 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._601__156
timestamp 1698175906
transform -1 0 58688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._601_
timestamp 1698175906
transform 1 0 58016 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._602__157
timestamp 1698175906
transform -1 0 38864 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._602_
timestamp 1698175906
transform 1 0 38304 0 1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._603_
timestamp 1698175906
transform 1 0 49392 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._603__158
timestamp 1698175906
transform 1 0 48944 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._604__159
timestamp 1698175906
transform -1 0 55328 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._604_
timestamp 1698175906
transform 1 0 54656 0 1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._605__160
timestamp 1698175906
transform -1 0 58240 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._605_
timestamp 1698175906
transform 1 0 56448 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._606__161
timestamp 1698175906
transform -1 0 58688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._606_
timestamp 1698175906
transform 1 0 58016 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._607__162
timestamp 1698175906
transform -1 0 31472 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._607_
timestamp 1698175906
transform 1 0 30800 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._608__163
timestamp 1698175906
transform -1 0 32032 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._608_
timestamp 1698175906
transform 1 0 31360 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._609__164
timestamp 1698175906
transform -1 0 31808 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._609_
timestamp 1698175906
transform 1 0 31136 0 1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._610__165
timestamp 1698175906
transform -1 0 32032 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._610_
timestamp 1698175906
transform 1 0 31360 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._611_
timestamp 1698175906
transform 1 0 60368 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._611__166
timestamp 1698175906
transform 1 0 59696 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._612_
timestamp 1698175906
transform 1 0 79856 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._612__167
timestamp 1698175906
transform -1 0 81312 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._613__168
timestamp 1698175906
transform 1 0 67312 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._613_
timestamp 1698175906
transform 1 0 68208 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._614_
timestamp 1698175906
transform 1 0 78736 0 1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._614__169
timestamp 1698175906
transform -1 0 79296 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._615__170
timestamp 1698175906
transform -1 0 61040 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._615_
timestamp 1698175906
transform 1 0 60368 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._616__171
timestamp 1698175906
transform 1 0 37184 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._616_
timestamp 1698175906
transform 1 0 37744 0 1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._617__172
timestamp 1698175906
transform 1 0 63504 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._617_
timestamp 1698175906
transform 1 0 63952 0 1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._618_
timestamp 1698175906
transform 1 0 38304 0 1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._618__173
timestamp 1698175906
transform -1 0 38864 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._619__174
timestamp 1698175906
transform -1 0 56784 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._619_
timestamp 1698175906
transform 1 0 55216 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._620__175
timestamp 1698175906
transform 1 0 48720 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._620_
timestamp 1698175906
transform 1 0 49168 0 -1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._621__176
timestamp 1698175906
transform -1 0 50512 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._621_
timestamp 1698175906
transform 1 0 49840 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._622__177
timestamp 1698175906
transform -1 0 49952 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._622_
timestamp 1698175906
transform 1 0 49392 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._623_
timestamp 1698175906
transform 1 0 25424 0 -1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._623__178
timestamp 1698175906
transform -1 0 25984 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._624__179
timestamp 1698175906
transform 1 0 25088 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._624_
timestamp 1698175906
transform 1 0 25536 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._625__180
timestamp 1698175906
transform -1 0 25760 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._625_
timestamp 1698175906
transform 1 0 25200 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._626__181
timestamp 1698175906
transform -1 0 26656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._626_
timestamp 1698175906
transform 1 0 25984 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._627__182
timestamp 1698175906
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._627_
timestamp 1698175906
transform 1 0 56448 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._628__183
timestamp 1698175906
transform -1 0 54544 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._628_
timestamp 1698175906
transform 1 0 53984 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._629__184
timestamp 1698175906
transform -1 0 35728 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._629_
timestamp 1698175906
transform 1 0 35056 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._630__185
timestamp 1698175906
transform 1 0 8624 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_adc_reg._630_
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_4  u_adc_reg._631_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._631__186
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._632__187
timestamp 1698175906
transform -1 0 26544 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_adc_reg._632_
timestamp 1698175906
transform 1 0 25872 0 -1 32928
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._633__188
timestamp 1698175906
transform -1 0 27776 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_adc_reg._633_
timestamp 1698175906
transform 1 0 27104 0 -1 34496
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._634__189
timestamp 1698175906
transform 1 0 5376 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._634_
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._635_
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._635__190
timestamp 1698175906
transform -1 0 2688 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._636__191
timestamp 1698175906
transform -1 0 2240 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._636_
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._637_
timestamp 1698175906
transform 1 0 6160 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._637__192
timestamp 1698175906
transform 1 0 5712 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._638__193
timestamp 1698175906
transform -1 0 12208 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._638_
timestamp 1698175906
transform 1 0 11536 0 -1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._639__194
timestamp 1698175906
transform -1 0 2240 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._639_
timestamp 1698175906
transform 1 0 1568 0 -1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._640_
timestamp 1698175906
transform 1 0 16688 0 1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._640__195
timestamp 1698175906
transform 1 0 16240 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._641__196
timestamp 1698175906
transform -1 0 5936 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._641_
timestamp 1698175906
transform 1 0 5264 0 -1 50176
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._642__197
timestamp 1698175906
transform -1 0 9856 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._642_
timestamp 1698175906
transform 1 0 8736 0 1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._643_
timestamp 1698175906
transform 1 0 2240 0 -1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._643__198
timestamp 1698175906
transform -1 0 2912 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._644__199
timestamp 1698175906
transform -1 0 3472 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._644_
timestamp 1698175906
transform 1 0 2800 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._645__200
timestamp 1698175906
transform -1 0 2912 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._645_
timestamp 1698175906
transform 1 0 2240 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._646__201
timestamp 1698175906
transform 1 0 8624 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._646_
timestamp 1698175906
transform 1 0 9408 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._647_
timestamp 1698175906
transform 1 0 2576 0 -1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._647__202
timestamp 1698175906
transform -1 0 3248 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._648_
timestamp 1698175906
transform 1 0 1568 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._648__203
timestamp 1698175906
transform -1 0 2688 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._649__204
timestamp 1698175906
transform -1 0 2688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._649_
timestamp 1698175906
transform 1 0 2128 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._650_
timestamp 1698175906
transform 1 0 5376 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._650__205
timestamp 1698175906
transform -1 0 5936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._651__206
timestamp 1698175906
transform -1 0 3024 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._651_
timestamp 1698175906
transform 1 0 2464 0 -1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._652__207
timestamp 1698175906
transform -1 0 2688 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._652_
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._653__208
timestamp 1698175906
transform -1 0 11648 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._653_
timestamp 1698175906
transform 1 0 11088 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._654__209
timestamp 1698175906
transform -1 0 2688 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._654_
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._655_
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._655__210
timestamp 1698175906
transform 1 0 4816 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._656_
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._656__211
timestamp 1698175906
transform 1 0 4816 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._657_
timestamp 1698175906
transform 1 0 2128 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._657__212
timestamp 1698175906
transform 1 0 1680 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._658_
timestamp 1698175906
transform 1 0 21056 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._658__213
timestamp 1698175906
transform 1 0 20608 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._659_
timestamp 1698175906
transform 1 0 8848 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._659__214
timestamp 1698175906
transform 1 0 8400 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._660_
timestamp 1698175906
transform 1 0 18368 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._660__215
timestamp 1698175906
transform 1 0 17920 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._661__216
timestamp 1698175906
transform 1 0 1680 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._661_
timestamp 1698175906
transform 1 0 2128 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._662__217
timestamp 1698175906
transform -1 0 7728 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._662_
timestamp 1698175906
transform 1 0 7056 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._663__218
timestamp 1698175906
transform 1 0 5040 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._663_
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._664__219
timestamp 1698175906
transform -1 0 2240 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._664_
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._665__220
timestamp 1698175906
transform -1 0 16912 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._665_
timestamp 1698175906
transform 1 0 15568 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._666__221
timestamp 1698175906
transform -1 0 27216 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._666_
timestamp 1698175906
transform 1 0 26544 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._667__222
timestamp 1698175906
transform -1 0 29456 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._667_
timestamp 1698175906
transform 1 0 28784 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._668_
timestamp 1698175906
transform 1 0 10080 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._668__223
timestamp 1698175906
transform 1 0 9632 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._669__224
timestamp 1698175906
transform -1 0 19376 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._669_
timestamp 1698175906
transform 1 0 18704 0 -1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._670_
timestamp 1698175906
transform 1 0 44688 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._670__225
timestamp 1698175906
transform 1 0 44016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._671__226
timestamp 1698175906
transform 1 0 49392 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._671_
timestamp 1698175906
transform 1 0 49840 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._672__227
timestamp 1698175906
transform -1 0 90720 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._672_
timestamp 1698175906
transform 1 0 90048 0 -1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._673__228
timestamp 1698175906
transform -1 0 87136 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._673_
timestamp 1698175906
transform 1 0 86464 0 1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._674_
timestamp 1698175906
transform 1 0 92512 0 1 48608
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._674__229
timestamp 1698175906
transform 1 0 92064 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._675__230
timestamp 1698175906
transform -1 0 86912 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._675_
timestamp 1698175906
transform 1 0 86352 0 1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._676__231
timestamp 1698175906
transform -1 0 87360 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._676_
timestamp 1698175906
transform 1 0 85904 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._677__232
timestamp 1698175906
transform -1 0 92848 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._677_
timestamp 1698175906
transform 1 0 91952 0 1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._678__233
timestamp 1698175906
transform 1 0 91168 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._678_
timestamp 1698175906
transform 1 0 91616 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._679_
timestamp 1698175906
transform 1 0 91616 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._679__234
timestamp 1698175906
transform -1 0 92400 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._680__235
timestamp 1698175906
transform -1 0 82880 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._680_
timestamp 1698175906
transform 1 0 82208 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._681_
timestamp 1698175906
transform 1 0 86576 0 1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._681__236
timestamp 1698175906
transform 1 0 86128 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._682__237
timestamp 1698175906
transform -1 0 85008 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._682_
timestamp 1698175906
transform 1 0 83776 0 -1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._683__238
timestamp 1698175906
transform -1 0 79408 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._683_
timestamp 1698175906
transform 1 0 77840 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._684__239
timestamp 1698175906
transform -1 0 85792 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._684_
timestamp 1698175906
transform 1 0 84448 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._685__240
timestamp 1698175906
transform -1 0 72688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._685_
timestamp 1698175906
transform 1 0 72016 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._686_
timestamp 1698175906
transform 1 0 69216 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._686__241
timestamp 1698175906
transform 1 0 68768 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._687__242
timestamp 1698175906
transform -1 0 66304 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._687_
timestamp 1698175906
transform 1 0 64848 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._688__243
timestamp 1698175906
transform 1 0 67536 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._688_
timestamp 1698175906
transform 1 0 68208 0 1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._689__244
timestamp 1698175906
transform -1 0 64176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._689_
timestamp 1698175906
transform 1 0 62496 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._690__245
timestamp 1698175906
transform -1 0 78064 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._690_
timestamp 1698175906
transform 1 0 75936 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._691_
timestamp 1698175906
transform 1 0 72016 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._691__246
timestamp 1698175906
transform 1 0 71568 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._692__247
timestamp 1698175906
transform -1 0 62160 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._692_
timestamp 1698175906
transform 1 0 61488 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._693__248
timestamp 1698175906
transform -1 0 66976 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._693_
timestamp 1698175906
transform 1 0 66528 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._694_
timestamp 1698175906
transform 1 0 78176 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._694__249
timestamp 1698175906
transform -1 0 78848 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._695__250
timestamp 1698175906
transform -1 0 62160 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._695_
timestamp 1698175906
transform 1 0 61488 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._696__251
timestamp 1698175906
transform -1 0 78960 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._696_
timestamp 1698175906
transform 1 0 77952 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._697_
timestamp 1698175906
transform 1 0 66864 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._697__252
timestamp 1698175906
transform -1 0 67424 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._698__253
timestamp 1698175906
transform -1 0 73248 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._698_
timestamp 1698175906
transform 1 0 72016 0 1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._699_
timestamp 1698175906
transform 1 0 82768 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._699__254
timestamp 1698175906
transform -1 0 83440 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._700__255
timestamp 1698175906
transform -1 0 86352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._700_
timestamp 1698175906
transform 1 0 85344 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._701__256
timestamp 1698175906
transform 1 0 75712 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._701_
timestamp 1698175906
transform 1 0 76048 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._702__257
timestamp 1698175906
transform -1 0 71344 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._702_
timestamp 1698175906
transform 1 0 70672 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg._703__258
timestamp 1698175906
transform -1 0 82208 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg._703_
timestamp 1698175906
transform 1 0 79856 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_adc_reg.u_reg_0._068_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._069_
timestamp 1698175906
transform -1 0 20832 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._070_
timestamp 1698175906
transform 1 0 19936 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._071_
timestamp 1698175906
transform -1 0 11088 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._072_
timestamp 1698175906
transform 1 0 8512 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._073_
timestamp 1698175906
transform -1 0 21728 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._074_
timestamp 1698175906
transform 1 0 20272 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._075_
timestamp 1698175906
transform 1 0 9184 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._076_
timestamp 1698175906
transform 1 0 8512 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._077_
timestamp 1698175906
transform -1 0 16128 0 -1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._078_
timestamp 1698175906
transform 1 0 13776 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._079_
timestamp 1698175906
transform -1 0 16800 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._080_
timestamp 1698175906
transform -1 0 15120 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._081_
timestamp 1698175906
transform -1 0 22848 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._082_
timestamp 1698175906
transform 1 0 19824 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._083_
timestamp 1698175906
transform -1 0 15008 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._084_
timestamp 1698175906
transform 1 0 12432 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_adc_reg.u_reg_0._085_
timestamp 1698175906
transform -1 0 11424 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._086_
timestamp 1698175906
transform -1 0 13104 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._087_
timestamp 1698175906
transform 1 0 13328 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._088_
timestamp 1698175906
transform -1 0 18928 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._089_
timestamp 1698175906
transform 1 0 18144 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._090_
timestamp 1698175906
transform -1 0 21952 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._091_
timestamp 1698175906
transform 1 0 20272 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._092_
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._093_
timestamp 1698175906
transform 1 0 8512 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._094_
timestamp 1698175906
transform -1 0 16800 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._095_
timestamp 1698175906
transform -1 0 15792 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._096_
timestamp 1698175906
transform -1 0 21616 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._097_
timestamp 1698175906
transform 1 0 21616 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._098_
timestamp 1698175906
transform -1 0 20944 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._099_
timestamp 1698175906
transform -1 0 21840 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._100_
timestamp 1698175906
transform -1 0 16464 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._101_
timestamp 1698175906
transform -1 0 15344 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_adc_reg.u_reg_0._102_
timestamp 1698175906
transform -1 0 11872 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._103_
timestamp 1698175906
transform -1 0 28560 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._104_
timestamp 1698175906
transform -1 0 27328 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._105_
timestamp 1698175906
transform -1 0 16576 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._106_
timestamp 1698175906
transform -1 0 14896 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._107_
timestamp 1698175906
transform -1 0 32368 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._108_
timestamp 1698175906
transform 1 0 31584 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._109_
timestamp 1698175906
transform -1 0 31808 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._110_
timestamp 1698175906
transform -1 0 30800 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._111_
timestamp 1698175906
transform -1 0 26544 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._112_
timestamp 1698175906
transform 1 0 24192 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._113_
timestamp 1698175906
transform -1 0 13664 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._114_
timestamp 1698175906
transform 1 0 13664 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._115_
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._116_
timestamp 1698175906
transform -1 0 20832 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._117_
timestamp 1698175906
transform -1 0 27552 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._118_
timestamp 1698175906
transform 1 0 26208 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  u_adc_reg.u_reg_0._119_
timestamp 1698175906
transform -1 0 12208 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._120_
timestamp 1698175906
transform -1 0 39872 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._121_
timestamp 1698175906
transform 1 0 38640 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._122_
timestamp 1698175906
transform -1 0 34496 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._123_
timestamp 1698175906
transform 1 0 32928 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._124_
timestamp 1698175906
transform -1 0 11984 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._125_
timestamp 1698175906
transform 1 0 11424 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._126_
timestamp 1698175906
transform -1 0 22848 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._127_
timestamp 1698175906
transform -1 0 21840 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._128_
timestamp 1698175906
transform -1 0 39984 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._129_
timestamp 1698175906
transform 1 0 38864 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._130_
timestamp 1698175906
transform -1 0 35056 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._131_
timestamp 1698175906
transform 1 0 33376 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._132_
timestamp 1698175906
transform -1 0 16464 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._133_
timestamp 1698175906
transform 1 0 14112 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  u_adc_reg.u_reg_0._134_
timestamp 1698175906
transform -1 0 24864 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  u_adc_reg.u_reg_0._135_
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_adc_reg.u_reg_0._136_
timestamp 1698175906
transform 1 0 20608 0 -1 42336
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._136__259
timestamp 1698175906
transform -1 0 21616 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_adc_reg.u_reg_0._137_
timestamp 1698175906
transform 1 0 9408 0 -1 47040
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._137__260
timestamp 1698175906
transform 1 0 8848 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._138__261
timestamp 1698175906
transform 1 0 20496 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._138_
timestamp 1698175906
transform 1 0 21168 0 1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._139__262
timestamp 1698175906
transform 1 0 8064 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  u_adc_reg.u_reg_0._139_
timestamp 1698175906
transform 1 0 9408 0 -1 43904
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._140__263
timestamp 1698175906
transform -1 0 14784 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._140_
timestamp 1698175906
transform 1 0 14112 0 1 47040
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._141__264
timestamp 1698175906
transform 1 0 14000 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._141_
timestamp 1698175906
transform 1 0 14224 0 1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._142__265
timestamp 1698175906
transform -1 0 21616 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._142_
timestamp 1698175906
transform 1 0 20496 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._143__266
timestamp 1698175906
transform -1 0 14224 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._143_
timestamp 1698175906
transform 1 0 13216 0 -1 42336
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._144__267
timestamp 1698175906
transform -1 0 14448 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._144_
timestamp 1698175906
transform 1 0 13104 0 -1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._145_
timestamp 1698175906
transform 1 0 18928 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._145__268
timestamp 1698175906
transform -1 0 19600 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._146_
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._146__269
timestamp 1698175906
transform -1 0 21952 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._147__270
timestamp 1698175906
transform 1 0 8064 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._147_
timestamp 1698175906
transform 1 0 8624 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._148__271
timestamp 1698175906
transform 1 0 14336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._148_
timestamp 1698175906
transform 1 0 14784 0 1 36064
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._149__272
timestamp 1698175906
transform -1 0 21616 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._149_
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._150__273
timestamp 1698175906
transform -1 0 21168 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._150_
timestamp 1698175906
transform 1 0 20496 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._151__274
timestamp 1698175906
transform -1 0 15792 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._151_
timestamp 1698175906
transform 1 0 14336 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._152__275
timestamp 1698175906
transform -1 0 27776 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._152_
timestamp 1698175906
transform 1 0 26208 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._153_
timestamp 1698175906
transform 1 0 13216 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._153__276
timestamp 1698175906
transform -1 0 14224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._154__277
timestamp 1698175906
transform 1 0 32480 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._154_
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._155__278
timestamp 1698175906
transform -1 0 31248 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._155_
timestamp 1698175906
transform 1 0 28896 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._156__279
timestamp 1698175906
transform 1 0 24416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._156_
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._157__280
timestamp 1698175906
transform -1 0 14784 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._157_
timestamp 1698175906
transform 1 0 13664 0 1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._158__281
timestamp 1698175906
transform -1 0 20048 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._158_
timestamp 1698175906
transform 1 0 19376 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._159_
timestamp 1698175906
transform 1 0 26432 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._159__282
timestamp 1698175906
transform -1 0 28000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._160__283
timestamp 1698175906
transform -1 0 39760 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._160_
timestamp 1698175906
transform 1 0 38640 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._161_
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._161__284
timestamp 1698175906
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._162_
timestamp 1698175906
transform 1 0 12656 0 -1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._162__285
timestamp 1698175906
transform 1 0 12208 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._163__286
timestamp 1698175906
transform -1 0 20944 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._163_
timestamp 1698175906
transform 1 0 20496 0 -1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._164__287
timestamp 1698175906
transform -1 0 40432 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._164_
timestamp 1698175906
transform 1 0 39200 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._165__288
timestamp 1698175906
transform -1 0 34496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._165_
timestamp 1698175906
transform 1 0 33264 0 -1 21952
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._166__289
timestamp 1698175906
transform -1 0 15232 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._166_
timestamp 1698175906
transform 1 0 14672 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  u_adc_reg.u_reg_0._167_
timestamp 1698175906
transform 1 0 24864 0 1 20384
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  u_adc_reg.u_reg_0._167__290
timestamp 1698175906
transform -1 0 25536 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_20  wire26
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 7030 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  wire114
timestamp 1698175906
transform 1 0 27216 0 -1 21952
box -86 -86 1654 870
<< labels >>
flabel metal4 s 4258 3076 4958 56508 0 FreeSans 5120 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 13258 3076 13958 56508 0 FreeSans 5120 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 22258 3076 22958 56508 0 FreeSans 5120 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 31258 3076 31958 56508 0 FreeSans 5120 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 40258 3076 40958 56508 0 FreeSans 5120 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 49258 3076 49958 56508 0 FreeSans 5120 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 58258 3076 58958 56508 0 FreeSans 5120 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 67258 3076 67958 56508 0 FreeSans 5120 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 76258 3076 76958 56508 0 FreeSans 5120 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 85258 3076 85958 56508 0 FreeSans 5120 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 94258 3076 94958 56508 0 FreeSans 5120 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 8758 3076 9458 56508 0 FreeSans 5120 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 17758 3076 18458 56508 0 FreeSans 5120 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 26758 3076 27458 56508 0 FreeSans 5120 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 35758 3076 36458 56508 0 FreeSans 5120 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 44758 3076 45458 56508 0 FreeSans 5120 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 53758 3076 54458 56508 0 FreeSans 5120 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 62758 3076 63458 56508 0 FreeSans 5120 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 71758 3076 72458 56508 0 FreeSans 5120 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 80758 3076 81458 56508 0 FreeSans 5120 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal4 s 89758 3076 90458 56508 0 FreeSans 5120 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal2 s 93856 0 93968 800 0 FreeSans 448 90 0 0 analog_dac_out
port 2 nsew signal input
flabel metal2 s 82880 0 82992 800 0 FreeSans 448 90 0 0 analog_din[0]
port 3 nsew signal input
flabel metal2 s 71904 0 72016 800 0 FreeSans 448 90 0 0 analog_din[1]
port 4 nsew signal input
flabel metal2 s 60928 0 61040 800 0 FreeSans 448 90 0 0 analog_din[2]
port 5 nsew signal input
flabel metal2 s 49952 0 50064 800 0 FreeSans 448 90 0 0 analog_din[3]
port 6 nsew signal input
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 analog_din[4]
port 7 nsew signal input
flabel metal2 s 28000 0 28112 800 0 FreeSans 448 90 0 0 analog_din[5]
port 8 nsew signal input
flabel metal3 s 0 4032 800 4144 0 FreeSans 448 0 0 0 clk
port 9 nsew signal input
flabel metal2 s 17024 0 17136 800 0 FreeSans 448 90 0 0 pulse1m_mclk
port 10 nsew signal input
flabel metal3 s 99200 58464 100000 58576 0 FreeSans 448 0 0 0 reg_ack
port 11 nsew signal tristate
flabel metal3 s 0 15232 800 15344 0 FreeSans 448 0 0 0 reg_addr[0]
port 12 nsew signal input
flabel metal3 s 0 14112 800 14224 0 FreeSans 448 0 0 0 reg_addr[1]
port 13 nsew signal input
flabel metal3 s 0 12992 800 13104 0 FreeSans 448 0 0 0 reg_addr[2]
port 14 nsew signal input
flabel metal3 s 0 11872 800 11984 0 FreeSans 448 0 0 0 reg_addr[3]
port 15 nsew signal input
flabel metal3 s 0 10752 800 10864 0 FreeSans 448 0 0 0 reg_addr[4]
port 16 nsew signal input
flabel metal3 s 0 9632 800 9744 0 FreeSans 448 0 0 0 reg_addr[5]
port 17 nsew signal input
flabel metal3 s 0 8512 800 8624 0 FreeSans 448 0 0 0 reg_addr[6]
port 18 nsew signal input
flabel metal3 s 0 7392 800 7504 0 FreeSans 448 0 0 0 reg_addr[7]
port 19 nsew signal input
flabel metal3 s 0 19712 800 19824 0 FreeSans 448 0 0 0 reg_be[0]
port 20 nsew signal input
flabel metal3 s 0 18592 800 18704 0 FreeSans 448 0 0 0 reg_be[1]
port 21 nsew signal input
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 reg_be[2]
port 22 nsew signal input
flabel metal3 s 0 16352 800 16464 0 FreeSans 448 0 0 0 reg_be[3]
port 23 nsew signal input
flabel metal3 s 0 5152 800 5264 0 FreeSans 448 0 0 0 reg_cs
port 24 nsew signal input
flabel metal3 s 99200 56672 100000 56784 0 FreeSans 448 0 0 0 reg_rdata[0]
port 25 nsew signal tristate
flabel metal3 s 99200 38752 100000 38864 0 FreeSans 448 0 0 0 reg_rdata[10]
port 26 nsew signal tristate
flabel metal3 s 99200 36960 100000 37072 0 FreeSans 448 0 0 0 reg_rdata[11]
port 27 nsew signal tristate
flabel metal3 s 99200 35168 100000 35280 0 FreeSans 448 0 0 0 reg_rdata[12]
port 28 nsew signal tristate
flabel metal3 s 99200 33376 100000 33488 0 FreeSans 448 0 0 0 reg_rdata[13]
port 29 nsew signal tristate
flabel metal3 s 99200 31584 100000 31696 0 FreeSans 448 0 0 0 reg_rdata[14]
port 30 nsew signal tristate
flabel metal3 s 99200 29792 100000 29904 0 FreeSans 448 0 0 0 reg_rdata[15]
port 31 nsew signal tristate
flabel metal3 s 99200 28000 100000 28112 0 FreeSans 448 0 0 0 reg_rdata[16]
port 32 nsew signal tristate
flabel metal3 s 99200 26208 100000 26320 0 FreeSans 448 0 0 0 reg_rdata[17]
port 33 nsew signal tristate
flabel metal3 s 99200 24416 100000 24528 0 FreeSans 448 0 0 0 reg_rdata[18]
port 34 nsew signal tristate
flabel metal3 s 99200 22624 100000 22736 0 FreeSans 448 0 0 0 reg_rdata[19]
port 35 nsew signal tristate
flabel metal3 s 99200 54880 100000 54992 0 FreeSans 448 0 0 0 reg_rdata[1]
port 36 nsew signal tristate
flabel metal3 s 99200 20832 100000 20944 0 FreeSans 448 0 0 0 reg_rdata[20]
port 37 nsew signal tristate
flabel metal3 s 99200 19040 100000 19152 0 FreeSans 448 0 0 0 reg_rdata[21]
port 38 nsew signal tristate
flabel metal3 s 99200 17248 100000 17360 0 FreeSans 448 0 0 0 reg_rdata[22]
port 39 nsew signal tristate
flabel metal3 s 99200 15456 100000 15568 0 FreeSans 448 0 0 0 reg_rdata[23]
port 40 nsew signal tristate
flabel metal3 s 99200 13664 100000 13776 0 FreeSans 448 0 0 0 reg_rdata[24]
port 41 nsew signal tristate
flabel metal3 s 99200 11872 100000 11984 0 FreeSans 448 0 0 0 reg_rdata[25]
port 42 nsew signal tristate
flabel metal3 s 99200 10080 100000 10192 0 FreeSans 448 0 0 0 reg_rdata[26]
port 43 nsew signal tristate
flabel metal3 s 99200 8288 100000 8400 0 FreeSans 448 0 0 0 reg_rdata[27]
port 44 nsew signal tristate
flabel metal3 s 99200 6496 100000 6608 0 FreeSans 448 0 0 0 reg_rdata[28]
port 45 nsew signal tristate
flabel metal3 s 99200 4704 100000 4816 0 FreeSans 448 0 0 0 reg_rdata[29]
port 46 nsew signal tristate
flabel metal3 s 99200 53088 100000 53200 0 FreeSans 448 0 0 0 reg_rdata[2]
port 47 nsew signal tristate
flabel metal3 s 99200 2912 100000 3024 0 FreeSans 448 0 0 0 reg_rdata[30]
port 48 nsew signal tristate
flabel metal3 s 99200 1120 100000 1232 0 FreeSans 448 0 0 0 reg_rdata[31]
port 49 nsew signal tristate
flabel metal3 s 99200 51296 100000 51408 0 FreeSans 448 0 0 0 reg_rdata[3]
port 50 nsew signal tristate
flabel metal3 s 99200 49504 100000 49616 0 FreeSans 448 0 0 0 reg_rdata[4]
port 51 nsew signal tristate
flabel metal3 s 99200 47712 100000 47824 0 FreeSans 448 0 0 0 reg_rdata[5]
port 52 nsew signal tristate
flabel metal3 s 99200 45920 100000 46032 0 FreeSans 448 0 0 0 reg_rdata[6]
port 53 nsew signal tristate
flabel metal3 s 99200 44128 100000 44240 0 FreeSans 448 0 0 0 reg_rdata[7]
port 54 nsew signal tristate
flabel metal3 s 99200 42336 100000 42448 0 FreeSans 448 0 0 0 reg_rdata[8]
port 55 nsew signal tristate
flabel metal3 s 99200 40544 100000 40656 0 FreeSans 448 0 0 0 reg_rdata[9]
port 56 nsew signal tristate
flabel metal3 s 0 55552 800 55664 0 FreeSans 448 0 0 0 reg_wdata[0]
port 57 nsew signal input
flabel metal3 s 0 44352 800 44464 0 FreeSans 448 0 0 0 reg_wdata[10]
port 58 nsew signal input
flabel metal3 s 0 43232 800 43344 0 FreeSans 448 0 0 0 reg_wdata[11]
port 59 nsew signal input
flabel metal3 s 0 42112 800 42224 0 FreeSans 448 0 0 0 reg_wdata[12]
port 60 nsew signal input
flabel metal3 s 0 40992 800 41104 0 FreeSans 448 0 0 0 reg_wdata[13]
port 61 nsew signal input
flabel metal3 s 0 39872 800 39984 0 FreeSans 448 0 0 0 reg_wdata[14]
port 62 nsew signal input
flabel metal3 s 0 38752 800 38864 0 FreeSans 448 0 0 0 reg_wdata[15]
port 63 nsew signal input
flabel metal3 s 0 37632 800 37744 0 FreeSans 448 0 0 0 reg_wdata[16]
port 64 nsew signal input
flabel metal3 s 0 36512 800 36624 0 FreeSans 448 0 0 0 reg_wdata[17]
port 65 nsew signal input
flabel metal3 s 0 35392 800 35504 0 FreeSans 448 0 0 0 reg_wdata[18]
port 66 nsew signal input
flabel metal3 s 0 34272 800 34384 0 FreeSans 448 0 0 0 reg_wdata[19]
port 67 nsew signal input
flabel metal3 s 0 54432 800 54544 0 FreeSans 448 0 0 0 reg_wdata[1]
port 68 nsew signal input
flabel metal3 s 0 33152 800 33264 0 FreeSans 448 0 0 0 reg_wdata[20]
port 69 nsew signal input
flabel metal3 s 0 32032 800 32144 0 FreeSans 448 0 0 0 reg_wdata[21]
port 70 nsew signal input
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 reg_wdata[22]
port 71 nsew signal input
flabel metal3 s 0 29792 800 29904 0 FreeSans 448 0 0 0 reg_wdata[23]
port 72 nsew signal input
flabel metal3 s 0 28672 800 28784 0 FreeSans 448 0 0 0 reg_wdata[24]
port 73 nsew signal input
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 reg_wdata[25]
port 74 nsew signal input
flabel metal3 s 0 26432 800 26544 0 FreeSans 448 0 0 0 reg_wdata[26]
port 75 nsew signal input
flabel metal3 s 0 25312 800 25424 0 FreeSans 448 0 0 0 reg_wdata[27]
port 76 nsew signal input
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 reg_wdata[28]
port 77 nsew signal input
flabel metal3 s 0 23072 800 23184 0 FreeSans 448 0 0 0 reg_wdata[29]
port 78 nsew signal input
flabel metal3 s 0 53312 800 53424 0 FreeSans 448 0 0 0 reg_wdata[2]
port 79 nsew signal input
flabel metal3 s 0 21952 800 22064 0 FreeSans 448 0 0 0 reg_wdata[30]
port 80 nsew signal input
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 reg_wdata[31]
port 81 nsew signal input
flabel metal3 s 0 52192 800 52304 0 FreeSans 448 0 0 0 reg_wdata[3]
port 82 nsew signal input
flabel metal3 s 0 51072 800 51184 0 FreeSans 448 0 0 0 reg_wdata[4]
port 83 nsew signal input
flabel metal3 s 0 49952 800 50064 0 FreeSans 448 0 0 0 reg_wdata[5]
port 84 nsew signal input
flabel metal3 s 0 48832 800 48944 0 FreeSans 448 0 0 0 reg_wdata[6]
port 85 nsew signal input
flabel metal3 s 0 47712 800 47824 0 FreeSans 448 0 0 0 reg_wdata[7]
port 86 nsew signal input
flabel metal3 s 0 46592 800 46704 0 FreeSans 448 0 0 0 reg_wdata[8]
port 87 nsew signal input
flabel metal3 s 0 45472 800 45584 0 FreeSans 448 0 0 0 reg_wdata[9]
port 88 nsew signal input
flabel metal3 s 0 6272 800 6384 0 FreeSans 448 0 0 0 reg_wr
port 89 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 reset_n
port 90 nsew signal input
flabel metal2 s 92960 59200 93072 60000 0 FreeSans 448 90 0 0 sar2dac[0]
port 91 nsew signal tristate
flabel metal2 s 80640 59200 80752 60000 0 FreeSans 448 90 0 0 sar2dac[1]
port 92 nsew signal tristate
flabel metal2 s 68320 59200 68432 60000 0 FreeSans 448 90 0 0 sar2dac[2]
port 93 nsew signal tristate
flabel metal2 s 56000 59200 56112 60000 0 FreeSans 448 90 0 0 sar2dac[3]
port 94 nsew signal tristate
flabel metal2 s 43680 59200 43792 60000 0 FreeSans 448 90 0 0 sar2dac[4]
port 95 nsew signal tristate
flabel metal2 s 31360 59200 31472 60000 0 FreeSans 448 90 0 0 sar2dac[5]
port 96 nsew signal tristate
flabel metal2 s 19040 59200 19152 60000 0 FreeSans 448 90 0 0 sar2dac[6]
port 97 nsew signal tristate
flabel metal2 s 6720 59200 6832 60000 0 FreeSans 448 90 0 0 sar2dac[7]
port 98 nsew signal tristate
rlabel metal1 49952 55664 49952 55664 0 VDD
rlabel metal1 49952 56448 49952 56448 0 VSS
rlabel metal2 76104 4592 76104 4592 0 COMP_0.Q
rlabel metal2 88200 10080 88200 10080 0 COMP_0.net1
rlabel metal3 83384 6664 83384 6664 0 COMP_0.net2
rlabel metal2 84112 10024 84112 10024 0 COMP_0.net3
rlabel metal2 78904 13104 78904 13104 0 COMP_0.net4
rlabel metal2 75880 3360 75880 3360 0 COMP_0.net7
rlabel metal2 72744 4984 72744 4984 0 COMP_1.Q
rlabel metal2 77112 5936 77112 5936 0 COMP_1.net1
rlabel metal2 81648 4312 81648 4312 0 COMP_1.net2
rlabel metal3 78960 5824 78960 5824 0 COMP_1.net3
rlabel metal2 70952 5096 70952 5096 0 COMP_1.net4
rlabel metal2 71848 3640 71848 3640 0 COMP_1.net7
rlabel metal2 61880 5096 61880 5096 0 COMP_2.Q
rlabel metal2 64456 6496 64456 6496 0 COMP_2.net1
rlabel metal3 59304 6664 59304 6664 0 COMP_2.net2
rlabel metal2 60088 4536 60088 4536 0 COMP_2.net3
rlabel metal3 63784 5096 63784 5096 0 COMP_2.net4
rlabel metal2 62440 6216 62440 6216 0 COMP_2.net7
rlabel metal2 50792 5376 50792 5376 0 COMP_3.Q
rlabel metal2 51352 8176 51352 8176 0 COMP_3.net1
rlabel metal2 47880 9688 47880 9688 0 COMP_3.net2
rlabel metal2 50344 4200 50344 4200 0 COMP_3.net3
rlabel metal2 49896 4816 49896 4816 0 COMP_3.net4
rlabel metal2 46312 5432 46312 5432 0 COMP_3.net7
rlabel metal2 44856 4144 44856 4144 0 COMP_4.Q
rlabel metal2 43904 15176 43904 15176 0 COMP_4.net1
rlabel metal3 43820 3304 43820 3304 0 COMP_4.net2
rlabel metal2 41944 4368 41944 4368 0 COMP_4.net3
rlabel metal2 42392 4368 42392 4368 0 COMP_4.net4
rlabel metal3 43960 3752 43960 3752 0 COMP_4.net7
rlabel metal2 37128 5768 37128 5768 0 COMP_5.Q
rlabel metal2 27608 6160 27608 6160 0 COMP_5.net1
rlabel metal2 34888 9912 34888 9912 0 COMP_5.net2
rlabel metal2 33432 3808 33432 3808 0 COMP_5.net3
rlabel metal2 34608 4536 34608 4536 0 COMP_5.net4
rlabel metal2 37016 5824 37016 5824 0 COMP_5.net7
rlabel metal2 50344 51352 50344 51352 0 CTRL._000_
rlabel metal3 68712 53592 68712 53592 0 CTRL._001_
rlabel metal2 66024 53256 66024 53256 0 CTRL._002_
rlabel metal2 57400 51296 57400 51296 0 CTRL._003_
rlabel metal2 41104 51688 41104 51688 0 CTRL._004_
rlabel metal2 32984 50512 32984 50512 0 CTRL._005_
rlabel metal2 29680 49896 29680 49896 0 CTRL._006_
rlabel metal2 26264 50904 26264 50904 0 CTRL._007_
rlabel metal2 48888 54936 48888 54936 0 CTRL._008_
rlabel metal2 51800 54824 51800 54824 0 CTRL._009_
rlabel metal2 60536 54824 60536 54824 0 CTRL._010_
rlabel metal2 62664 52472 62664 52472 0 CTRL._011_
rlabel metal2 41384 54936 41384 54936 0 CTRL._012_
rlabel metal2 34552 54488 34552 54488 0 CTRL._013_
rlabel metal2 30072 54488 30072 54488 0 CTRL._014_
rlabel metal2 25144 52528 25144 52528 0 CTRL._015_
rlabel metal2 30072 52472 30072 52472 0 CTRL._016_
rlabel metal2 27944 52752 27944 52752 0 CTRL._017_
rlabel metal3 27384 52024 27384 52024 0 CTRL._018_
rlabel metal2 27720 52976 27720 52976 0 CTRL._019_
rlabel metal2 50792 52360 50792 52360 0 CTRL._020_
rlabel metal2 52696 54768 52696 54768 0 CTRL._021_
rlabel metal2 50792 53256 50792 53256 0 CTRL._022_
rlabel metal2 43960 52024 43960 52024 0 CTRL._023_
rlabel metal2 43736 52808 43736 52808 0 CTRL._024_
rlabel metal2 52920 54712 52920 54712 0 CTRL._025_
rlabel metal2 47768 54656 47768 54656 0 CTRL._026_
rlabel metal2 47320 53816 47320 53816 0 CTRL._027_
rlabel metal2 46424 51688 46424 51688 0 CTRL._028_
rlabel metal2 49168 52248 49168 52248 0 CTRL._029_
rlabel metal2 41384 51352 41384 51352 0 CTRL._030_
rlabel metal2 46760 53088 46760 53088 0 CTRL._031_
rlabel metal3 47096 51352 47096 51352 0 CTRL._032_
rlabel metal2 50232 53592 50232 53592 0 CTRL._033_
rlabel metal2 48944 54488 48944 54488 0 CTRL._034_
rlabel metal2 49336 53144 49336 53144 0 CTRL._035_
rlabel metal3 54292 55048 54292 55048 0 CTRL._036_
rlabel metal3 61376 53480 61376 53480 0 CTRL._037_
rlabel metal2 57848 52976 57848 52976 0 CTRL._038_
rlabel metal2 58408 54824 58408 54824 0 CTRL._039_
rlabel metal3 62776 53816 62776 53816 0 CTRL._040_
rlabel metal2 56840 53984 56840 53984 0 CTRL._041_
rlabel metal2 57288 52920 57288 52920 0 CTRL._042_
rlabel metal2 55720 52192 55720 52192 0 CTRL._043_
rlabel metal2 40936 53200 40936 53200 0 CTRL._044_
rlabel metal2 40824 54712 40824 54712 0 CTRL._045_
rlabel metal2 41328 52920 41328 52920 0 CTRL._046_
rlabel metal2 35112 53760 35112 53760 0 CTRL._047_
rlabel metal2 35224 53256 35224 53256 0 CTRL._048_
rlabel metal2 33320 52472 33320 52472 0 CTRL._049_
rlabel metal2 29624 53088 29624 53088 0 CTRL._050_
rlabel metal3 30352 53480 30352 53480 0 CTRL._051_
rlabel metal3 48160 52136 48160 52136 0 CTRL.cmp
rlabel metal2 39928 51240 39928 51240 0 CTRL.done
rlabel metal2 53928 54040 53928 54040 0 CTRL.next\[0\]
rlabel metal2 58408 54320 58408 54320 0 CTRL.next\[1\]
rlabel metal3 59584 52248 59584 52248 0 CTRL.next\[2\]
rlabel metal3 44632 54544 44632 54544 0 CTRL.next\[3\]
rlabel metal2 39256 53424 39256 53424 0 CTRL.next\[4\]
rlabel metal2 35448 53200 35448 53200 0 CTRL.next\[5\]
rlabel metal3 24948 52248 24948 52248 0 CTRL.next\[6\]
rlabel metal2 41272 50848 41272 50848 0 CTRL.nstate\[0\]
rlabel metal2 46872 51016 46872 51016 0 CTRL.nstate\[1\]
rlabel metal2 55328 37464 55328 37464 0 CTRL.out\[0\]
rlabel metal2 67256 53368 67256 53368 0 CTRL.out\[1\]
rlabel metal2 68152 52752 68152 52752 0 CTRL.out\[2\]
rlabel metal2 55496 50960 55496 50960 0 CTRL.out\[3\]
rlabel metal2 42616 49784 42616 49784 0 CTRL.out\[4\]
rlabel metal2 39424 46424 39424 46424 0 CTRL.out\[5\]
rlabel metal2 66136 39200 66136 39200 0 CTRL.out\[6\]
rlabel metal2 44800 40264 44800 40264 0 CTRL.out\[7\]
rlabel metal2 51688 53368 51688 53368 0 CTRL.outn\[0\]
rlabel metal2 68376 54544 68376 54544 0 CTRL.outn\[1\]
rlabel metal3 66080 53704 66080 53704 0 CTRL.outn\[2\]
rlabel metal2 55832 53424 55832 53424 0 CTRL.outn\[3\]
rlabel metal2 42728 53368 42728 53368 0 CTRL.outn\[4\]
rlabel metal2 33264 52136 33264 52136 0 CTRL.outn\[5\]
rlabel metal2 25816 54096 25816 54096 0 CTRL.outn\[6\]
rlabel metal2 26600 54152 26600 54152 0 CTRL.outn\[7\]
rlabel metal3 48888 54600 48888 54600 0 CTRL.shift\[0\]
rlabel metal2 41048 51128 41048 51128 0 CTRL.start
rlabel metal2 44296 51072 44296 51072 0 CTRL.state\[0\]
rlabel metal2 50008 51688 50008 51688 0 CTRL.state\[1\]
rlabel metal2 46088 11760 46088 11760 0 _00_
rlabel metal2 45640 8904 45640 8904 0 _02_
rlabel metal2 45416 8736 45416 8736 0 _03_
rlabel metal3 47544 8232 47544 8232 0 _04_
rlabel metal2 45752 9912 45752 9912 0 _05_
rlabel metal2 94080 3640 94080 3640 0 analog_dac_out
rlabel metal2 82936 2142 82936 2142 0 analog_din[0]
rlabel metal2 74424 4256 74424 4256 0 analog_din[1]
rlabel metal2 60984 2058 60984 2058 0 analog_din[2]
rlabel metal2 50176 2184 50176 2184 0 analog_din[3]
rlabel metal3 39424 3416 39424 3416 0 analog_din[4]
rlabel metal2 28224 3416 28224 3416 0 analog_din[5]
rlabel metal3 21112 14504 21112 14504 0 clk
rlabel metal2 76216 6328 76216 6328 0 clknet_0_COMP_0.Q
rlabel metal2 82264 11648 82264 11648 0 clknet_0_COMP_0.net1
rlabel metal2 81704 7588 81704 7588 0 clknet_0_COMP_0.net2
rlabel metal3 82992 9016 82992 9016 0 clknet_0_COMP_0.net3
rlabel metal2 85176 10248 85176 10248 0 clknet_0_COMP_0.net4
rlabel metal3 67256 6552 67256 6552 0 clknet_0_COMP_1.Q
rlabel metal3 77616 9016 77616 9016 0 clknet_0_COMP_1.net1
rlabel metal2 81984 8008 81984 8008 0 clknet_0_COMP_1.net2
rlabel metal2 84000 7448 84000 7448 0 clknet_0_COMP_1.net3
rlabel metal2 76104 11424 76104 11424 0 clknet_0_COMP_1.net4
rlabel metal2 64680 6384 64680 6384 0 clknet_0_COMP_2.Q
rlabel metal2 68880 5992 68880 5992 0 clknet_0_COMP_2.net1
rlabel metal2 64344 8288 64344 8288 0 clknet_0_COMP_2.net2
rlabel metal2 63112 8512 63112 8512 0 clknet_0_COMP_2.net3
rlabel metal2 66248 7952 66248 7952 0 clknet_0_COMP_2.net4
rlabel metal2 55384 6720 55384 6720 0 clknet_0_COMP_3.Q
rlabel metal3 52808 4368 52808 4368 0 clknet_0_COMP_3.net1
rlabel metal3 52416 7448 52416 7448 0 clknet_0_COMP_3.net2
rlabel metal2 54488 6664 54488 6664 0 clknet_0_COMP_3.net3
rlabel metal3 54488 5208 54488 5208 0 clknet_0_COMP_3.net4
rlabel metal2 41944 6664 41944 6664 0 clknet_0_COMP_4.Q
rlabel metal2 43176 6720 43176 6720 0 clknet_0_COMP_4.net1
rlabel metal2 47208 11312 47208 11312 0 clknet_0_COMP_4.net2
rlabel metal3 42616 5208 42616 5208 0 clknet_0_COMP_4.net3
rlabel metal2 46424 8680 46424 8680 0 clknet_0_COMP_4.net4
rlabel metal2 40040 8960 40040 8960 0 clknet_0_COMP_5.Q
rlabel metal2 31136 11368 31136 11368 0 clknet_0_COMP_5.net1
rlabel metal2 37240 11088 37240 11088 0 clknet_0_COMP_5.net2
rlabel metal3 30240 9688 30240 9688 0 clknet_0_COMP_5.net3
rlabel metal3 33600 9016 33600 9016 0 clknet_0_COMP_5.net4
rlabel metal3 45808 53032 45808 53032 0 clknet_0_CTRL.cmp
rlabel metal2 44184 20160 44184 20160 0 clknet_0_clk
rlabel metal2 65576 12264 65576 12264 0 clknet_1_0__leaf_COMP_0.Q
rlabel metal2 80472 13384 80472 13384 0 clknet_1_0__leaf_COMP_0.net1
rlabel metal2 77280 5880 77280 5880 0 clknet_1_0__leaf_COMP_0.net2
rlabel metal2 78288 11144 78288 11144 0 clknet_1_0__leaf_COMP_0.net3
rlabel metal2 91224 8344 91224 8344 0 clknet_1_0__leaf_COMP_0.net4
rlabel metal2 53480 9520 53480 9520 0 clknet_1_0__leaf_COMP_1.Q
rlabel metal2 71456 14504 71456 14504 0 clknet_1_0__leaf_COMP_1.net1
rlabel metal2 69720 12488 69720 12488 0 clknet_1_0__leaf_COMP_1.net2
rlabel metal2 74088 7000 74088 7000 0 clknet_1_0__leaf_COMP_1.net3
rlabel metal2 71288 9072 71288 9072 0 clknet_1_0__leaf_COMP_1.net4
rlabel metal2 51240 10640 51240 10640 0 clknet_1_0__leaf_COMP_2.Q
rlabel metal2 65800 7896 65800 7896 0 clknet_1_0__leaf_COMP_2.net1
rlabel metal2 60480 13720 60480 13720 0 clknet_1_0__leaf_COMP_2.net2
rlabel metal2 59864 7784 59864 7784 0 clknet_1_0__leaf_COMP_2.net3
rlabel metal2 60536 4704 60536 4704 0 clknet_1_0__leaf_COMP_2.net4
rlabel metal2 49112 6384 49112 6384 0 clknet_1_0__leaf_COMP_3.Q
rlabel metal2 48104 10136 48104 10136 0 clknet_1_0__leaf_COMP_3.net1
rlabel metal2 51128 11144 51128 11144 0 clknet_1_0__leaf_COMP_3.net2
rlabel metal2 49448 4704 49448 4704 0 clknet_1_0__leaf_COMP_3.net3
rlabel metal2 50120 4928 50120 4928 0 clknet_1_0__leaf_COMP_3.net4
rlabel metal3 40404 7448 40404 7448 0 clknet_1_0__leaf_COMP_4.Q
rlabel metal2 44072 5656 44072 5656 0 clknet_1_0__leaf_COMP_4.net1
rlabel metal2 41216 15176 41216 15176 0 clknet_1_0__leaf_COMP_4.net2
rlabel metal2 41720 4816 41720 4816 0 clknet_1_0__leaf_COMP_4.net3
rlabel metal2 41272 4984 41272 4984 0 clknet_1_0__leaf_COMP_4.net4
rlabel metal2 37128 8120 37128 8120 0 clknet_1_0__leaf_COMP_5.Q
rlabel metal2 34216 5656 34216 5656 0 clknet_1_0__leaf_COMP_5.net1
rlabel metal2 26824 6552 26824 6552 0 clknet_1_0__leaf_COMP_5.net2
rlabel metal2 34104 4816 34104 4816 0 clknet_1_0__leaf_COMP_5.net3
rlabel metal2 33992 4200 33992 4200 0 clknet_1_0__leaf_COMP_5.net4
rlabel metal2 41944 52976 41944 52976 0 clknet_1_0__leaf_CTRL.cmp
rlabel metal2 75544 5096 75544 5096 0 clknet_1_1__leaf_COMP_0.Q
rlabel metal3 83608 9688 83608 9688 0 clknet_1_1__leaf_COMP_0.net1
rlabel metal2 82880 15176 82880 15176 0 clknet_1_1__leaf_COMP_0.net2
rlabel metal2 77056 13720 77056 13720 0 clknet_1_1__leaf_COMP_0.net3
rlabel metal2 86184 7336 86184 7336 0 clknet_1_1__leaf_COMP_0.net4
rlabel metal2 71400 7784 71400 7784 0 clknet_1_1__leaf_COMP_1.Q
rlabel metal2 71232 3528 71232 3528 0 clknet_1_1__leaf_COMP_1.net1
rlabel metal2 71064 7784 71064 7784 0 clknet_1_1__leaf_COMP_1.net2
rlabel metal2 81592 6328 81592 6328 0 clknet_1_1__leaf_COMP_1.net3
rlabel metal2 70280 6272 70280 6272 0 clknet_1_1__leaf_COMP_1.net4
rlabel metal2 59192 7896 59192 7896 0 clknet_1_1__leaf_COMP_2.Q
rlabel metal2 62552 6272 62552 6272 0 clknet_1_1__leaf_COMP_2.net1
rlabel metal2 62440 9016 62440 9016 0 clknet_1_1__leaf_COMP_2.net2
rlabel metal4 75656 4687 75656 4687 0 clknet_1_1__leaf_COMP_2.net3
rlabel metal2 63896 7056 63896 7056 0 clknet_1_1__leaf_COMP_2.net4
rlabel metal2 52136 11872 52136 11872 0 clknet_1_1__leaf_COMP_3.Q
rlabel metal2 46200 6608 46200 6608 0 clknet_1_1__leaf_COMP_3.net1
rlabel metal2 49336 5656 49336 5656 0 clknet_1_1__leaf_COMP_3.net2
rlabel metal2 50008 6272 50008 6272 0 clknet_1_1__leaf_COMP_3.net3
rlabel metal2 50232 8400 50232 8400 0 clknet_1_1__leaf_COMP_3.net4
rlabel metal2 46312 7392 46312 7392 0 clknet_1_1__leaf_COMP_4.Q
rlabel metal2 45192 4144 45192 4144 0 clknet_1_1__leaf_COMP_4.net1
rlabel metal2 42448 7448 42448 7448 0 clknet_1_1__leaf_COMP_4.net2
rlabel metal2 40936 6328 40936 6328 0 clknet_1_1__leaf_COMP_4.net3
rlabel metal2 42952 4256 42952 4256 0 clknet_1_1__leaf_COMP_4.net4
rlabel metal3 44464 8120 44464 8120 0 clknet_1_1__leaf_COMP_5.Q
rlabel metal2 37408 5320 37408 5320 0 clknet_1_1__leaf_COMP_5.net1
rlabel metal2 37464 7504 37464 7504 0 clknet_1_1__leaf_COMP_5.net2
rlabel metal3 35952 7560 35952 7560 0 clknet_1_1__leaf_COMP_5.net3
rlabel metal2 38080 5096 38080 5096 0 clknet_1_1__leaf_COMP_5.net4
rlabel metal2 48944 52920 48944 52920 0 clknet_1_1__leaf_CTRL.cmp
rlabel metal3 40656 49672 40656 49672 0 clknet_2_0__leaf_clk
rlabel metal2 26152 52136 26152 52136 0 clknet_2_1__leaf_clk
rlabel metal2 78120 3752 78120 3752 0 clknet_2_2__leaf_clk
rlabel metal2 69608 53200 69608 53200 0 clknet_2_3__leaf_clk
rlabel metal2 83272 4368 83272 4368 0 net1
rlabel metal3 17696 12264 17696 12264 0 net10
rlabel metal2 5768 26152 5768 26152 0 net100
rlabel metal3 29960 24808 29960 24808 0 net101
rlabel metal2 29736 21560 29736 21560 0 net102
rlabel metal3 47600 50456 47600 50456 0 net103
rlabel metal3 40488 48440 40488 48440 0 net104
rlabel metal2 69496 24080 69496 24080 0 net105
rlabel metal2 53200 29624 53200 29624 0 net106
rlabel metal2 56728 38360 56728 38360 0 net107
rlabel metal3 65884 50456 65884 50456 0 net108
rlabel metal2 76160 25480 76160 25480 0 net109
rlabel metal2 25816 32368 25816 32368 0 net11
rlabel metal2 74312 50960 74312 50960 0 net110
rlabel metal3 93968 49672 93968 49672 0 net111
rlabel metal2 74872 21504 74872 21504 0 net112
rlabel metal2 5880 21168 5880 21168 0 net113
rlabel metal2 28392 21616 28392 21616 0 net114
rlabel metal2 44968 5656 44968 5656 0 net115
rlabel metal2 75544 13664 75544 13664 0 net116
rlabel metal2 74536 5936 74536 5936 0 net117
rlabel metal3 78764 6104 78764 6104 0 net118
rlabel metal2 78232 6104 78232 6104 0 net119
rlabel metal2 27944 26040 27944 26040 0 net12
rlabel metal2 74872 6272 74872 6272 0 net120
rlabel metal2 75320 4536 75320 4536 0 net121
rlabel metal2 63560 4088 63560 4088 0 net122
rlabel metal2 62216 6944 62216 6944 0 net123
rlabel metal3 47880 3528 47880 3528 0 net124
rlabel metal2 49112 4872 49112 4872 0 net125
rlabel metal3 39816 3640 39816 3640 0 net126
rlabel metal2 41384 5936 41384 5936 0 net127
rlabel metal2 34328 4592 34328 4592 0 net128
rlabel metal2 33768 4200 33768 4200 0 net129
rlabel metal3 4480 22344 4480 22344 0 net13
rlabel metal2 48608 28392 48608 28392 0 net130
rlabel metal2 50232 29680 50232 29680 0 net131
rlabel metal2 40376 27888 40376 27888 0 net132
rlabel metal2 38920 33600 38920 33600 0 net133
rlabel metal2 55048 34832 55048 34832 0 net134
rlabel metal2 80808 43624 80808 43624 0 net135
rlabel metal2 69888 42728 69888 42728 0 net136
rlabel metal3 72296 37800 72296 37800 0 net137
rlabel metal2 62384 42728 62384 42728 0 net138
rlabel metal2 43624 44352 43624 44352 0 net139
rlabel metal2 2576 21224 2576 21224 0 net14
rlabel metal2 63112 37968 63112 37968 0 net140
rlabel metal3 43736 38920 43736 38920 0 net141
rlabel metal2 63224 33712 63224 33712 0 net142
rlabel metal2 80248 48496 80248 48496 0 net143
rlabel metal2 71064 47880 71064 47880 0 net144
rlabel metal2 78008 41608 78008 41608 0 net145
rlabel metal2 65464 50064 65464 50064 0 net146
rlabel metal2 43512 47488 43512 47488 0 net147
rlabel metal2 68488 35336 68488 35336 0 net148
rlabel metal2 44072 41832 44072 41832 0 net149
rlabel metal2 2072 18088 2072 18088 0 net15
rlabel metal3 53312 38920 53312 38920 0 net150
rlabel metal2 77056 50568 77056 50568 0 net151
rlabel metal2 70560 50568 70560 50568 0 net152
rlabel metal2 70840 41104 70840 41104 0 net153
rlabel metal2 60200 50568 60200 50568 0 net154
rlabel metal2 36456 47768 36456 47768 0 net155
rlabel metal2 58184 37940 58184 37940 0 net156
rlabel metal2 38584 41608 38584 41608 0 net157
rlabel metal2 49224 32592 49224 32592 0 net158
rlabel metal2 54936 48104 54936 48104 0 net159
rlabel metal3 4424 20776 4424 20776 0 net16
rlabel metal2 56728 43792 56728 43792 0 net160
rlabel metal2 58184 41216 58184 41216 0 net161
rlabel metal2 30968 46256 30968 46256 0 net162
rlabel metal2 31640 42840 31640 42840 0 net163
rlabel metal2 31136 39592 31136 39592 0 net164
rlabel metal2 31640 36568 31640 36568 0 net165
rlabel metal2 59976 31696 59976 31696 0 net166
rlabel metal3 80248 45864 80248 45864 0 net167
rlabel metal2 67592 46648 67592 46648 0 net168
rlabel metal2 79016 38780 79016 38780 0 net169
rlabel metal3 44576 25368 44576 25368 0 net17
rlabel metal2 60648 46536 60648 46536 0 net170
rlabel metal2 37464 44744 37464 44744 0 net171
rlabel metal2 63784 41104 63784 41104 0 net172
rlabel metal2 38584 38472 38584 38472 0 net173
rlabel metal2 55384 30072 55384 30072 0 net174
rlabel metal2 49000 48272 49000 48272 0 net175
rlabel metal2 50176 43512 50176 43512 0 net176
rlabel metal3 49280 40376 49280 40376 0 net177
rlabel metal2 25704 46200 25704 46200 0 net178
rlabel metal2 25368 43568 25368 43568 0 net179
rlabel metal3 7112 56168 7112 56168 0 net18
rlabel metal2 25480 40656 25480 40656 0 net180
rlabel metal2 26320 37240 26320 37240 0 net181
rlabel metal2 56112 29512 56112 29512 0 net182
rlabel metal2 54264 25872 54264 25872 0 net183
rlabel metal2 35336 28112 35336 28112 0 net184
rlabel metal2 9240 33096 9240 33096 0 net185
rlabel metal2 32536 34160 32536 34160 0 net186
rlabel metal2 26208 32536 26208 32536 0 net187
rlabel metal2 27384 34216 27384 34216 0 net188
rlabel metal2 5656 22792 5656 22792 0 net189
rlabel metal2 2016 45192 2016 45192 0 net19
rlabel metal2 1848 22904 1848 22904 0 net190
rlabel metal2 1904 19992 1904 19992 0 net191
rlabel metal2 5992 20720 5992 20720 0 net192
rlabel metal2 11704 50624 11704 50624 0 net193
rlabel metal2 1848 49056 1848 49056 0 net194
rlabel metal2 16632 50568 16632 50568 0 net195
rlabel metal2 5600 49784 5600 49784 0 net196
rlabel metal2 9072 49000 9072 49000 0 net197
rlabel metal2 2520 46928 2520 46928 0 net198
rlabel metal2 3080 45360 3080 45360 0 net199
rlabel metal2 83496 12096 83496 12096 0 net2
rlabel metal2 2072 43232 2072 43232 0 net20
rlabel metal2 2576 43512 2576 43512 0 net200
rlabel metal2 8904 41104 8904 41104 0 net201
rlabel metal2 2856 42224 2856 42224 0 net202
rlabel metal2 1848 40096 1848 40096 0 net203
rlabel metal2 2408 38080 2408 38080 0 net204
rlabel metal2 5656 39928 5656 39928 0 net205
rlabel metal2 2744 35952 2744 35952 0 net206
rlabel metal2 1848 34272 1848 34272 0 net207
rlabel metal2 11368 34384 11368 34384 0 net208
rlabel metal2 1848 31080 1848 31080 0 net209
rlabel metal2 2072 41944 2072 41944 0 net21
rlabel metal2 5096 34832 5096 34832 0 net210
rlabel metal2 5096 31696 5096 31696 0 net211
rlabel metal2 1960 29456 1960 29456 0 net212
rlabel metal2 20888 31024 20888 31024 0 net213
rlabel metal2 8680 30128 8680 30128 0 net214
rlabel metal2 18200 29456 18200 29456 0 net215
rlabel metal2 1960 27888 1960 27888 0 net216
rlabel metal2 7336 27720 7336 27720 0 net217
rlabel metal2 5320 25928 5320 25928 0 net218
rlabel metal2 1904 24696 1904 24696 0 net219
rlabel metal2 2800 40936 2800 40936 0 net22
rlabel metal2 15848 23800 15848 23800 0 net220
rlabel metal2 26600 23408 26600 23408 0 net221
rlabel metal2 29120 21560 29120 21560 0 net222
rlabel metal2 9912 21616 9912 21616 0 net223
rlabel metal2 19040 19992 19040 19992 0 net224
rlabel metal2 44296 25480 44296 25480 0 net225
rlabel metal2 49672 26320 49672 26320 0 net226
rlabel metal2 90496 35672 90496 35672 0 net227
rlabel metal2 86744 49672 86744 49672 0 net228
rlabel metal2 92344 48944 92344 48944 0 net229
rlabel metal2 2072 40768 2072 40768 0 net23
rlabel metal2 86632 43176 86632 43176 0 net230
rlabel metal2 86240 45864 86240 45864 0 net231
rlabel metal2 92008 46312 92008 46312 0 net232
rlabel metal2 91448 43568 91448 43568 0 net233
rlabel metal2 91896 39928 91896 39928 0 net234
rlabel metal2 82488 40656 82488 40656 0 net235
rlabel metal2 86408 39536 86408 39536 0 net236
rlabel metal3 84336 38920 84336 38920 0 net237
rlabel metal2 78120 35112 78120 35112 0 net238
rlabel metal2 84616 35280 84616 35280 0 net239
rlabel metal2 11816 36736 11816 36736 0 net24
rlabel metal2 72184 35336 72184 35336 0 net240
rlabel metal2 69048 31696 69048 31696 0 net241
rlabel metal2 65128 31080 65128 31080 0 net242
rlabel metal2 67816 28560 67816 28560 0 net243
rlabel metal3 63336 27048 63336 27048 0 net244
rlabel metal2 76216 28112 76216 28112 0 net245
rlabel metal2 71848 25424 71848 25424 0 net246
rlabel metal2 61768 24584 61768 24584 0 net247
rlabel metal2 66696 25536 66696 25536 0 net248
rlabel metal2 78512 25480 78512 25480 0 net249
rlabel metal2 2072 30968 2072 30968 0 net25
rlabel metal2 61768 21448 61768 21448 0 net250
rlabel metal2 78232 22232 78232 22232 0 net251
rlabel metal2 67144 22680 67144 22680 0 net252
rlabel metal2 72184 22792 72184 22792 0 net253
rlabel metal2 83048 22680 83048 22680 0 net254
rlabel metal2 85624 19320 85624 19320 0 net255
rlabel metal2 75992 19656 75992 19656 0 net256
rlabel metal2 71008 19208 71008 19208 0 net257
rlabel metal3 81032 20216 81032 20216 0 net258
rlabel metal2 20664 42224 20664 42224 0 net259
rlabel metal2 2128 36232 2128 36232 0 net26
rlabel metal2 9352 47208 9352 47208 0 net260
rlabel metal2 20832 48776 20832 48776 0 net261
rlabel metal2 8344 43904 8344 43904 0 net262
rlabel metal2 14168 48104 14168 48104 0 net263
rlabel metal2 14280 44744 14280 44744 0 net264
rlabel metal2 20776 44968 20776 44968 0 net265
rlabel metal2 13272 42392 13272 42392 0 net266
rlabel metal2 13384 39088 13384 39088 0 net267
rlabel metal2 19264 40376 19264 40376 0 net268
rlabel metal2 21616 38024 21616 38024 0 net269
rlabel metal3 4368 31752 4368 31752 0 net27
rlabel metal2 8456 36904 8456 36904 0 net270
rlabel metal2 14616 36400 14616 36400 0 net271
rlabel metal2 21224 35560 21224 35560 0 net272
rlabel metal2 20552 33376 20552 33376 0 net273
rlabel metal3 15064 32312 15064 32312 0 net274
rlabel metal2 26488 31248 26488 31248 0 net275
rlabel metal2 13496 29680 13496 29680 0 net276
rlabel metal2 32760 31248 32760 31248 0 net277
rlabel metal2 29176 28112 29176 28112 0 net278
rlabel metal2 24752 28392 24752 28392 0 net279
rlabel metal3 2408 34664 2408 34664 0 net28
rlabel metal2 14000 27048 14000 27048 0 net280
rlabel metal2 19712 26264 19712 26264 0 net281
rlabel metal2 26488 24976 26488 24976 0 net282
rlabel metal2 38920 23800 38920 23800 0 net283
rlabel metal2 32536 24752 32536 24752 0 net284
rlabel metal2 12488 24752 12488 24752 0 net285
rlabel metal2 20664 23408 20664 23408 0 net286
rlabel metal3 39704 20776 39704 20776 0 net287
rlabel metal2 33432 21840 33432 21840 0 net288
rlabel metal2 14952 21448 14952 21448 0 net289
rlabel metal2 2072 54376 2072 54376 0 net29
rlabel metal2 25200 20776 25200 20776 0 net290
rlabel metal2 77728 14056 77728 14056 0 net291
rlabel metal2 78288 4200 78288 4200 0 net292
rlabel metal2 74816 5320 74816 5320 0 net293
rlabel metal2 67984 5320 67984 5320 0 net294
rlabel metal2 58856 13608 58856 13608 0 net295
rlabel metal2 58184 5320 58184 5320 0 net296
rlabel metal2 45976 4312 45976 4312 0 net297
rlabel metal2 49784 9464 49784 9464 0 net298
rlabel metal2 41776 15288 41776 15288 0 net299
rlabel metal2 73976 5824 73976 5824 0 net3
rlabel metal3 2744 31864 2744 31864 0 net30
rlabel metal2 43512 4200 43512 4200 0 net300
rlabel metal2 30744 5992 30744 5992 0 net301
rlabel metal2 33432 5040 33432 5040 0 net302
rlabel metal2 77896 3752 77896 3752 0 net303
rlabel metal2 78400 11368 78400 11368 0 net304
rlabel metal2 70168 5600 70168 5600 0 net305
rlabel metal3 69048 3752 69048 3752 0 net306
rlabel metal2 59080 3696 59080 3696 0 net307
rlabel metal2 58240 3752 58240 3752 0 net308
rlabel metal2 47768 8232 47768 8232 0 net309
rlabel metal2 2184 31864 2184 31864 0 net31
rlabel metal2 46872 8008 46872 8008 0 net310
rlabel metal3 43176 3304 43176 3304 0 net311
rlabel metal2 42224 15400 42224 15400 0 net312
rlabel metal2 34216 6552 34216 6552 0 net313
rlabel metal2 27944 5824 27944 5824 0 net314
rlabel metal3 70728 3640 70728 3640 0 net315
rlabel metal2 45864 5880 45864 5880 0 net316
rlabel metal2 82488 4368 82488 4368 0 net317
rlabel metal2 71176 6944 71176 6944 0 net318
rlabel metal2 62888 5936 62888 5936 0 net319
rlabel metal2 2408 29568 2408 29568 0 net32
rlabel metal2 49616 5880 49616 5880 0 net320
rlabel metal3 44016 3528 44016 3528 0 net321
rlabel metal2 37688 5096 37688 5096 0 net322
rlabel metal2 77336 4480 77336 4480 0 net323
rlabel metal2 59640 6888 59640 6888 0 net324
rlabel metal2 41048 6664 41048 6664 0 net325
rlabel metal3 36064 6888 36064 6888 0 net326
rlabel metal2 45976 12040 45976 12040 0 net327
rlabel metal2 52696 30072 52696 30072 0 net328
rlabel metal3 78624 4424 78624 4424 0 net329
rlabel metal2 2072 29792 2072 29792 0 net33
rlabel metal2 2072 28560 2072 28560 0 net34
rlabel metal2 2128 26936 2128 26936 0 net35
rlabel metal2 2296 25760 2296 25760 0 net36
rlabel metal2 2072 25536 2072 25536 0 net37
rlabel metal2 2072 23520 2072 23520 0 net38
rlabel metal2 2744 22568 2744 22568 0 net39
rlabel metal2 61936 13832 61936 13832 0 net4
rlabel metal2 1960 51968 1960 51968 0 net40
rlabel metal2 1960 21840 1960 21840 0 net41
rlabel metal2 2240 21672 2240 21672 0 net42
rlabel metal2 2072 52360 2072 52360 0 net43
rlabel metal2 2296 50232 2296 50232 0 net44
rlabel metal2 2072 50400 2072 50400 0 net45
rlabel metal2 2744 46928 2744 46928 0 net46
rlabel metal2 2688 44744 2688 44744 0 net47
rlabel metal3 5236 47320 5236 47320 0 net48
rlabel metal2 2128 45640 2128 45640 0 net49
rlabel metal2 50232 3640 50232 3640 0 net5
rlabel metal2 2296 6384 2296 6384 0 net50
rlabel metal2 6440 21504 6440 21504 0 net51
rlabel metal2 96544 55048 96544 55048 0 net52
rlabel metal2 96488 38920 96488 38920 0 net53
rlabel metal2 96600 38752 96600 38752 0 net54
rlabel metal2 96600 36792 96600 36792 0 net55
rlabel metal2 96600 35224 96600 35224 0 net56
rlabel metal3 96824 34104 96824 34104 0 net57
rlabel metal2 96936 31640 96936 31640 0 net58
rlabel metal2 96936 30128 96936 30128 0 net59
rlabel metal2 44576 15400 44576 15400 0 net6
rlabel metal3 96824 28616 96824 28616 0 net60
rlabel metal2 96600 27216 96600 27216 0 net61
rlabel metal2 96936 25536 96936 25536 0 net62
rlabel metal2 76664 23520 76664 23520 0 net63
rlabel metal3 94024 51576 94024 51576 0 net64
rlabel metal2 96936 21672 96936 21672 0 net65
rlabel metal2 71512 21392 71512 21392 0 net66
rlabel metal2 96936 17528 96936 17528 0 net67
rlabel metal2 96824 16072 96824 16072 0 net68
rlabel metal3 96936 14448 96936 14448 0 net69
rlabel metal2 25928 5208 25928 5208 0 net7
rlabel metal3 81368 12208 81368 12208 0 net70
rlabel metal2 96936 10640 96936 10640 0 net71
rlabel metal3 92064 9240 92064 9240 0 net72
rlabel metal2 90440 17416 90440 17416 0 net73
rlabel metal3 81536 5432 81536 5432 0 net74
rlabel metal2 96600 52080 96600 52080 0 net75
rlabel metal2 75264 13944 75264 13944 0 net76
rlabel metal2 86072 16268 86072 16268 0 net77
rlabel metal2 96600 45304 96600 45304 0 net78
rlabel metal2 96600 49112 96600 49112 0 net79
rlabel metal2 38640 25032 38640 25032 0 net8
rlabel metal2 96600 47544 96600 47544 0 net80
rlabel metal2 95928 45416 95928 45416 0 net81
rlabel metal2 96936 43988 96936 43988 0 net82
rlabel metal2 96600 41440 96600 41440 0 net83
rlabel metal2 96656 40600 96656 40600 0 net84
rlabel metal2 82152 55384 82152 55384 0 net85
rlabel metal3 75208 55048 75208 55048 0 net86
rlabel metal2 67144 55608 67144 55608 0 net87
rlabel metal2 56056 55300 56056 55300 0 net88
rlabel metal2 43288 55608 43288 55608 0 net89
rlabel metal2 9800 23464 9800 23464 0 net9
rlabel metal2 32424 55608 32424 55608 0 net90
rlabel metal2 25480 55608 25480 55608 0 net91
rlabel metal2 8232 56000 8232 56000 0 net92
rlabel metal2 5656 24752 5656 24752 0 net93
rlabel metal2 5096 30408 5096 30408 0 net94
rlabel metal2 21784 21728 21784 21728 0 net95
rlabel metal2 5656 47992 5656 47992 0 net96
rlabel metal2 5768 46088 5768 46088 0 net97
rlabel metal2 24248 36232 24248 36232 0 net98
rlabel metal2 7000 43624 7000 43624 0 net99
rlabel metal2 17304 3360 17304 3360 0 pulse1m_mclk
rlabel metal2 97720 57400 97720 57400 0 reg_ack
rlabel metal2 1736 13384 1736 13384 0 reg_addr[2]
rlabel metal2 1736 12040 1736 12040 0 reg_addr[3]
rlabel metal2 1736 11032 1736 11032 0 reg_addr[4]
rlabel metal3 1246 9688 1246 9688 0 reg_addr[5]
rlabel metal2 1736 19488 1736 19488 0 reg_be[0]
rlabel metal2 2240 18424 2240 18424 0 reg_be[1]
rlabel metal3 1246 17528 1246 17528 0 reg_be[2]
rlabel metal2 1736 16632 1736 16632 0 reg_be[3]
rlabel metal3 1302 5208 1302 5208 0 reg_cs
rlabel metal2 95928 56336 95928 56336 0 reg_rdata[0]
rlabel metal2 98056 39144 98056 39144 0 reg_rdata[10]
rlabel metal2 98056 37072 98056 37072 0 reg_rdata[11]
rlabel metal2 97720 35336 97720 35336 0 reg_rdata[12]
rlabel metal2 97720 33656 97720 33656 0 reg_rdata[13]
rlabel metal3 98658 31640 98658 31640 0 reg_rdata[14]
rlabel metal2 98056 29960 98056 29960 0 reg_rdata[15]
rlabel metal2 97720 28336 97720 28336 0 reg_rdata[16]
rlabel metal2 97720 26600 97720 26600 0 reg_rdata[17]
rlabel metal2 98056 24528 98056 24528 0 reg_rdata[18]
rlabel metal2 98056 22848 98056 22848 0 reg_rdata[19]
rlabel metal2 98056 55048 98056 55048 0 reg_rdata[1]
rlabel metal2 98056 21168 98056 21168 0 reg_rdata[20]
rlabel metal3 98658 19096 98658 19096 0 reg_rdata[21]
rlabel metal2 98056 17416 98056 17416 0 reg_rdata[22]
rlabel metal2 98056 15736 98056 15736 0 reg_rdata[23]
rlabel metal2 98056 14056 98056 14056 0 reg_rdata[24]
rlabel metal2 98056 11984 98056 11984 0 reg_rdata[25]
rlabel metal2 98056 10304 98056 10304 0 reg_rdata[26]
rlabel metal3 98490 8344 98490 8344 0 reg_rdata[27]
rlabel metal3 98658 6552 98658 6552 0 reg_rdata[28]
rlabel metal2 97720 4928 97720 4928 0 reg_rdata[29]
rlabel metal2 98056 53368 98056 53368 0 reg_rdata[2]
rlabel metal2 97720 3192 97720 3192 0 reg_rdata[30]
rlabel metal2 97776 4088 97776 4088 0 reg_rdata[31]
rlabel metal2 97720 51744 97720 51744 0 reg_rdata[3]
rlabel metal2 98056 49616 98056 49616 0 reg_rdata[4]
rlabel metal2 98056 47936 98056 47936 0 reg_rdata[5]
rlabel metal2 98056 46256 98056 46256 0 reg_rdata[6]
rlabel metal3 98658 44184 98658 44184 0 reg_rdata[7]
rlabel metal2 98056 42504 98056 42504 0 reg_rdata[8]
rlabel metal2 98056 40824 98056 40824 0 reg_rdata[9]
rlabel metal2 1736 55832 1736 55832 0 reg_wdata[0]
rlabel metal2 1736 44744 1736 44744 0 reg_wdata[10]
rlabel metal3 1302 43288 1302 43288 0 reg_wdata[11]
rlabel metal2 1736 42392 1736 42392 0 reg_wdata[12]
rlabel metal3 1582 41048 1582 41048 0 reg_wdata[13]
rlabel metal2 1736 40488 1736 40488 0 reg_wdata[14]
rlabel metal3 1302 38808 1302 38808 0 reg_wdata[15]
rlabel metal2 1736 37800 1736 37800 0 reg_wdata[16]
rlabel metal2 1736 36512 1736 36512 0 reg_wdata[17]
rlabel metal2 1736 35560 1736 35560 0 reg_wdata[18]
rlabel metal2 1736 34552 1736 34552 0 reg_wdata[19]
rlabel metal2 1736 54824 1736 54824 0 reg_wdata[1]
rlabel metal3 1246 33208 1246 33208 0 reg_wdata[20]
rlabel metal2 1736 32312 1736 32312 0 reg_wdata[21]
rlabel metal2 1736 31304 1736 31304 0 reg_wdata[22]
rlabel metal2 1736 29960 1736 29960 0 reg_wdata[23]
rlabel metal2 1736 28672 1736 28672 0 reg_wdata[24]
rlabel metal2 1736 27328 1736 27328 0 reg_wdata[25]
rlabel metal2 2632 26768 2632 26768 0 reg_wdata[26]
rlabel metal3 1246 25368 1246 25368 0 reg_wdata[27]
rlabel metal2 1736 24080 1736 24080 0 reg_wdata[28]
rlabel metal2 2408 23660 2408 23660 0 reg_wdata[29]
rlabel metal2 1736 53480 1736 53480 0 reg_wdata[2]
rlabel metal2 1736 22120 1736 22120 0 reg_wdata[30]
rlabel metal2 1736 21224 1736 21224 0 reg_wdata[31]
rlabel metal2 1736 52584 1736 52584 0 reg_wdata[3]
rlabel metal2 1736 51240 1736 51240 0 reg_wdata[4]
rlabel metal2 1736 50232 1736 50232 0 reg_wdata[5]
rlabel metal3 1582 48888 1582 48888 0 reg_wdata[6]
rlabel metal2 1736 48328 1736 48328 0 reg_wdata[7]
rlabel metal3 1302 46648 1302 46648 0 reg_wdata[8]
rlabel metal2 1736 45640 1736 45640 0 reg_wdata[9]
rlabel metal2 1736 6384 1736 6384 0 reg_wr
rlabel metal2 6104 2086 6104 2086 0 reset_n
rlabel metal2 94024 56448 94024 56448 0 sar2dac[0]
rlabel metal2 82264 56280 82264 56280 0 sar2dac[1]
rlabel metal2 69048 56112 69048 56112 0 sar2dac[2]
rlabel metal2 57064 56448 57064 56448 0 sar2dac[3]
rlabel metal2 44408 56280 44408 56280 0 sar2dac[4]
rlabel metal3 31808 56280 31808 56280 0 sar2dac[5]
rlabel metal2 19152 55944 19152 55944 0 sar2dac[6]
rlabel metal2 7336 56392 7336 56392 0 sar2dac[7]
rlabel metal2 57176 28616 57176 28616 0 u_adc_reg._000_
rlabel metal3 48888 25480 48888 25480 0 u_adc_reg._001_
rlabel metal2 35672 27384 35672 27384 0 u_adc_reg._002_
rlabel metal2 48104 28112 48104 28112 0 u_adc_reg._003_
rlabel metal2 50568 29568 50568 29568 0 u_adc_reg._004_
rlabel metal2 41384 28112 41384 28112 0 u_adc_reg._005_
rlabel metal2 39424 33320 39424 33320 0 u_adc_reg._006_
rlabel metal2 55720 34608 55720 34608 0 u_adc_reg._007_
rlabel metal2 80136 43904 80136 43904 0 u_adc_reg._008_
rlabel metal2 70280 43176 70280 43176 0 u_adc_reg._009_
rlabel metal2 72744 37520 72744 37520 0 u_adc_reg._010_
rlabel metal2 62776 43176 62776 43176 0 u_adc_reg._011_
rlabel metal2 43960 43792 43960 43792 0 u_adc_reg._012_
rlabel metal2 64456 37744 64456 37744 0 u_adc_reg._013_
rlabel metal2 43960 37520 43960 37520 0 u_adc_reg._014_
rlabel metal2 63000 35224 63000 35224 0 u_adc_reg._015_
rlabel metal2 79576 47768 79576 47768 0 u_adc_reg._016_
rlabel metal2 71400 47880 71400 47880 0 u_adc_reg._017_
rlabel metal2 78120 41832 78120 41832 0 u_adc_reg._018_
rlabel metal2 65016 49840 65016 49840 0 u_adc_reg._019_
rlabel metal2 43960 47488 43960 47488 0 u_adc_reg._020_
rlabel metal2 68376 35588 68376 35588 0 u_adc_reg._021_
rlabel metal2 44296 41104 44296 41104 0 u_adc_reg._022_
rlabel metal2 53256 38472 53256 38472 0 u_adc_reg._023_
rlabel metal2 76552 50512 76552 50512 0 u_adc_reg._024_
rlabel metal2 70952 51016 70952 51016 0 u_adc_reg._025_
rlabel metal3 71960 40600 71960 40600 0 u_adc_reg._026_
rlabel metal2 60984 50288 60984 50288 0 u_adc_reg._027_
rlabel metal2 37352 47768 37352 47768 0 u_adc_reg._028_
rlabel metal2 58744 37520 58744 37520 0 u_adc_reg._029_
rlabel metal2 39032 41384 39032 41384 0 u_adc_reg._030_
rlabel metal2 50904 32088 50904 32088 0 u_adc_reg._031_
rlabel metal2 55384 47880 55384 47880 0 u_adc_reg._032_
rlabel metal2 57064 45192 57064 45192 0 u_adc_reg._033_
rlabel metal2 57400 40432 57400 40432 0 u_adc_reg._034_
rlabel metal2 31528 45976 31528 45976 0 u_adc_reg._035_
rlabel metal2 32088 43176 32088 43176 0 u_adc_reg._036_
rlabel metal2 31864 39704 31864 39704 0 u_adc_reg._037_
rlabel metal2 32088 36904 32088 36904 0 u_adc_reg._038_
rlabel metal2 61208 31472 61208 31472 0 u_adc_reg._039_
rlabel metal2 79856 45640 79856 45640 0 u_adc_reg._040_
rlabel metal2 68600 45584 68600 45584 0 u_adc_reg._041_
rlabel metal2 78568 37968 78568 37968 0 u_adc_reg._042_
rlabel metal2 61096 46088 61096 46088 0 u_adc_reg._043_
rlabel metal2 38472 44968 38472 44968 0 u_adc_reg._044_
rlabel metal2 65240 40880 65240 40880 0 u_adc_reg._045_
rlabel metal2 39480 37744 39480 37744 0 u_adc_reg._046_
rlabel metal2 55832 30072 55832 30072 0 u_adc_reg._047_
rlabel metal2 50568 47768 50568 47768 0 u_adc_reg._048_
rlabel metal2 50568 43792 50568 43792 0 u_adc_reg._049_
rlabel metal2 50680 40656 50680 40656 0 u_adc_reg._050_
rlabel metal2 26936 46200 26936 46200 0 u_adc_reg._051_
rlabel metal2 26264 43064 26264 43064 0 u_adc_reg._052_
rlabel metal2 26600 39928 26600 39928 0 u_adc_reg._053_
rlabel metal2 27160 36792 27160 36792 0 u_adc_reg._054_
rlabel metal2 90832 35672 90832 35672 0 u_adc_reg._055_
rlabel metal2 86296 49336 86296 49336 0 u_adc_reg._056_
rlabel metal2 92904 48160 92904 48160 0 u_adc_reg._057_
rlabel metal2 86856 42448 86856 42448 0 u_adc_reg._058_
rlabel metal2 86464 47208 86464 47208 0 u_adc_reg._059_
rlabel metal2 92232 46312 92232 46312 0 u_adc_reg._060_
rlabel metal2 92064 42168 92064 42168 0 u_adc_reg._061_
rlabel metal2 91840 40600 91840 40600 0 u_adc_reg._062_
rlabel metal2 82600 40040 82600 40040 0 u_adc_reg._063_
rlabel metal3 86072 39592 86072 39592 0 u_adc_reg._064_
rlabel metal2 84392 37520 84392 37520 0 u_adc_reg._065_
rlabel metal2 78400 34888 78400 34888 0 u_adc_reg._066_
rlabel metal2 84896 34888 84896 34888 0 u_adc_reg._067_
rlabel metal2 72800 34328 72800 34328 0 u_adc_reg._068_
rlabel metal2 69832 31472 69832 31472 0 u_adc_reg._069_
rlabel metal3 65352 30968 65352 30968 0 u_adc_reg._070_
rlabel metal2 68768 28616 68768 28616 0 u_adc_reg._071_
rlabel metal2 63112 27384 63112 27384 0 u_adc_reg._072_
rlabel metal3 76216 27160 76216 27160 0 u_adc_reg._073_
rlabel metal2 72632 25816 72632 25816 0 u_adc_reg._074_
rlabel metal2 62328 23912 62328 23912 0 u_adc_reg._075_
rlabel metal2 67256 26096 67256 26096 0 u_adc_reg._076_
rlabel metal3 78120 25480 78120 25480 0 u_adc_reg._077_
rlabel metal2 62328 20776 62328 20776 0 u_adc_reg._078_
rlabel metal2 78568 22512 78568 22512 0 u_adc_reg._079_
rlabel metal2 68488 22792 68488 22792 0 u_adc_reg._080_
rlabel metal2 72744 22512 72744 22512 0 u_adc_reg._081_
rlabel metal3 82768 23128 82768 23128 0 u_adc_reg._082_
rlabel metal3 85624 20552 85624 20552 0 u_adc_reg._083_
rlabel metal2 76664 19320 76664 19320 0 u_adc_reg._084_
rlabel metal3 71792 20552 71792 20552 0 u_adc_reg._085_
rlabel metal2 80584 19376 80584 19376 0 u_adc_reg._086_
rlabel metal2 43400 25200 43400 25200 0 u_adc_reg._087_
rlabel metal2 35448 26376 35448 26376 0 u_adc_reg._088_
rlabel metal2 39032 35336 39032 35336 0 u_adc_reg._089_
rlabel metal2 43736 21112 43736 21112 0 u_adc_reg._090_
rlabel metal2 38808 29848 38808 29848 0 u_adc_reg._091_
rlabel metal2 12040 26656 12040 26656 0 u_adc_reg._092_
rlabel metal2 56952 27888 56952 27888 0 u_adc_reg._093_
rlabel metal2 75096 26376 75096 26376 0 u_adc_reg._094_
rlabel metal3 91784 48216 91784 48216 0 u_adc_reg._095_
rlabel metal3 57288 29512 57288 29512 0 u_adc_reg._096_
rlabel metal2 54936 29120 54936 29120 0 u_adc_reg._097_
rlabel metal2 44072 30576 44072 30576 0 u_adc_reg._098_
rlabel metal2 44184 29624 44184 29624 0 u_adc_reg._099_
rlabel metal2 47600 28616 47600 28616 0 u_adc_reg._100_
rlabel metal2 44072 29232 44072 29232 0 u_adc_reg._101_
rlabel metal2 47208 30520 47208 30520 0 u_adc_reg._102_
rlabel metal2 46424 31808 46424 31808 0 u_adc_reg._103_
rlabel metal2 46200 33040 46200 33040 0 u_adc_reg._104_
rlabel metal2 46312 30240 46312 30240 0 u_adc_reg._105_
rlabel metal2 46200 29848 46200 29848 0 u_adc_reg._106_
rlabel metal2 43400 31864 43400 31864 0 u_adc_reg._107_
rlabel metal2 41720 28896 41720 28896 0 u_adc_reg._108_
rlabel metal2 39984 34104 39984 34104 0 u_adc_reg._109_
rlabel metal2 45080 33208 45080 33208 0 u_adc_reg._110_
rlabel metal2 46872 33152 46872 33152 0 u_adc_reg._111_
rlabel metal2 57512 35672 57512 35672 0 u_adc_reg._112_
rlabel metal2 56448 34104 56448 34104 0 u_adc_reg._113_
rlabel metal3 79072 44184 79072 44184 0 u_adc_reg._114_
rlabel metal3 71568 43512 71568 43512 0 u_adc_reg._115_
rlabel metal2 72856 38024 72856 38024 0 u_adc_reg._116_
rlabel metal2 63448 43680 63448 43680 0 u_adc_reg._117_
rlabel metal2 44632 44184 44632 44184 0 u_adc_reg._118_
rlabel metal2 65016 37240 65016 37240 0 u_adc_reg._119_
rlabel metal2 44632 37912 44632 37912 0 u_adc_reg._120_
rlabel metal2 45584 33544 45584 33544 0 u_adc_reg._121_
rlabel metal2 61600 34328 61600 34328 0 u_adc_reg._122_
rlabel metal2 62216 35000 62216 35000 0 u_adc_reg._123_
rlabel metal2 79240 47712 79240 47712 0 u_adc_reg._124_
rlabel metal3 72072 48216 72072 48216 0 u_adc_reg._125_
rlabel metal2 77560 42392 77560 42392 0 u_adc_reg._126_
rlabel metal2 64792 49504 64792 49504 0 u_adc_reg._127_
rlabel metal2 44968 47936 44968 47936 0 u_adc_reg._128_
rlabel metal2 68152 35840 68152 35840 0 u_adc_reg._129_
rlabel metal2 44744 40600 44744 40600 0 u_adc_reg._130_
rlabel metal2 43064 32536 43064 32536 0 u_adc_reg._131_
rlabel metal2 54096 37352 54096 37352 0 u_adc_reg._132_
rlabel metal2 53648 37464 53648 37464 0 u_adc_reg._133_
rlabel metal2 76384 50568 76384 50568 0 u_adc_reg._134_
rlabel metal2 72576 51464 72576 51464 0 u_adc_reg._135_
rlabel metal2 72912 40376 72912 40376 0 u_adc_reg._136_
rlabel metal2 61544 49784 61544 49784 0 u_adc_reg._137_
rlabel metal2 39144 47096 39144 47096 0 u_adc_reg._138_
rlabel metal3 59976 37912 59976 37912 0 u_adc_reg._139_
rlabel metal2 41048 41272 41048 41272 0 u_adc_reg._140_
rlabel metal3 42056 32536 42056 32536 0 u_adc_reg._141_
rlabel metal2 54488 32480 54488 32480 0 u_adc_reg._142_
rlabel metal3 52360 32312 52360 32312 0 u_adc_reg._143_
rlabel metal2 56392 48216 56392 48216 0 u_adc_reg._144_
rlabel metal2 56392 44800 56392 44800 0 u_adc_reg._145_
rlabel metal2 57008 40488 57008 40488 0 u_adc_reg._146_
rlabel metal2 32536 46984 32536 46984 0 u_adc_reg._147_
rlabel metal2 33432 43848 33432 43848 0 u_adc_reg._148_
rlabel metal2 33432 40712 33432 40712 0 u_adc_reg._149_
rlabel metal2 33488 37352 33488 37352 0 u_adc_reg._150_
rlabel metal2 44072 32872 44072 32872 0 u_adc_reg._151_
rlabel metal2 62104 33320 62104 33320 0 u_adc_reg._152_
rlabel metal2 61544 32032 61544 32032 0 u_adc_reg._153_
rlabel metal2 78680 45528 78680 45528 0 u_adc_reg._154_
rlabel metal3 69552 45080 69552 45080 0 u_adc_reg._155_
rlabel metal2 78680 37520 78680 37520 0 u_adc_reg._156_
rlabel metal2 62440 45976 62440 45976 0 u_adc_reg._157_
rlabel metal2 41048 45528 41048 45528 0 u_adc_reg._158_
rlabel metal3 66080 40376 66080 40376 0 u_adc_reg._159_
rlabel metal3 40432 37240 40432 37240 0 u_adc_reg._160_
rlabel metal2 53200 36232 53200 36232 0 u_adc_reg._161_
rlabel metal2 56168 31836 56168 31836 0 u_adc_reg._162_
rlabel metal2 51912 47096 51912 47096 0 u_adc_reg._163_
rlabel metal3 53312 44184 53312 44184 0 u_adc_reg._164_
rlabel metal2 53648 40600 53648 40600 0 u_adc_reg._165_
rlabel metal2 27272 46144 27272 46144 0 u_adc_reg._166_
rlabel metal2 27272 43008 27272 43008 0 u_adc_reg._167_
rlabel metal2 26824 39872 26824 39872 0 u_adc_reg._168_
rlabel metal2 27552 36456 27552 36456 0 u_adc_reg._169_
rlabel metal2 89320 36008 89320 36008 0 u_adc_reg._170_
rlabel metal2 47320 33656 47320 33656 0 u_adc_reg._171_
rlabel metal2 47208 35392 47208 35392 0 u_adc_reg._172_
rlabel metal2 47992 35392 47992 35392 0 u_adc_reg._173_
rlabel metal2 59864 32984 59864 32984 0 u_adc_reg._174_
rlabel metal3 48776 34776 48776 34776 0 u_adc_reg._175_
rlabel metal3 50456 33040 50456 33040 0 u_adc_reg._176_
rlabel metal2 51688 35672 51688 35672 0 u_adc_reg._177_
rlabel metal2 60760 33656 60760 33656 0 u_adc_reg._178_
rlabel metal2 63392 32424 63392 32424 0 u_adc_reg._179_
rlabel metal2 52472 34888 52472 34888 0 u_adc_reg._180_
rlabel metal2 52808 35392 52808 35392 0 u_adc_reg._181_
rlabel metal2 50624 37352 50624 37352 0 u_adc_reg._182_
rlabel metal2 51520 36456 51520 36456 0 u_adc_reg._183_
rlabel metal2 53368 36232 53368 36232 0 u_adc_reg._184_
rlabel metal2 53592 35840 53592 35840 0 u_adc_reg._185_
rlabel metal3 46592 35672 46592 35672 0 u_adc_reg._186_
rlabel metal2 54152 35224 54152 35224 0 u_adc_reg._187_
rlabel metal2 69496 21952 69496 21952 0 u_adc_reg._188_
rlabel metal2 89096 35224 89096 35224 0 u_adc_reg._189_
rlabel metal2 90216 35896 90216 35896 0 u_adc_reg._190_
rlabel metal2 77168 46648 77168 46648 0 u_adc_reg._191_
rlabel metal2 77672 46256 77672 46256 0 u_adc_reg._192_
rlabel metal2 51576 34720 51576 34720 0 u_adc_reg._193_
rlabel metal2 76776 46760 76776 46760 0 u_adc_reg._194_
rlabel metal2 50120 40936 50120 40936 0 u_adc_reg._195_
rlabel metal2 78120 46984 78120 46984 0 u_adc_reg._196_
rlabel metal2 78456 47824 78456 47824 0 u_adc_reg._197_
rlabel metal2 86128 49224 86128 49224 0 u_adc_reg._198_
rlabel metal2 74032 46648 74032 46648 0 u_adc_reg._199_
rlabel metal2 73080 46368 73080 46368 0 u_adc_reg._200_
rlabel metal2 73416 46144 73416 46144 0 u_adc_reg._201_
rlabel metal2 74984 46816 74984 46816 0 u_adc_reg._202_
rlabel metal2 91672 47880 91672 47880 0 u_adc_reg._203_
rlabel metal3 93072 47432 93072 47432 0 u_adc_reg._204_
rlabel metal2 76384 40264 76384 40264 0 u_adc_reg._205_
rlabel metal2 77616 38920 77616 38920 0 u_adc_reg._206_
rlabel metal2 59304 41160 59304 41160 0 u_adc_reg._207_
rlabel metal3 77392 40376 77392 40376 0 u_adc_reg._208_
rlabel metal2 87528 41216 87528 41216 0 u_adc_reg._209_
rlabel metal3 88200 41944 88200 41944 0 u_adc_reg._210_
rlabel metal2 66472 44968 66472 44968 0 u_adc_reg._211_
rlabel metal2 64904 46256 64904 46256 0 u_adc_reg._212_
rlabel metal3 65240 46760 65240 46760 0 u_adc_reg._213_
rlabel metal2 65240 47376 65240 47376 0 u_adc_reg._214_
rlabel metal2 86408 46592 86408 46592 0 u_adc_reg._215_
rlabel metal2 87304 46928 87304 46928 0 u_adc_reg._216_
rlabel metal2 49112 45080 49112 45080 0 u_adc_reg._217_
rlabel metal2 47320 45584 47320 45584 0 u_adc_reg._218_
rlabel metal3 43064 45528 43064 45528 0 u_adc_reg._219_
rlabel metal2 48048 45752 48048 45752 0 u_adc_reg._220_
rlabel metal2 92008 45248 92008 45248 0 u_adc_reg._221_
rlabel metal2 92904 45976 92904 45976 0 u_adc_reg._222_
rlabel metal2 67928 39256 67928 39256 0 u_adc_reg._223_
rlabel metal2 68712 39984 68712 39984 0 u_adc_reg._224_
rlabel metal2 68152 40544 68152 40544 0 u_adc_reg._225_
rlabel metal2 68936 40152 68936 40152 0 u_adc_reg._226_
rlabel metal2 91448 42112 91448 42112 0 u_adc_reg._227_
rlabel metal2 92344 42224 92344 42224 0 u_adc_reg._228_
rlabel metal2 50064 37912 50064 37912 0 u_adc_reg._229_
rlabel metal2 48328 38724 48328 38724 0 u_adc_reg._230_
rlabel metal2 38528 37464 38528 37464 0 u_adc_reg._231_
rlabel metal2 49000 39424 49000 39424 0 u_adc_reg._232_
rlabel metal2 89096 38528 89096 38528 0 u_adc_reg._233_
rlabel metal2 92008 39200 92008 39200 0 u_adc_reg._234_
rlabel metal3 36568 39648 36568 39648 0 u_adc_reg._235_
rlabel metal2 75040 21560 75040 21560 0 u_adc_reg._236_
rlabel metal3 83496 39592 83496 39592 0 u_adc_reg._237_
rlabel metal3 55636 39592 55636 39592 0 u_adc_reg._238_
rlabel metal2 85512 39592 85512 39592 0 u_adc_reg._239_
rlabel metal2 37352 37632 37352 37632 0 u_adc_reg._240_
rlabel metal2 85064 38024 85064 38024 0 u_adc_reg._241_
rlabel metal2 78008 36176 78008 36176 0 u_adc_reg._242_
rlabel metal3 79464 35672 79464 35672 0 u_adc_reg._243_
rlabel metal2 36848 35448 36848 35448 0 u_adc_reg._244_
rlabel metal2 86016 33880 86016 33880 0 u_adc_reg._245_
rlabel metal2 72632 34104 72632 34104 0 u_adc_reg._246_
rlabel metal2 68936 26096 68936 26096 0 u_adc_reg._247_
rlabel metal3 73864 34104 73864 34104 0 u_adc_reg._248_
rlabel metal3 55440 31136 55440 31136 0 u_adc_reg._249_
rlabel metal2 72352 30744 72352 30744 0 u_adc_reg._250_
rlabel metal2 64904 32032 64904 32032 0 u_adc_reg._251_
rlabel metal2 66472 30968 66472 30968 0 u_adc_reg._252_
rlabel metal2 68376 29008 68376 29008 0 u_adc_reg._253_
rlabel metal2 70504 28728 70504 28728 0 u_adc_reg._254_
rlabel metal3 67760 26376 67760 26376 0 u_adc_reg._255_
rlabel metal2 61096 28448 61096 28448 0 u_adc_reg._256_
rlabel metal2 61320 28728 61320 28728 0 u_adc_reg._257_
rlabel metal3 64680 27608 64680 27608 0 u_adc_reg._258_
rlabel metal2 76216 27048 76216 27048 0 u_adc_reg._259_
rlabel metal2 77168 27048 77168 27048 0 u_adc_reg._260_
rlabel metal2 72576 26488 72576 26488 0 u_adc_reg._261_
rlabel metal2 74200 25592 74200 25592 0 u_adc_reg._262_
rlabel metal2 62272 25480 62272 25480 0 u_adc_reg._263_
rlabel metal3 64008 25480 64008 25480 0 u_adc_reg._264_
rlabel metal2 67144 26656 67144 26656 0 u_adc_reg._265_
rlabel metal2 68600 25648 68600 25648 0 u_adc_reg._266_
rlabel metal2 76776 25648 76776 25648 0 u_adc_reg._267_
rlabel metal2 77896 25200 77896 25200 0 u_adc_reg._268_
rlabel metal2 62328 23520 62328 23520 0 u_adc_reg._269_
rlabel metal2 64288 21784 64288 21784 0 u_adc_reg._270_
rlabel metal3 77784 23184 77784 23184 0 u_adc_reg._271_
rlabel metal2 80248 22456 80248 22456 0 u_adc_reg._272_
rlabel metal2 60088 23016 60088 23016 0 u_adc_reg._273_
rlabel metal2 69048 22344 69048 22344 0 u_adc_reg._274_
rlabel metal2 73528 23520 73528 23520 0 u_adc_reg._275_
rlabel metal2 74984 22064 74984 22064 0 u_adc_reg._276_
rlabel metal2 46312 22848 46312 22848 0 u_adc_reg._277_
rlabel metal3 83664 22232 83664 22232 0 u_adc_reg._278_
rlabel metal2 84392 21112 84392 21112 0 u_adc_reg._279_
rlabel metal2 85736 20776 85736 20776 0 u_adc_reg._280_
rlabel metal2 76328 20384 76328 20384 0 u_adc_reg._281_
rlabel metal2 78064 19768 78064 19768 0 u_adc_reg._282_
rlabel metal3 64232 20776 64232 20776 0 u_adc_reg._283_
rlabel metal2 73192 20496 73192 20496 0 u_adc_reg._284_
rlabel metal3 43680 19880 43680 19880 0 u_adc_reg._285_
rlabel metal3 82376 19992 82376 19992 0 u_adc_reg._286_
rlabel metal2 45416 13384 45416 13384 0 u_adc_reg.adc_ch_no\[0\]
rlabel metal2 53704 28952 53704 28952 0 u_adc_reg.adc_ch_no\[1\]
rlabel metal2 44352 26152 44352 26152 0 u_adc_reg.adc_ch_no\[2\]
rlabel metal2 21896 42280 21896 42280 0 u_adc_reg.reg_0\[0\]
rlabel metal3 23184 37240 23184 37240 0 u_adc_reg.reg_0\[10\]
rlabel metal2 11928 36792 11928 36792 0 u_adc_reg.reg_0\[11\]
rlabel metal2 17528 36120 17528 36120 0 u_adc_reg.reg_0\[12\]
rlabel metal2 21000 35112 21000 35112 0 u_adc_reg.reg_0\[13\]
rlabel metal2 20384 33320 20384 33320 0 u_adc_reg.reg_0\[14\]
rlabel metal3 17416 31640 17416 31640 0 u_adc_reg.reg_0\[15\]
rlabel metal3 33544 30744 33544 30744 0 u_adc_reg.reg_0\[16\]
rlabel metal2 16968 29008 16968 29008 0 u_adc_reg.reg_0\[17\]
rlabel metal2 61768 28560 61768 28560 0 u_adc_reg.reg_0\[18\]
rlabel metal2 59976 27216 59976 27216 0 u_adc_reg.reg_0\[19\]
rlabel metal2 13160 46200 13160 46200 0 u_adc_reg.reg_0\[1\]
rlabel metal3 26376 28728 26376 28728 0 u_adc_reg.reg_0\[20\]
rlabel metal2 17416 27664 17416 27664 0 u_adc_reg.reg_0\[21\]
rlabel metal2 23128 26656 23128 26656 0 u_adc_reg.reg_0\[22\]
rlabel metal2 28448 25256 28448 25256 0 u_adc_reg.reg_0\[23\]
rlabel metal2 40208 24584 40208 24584 0 u_adc_reg.reg_0\[24\]
rlabel metal2 34776 24360 34776 24360 0 u_adc_reg.reg_0\[25\]
rlabel metal2 16408 24248 16408 24248 0 u_adc_reg.reg_0\[26\]
rlabel metal2 23128 23408 23128 23408 0 u_adc_reg.reg_0\[27\]
rlabel metal3 43764 21784 43764 21784 0 u_adc_reg.reg_0\[28\]
rlabel metal2 37016 21000 37016 21000 0 u_adc_reg.reg_0\[29\]
rlabel metal2 24920 47040 24920 47040 0 u_adc_reg.reg_0\[2\]
rlabel metal2 16856 21168 16856 21168 0 u_adc_reg.reg_0\[30\]
rlabel metal3 26432 20776 26432 20776 0 u_adc_reg.reg_0\[31\]
rlabel metal3 10696 44296 10696 44296 0 u_adc_reg.reg_0\[3\]
rlabel metal2 17752 47208 17752 47208 0 u_adc_reg.reg_0\[4\]
rlabel metal3 18872 44072 18872 44072 0 u_adc_reg.reg_0\[5\]
rlabel metal2 24248 44464 24248 44464 0 u_adc_reg.reg_0\[6\]
rlabel metal2 14392 42616 14392 42616 0 u_adc_reg.reg_0\[7\]
rlabel metal2 13608 40264 13608 40264 0 u_adc_reg.reg_0\[8\]
rlabel metal2 22680 40824 22680 40824 0 u_adc_reg.reg_0\[9\]
rlabel metal2 57736 34944 57736 34944 0 u_adc_reg.reg_1\[0\]
rlabel metal3 80752 43624 80752 43624 0 u_adc_reg.reg_1\[1\]
rlabel metal2 73528 43652 73528 43652 0 u_adc_reg.reg_1\[2\]
rlabel metal2 76104 37464 76104 37464 0 u_adc_reg.reg_1\[3\]
rlabel metal2 65856 42952 65856 42952 0 u_adc_reg.reg_1\[4\]
rlabel metal2 47208 43960 47208 43960 0 u_adc_reg.reg_1\[5\]
rlabel metal3 67536 38920 67536 38920 0 u_adc_reg.reg_1\[6\]
rlabel metal2 47208 37632 47208 37632 0 u_adc_reg.reg_1\[7\]
rlabel metal2 63784 32928 63784 32928 0 u_adc_reg.reg_2\[0\]
rlabel metal3 81032 48328 81032 48328 0 u_adc_reg.reg_2\[1\]
rlabel metal2 73528 48272 73528 48272 0 u_adc_reg.reg_2\[2\]
rlabel metal2 78680 41720 78680 41720 0 u_adc_reg.reg_2\[3\]
rlabel metal2 65912 49224 65912 49224 0 u_adc_reg.reg_2\[4\]
rlabel metal2 46984 47096 46984 47096 0 u_adc_reg.reg_2\[5\]
rlabel metal2 69608 36120 69608 36120 0 u_adc_reg.reg_2\[6\]
rlabel metal2 48440 40712 48440 40712 0 u_adc_reg.reg_2\[7\]
rlabel metal3 53928 37352 53928 37352 0 u_adc_reg.reg_3\[0\]
rlabel metal3 79240 50456 79240 50456 0 u_adc_reg.reg_3\[1\]
rlabel metal2 73864 49672 73864 49672 0 u_adc_reg.reg_3\[2\]
rlabel metal3 75544 41048 75544 41048 0 u_adc_reg.reg_3\[3\]
rlabel metal3 64512 49560 64512 49560 0 u_adc_reg.reg_3\[4\]
rlabel metal3 44128 47992 44128 47992 0 u_adc_reg.reg_3\[5\]
rlabel metal2 61768 37688 61768 37688 0 u_adc_reg.reg_3\[6\]
rlabel metal3 45808 41048 45808 41048 0 u_adc_reg.reg_3\[7\]
rlabel metal2 53088 32760 53088 32760 0 u_adc_reg.reg_4\[0\]
rlabel metal2 58464 47208 58464 47208 0 u_adc_reg.reg_4\[1\]
rlabel metal2 56784 44296 56784 44296 0 u_adc_reg.reg_4\[2\]
rlabel metal3 59416 41160 59416 41160 0 u_adc_reg.reg_4\[3\]
rlabel metal2 34552 46368 34552 46368 0 u_adc_reg.reg_4\[4\]
rlabel metal3 34664 42952 34664 42952 0 u_adc_reg.reg_4\[5\]
rlabel metal2 34888 40152 34888 40152 0 u_adc_reg.reg_4\[6\]
rlabel metal2 35112 36848 35112 36848 0 u_adc_reg.reg_4\[7\]
rlabel metal2 62552 32256 62552 32256 0 u_adc_reg.reg_5\[0\]
rlabel metal2 78344 45360 78344 45360 0 u_adc_reg.reg_5\[1\]
rlabel metal3 71232 45640 71232 45640 0 u_adc_reg.reg_5\[2\]
rlabel metal2 78344 37520 78344 37520 0 u_adc_reg.reg_5\[3\]
rlabel metal3 63392 45640 63392 45640 0 u_adc_reg.reg_5\[4\]
rlabel metal3 44464 45080 44464 45080 0 u_adc_reg.reg_5\[5\]
rlabel metal2 66920 39816 66920 39816 0 u_adc_reg.reg_5\[6\]
rlabel metal3 45080 38248 45080 38248 0 u_adc_reg.reg_5\[7\]
rlabel metal2 59024 28840 59024 28840 0 u_adc_reg.reg_6\[0\]
rlabel metal3 56168 46424 56168 46424 0 u_adc_reg.reg_6\[1\]
rlabel metal2 54936 44688 54936 44688 0 u_adc_reg.reg_6\[2\]
rlabel metal2 54040 40320 54040 40320 0 u_adc_reg.reg_6\[3\]
rlabel metal3 32424 46536 32424 46536 0 u_adc_reg.reg_6\[4\]
rlabel metal3 32592 43512 32592 43512 0 u_adc_reg.reg_6\[5\]
rlabel metal3 32536 40376 32536 40376 0 u_adc_reg.reg_6\[6\]
rlabel metal3 32424 37240 32424 37240 0 u_adc_reg.reg_6\[7\]
rlabel metal2 53592 26656 53592 26656 0 u_adc_reg.reg_cs_2l
rlabel metal2 48440 25984 48440 25984 0 u_adc_reg.reg_cs_l
rlabel metal3 94976 35896 94976 35896 0 u_adc_reg.reg_rdata\[0\]
rlabel metal2 96264 37464 96264 37464 0 u_adc_reg.reg_rdata\[10\]
rlabel metal2 81592 35728 81592 35728 0 u_adc_reg.reg_rdata\[11\]
rlabel metal2 85848 34552 85848 34552 0 u_adc_reg.reg_rdata\[12\]
rlabel metal2 75768 34496 75768 34496 0 u_adc_reg.reg_rdata\[13\]
rlabel metal2 72520 31192 72520 31192 0 u_adc_reg.reg_rdata\[14\]
rlabel metal2 68600 30464 68600 30464 0 u_adc_reg.reg_rdata\[15\]
rlabel metal3 71344 28616 71344 28616 0 u_adc_reg.reg_rdata\[16\]
rlabel metal2 66304 27272 66304 27272 0 u_adc_reg.reg_rdata\[17\]
rlabel metal3 81872 27608 81872 27608 0 u_adc_reg.reg_rdata\[18\]
rlabel metal2 75768 24584 75768 24584 0 u_adc_reg.reg_rdata\[19\]
rlabel metal2 90776 50288 90776 50288 0 u_adc_reg.reg_rdata\[1\]
rlabel metal2 65240 23632 65240 23632 0 u_adc_reg.reg_rdata\[20\]
rlabel metal3 69552 24920 69552 24920 0 u_adc_reg.reg_rdata\[21\]
rlabel metal2 81928 25088 81928 25088 0 u_adc_reg.reg_rdata\[22\]
rlabel metal3 64904 21000 64904 21000 0 u_adc_reg.reg_rdata\[23\]
rlabel metal2 81704 21672 81704 21672 0 u_adc_reg.reg_rdata\[24\]
rlabel metal2 69384 22568 69384 22568 0 u_adc_reg.reg_rdata\[25\]
rlabel metal2 75768 21896 75768 21896 0 u_adc_reg.reg_rdata\[26\]
rlabel metal2 86520 22288 86520 22288 0 u_adc_reg.reg_rdata\[27\]
rlabel metal2 89096 19768 89096 19768 0 u_adc_reg.reg_rdata\[28\]
rlabel metal2 79800 19768 79800 19768 0 u_adc_reg.reg_rdata\[29\]
rlabel metal2 96264 48720 96264 48720 0 u_adc_reg.reg_rdata\[2\]
rlabel metal2 74424 19768 74424 19768 0 u_adc_reg.reg_rdata\[30\]
rlabel metal2 83608 18312 83608 18312 0 u_adc_reg.reg_rdata\[31\]
rlabel metal2 96264 43512 96264 43512 0 u_adc_reg.reg_rdata\[3\]
rlabel metal2 96152 46984 96152 46984 0 u_adc_reg.reg_rdata\[4\]
rlabel metal3 94136 45640 94136 45640 0 u_adc_reg.reg_rdata\[5\]
rlabel metal2 95592 43932 95592 43932 0 u_adc_reg.reg_rdata\[6\]
rlabel metal3 93520 40376 93520 40376 0 u_adc_reg.reg_rdata\[7\]
rlabel metal2 96264 40824 96264 40824 0 u_adc_reg.reg_rdata\[8\]
rlabel metal2 96264 39872 96264 39872 0 u_adc_reg.reg_rdata\[9\]
rlabel metal2 50456 34496 50456 34496 0 u_adc_reg.sw_addr\[0\]
rlabel metal2 50456 37184 50456 37184 0 u_adc_reg.sw_addr\[1\]
rlabel metal2 51016 34664 51016 34664 0 u_adc_reg.sw_addr\[2\]
rlabel metal2 39144 34832 39144 34832 0 u_adc_reg.sw_addr\[3\]
rlabel metal2 57736 26096 57736 26096 0 u_adc_reg.sw_rd_en
rlabel metal3 17528 42616 17528 42616 0 u_adc_reg.sw_reg_wdata\[0\]
rlabel metal2 5320 38976 5320 38976 0 u_adc_reg.sw_reg_wdata\[10\]
rlabel metal3 7140 37352 7140 37352 0 u_adc_reg.sw_reg_wdata\[11\]
rlabel metal2 9128 39872 9128 39872 0 u_adc_reg.sw_reg_wdata\[12\]
rlabel metal3 7308 35672 7308 35672 0 u_adc_reg.sw_reg_wdata\[13\]
rlabel metal2 19544 33600 19544 33600 0 u_adc_reg.sw_reg_wdata\[14\]
rlabel metal2 15176 33544 15176 33544 0 u_adc_reg.sw_reg_wdata\[15\]
rlabel metal2 5320 30184 5320 30184 0 u_adc_reg.sw_reg_wdata\[16\]
rlabel metal3 12488 33320 12488 33320 0 u_adc_reg.sw_reg_wdata\[17\]
rlabel metal2 30632 31528 30632 31528 0 u_adc_reg.sw_reg_wdata\[18\]
rlabel metal2 5656 28224 5656 28224 0 u_adc_reg.sw_reg_wdata\[19\]
rlabel metal2 9688 47656 9688 47656 0 u_adc_reg.sw_reg_wdata\[1\]
rlabel metal2 25200 28504 25200 28504 0 u_adc_reg.sw_reg_wdata\[20\]
rlabel metal2 12544 27944 12544 27944 0 u_adc_reg.sw_reg_wdata\[21\]
rlabel metal2 22232 26936 22232 26936 0 u_adc_reg.sw_reg_wdata\[22\]
rlabel metal2 5880 26600 5880 26600 0 u_adc_reg.sw_reg_wdata\[23\]
rlabel metal2 10808 25480 10808 25480 0 u_adc_reg.sw_reg_wdata\[24\]
rlabel metal2 9688 24640 9688 24640 0 u_adc_reg.sw_reg_wdata\[25\]
rlabel metal2 10584 25144 10584 25144 0 u_adc_reg.sw_reg_wdata\[26\]
rlabel metal2 21448 23744 21448 23744 0 u_adc_reg.sw_reg_wdata\[27\]
rlabel metal2 38696 22568 38696 22568 0 u_adc_reg.sw_reg_wdata\[28\]
rlabel metal2 33656 21000 33656 21000 0 u_adc_reg.sw_reg_wdata\[29\]
rlabel metal2 20440 49336 20440 49336 0 u_adc_reg.sw_reg_wdata\[2\]
rlabel metal3 14504 21672 14504 21672 0 u_adc_reg.sw_reg_wdata\[30\]
rlabel metal3 22960 20664 22960 20664 0 u_adc_reg.sw_reg_wdata\[31\]
rlabel metal2 10360 45528 10360 45528 0 u_adc_reg.sw_reg_wdata\[3\]
rlabel metal2 14952 48552 14952 48552 0 u_adc_reg.sw_reg_wdata\[4\]
rlabel metal2 5992 45808 5992 45808 0 u_adc_reg.sw_reg_wdata\[5\]
rlabel metal2 6552 44688 6552 44688 0 u_adc_reg.sw_reg_wdata\[6\]
rlabel metal3 7196 43288 7196 43288 0 u_adc_reg.sw_reg_wdata\[7\]
rlabel metal2 11928 39816 11928 39816 0 u_adc_reg.sw_reg_wdata\[8\]
rlabel metal2 17640 41104 17640 41104 0 u_adc_reg.sw_reg_wdata\[9\]
rlabel metal2 54600 27776 54600 27776 0 u_adc_reg.sw_wr_en
rlabel metal2 10920 22736 10920 22736 0 u_adc_reg.sw_wr_en_0
rlabel metal2 20440 41888 20440 41888 0 u_adc_reg.u_reg_0._000_
rlabel metal2 9016 46704 9016 46704 0 u_adc_reg.u_reg_0._001_
rlabel metal2 20776 47376 20776 47376 0 u_adc_reg.u_reg_0._002_
rlabel metal3 9408 44072 9408 44072 0 u_adc_reg.u_reg_0._003_
rlabel metal2 14280 47880 14280 47880 0 u_adc_reg.u_reg_0._004_
rlabel metal2 14616 44744 14616 44744 0 u_adc_reg.u_reg_0._005_
rlabel metal2 20720 45304 20720 45304 0 u_adc_reg.u_reg_0._006_
rlabel metal3 13384 42504 13384 42504 0 u_adc_reg.u_reg_0._007_
rlabel metal2 13832 39088 13832 39088 0 u_adc_reg.u_reg_0._008_
rlabel metal2 18648 39312 18648 39312 0 u_adc_reg.u_reg_0._009_
rlabel metal2 20776 37968 20776 37968 0 u_adc_reg.u_reg_0._010_
rlabel metal2 9016 36904 9016 36904 0 u_adc_reg.u_reg_0._011_
rlabel metal2 15288 36904 15288 36904 0 u_adc_reg.u_reg_0._012_
rlabel metal2 21896 35336 21896 35336 0 u_adc_reg.u_reg_0._013_
rlabel metal2 21280 32536 21280 32536 0 u_adc_reg.u_reg_0._014_
rlabel metal2 14952 31836 14952 31836 0 u_adc_reg.u_reg_0._015_
rlabel metal2 26712 31528 26712 31528 0 u_adc_reg.u_reg_0._016_
rlabel metal2 14000 29400 14000 29400 0 u_adc_reg.u_reg_0._017_
rlabel metal2 32088 30184 32088 30184 0 u_adc_reg.u_reg_0._018_
rlabel metal2 29624 28280 29624 28280 0 u_adc_reg.u_reg_0._019_
rlabel metal2 24696 27888 24696 27888 0 u_adc_reg.u_reg_0._020_
rlabel metal2 14168 27496 14168 27496 0 u_adc_reg.u_reg_0._021_
rlabel metal2 20328 25816 20328 25816 0 u_adc_reg.u_reg_0._022_
rlabel metal2 26656 26376 26656 26376 0 u_adc_reg.u_reg_0._023_
rlabel metal2 39144 24584 39144 24584 0 u_adc_reg.u_reg_0._024_
rlabel metal2 33544 25256 33544 25256 0 u_adc_reg.u_reg_0._025_
rlabel metal3 12600 24920 12600 24920 0 u_adc_reg.u_reg_0._026_
rlabel metal2 21336 22680 21336 22680 0 u_adc_reg.u_reg_0._027_
rlabel metal2 39368 21224 39368 21224 0 u_adc_reg.u_reg_0._028_
rlabel metal2 33880 21840 33880 21840 0 u_adc_reg.u_reg_0._029_
rlabel metal2 14616 21224 14616 21224 0 u_adc_reg.u_reg_0._030_
rlabel metal2 25592 20496 25592 20496 0 u_adc_reg.u_reg_0._031_
rlabel metal3 10808 47320 10808 47320 0 u_adc_reg.u_reg_0._032_
rlabel metal2 20216 42224 20216 42224 0 u_adc_reg.u_reg_0._033_
rlabel metal2 8680 46984 8680 46984 0 u_adc_reg.u_reg_0._034_
rlabel metal2 20552 47712 20552 47712 0 u_adc_reg.u_reg_0._035_
rlabel metal2 9128 44296 9128 44296 0 u_adc_reg.u_reg_0._036_
rlabel metal3 14952 48216 14952 48216 0 u_adc_reg.u_reg_0._037_
rlabel metal3 15736 45080 15736 45080 0 u_adc_reg.u_reg_0._038_
rlabel metal3 21336 44408 21336 44408 0 u_adc_reg.u_reg_0._039_
rlabel metal2 12712 42672 12712 42672 0 u_adc_reg.u_reg_0._040_
rlabel metal2 20216 35616 20216 35616 0 u_adc_reg.u_reg_0._041_
rlabel metal3 13160 39480 13160 39480 0 u_adc_reg.u_reg_0._042_
rlabel metal2 18424 39984 18424 39984 0 u_adc_reg.u_reg_0._043_
rlabel metal2 21672 37576 21672 37576 0 u_adc_reg.u_reg_0._044_
rlabel metal3 9184 37352 9184 37352 0 u_adc_reg.u_reg_0._045_
rlabel metal2 16520 36568 16520 36568 0 u_adc_reg.u_reg_0._046_
rlabel metal2 21560 35672 21560 35672 0 u_adc_reg.u_reg_0._047_
rlabel metal2 21112 33320 21112 33320 0 u_adc_reg.u_reg_0._048_
rlabel metal3 15680 32648 15680 32648 0 u_adc_reg.u_reg_0._049_
rlabel metal2 25480 29400 25480 29400 0 u_adc_reg.u_reg_0._050_
rlabel metal2 28280 31080 28280 31080 0 u_adc_reg.u_reg_0._051_
rlabel metal3 15512 30072 15512 30072 0 u_adc_reg.u_reg_0._052_
rlabel metal2 31864 30296 31864 30296 0 u_adc_reg.u_reg_0._053_
rlabel metal2 31304 27272 31304 27272 0 u_adc_reg.u_reg_0._054_
rlabel metal2 24472 28224 24472 28224 0 u_adc_reg.u_reg_0._055_
rlabel metal2 13608 27832 13608 27832 0 u_adc_reg.u_reg_0._056_
rlabel metal2 20664 25760 20664 25760 0 u_adc_reg.u_reg_0._057_
rlabel metal2 27272 25984 27272 25984 0 u_adc_reg.u_reg_0._058_
rlabel metal2 20272 24024 20272 24024 0 u_adc_reg.u_reg_0._059_
rlabel metal2 39592 25200 39592 25200 0 u_adc_reg.u_reg_0._060_
rlabel metal2 34216 24752 34216 24752 0 u_adc_reg.u_reg_0._061_
rlabel metal2 11704 24976 11704 24976 0 u_adc_reg.u_reg_0._062_
rlabel metal2 21672 23016 21672 23016 0 u_adc_reg.u_reg_0._063_
rlabel metal2 39144 21840 39144 21840 0 u_adc_reg.u_reg_0._064_
rlabel metal2 34776 21672 34776 21672 0 u_adc_reg.u_reg_0._065_
rlabel metal3 15288 21560 15288 21560 0 u_adc_reg.u_reg_0._066_
rlabel metal3 24976 20552 24976 20552 0 u_adc_reg.u_reg_0._067_
rlabel metal2 9240 22960 9240 22960 0 u_adc_reg.u_reg_0.we\[0\]
rlabel metal3 7784 23240 7784 23240 0 u_adc_reg.u_reg_0.we\[1\]
rlabel metal3 7896 20104 7896 20104 0 u_adc_reg.u_reg_0.we\[2\]
rlabel metal2 9856 21000 9856 21000 0 u_adc_reg.u_reg_0.we\[3\]
<< properties >>
string FIXED_BBOX 0 0 100000 60000
<< end >>
