* NGSPICE file created from temp_sensor.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_3 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_1 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_4 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__invz_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__invz_4 EN I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_8 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

.subckt temp_sensor clk i_wb_addr[0] i_wb_addr[10] i_wb_addr[11] i_wb_addr[12] i_wb_addr[13]
+ i_wb_addr[14] i_wb_addr[15] i_wb_addr[16] i_wb_addr[17] i_wb_addr[18] i_wb_addr[19]
+ i_wb_addr[1] i_wb_addr[20] i_wb_addr[21] i_wb_addr[22] i_wb_addr[23] i_wb_addr[24]
+ i_wb_addr[25] i_wb_addr[26] i_wb_addr[27] i_wb_addr[28] i_wb_addr[29] i_wb_addr[2]
+ i_wb_addr[30] i_wb_addr[31] i_wb_addr[3] i_wb_addr[4] i_wb_addr[5] i_wb_addr[6]
+ i_wb_addr[7] i_wb_addr[8] i_wb_addr[9] i_wb_cyc i_wb_data[0] i_wb_data[10] i_wb_data[11]
+ i_wb_data[12] i_wb_data[13] i_wb_data[14] i_wb_data[15] i_wb_data[16] i_wb_data[17]
+ i_wb_data[18] i_wb_data[19] i_wb_data[1] i_wb_data[20] i_wb_data[21] i_wb_data[22]
+ i_wb_data[23] i_wb_data[24] i_wb_data[25] i_wb_data[26] i_wb_data[27] i_wb_data[28]
+ i_wb_data[29] i_wb_data[2] i_wb_data[30] i_wb_data[31] i_wb_data[3] i_wb_data[4]
+ i_wb_data[5] i_wb_data[6] i_wb_data[7] i_wb_data[8] i_wb_data[9] i_wb_stb i_wb_we
+ io_oeb[0] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_out[0] io_out[1]
+ io_out[2] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] o_wb_ack o_wb_data[0]
+ o_wb_data[1] o_wb_data[2] o_wb_data[3] o_wb_data[4] o_wb_data[5] o_wb_data[6] o_wb_data[7]
+ o_wb_stall reset vdd vss io_oeb[2] io_oeb[1]
XTAP_TAPCELL_ROW_136_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2106_ _0124_ clknet_leaf_0_clk cal_lut\[143\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2037_ _0055_ clknet_leaf_13_clk cal_lut\[120\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1454__A1 _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1206__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1221__A4 _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_83_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1700__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1445__A1 _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._061_ dec1.i_bin\[6\] dec1._002_ dec1._012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1748__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1428__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1920__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1270_ _0834_ _0835_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_133_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1684__A1 _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1436__A1 _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0985_ ctr\[2\] ctr\[3\] _0565_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1739__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1606_ temp1.dac.i_enable _0333_ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1911__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1537_ _0239_ _0282_ _0297_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_38_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1468_ cal_lut\[52\] _0231_ _0977_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1399_ net28 _0955_ _0956_ _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_49_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_80_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1902__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1666__A1 _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1418__A1 _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2052__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1197__A3 _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1322_ _0590_ _0842_ _0840_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1253_ cal_lut\[144\] _0650_ _0628_ cal_lut\[126\] _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1106__B1 _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1184_ _0744_ _0746_ _0749_ _0752_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_148_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1409__A1 _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1896__A1 _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input36_I i_wb_data[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1648__A1 _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2075__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1820__A1 _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_137_Right_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1639__A1 _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1441__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1940_ _0348_ _0536_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_138_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1871_ cal_lut\[2\] _0497_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1878__A1 _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1305_ _0869_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1236_ cal_lut\[84\] _0679_ _0618_ cal_lut\[12\] _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1167_ _0734_ _0735_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2098__CLK clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1098_ _0598_ cal_lut\[32\] _0612_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_19_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1030__A2 _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1097__A2 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2070_ _0088_ clknet_leaf_0_clk cal_lut\[171\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1088__A2 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1021_ _0587_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_72_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1923_ cal_lut\[27\] _0506_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1260__A2 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1854_ _0278_ _0451_ _0485_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1785_ _0745_ _0386_ _0448_ _0430_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_97_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1079__A2 _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1219_ _0598_ cal_lut\[41\] _0766_ _0787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2199_ _0217_ clknet_leaf_7_clk en_dbg\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp_sensor_69 io_oeb[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__1251__A2 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2113__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1703__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1490__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1242__A2 _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1570_ _0272_ _0283_ _0314_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2122_ _0140_ clknet_leaf_5_clk cal_lut\[159\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_108_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
Xtemp1.dac.parallel_cells\[2\].vdac_batch._4_ temp1.dac.i_data\[2\] temp1.dac.i_data\[5\]
+ temp1.dac.parallel_cells\[2\].vdac_batch._1_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_116_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2053_ _0071_ clknet_leaf_6_clk ctr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1004_ ctr\[0\] _0564_ clknet_leaf_6_clk _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_29_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1481__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2136__CLK clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1906_ _0249_ _0496_ _0517_ _0508_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1233__A2 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1837_ cal_lut\[88\] _0461_ _0976_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1768_ _0437_ _0386_ _0438_ _0430_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1699_ net56 _0386_ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_139_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1804__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1472__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1224__A2 cal_lut\[155\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2009__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1160__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2159__CLK clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1463__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.vdac_single._4_ net79 net80 temp1.dac.vdac_single._1_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_143_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1215__A2 _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1622_ _0940_ _0345_ _0347_ _0348_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_111_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1553_ cal_lut\[117\] _0292_ _0298_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1484_ _0263_ _0962_ _0264_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_136_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2105_ _0123_ clknet_leaf_1_clk cal_lut\[142\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2036_ _0054_ clknet_leaf_12_clk cal_lut\[119\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1454__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.vdac_single.einvp_batch\[0\].pupd temp1.dac.vdac_single.en_pupd temp1.dac.vdac_single.npu_pd
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XTAP_TAPCELL_ROW_60_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input66_I i_wb_stb vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1534__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1445__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._060_ dec1.i_bin\[3\] dec1._008_ dec1._010_ dec1._011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_110_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_11_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Left_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_39_Left_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1381__A1 _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1444__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1133__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1684__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1436__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0984_ _0563_ _0564_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_13_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_120_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1605_ _0332_ _0330_ dec1.i_tens _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1536_ cal_lut\[109\] _0292_ _0266_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1467_ net44 _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1398_ net30 net29 _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1675__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2019_ _0037_ clknet_leaf_18_clk cal_lut\[102\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1060__B1 _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1363__A1 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1666__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1418__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1991__CLK clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1321_ _0856_ _0882_ _0883_ _0884_ _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1252_ cal_lut\[174\] _0655_ _0626_ cal_lut\[168\] _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1657__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_56_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1183_ _0750_ _0645_ _0751_ _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1409__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_65_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_10_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1345__A1 ctr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1519_ cal_lut\[101\] _0283_ _0266_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1896__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input29_I i_wb_addr[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_74_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1648__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_83_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1820__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1584__A1 ctr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1706__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_92_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1639__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1811__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1870_ _0940_ _0496_ _0498_ _0430_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_9_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1878__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1304_ _0833_ _0839_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1235_ _0802_ dec1.i_bin\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1166_ _0593_ cal_lut\[130\] _0612_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1097_ cal_lut\[68\] _0608_ _0610_ cal_lut\[74\] _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__1802__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1079__B _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_1_0__f_net81 clknet_0_net81 clknet_1_0__leaf_net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1999_ _0017_ clknet_leaf_16_clk cal_lut\[50\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1566__A1 _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1807__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1869__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2042__CLK clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2192__CLK clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1008__I _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1020_ _0588_ _0591_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_72_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1922_ _0265_ _0497_ _0525_ _0508_ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1853_ cal_lut\[96\] _0449_ _0976_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1548__A1 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1784_ net58 _0384_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2065__CLK clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1218_ _0646_ _0644_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2198_ _0216_ clknet_leaf_7_clk en_dbg\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1149_ _0594_ _0590_ cal_lut\[27\] _0646_ _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_62_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1236__B1 _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_20_Left_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1447__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2088__CLK clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2121_ _0139_ clknet_leaf_5_clk cal_lut\[158\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2052_ _0070_ clknet_leaf_5_clk ctr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xtemp1.dac.parallel_cells\[2\].vdac_batch._3_ temp1.dac.i_data\[2\] temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1003_ ctr\[7\] _0564_ _0577_ temp1.dac.i_data\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XTAP_TAPCELL_ROW_116_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1905_ cal_lut\[18\] _0506_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1836_ _0259_ _0451_ _0476_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1767_ net50 _0404_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1698_ cal_lut\[131\] _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_148_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input11_I i_wb_addr[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XTAP_TAPCELL_ROW_63_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1224__A3 _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1932__A1 _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1160__A2 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.vdac_single._3_ net78 temp1.dac.vdac_single.npu_pd vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_14_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1021__I _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1621_ _0963_ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1552_ _0253_ _0282_ _0305_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1483_ cal_lut\[57\] _0231_ _0977_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1691__I _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1624__C _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I i_wb_addr[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2104_ _0122_ clknet_leaf_1_clk cal_lut\[141\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2103__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2035_ _0053_ clknet_leaf_1_clk cal_lut\[118\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1206__A3 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1819_ cal_lut\[79\] _0461_ _0453_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1914__A1 _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1815__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input59_I i_wb_data[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1709__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.vdac_single.einvp_batch\[0\].vref temp1.dac.vdac_single.en_vref temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XANTENNA__2126__CLK clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1133__A2 cal_lut\[129\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_103_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0983_ ctr\[1\] _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_14_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1604_ ctr\[12\] _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_112_Left_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1535_ _0237_ _0282_ _0296_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1372__A2 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1466_ _0251_ _0961_ _0252_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1397_ net27 _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1124__A2 _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_121_Left_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2018_ _0036_ clknet_leaf_18_clk cal_lut\[101\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_72_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1545__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2149__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1051__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1320_ _0833_ _0841_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_1251_ cal_lut\[180\] _0658_ _0630_ cal_lut\[186\] _0818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1106__A2 _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1902__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1182_ _0594_ _0590_ cal_lut\[28\] _0646_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_91_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1042__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1518_ _0971_ _0282_ _0287_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1449_ net38 _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_65_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1033__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.vdac_single.einvp_batch\[0\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1336__A2 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1722__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1024__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1575__A2 _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1185__B _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1303_ _0583_ _0842_ _0840_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1632__C _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1234_ _0800_ _0801_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1165_ _0598_ cal_lut\[34\] _0612_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_126_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1096_ cal_lut\[56\] _0602_ _0605_ cal_lut\[62\] _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1998_ _0016_ clknet_leaf_16_clk cal_lut\[49\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1566__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input41_I i_wb_data[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1823__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1557__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1245__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1921_ cal_lut\[26\] _0506_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1796__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1852_ _0276_ _0451_ _0484_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1548__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1783_ _0713_ _0386_ _0447_ _0430_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2197_ _0215_ clknet_leaf_6_clk o_wb_data[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1217_ _0782_ _0645_ _0783_ _0784_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__1484__A1 _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1148_ cal_lut\[111\] _0718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1079_ cal_lut\[139\] _0650_ _0592_ _0651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_62_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1539__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1553__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1172__B1 _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1711__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1475__A1 _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1227__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1778__A2 _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1950__A2 _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1163__B1 _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1702__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2120_ _0138_ clknet_leaf_4_clk cal_lut\[157\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2051_ _0069_ clknet_leaf_5_clk ctr\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1002_ ctr\[6\] _0564_ _0577_ temp1.dac.i_data\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_16_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1910__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1466__A1 _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_116_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1218__A1 _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1904_ _0247_ _0496_ _0516_ _0508_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_89_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1835_ cal_lut\[87\] _0461_ _0976_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2032__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1766_ cal_lut\[153\] _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1941__A2 _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1697_ _0389_ _0385_ _0390_ _0388_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_148_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1154__B1 _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2182__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1457__A1 _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1209__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1932__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1448__A1 _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_14_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1620_ cal_lut\[161\] _0346_ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1551_ cal_lut\[116\] _0292_ _0298_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1923__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1482_ net50 _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__1136__B1 _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2103_ _0121_ clknet_leaf_1_clk cal_lut\[140\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_37_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2034_ _0052_ clknet_leaf_1_clk cal_lut\[117\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1439__A1 _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1818_ _0241_ _0450_ _0467_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1749_ _0424_ _0385_ _0425_ _0388_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_68_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1914__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1678__A1 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1831__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2078__CLK clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1850__A1 _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1725__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1905__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1133__A3 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._4__A2 temp1.dac.i_data\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0982_ ctr\[0\] _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_104_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_132_Right_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1603_ _0965_ _0331_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1534_ cal_lut\[108\] _0292_ _0266_ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1465_ cal_lut\[51\] _0231_ _0977_ _0252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1396_ net67 net33 net66 _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2017_ _0035_ clknet_leaf_18_clk cal_lut\[100\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1832__A1 _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1060__A2 _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1561__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1787__I _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1051__A2 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1250_ cal_lut\[42\] _0816_ _0656_ cal_lut\[18\] _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1471__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1181_ cal_lut\[112\] _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].pupd temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_115_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1814__A1 _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_24_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1517_ cal_lut\[100\] _0283_ _0266_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1448_ _0239_ _0961_ _0240_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1379_ temp1.dac.i_enable _0870_ _0937_ _0938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1805__A1 _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2116__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1291__B _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_140_Left_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_138_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1024__A2 _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1302_ _0856_ _0865_ _0866_ _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1233_ dbg3\[5\] _0585_ _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1164_ cal_lut\[70\] _0608_ _0610_ cal_lut\[76\] _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1095_ cal_lut\[152\] _0596_ _0600_ cal_lut\[134\] _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_35_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2139__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1997_ _0015_ clknet_leaf_2_clk cal_lut\[48\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input34_I i_wb_data[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1493__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1245__A2 cal_lut\[156\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1920_ _0263_ _0497_ _0524_ _0508_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1851_ cal_lut\[95\] _0449_ _0976_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1908__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1782_ net57 _0384_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1953__B1 _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1643__C _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2196_ _0214_ clknet_leaf_5_clk o_wb_data[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_119_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1216_ cal_lut\[71\] _0608_ _0621_ cal_lut\[107\] _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_46_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1147_ _0593_ _0715_ _0599_ _0640_ _0716_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__1484__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1078_ _0597_ _0589_ _0603_ _0607_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__1885__I _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0995__A1 dec1.i_ones vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1475__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._7__I temp1.dac.i_enable vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1227__A2 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0986__A1 ctr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1728__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac._5_ temp1.dac._1_ temp1.dac.i_data\[5\] temp1.dac._0_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_107_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2050_ _0068_ clknet_leaf_5_clk ctr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1001_ _0562_ _0564_ _0577_ temp1.dac.i_data\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_88_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1466__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1903_ cal_lut\[17\] _0506_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xtemp1.dac.parallel_cells\[0\].vdac_batch._8_ temp1.dac.parallel_cells\[0\].vdac_batch._0_
+ temp1.dac.parallel_cells\[0\].vdac_batch._1_ temp1.dac.parallel_cells\[0\].vdac_batch.en_vref
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1834_ _0257_ _0451_ _0475_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1765_ _0435_ _0386_ _0436_ _0430_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1696_ net45 _0386_ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_148_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1457__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2179_ _0197_ clknet_leaf_11_clk cal_lut\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_146_Right_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1829__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1696__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1448__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1994__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_9_clk_I clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1620__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1550_ _0251_ _0282_ _0304_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1474__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1481_ _0261_ _0962_ _0262_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._5__A1 temp1.dac.i_enable vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2102_ _0120_ clknet_leaf_0_clk cal_lut\[139\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2033_ _0051_ clknet_leaf_16_clk cal_lut\[116\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1439__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1817_ cal_lut\[78\] _0461_ _0453_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1748_ net43 _0404_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1679_ cal_lut\[189\] _0344_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1127__A1 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1678__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1403__I _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1559__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1850__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1669__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1313__I _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2022__CLK clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1841__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_17_Left_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2172__CLK clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0981_ ctr\[5\] _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_13_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1602_ ctr\[12\] _0330_ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_22_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1916__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1533_ _0235_ _0282_ _0295_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1464_ net43 _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XPHY_EDGE_ROW_26_Left_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1395_ _0949_ _0951_ _0952_ _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_38_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1124__A4 _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2016_ _0034_ clknet_leaf_18_clk cal_lut\[99\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_35_Left_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1832__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input64_I i_wb_data[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1899__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_44_Left_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1520__A1 _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2045__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2195__CLK clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1823__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1587__A1 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1051__A3 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1339__A1 clknet_leaf_8_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1180_ _0593_ _0747_ _0599_ _0640_ _0748_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__1511__A1 cal_lut\[97\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1814__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1578__A1 _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_12_clk clknet_1_0__leaf_clk clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1042__A3 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2068__CLK clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1516_ _0969_ _0282_ _0286_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1447_ cal_lut\[45\] _0231_ _0977_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1378_ _0842_ _0935_ _0936_ _0870_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1805__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_92_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1837__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_61_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xtemp1.dac.vdac_single._3__78 net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_36_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1301_ _0564_ _0856_ _0842_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_19_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_1_clk clknet_1_0__leaf_clk clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1232_ _0762_ _0592_ _0781_ _0799_ _0585_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1163_ cal_lut\[58\] _0602_ _0605_ cal_lut\[64\] _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_126_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1094_ cal_lut\[2\] _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1501__I net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1799__A1 _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1996_ _0014_ clknet_leaf_2_clk cal_lut\[47\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1971__A1 ctr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input27_I i_wb_addr[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1239__B1 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1567__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1962__A1 _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1190__A2 _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1245__A3 _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1850_ _0274_ _0451_ _0483_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1477__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1781_ _0681_ _0386_ _0446_ _0430_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_112_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1924__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_127_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2195_ _0213_ clknet_leaf_6_clk o_wb_data[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2106__CLK clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1215_ cal_lut\[17\] _0656_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1146_ cal_lut\[87\] _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_9_Left_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1077_ _0638_ _0642_ _0648_ _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_62_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1979_ ctr\[7\] clknet_1_1__leaf__0553_ _0559_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_30_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1172__A2 _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1406__I _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1227__A3 _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0980__I ctr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2129__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac._4_ temp1.dac.i_enable temp1.dac._1_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1000_ ctr\[4\] _0564_ _0577_ temp1.dac.i_data\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_29_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1902_ _0245_ _0496_ _0515_ _0508_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_44_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[0\].vdac_batch._7_ temp1.dac.i_enable temp1.dac.parallel_cells\[0\].vdac_batch._0_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1833_ cal_lut\[86\] _0461_ _0976_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1764_ net49 _0404_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1926__A1 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1695_ cal_lut\[130\] _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1654__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1154__A2 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2178_ _0196_ clknet_leaf_1_clk cal_lut\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1129_ cal_lut\[153\] _0596_ _0600_ cal_lut\[135\] _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_79_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1209__A3 _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1845__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_128_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1081__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1908__A1 _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1480_ cal_lut\[56\] _0231_ _0977_ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_69_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1136__A2 _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2101_ _0119_ clknet_leaf_0_clk cal_lut\[138\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1490__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2032_ _0050_ clknet_leaf_17_clk cal_lut\[115\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_99_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1072__A1 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1816_ _0239_ _0450_ _0466_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_32_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1747_ cal_lut\[147\] _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1678_ _0270_ _0346_ _0377_ _0362_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_68_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1127__A2 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_84_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1063__A1 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1575__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0980_ ctr\[7\] _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1601_ ctr\[11\] _0571_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1532_ cal_lut\[107\] _0292_ _0266_ _0295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1463_ _0249_ _0961_ _0250_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1932__C _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1394_ net18 net17 net20 net19 _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA_input1_I i_wb_addr[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1504__I net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2015_ _0033_ clknet_leaf_18_clk cal_lut\[98\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1045__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input57_I i_wb_data[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1984__CLK clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_8_clk_I clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1520__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1036__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1752__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1511__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1027__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._099_ dec1._009_ dec1._034_ dec1._047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1943__B _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1515_ cal_lut\[99\] _0283_ _0266_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1662__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1446_ net37 _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_1377_ ctr\[1\] _0842_ _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1502__A2 _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1569__A2 _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2012__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1853__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2162__CLK clknet_leaf_8_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1257__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1009__A1 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1300_ ctr\[9\] _0864_ _0843_ _0865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1231_ _0785_ _0790_ _0794_ _0798_ _0799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_126_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1162_ cal_lut\[154\] _0596_ _0600_ cal_lut\[136\] _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1093_ _0584_ _0585_ _0664_ dec1.i_bin\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_143_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1799__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1995_ _0013_ clknet_leaf_16_clk cal_lut\[46\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2035__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2185__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1429_ _0226_ _0961_ _0227_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_temp1.dcdc_EN temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1962__A2 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1583__B _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1714__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1478__A1 _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1650__A1 _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1780_ net55 _0384_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_115_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1953__A2 _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_1__f_temp1.i_precharge_n clknet_0_temp1.i_precharge_n clknet_1_1__leaf_temp1.i_precharge_n
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1493__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1705__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2194_ _0212_ clknet_leaf_5_clk o_wb_data[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1469__A1 _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1214_ cal_lut\[113\] _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1145_ cal_lut\[39\] _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1076_ _0643_ _0645_ _0647_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1641__A1 _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1978_ dbg3\[5\] clknet_1_1__leaf__0553_ _0976_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1944__A2 _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2200__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1880__A1 _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_119_Left_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1578__B _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1632__A1 _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XPHY_EDGE_ROW_128_Left_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_137_Left_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_88_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_29_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1901_ cal_lut\[16\] _0506_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1832_ _0255_ _0451_ _0474_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xtemp1.dac.parallel_cells\[0\].vdac_batch._6_ temp1.dac.parallel_cells\[0\].vdac_batch._2_
+ temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_146_Left_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1763_ cal_lut\[152\] _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_106_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1694_ _0382_ _0385_ _0387_ _0388_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1926__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1139__B1 _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1951__B _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1670__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2177_ _0195_ clknet_leaf_1_clk cal_lut\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_95_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1862__A1 _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1128_ cal_lut\[3\] _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1059_ _0594_ _0590_ _0588_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_87_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1090__A2 _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1917__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_145_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1081__A2 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1908__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2100_ _0118_ clknet_leaf_0_clk cal_lut\[137\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2031_ _0049_ clknet_leaf_1_clk cal_lut\[114\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1844__A1 _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1072__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1946__B _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1815_ cal_lut\[77\] _0461_ _0453_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1746_ _0422_ _0385_ _0423_ _0388_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1677_ cal_lut\[188\] _0356_ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_7_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2119__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1063__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1826__A1 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1054__A2 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1600_ _0965_ _0329_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1531_ _0233_ _0282_ _0294_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1462_ cal_lut\[50\] _0231_ _0977_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1393_ net25 net24 _0950_ _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_2_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2014_ _0032_ clknet_leaf_18_clk cal_lut\[97\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1729_ cal_lut\[141\] _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1808__A1 _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2091__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1036__A2 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1027__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1496__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._098_ dec1._001_ dec1._045_ dec1._025_ dec1._046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_40_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1514_ _0967_ _0282_ _0285_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1445_ _0237_ _0961_ _0238_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1376_ ctr\[7\] _0856_ _0934_ _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_dec1._078__A1 dec1.i_ones vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_100_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1193__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1230_ _0796_ _0797_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1161_ cal_lut\[4\] _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_126_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1496__A2 _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1092_ _0585_ _0663_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_142_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1994_ _0012_ clknet_leaf_2_clk cal_lut\[45\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_7_clk_I clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1420__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1428_ cal_lut\[39\] _0962_ _0977_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1487__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1359_ _0917_ _0918_ _0919_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0998__A1 ctr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1411__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1190__A4 _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1478__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_141_Right_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1997__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1650__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1166__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1213_ _0768_ _0771_ _0776_ _0780_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_46_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2193_ _0211_ clknet_leaf_5_clk o_wb_data[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1469__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1144_ _0598_ _0713_ _0604_ _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1075_ _0594_ _0590_ cal_lut\[25\] _0646_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__1949__B _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2002__CLK clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1641__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1668__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2152__CLK clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1977_ ctr\[6\] clknet_1_0__leaf__0553_ _0558_ _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input32_I i_wb_addr[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_125_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1880__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1632__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1699__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2025__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1871__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2175__CLK clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1623__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1900_ _0243_ _0496_ _0514_ _0508_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1831_ cal_lut\[85\] _0461_ _0453_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xtemp1.dac.parallel_cells\[0\].vdac_batch._5_ temp1.dac.i_enable temp1.dac.parallel_cells\[0\].vdac_batch._1_
+ temp1.dac.parallel_cells\[0\].vdac_batch._2_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1762_ _0433_ _0386_ _0434_ _0430_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1693_ _0963_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_122_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2176_ _0194_ clknet_leaf_1_clk cal_lut\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_107_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1127_ _0603_ _0585_ _0697_ dec1.i_bin\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1058_ _0597_ _0584_ _0580_ _0609_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_130_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref temp1.dac.parallel_cells\[1\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1378__A1 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_113_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2048__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1550__A1 _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2198__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1853__A2 _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1081__A3 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._58_ seg1._22_ seg1._24_ seg1._25_ seg1.o_segments\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_104_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1771__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2030_ _0048_ clknet_leaf_2_clk cal_lut\[113\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1844__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1499__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1057__B1 _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1814_ _0237_ _0450_ _0465_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1745_ net42 _0404_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1676_ _0268_ _0346_ _0376_ _0362_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_68_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2159_ _0177_ clknet_leaf_3_clk cal_lut\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1835__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1826__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1039__B1 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1054__A3 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1211__B1 _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1530_ cal_lut\[106\] _0292_ _0266_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1461_ net42 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1392_ net22 net21 _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1514__A1 _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1817__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2013_ _0031_ clknet_leaf_12_clk cal_lut\[64\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_clk clknet_1_0__leaf_clk clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1676__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1728_ _0410_ _0385_ _0411_ _0388_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1202__B1 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1659_ cal_lut\[179\] _0356_ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Left_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1808__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_22_Left_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1036__A3 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_31_Left_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1621__I _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1027__A3 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xdec1._097_ dec1._027_ dec1._045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xtemp1.inv2_2 clknet_1_0__leaf_net81 net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1513_ cal_lut\[98\] _0283_ _0266_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2109__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1444_ cal_lut\[44\] _0231_ _0977_ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_4_clk clknet_1_1__leaf_clk clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1375_ _0833_ _0838_ _0849_ dec1.i_tens _0933_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_65_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1974__A1 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input62_I i_wb_data[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_138_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1193__A2 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1160_ _0594_ _0585_ _0729_ dec1.i_bin\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1091_ _0586_ _0592_ _0616_ _0662_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__1248__A3 _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1993_ _0011_ clknet_leaf_2_clk cal_lut\[44\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1956__A1 _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1427_ net62 _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__1970__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2081__CLK clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1358_ dec1.i_ones _0835_ _0855_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1289_ _0833_ _0834_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_135_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_128_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1938__A1 _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1774__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1166__A2 cal_lut\[130\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1212_ _0777_ _0778_ _0779_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2192_ _0210_ clknet_leaf_6_clk o_wb_data[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1143_ cal_lut\[159\] _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1074_ _0587_ _0583_ _0580_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1976_ _0593_ clknet_1_0__leaf__0553_ _0976_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1684__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1157__A2 _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input25_I i_wb_addr[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XTAP_TAPCELL_ROW_125_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1093__A1 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_148_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_6_clk_I clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1084__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1830_ _0253_ _0450_ _0473_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xtemp1.dac.parallel_cells\[0\].vdac_batch._4_ temp1.dac.i_data\[0\] temp1.dac.i_data\[5\]
+ temp1.dac.parallel_cells\[0\].vdac_batch._1_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1761_ net48 _0404_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1692_ net34 _0386_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1139__A2 _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2175_ _0193_ clknet_leaf_3_clk cal_lut\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_107_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1126_ _0585_ _0696_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1057_ cal_lut\[163\] _0626_ _0628_ cal_lut\[121\] _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_87_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1075__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1090__A4 _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1959_ _0835_ _0493_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_8_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1987__CLK clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1550__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1066__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xseg1._57_ seg1._11_ seg1._04_ seg1._06_ seg1._25_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_27_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1541__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2142__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_59_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_104_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1057__A1 cal_lut\[163\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_0_clk net84 clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_84_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1813_ cal_lut\[76\] _0461_ _0453_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1744_ cal_lut\[146\] _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_68_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1675_ cal_lut\[187\] _0356_ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1780__A2 _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_5_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1532__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_77_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2158_ _0176_ clknet_leaf_8_clk cal_lut\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1296__A1 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2089_ _0107_ clknet_leaf_13_clk cal_lut\[190\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1109_ cal_lut\[80\] _0679_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_51_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_86_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2015__CLK clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1771__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1872__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2165__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1523__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_95_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_74_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_0_net81 net81 clknet_0_net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_13_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1619__I _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_136_Right_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1762__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1460_ _0247_ _0961_ _0248_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1391_ _0947_ _0948_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1514__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2012_ _0030_ clknet_leaf_12_clk cal_lut\[63\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_132_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2038__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1202__A1 cal_lut\[101\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1727_ net36 _0404_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1202__B2 cal_lut\[149\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2188__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1658_ _0249_ _0345_ _0367_ _0362_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1505__A2 _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1589_ ctr\[6\] _0323_ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_48_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1680__A1 _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1027__A4 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1777__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1432__A1 _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._096_ dec1._025_ dec1._028_ dec1._044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xtemp1.inv2_3 clknet_1_1__leaf_net81 net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1512_ _0940_ _0282_ _0284_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_10_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1443_ net36 _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_1374_ cal_ena _0849_ _0933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1120__B1 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1968__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1187__B1 _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input55_I i_wb_data[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2203__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1662__A1 _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1965__A2 _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1090_ _0619_ _0633_ _0649_ _0661_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1102__B1 _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1992_ _0010_ clknet_leaf_2_clk cal_lut\[43\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xdec1._079_ dec1.i_bin\[0\] dec1._030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1708__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1169__B1 _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1426_ _0975_ _0961_ _0978_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1357_ _0561_ _0846_ _0844_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_50_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1892__A1 _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1288_ _0844_ _0851_ _0852_ _0853_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1644__A1 cal_lut\[172\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1947__A2 _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1717__I _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1880__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_56_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1938__A2 _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1166__A3 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1211_ cal_lut\[53\] _0631_ _0628_ cal_lut\[125\] _0779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2191_ _0209_ clknet_leaf_6_clk o_wb_data[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1142_ cal_lut\[81\] _0679_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1874__A1 _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1073_ _0587_ _0583_ _0581_ _0644_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__1626__A1 _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1975_ _0562_ clknet_1_1__leaf__0553_ _0557_ _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1929__A2 _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1409_ _0940_ _0961_ _0966_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1865__A1 _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input18_I i_wb_addr[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1093__A2 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1084__A2 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_106_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
Xtemp1.dac.parallel_cells\[0\].vdac_batch._3_ temp1.dac.i_data\[0\] temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1760_ cal_lut\[151\] _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1785__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2071__CLK clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1691_ _0384_ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_122_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_115_Left_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2174_ _0192_ clknet_leaf_3_clk cal_lut\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._7__I temp1.dac.i_enable vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1125_ _0665_ _0592_ _0672_ _0695_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_107_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_124_Left_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1056_ _0587_ _0594_ _0590_ _0627_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA__1075__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1976__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1958_ _0348_ _0547_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_31_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1889_ cal_lut\[10\] _0506_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_133_Left_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1838__A1 _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_142_Left_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._56_ dec1.o_dec\[1\] seg1._03_ seg1._00_ seg1._24_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_118_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1057__A2 _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1796__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1812_ _0235_ _0450_ _0464_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1743_ _0420_ _0385_ _0421_ _0388_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1674_ _0265_ _0346_ _0375_ _0362_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_68_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2157_ _0175_ clknet_leaf_7_clk cal_ena vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_108_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1296__A2 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2088_ _0106_ clknet_leaf_13_clk cal_lut\[189\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1108_ _0587_ _0583_ _0581_ _0609_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_1039_ cal_lut\[67\] _0608_ _0610_ cal_lut\[73\] _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_51_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_5_clk_I clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1220__A2 _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1039__A2 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1211__A2 _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._39_ dec1.o_dec\[1\] dec1.o_dec\[0\] seg1._12_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1390_ net9 net8 net11 net10 _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_54_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2011_ _0029_ clknet_leaf_12_clk cal_lut\[62\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1450__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1202__A2 _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1726_ cal_lut\[140\] _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1657_ cal_lut\[178\] _0356_ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_95_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1588_ _0562_ _0567_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1441__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2132__CLK clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1680__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1432__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._095_ dec1._000_ dec1._008_ dec1._035_ dec1._043_ dec1._029_ dec1.o_dec\[2\]
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_4
X_1511_ cal_lut\[97\] _0283_ _0266_ _0284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1442_ _0235_ _0961_ _0236_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1373_ temp1.dac.i_enable _0872_ _0932_ io_out[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1499__A2 _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2005__CLK clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1671__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2155__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1187__A1 cal_lut\[172\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1709_ _0397_ _0385_ _0398_ _0388_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_input48_I i_wb_data[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1111__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1662__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1878__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1414__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1965__A3 _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2028__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1350__A1 temp1.dac.i_data\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2178__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1653__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1991_ _0009_ clknet_leaf_3_clk cal_lut\[42\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._078_ dec1.i_ones dec1._000_ dec1._029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_50_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1425_ cal_lut\[38\] _0962_ _0977_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1356_ _0800_ _0801_ _0849_ _0916_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1892__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1287_ _0833_ _0834_ _0838_ _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_92_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1644__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._4__A2 temp1.dac.i_data\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1580__A1 _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1883__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1635__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1096__B1 _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1210_ _0593_ cal_lut\[131\] _0612_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_46_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2190_ _0208_ clknet_leaf_5_clk o_wb_data[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1141_ _0707_ _0708_ _0709_ _0710_ _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1874__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1072_ _0589_ _0590_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__1626__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1974_ _0589_ clknet_1_1__leaf__0553_ _0976_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1562__A1 _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1157__A4 _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1408_ cal_lut\[33\] _0962_ _0965_ _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1314__A1 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1339_ clknet_leaf_8_clk _0901_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1865__A2 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1502__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1250__B1 _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1084__A3 _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1241__B1 _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1690_ _0384_ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_106_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1544__A1 _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2173_ _0191_ clknet_leaf_1_clk cal_lut\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1847__A2 _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1124_ _0673_ _0678_ _0689_ _0694_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1055_ _0583_ _0580_ _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_145_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_113_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1957_ o_wb_data[7] _0533_ _0535_ io_out[7] _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1232__B1 _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1888_ _0230_ _0496_ _0507_ _0508_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1535__A1 _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input30_I i_wb_addr[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1838__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._55_ seg1._00_ seg1._23_ seg1._10_ seg1.o_segments\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1526__A1 _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1829__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1811_ cal_lut\[75\] _0461_ _0453_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1742_ net41 _0404_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1673_ cal_lut\[186\] _0356_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1517__A1 cal_lut\[100\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2156_ _0174_ clknet_leaf_5_clk o_wb_ack vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2087_ _0105_ clknet_leaf_13_clk cal_lut\[188\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_18_clk clknet_1_0__leaf_clk clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1107_ _0674_ _0675_ _0676_ _0677_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1038_ _0588_ _0609_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_75_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2061__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_1__f__0553_ clknet_0__0553_ clknet_1_1__leaf__0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xseg1._38_ seg1._00_ seg1._11_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2010_ _0028_ clknet_leaf_10_clk cal_lut\[61\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_33_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1725_ _0408_ _0385_ _0409_ _0388_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_79_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1656_ _0247_ _0345_ _0366_ _0362_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xclkbuf_leaf_7_clk clknet_1_1__leaf_clk clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1587_ _0965_ _0322_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2084__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1910__A1 _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2139_ _0157_ clknet_leaf_2_clk cal_lut\[80\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1977__A1 ctr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1420__B _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1968__A1 _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._094_ dec1._027_ dec1._042_ dec1._038_ dec1._041_ dec1._043_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__1196__A2 _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1510_ _0281_ _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_120_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1441_ cal_lut\[43\] _0231_ _0977_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1372_ clknet_1_1__leaf_temp1.i_precharge_n _0870_ _0931_ _0872_ _0932_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_4_clk_I clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1120__A2 _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1187__A2 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1708_ net61 _0386_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1639_ _0230_ _0345_ _0357_ _0348_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1505__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1894__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1350__A2 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1102__A2 _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1990_ _0008_ clknet_leaf_10_clk cal_lut\[41\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._077_ dec1._024_ dec1._025_ dec1._027_ dec1._028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_27_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1169__A2 _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1424_ _0976_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1355_ _0846_ _0915_ _0916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_92_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1286_ ctr\[8\] _0843_ _0852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_92_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2122__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input60_I i_wb_data[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1571__A2 _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2145__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1323__A2 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1140_ cal_lut\[183\] _0630_ _0631_ cal_lut\[51\] _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1071_ cal_lut\[109\] _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1087__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1973_ ctr\[4\] clknet_1_0__leaf__0553_ _0556_ _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_70_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1562__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1407_ _0964_ _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__1314__A2 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1338_ _0563_ ctr\[1\] _0875_ _0901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1269_ en_dbg\[0\] _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2018__CLK clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1002__A1 ctr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2168__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1553__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1792__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1544__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Left_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2172_ _0190_ clknet_leaf_0_clk cal_lut\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1123_ _0690_ _0691_ _0692_ _0693_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_73_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1054_ _0597_ _0594_ _0590_ _0607_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_73_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1075__A4 _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Left_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_38_Left_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1956_ _0348_ _0546_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_31_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1887_ _0963_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_98_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1783__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_131_Right_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1535__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input23_I i_wb_addr[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1299__A1 ctr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1513__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1232__C _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1774__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xseg1._54_ seg1._12_ seg1._22_ seg1._23_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1526__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1810_ _0233_ _0450_ _0463_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_13_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1741_ cal_lut\[145\] _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1672_ _0263_ _0346_ _0374_ _0362_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1765__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1517__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2155_ _0173_ clknet_leaf_11_clk cal_lut\[96\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1106_ cal_lut\[182\] _0630_ _0631_ cal_lut\[50\] _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2086_ _0104_ clknet_leaf_13_clk cal_lut\[187\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_36_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1037_ _0589_ _0590_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_133_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1205__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1939_ o_wb_data[0] _0533_ _0535_ io_out[0] _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1756__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2206__CLK clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_64_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_66_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_73_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xseg1._37_ seg1._00_ seg1._09_ seg1._10_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_82_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_91_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1724_ net35 _0404_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_110_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1655_ cal_lut\[177\] _0356_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1586_ _0562_ _0567_ _0322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1910__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2207_ _0225_ clknet_leaf_6_clk temp_delay_last vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1674__A1 _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2138_ _0156_ clknet_leaf_3_clk cal_lut\[79\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2069_ _0087_ clknet_leaf_17_clk cal_lut\[170\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1426__A1 _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1901__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._093_ dec1.i_bin\[1\] dec1._041_ dec1._042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xtemp1.dac.parallel_cells\[3\].vdac_batch._8_ temp1.dac.parallel_cells\[3\].vdac_batch._0_
+ temp1.dac.parallel_cells\[3\].vdac_batch._1_ temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1440_ net35 _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_1371_ _0563_ _0884_ _0929_ _0930_ _0870_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__1105__B1 _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1656__A1 _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1959__A2 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2051__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1707_ cal_lut\[134\] _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1638_ cal_lut\[169\] _0356_ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1569_ cal_lut\[125\] _0281_ _0298_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1521__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1431__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2074__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1810__A1 _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._076_ dec1._017_ dec1._026_ dec1._027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_50_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1423_ _0964_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_10_Left_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1354_ seg1.o_segments\[5\] _0847_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1285_ ctr\[2\] _0846_ _0848_ _0850_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._3__I temp1.dac.i_data\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1801__A1 _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input53_I i_wb_data[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2097__CLK clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_145_Right_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_clk_I clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1070_ _0593_ _0639_ _0599_ _0640_ _0641_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_99_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1972_ _0590_ clknet_1_0__leaf__0553_ _0976_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xdec1._059_ dec1._003_ dec1._009_ dec1._010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_70_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_140_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1336__B _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1406_ _0963_ _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1337_ _0897_ _0898_ _0899_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_127_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1268_ en_dbg\[1\] _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_36_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1199_ _0593_ cal_lut\[137\] _0766_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1078__A2 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1241__A2 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2112__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2171_ _0189_ clknet_leaf_0_clk cal_lut\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1122_ cal_lut\[176\] _0658_ _0659_ cal_lut\[116\] _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1053_ cal_lut\[43\] _0623_ _0624_ cal_lut\[19\] _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1480__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1955_ o_wb_data[6] _0533_ _0535_ io_out[6] _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1232__A2 _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1886_ cal_lut\[9\] _0506_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__0991__A1 dec1.i_ones vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_102_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input16_I i_wb_addr[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1471__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_111_Left_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_62_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1223__A2 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2135__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1755__I _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._53_ dec1.o_dec\[2\] seg1._13_ seg1._22_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1462__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1740_ _0418_ _0385_ _0419_ _0388_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_40_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1671_ cal_lut\[185\] _0356_ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I i_wb_addr[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2008__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2154_ _0172_ clknet_leaf_10_clk cal_lut\[95\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1105_ cal_lut\[164\] _0626_ _0628_ cal_lut\[122\] _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2085_ _0103_ clknet_leaf_16_clk cal_lut\[186\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1036_ _0587_ _0594_ _0590_ _0607_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__2158__CLK clknet_leaf_8_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1453__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1938_ _0534_ _0533_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1869_ cal_lut\[1\] _0497_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_98_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1692__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_1_1__f__0551_ clknet_0__0551_ clknet_1_1__leaf__0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1444__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._36_ seg1._08_ seg1._09_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_129_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1132__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1683__A2 _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1435__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1199__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1723_ cal_lut\[139\] _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
X_1654_ _0245_ _0345_ _0365_ _0362_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_110_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1585_ _0567_ _0321_ _0965_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2206_ _0224_ clknet_leaf_6_clk dbg3\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2137_ _0155_ clknet_leaf_17_clk cal_lut\[78\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1674__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
X_2068_ _0086_ clknet_leaf_0_clk cal_lut\[169\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1019_ _0589_ _0590_ _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
XANTENNA__1426__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1519__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1114__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1665__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1417__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xdec1._092_ dec1._021_ dec1._023_ dec1._041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[3\].vdac_batch._7_ temp1.dac.i_enable temp1.dac.parallel_cells\[3\].vdac_batch._0_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1050__B1 _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1370_ ctr\[6\] _0853_ _0884_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1656__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1408__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1990__CLK clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1592__A1 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1706_ _0395_ _0385_ _0396_ _0388_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xclkbuf_0__0553_ _0553_ clknet_0__0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_111_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1637_ _0344_ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1568_ _0270_ _0283_ _0313_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1895__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1499_ cal_lut\[62\] _0960_ _0266_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1802__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1335__A1 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1886__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1638__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xdec1._075_ dec1._011_ dec1._014_ dec1._020_ dec1._026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1810__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1574__A1 _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1422_ net61 _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_76_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1353_ _0914_ io_out[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1877__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1284_ seg1.o_segments\[0\] _0849_ _0846_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1629__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1801__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0999_ ctr\[3\] _0564_ _0577_ temp1.dac.i_data\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_26_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input46_I i_wb_data[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1317__A1 ctr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1532__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1253__B1 _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1556__A1 _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2041__CLK clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2191__CLK clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1971_ ctr\[3\] clknet_1_1__leaf__0553_ _0555_ _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1795__A1 _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._058_ dec1.i_bin\[5\] dec1.i_bin\[4\] dec1.i_bin\[6\] dec1._009_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_0_102_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1405_ net68 _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1336_ temp1.dac.i_data\[3\] _0870_ _0872_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput1 i_wb_addr[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1267_ en_dbg\[2\] _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__1078__A3 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1198_ _0589_ _0603_ _0584_ _0580_ _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_19_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2064__CLK clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_clk_I net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1529__A1 _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2170_ _0188_ clknet_leaf_0_clk cal_lut\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1121_ cal_lut\[170\] _0655_ _0656_ cal_lut\[14\] _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_73_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1052_ _0587_ _0591_ _0607_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_73_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1954_ _0348_ _0545_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_22_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1885_ _0495_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_98_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2087__CLK clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1940__A1 _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1319_ ctr\[2\] _0853_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_clkbuf_leaf_2_clk_I clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xseg1._52_ seg1._20_ seg1._21_ seg1.o_segments\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1670_ _0261_ _0346_ _0373_ _0362_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_7_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1922__A1 _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2153_ _0171_ clknet_leaf_10_clk cal_lut\[94\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1104_ cal_lut\[44\] _0623_ _0624_ cal_lut\[20\] _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2084_ _0102_ clknet_leaf_12_clk cal_lut\[185\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1035_ _0583_ _0580_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_91_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1937_ _0946_ _0488_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__1205__A3 _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1868_ _0495_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_31_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1799_ _0973_ _0450_ _0457_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1141__A2 _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2102__CLK clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1766__I cal_lut\[153\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xseg1._35_ dec1.o_dec\[1\] dec1.o_dec\[2\] dec1.o_dec\[0\] seg1._08_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1904__A1 _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1380__A2 _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1450__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1199__A2 cal_lut\[137\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_130_Left_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1722_ _0406_ _0385_ _0407_ _0388_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_13_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1653_ cal_lut\[176\] _0356_ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1584_ ctr\[4\] _0566_ _0321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_119_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2125__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2205_ _0223_ clknet_leaf_7_clk dbg3\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2136_ _0154_ clknet_leaf_18_clk cal_lut\[77\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2067_ _0085_ clknet_leaf_17_clk cal_lut\[168\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1018_ dbg3\[2\] _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_39_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._091_ dec1.i_tens dec1._037_ dec1._038_ dec1._040_ dec1.o_dec\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_54_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref temp1.dac.parallel_cells\[1\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_4
XFILLER_0_40_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[3\].vdac_batch._6_ temp1.dac.parallel_cells\[3\].vdac_batch._2_
+ temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_105_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2148__CLK clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1105__A2 _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1705_ net60 _0386_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1041__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1636_ _0228_ _0345_ _0355_ _0348_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1567_ cal_lut\[124\] _0292_ _0298_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1498_ net55 _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_55_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2119_ _0137_ clknet_leaf_4_clk cal_lut\[156\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1032__A1 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1335__A2 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1712__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1099__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._074_ dec1._018_ dec1._021_ dec1._025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1023__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1574__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1421_ _0973_ _0961_ _0974_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1352_ _0901_ _0913_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1283_ _0833_ en_dbg\[1\] _0835_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__1622__C _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0998_ ctr\[2\] _0564_ _0577_ temp1.dac.i_data\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_26_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1565__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1619_ _0344_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1813__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input39_I i_wb_data[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1556__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1308__A2 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1970_ _0583_ clknet_1_1__leaf__0553_ _0976_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1244__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1795__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._057_ dec1.i_bin\[6\] dec1._002_ dec1._005_ dec1._007_ dec1._008_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_102_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1547__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1404_ _0960_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1335_ _0589_ _0842_ _0840_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput2 i_wb_addr[10] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1266_ _0832_ dec1.i_bin\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_36_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1197_ _0598_ cal_lut\[59\] _0595_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_19_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1859__I _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1543__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1171__B1 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1769__I cal_lut\[154\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1226__A1 _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1777__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1529__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1453__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1120_ cal_lut\[98\] _0652_ _0653_ cal_lut\[146\] _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1162__B1 _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1051_ _0587_ _0589_ _0603_ _0607_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_73_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1900__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1953_ o_wb_data[5] _0533_ _0535_ io_out[5] _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_125_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1768__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1884_ _0228_ _0496_ _0505_ _0430_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1153__B1 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1318_ ctr\[10\] _0881_ _0843_ _0882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_16_Left_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1249_ _0593_ _0599_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_78_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1759__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_25_Left_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xseg1._51_ dec1.o_dec\[1\] seg1._03_ seg1._11_ seg1._01_ seg1._21_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2031__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1931__A2 _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_1_1__f__0902_ clknet_0__0902_ clknet_1_1__leaf__0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2181__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_34_Left_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_144_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_43_Left_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1922__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1686__A1 _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2152_ _0170_ clknet_leaf_10_clk cal_lut\[93\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1103_ cal_lut\[188\] _0620_ _0621_ cal_lut\[104\] _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_2083_ _0101_ clknet_leaf_12_clk cal_lut\[184\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1630__C _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1034_ cal_lut\[55\] _0602_ _0605_ cal_lut\[61\] _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_124_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2054__CLK clknet_leaf_8_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1936_ _0532_ net33 net66 _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_1867_ _0495_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xinput60 i_wb_data[4] net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1798_ cal_lut\[69\] _0451_ _0453_ _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1913__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input21_I i_wb_addr[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1821__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1429__A1 _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._34_ seg1._00_ seg1._02_ seg1._04_ seg1._07_ seg1.o_segments\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1904__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1715__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1668__A1 _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1132__A3 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XTAP_TAPCELL_ROW_73_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._5__A1 temp1.dac.i_enable vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2077__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_51_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1022__I _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1840__A1 _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1721_ net65 _0404_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1199__A3 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1652_ _0243_ _0345_ _0364_ _0362_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_79_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_1_clk_I clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1583_ _0566_ _0320_ _0965_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2204_ _0222_ clknet_leaf_6_clk dbg3\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2135_ _0153_ clknet_leaf_17_clk cal_lut\[76\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_1_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2066_ _0084_ clknet_leaf_13_clk cal_lut\[167\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1017_ dbg3\[3\] _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_48_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1867__I _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1919_ cal_lut\[25\] _0506_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_71_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1898__A1 _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1551__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1114__A3 _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._090_ dec1._029_ dec1._039_ dec1._040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_54_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1822__A1 _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[3\].vdac_batch._5_ temp1.dac.i_enable temp1.dac.parallel_cells\[3\].vdac_batch._1_
+ temp1.dac.parallel_cells\[3\].vdac_batch._2_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1050__A2 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1687__I cal_lut\[129\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_140_Right_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1704_ cal_lut\[133\] _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_53_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0__0551_ _0551_ clknet_0__0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1635_ cal_lut\[168\] _0346_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1566_ _0268_ _0283_ _0312_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1497_ _0272_ _0962_ _0273_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2118_ _0136_ clknet_leaf_4_clk cal_lut\[155\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2049_ _0067_ clknet_leaf_5_clk ctr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_44_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1032__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_8_Left_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._073_ dec1._001_ dec1._021_ dec1._023_ dec1._024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_137_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2115__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1023__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1456__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1420_ cal_lut\[37\] _0962_ _0965_ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1351_ _0910_ _0911_ _0912_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1282_ dec1.i_bin\[0\] _0847_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1262__A2 _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0997_ _0573_ _0576_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_26_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1618_ _0344_ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_41_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1549_ cal_lut\[115\] _0292_ _0298_ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2138__CLK clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1253__A2 _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._056_ dec1.i_bin\[6\] dec1._003_ dec1._006_ dec1._007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_70_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1403_ _0960_ _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1334_ _0856_ _0895_ _0896_ _0884_ _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_127_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1180__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1265_ _0830_ _0831_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xinput3 i_wb_addr[11] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1196_ cal_lut\[167\] _0626_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1483__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_89_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input51_I i_wb_data[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_98_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1474__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0985__A1 ctr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1162__B2 cal_lut\[136\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1162__A1 cal_lut\[154\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1025__I _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1050_ cal_lut\[187\] _0620_ _0621_ cal_lut\[103\] _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_48_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1465__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1952_ _0543_ _0544_ _0348_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_22_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1695__I cal_lut\[130\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1883_ cal_lut\[8\] _0497_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1628__C _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1153__A1 cal_lut\[99\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1317_ ctr\[4\] _0846_ _0879_ _0880_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1248_ _0808_ _0809_ _0814_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_106_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1456__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1179_ cal_lut\[88\] _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_93_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1819__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xseg1._50_ seg1._00_ seg1._19_ seg1._20_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1144__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1447__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._4__A1 temp1.dac.i_data\[4\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1686__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2151_ _0169_ clknet_leaf_10_clk cal_lut\[92\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2082_ _0100_ clknet_leaf_13_clk cal_lut\[183\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1102_ cal_lut\[92\] _0617_ _0618_ cal_lut\[8\] _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1033_ _0587_ _0604_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1438__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1935_ net67 _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_33_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1993__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1866_ _0343_ _0491_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_31_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput61 i_wb_data[5] net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1797_ _0971_ _0450_ _0456_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput50 i_wb_data[24] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_99_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1126__A1 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1677__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input14_I i_wb_addr[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1429__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1549__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._33_ seg1._05_ seg1._06_ seg1._00_ seg1._07_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1668__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1731__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_73_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1459__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1840__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1720_ cal_lut\[138\] _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1053__B1 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1651_ cal_lut\[175\] _0356_ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_21_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1906__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1582_ ctr\[2\] _0565_ ctr\[3\] _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1108__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input6_I i_wb_addr[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1659__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2203_ _0221_ clknet_leaf_5_clk dbg3\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1641__C _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2134_ _0152_ clknet_leaf_17_clk cal_lut\[75\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2065_ _0083_ clknet_leaf_15_clk cal_lut\[166\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2021__CLK clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1016_ _0587_ _0583_ _0580_ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_0_48_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_8_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1831__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2171__CLK clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1918_ _0261_ _0497_ _0523_ _0508_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1849_ cal_lut\[94\] _0449_ _0976_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1347__A1 ctr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1898__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_70_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1822__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[3\].vdac_batch._4_ temp1.dac.i_data\[3\] temp1.dac.i_data\[5\]
+ temp1.dac.parallel_cells\[3\].vdac_batch._1_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_62_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1586__A1 _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1889__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2044__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2194__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1813__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11_clk clknet_1_1__leaf_clk clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1703_ _0393_ _0385_ _0394_ _0388_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_53_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1041__A3 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1634_ _0226_ _0345_ _0354_ _0348_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1636__C _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1329__A1 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1565_ cal_lut\[123\] _0292_ _0298_ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1496_ cal_lut\[61\] _0960_ _0266_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1371__C _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2117_ _0135_ clknet_leaf_4_clk cal_lut\[154\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2048_ _0066_ clknet_leaf_5_clk ctr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__1804__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1568__A1 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_70_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1827__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1032__A3 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2067__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1099__A3 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1788__I _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_0_clk_I clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._072_ dec1._019_ dec1._022_ dec1._017_ dec1._023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_137_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_109_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1023__A3 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1350_ temp1.dac.i_data\[4\] _0870_ _0872_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_118_Left_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1281_ _0833_ en_dbg\[1\] _0835_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
Xclkbuf_leaf_0_clk clknet_1_0__leaf_clk clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1698__I cal_lut\[131\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_127_Left_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0996_ _0575_ _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_41_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1617_ _0337_ _0343_ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_41_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1970__A1 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_136_Left_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1548_ _0249_ _0282_ _0303_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1479_ net49 _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XPHY_EDGE_ROW_145_Left_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1238__B1 _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1557__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1229__B1 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1244__A3 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._055_ dec1.i_bin\[5\] dec1._006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1402_ _0959_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__1914__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1333_ ctr\[3\] _0853_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1264_ cal_lut\[6\] _0786_ cal_ena _0831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput4 i_wb_addr[12] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1195_ cal_lut\[179\] _0658_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0979_ dec1.i_ones dec1.i_tens vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_14_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input44_I i_wb_data[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2105__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0985__A2 ctr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1934__A1 _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1734__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1951_ _0901_ _0913_ _0535_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1882_ _0226_ _0496_ _0504_ _0430_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_22_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_135_Right_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2128__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1153__A2 _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1316_ seg1.o_segments\[2\] _0849_ _0846_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1247_ _0810_ _0811_ _0812_ _0813_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_2_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1178_ cal_lut\[40\] _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_94_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1916__A1 _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1835__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_45_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1080__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._4__A2 temp1.dac.i_data\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1480__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2150_ _0168_ clknet_leaf_10_clk cal_lut\[91\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2081_ _0099_ clknet_leaf_16_clk cal_lut\[182\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1101_ _0666_ _0667_ _0668_ _0671_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1032_ _0589_ _0603_ _0583_ _0581_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_33_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1639__C _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1934_ _0278_ _0497_ _0531_ _0963_ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_16_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput40 i_wb_data[15] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1865_ _0971_ _0493_ _0494_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput62 i_wb_data[6] net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1796_ cal_lut\[68\] _0451_ _0453_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput51 i_wb_data[25] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XTAP_TAPCELL_ROW_50_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xseg1._32_ dec1.o_dec\[1\] seg1._01_ dec1.o_dec\[2\] seg1._06_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1565__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1650_ _0241_ _0345_ _0363_ _0362_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_79_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1581_ _0319_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1108__A2 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1922__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2202_ _0220_ clknet_leaf_6_clk dbg3\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2133_ _0151_ clknet_leaf_14_clk cal_lut\[74\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_1_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2064_ _0082_ clknet_leaf_15_clk cal_lut\[165\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1015_ dbg3\[4\] _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
Xclkbuf_0__0902_ _0902_ clknet_0__0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1292__A1 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1917_ cal_lut\[24\] _0506_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1848_ _0272_ _0451_ _0482_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1779_ _0634_ _0386_ _0445_ _0430_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1404__I _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[3\].vdac_batch._3_ temp1.dac.i_data\[3\] temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__1035__A1 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1983__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1577__A2 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1702_ net59 _0386_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1633_ cal_lut\[167\] _0346_ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1564_ _0265_ _0283_ _0311_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_69_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1495_ net54 _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_39_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1652__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2116_ _0134_ clknet_leaf_4_clk cal_lut\[153\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2047_ _0065_ clknet_leaf_6_clk ctr\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_12_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1265__A1 _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1568__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1032__A4 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1843__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1740__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1256__A1 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._071_ dec1._011_ dec1._014_ dec1._022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1737__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1559__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1023__A4 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2011__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1731__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1280_ _0845_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_92_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2161__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1798__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1262__A4 _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0995_ dec1.i_ones ctr\[9\] _0574_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_26_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1616_ _0338_ _0941_ _0340_ _0342_ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__1722__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1547_ cal_lut\[114\] _0292_ _0298_ _0303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1478_ _0259_ _0962_ _0260_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1238__B2 cal_lut\[102\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1238__A1 cal_lut\[138\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1789__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2034__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1961__A2 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1573__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2184__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xdec1._054_ dec1.i_bin\[6\] dec1._003_ dec1._004_ dec1._005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_11_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1952__A2 _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1401_ _0946_ _0958_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1483__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1332_ ctr\[11\] _0894_ _0843_ _0895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1263_ _0807_ _0815_ _0829_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__1180__A3 _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 i_wb_addr[13] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1930__C _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1194_ cal_lut\[5\] _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_52_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input37_I i_wb_data[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0985__A3 _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1934__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1870__A1 _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1950_ o_wb_data[4] _0533_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1622__A1 _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1881_ cal_lut\[7\] _0497_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1925__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1138__B1 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1315_ _0585_ _0696_ _0847_ _0878_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__1660__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1246_ _0593_ cal_lut\[162\] _0772_ _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_2_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1177_ _0598_ _0745_ _0604_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_106_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1916__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1129__B1 _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1851__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1852__A1 _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_12_Left_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1907__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1135__A3 _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1100_ _0669_ _0670_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_84_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_21_Left_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2080_ _0098_ clknet_leaf_12_clk cal_lut\[181\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_76_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1031_ _0590_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_33_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1933_ cal_lut\[32\] _0495_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_83_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput30 i_wb_addr[7] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1864_ cal_ena _0493_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput63 i_wb_data[7] net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1795_ _0969_ _0450_ _0455_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput41 i_wb_data[16] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput52 i_wb_data[26] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1229_ cal_lut\[83\] _0679_ _0624_ cal_lut\[23\] _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1834__A1 _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._31_ dec1.o_dec\[1\] seg1._01_ seg1._05_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2118__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1580_ _0963_ _0318_ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_95_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1108__A3 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2201_ _0219_ clknet_leaf_5_clk dbg3\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2132_ _0150_ clknet_leaf_14_clk cal_lut\[73\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2063_ _0081_ clknet_leaf_15_clk cal_lut\[164\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1816__A1 _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1014_ cal_lut\[1\] _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1510__I _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1292__A2 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1916_ _0259_ _0497_ _0522_ _0508_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1847_ cal_lut\[93\] _0449_ _0976_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1778_ net54 _0384_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_85_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1035__A2 _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2090__CLK clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1701_ cal_lut\[132\] _0393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1632_ _0975_ _0345_ _0353_ _0348_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1563_ cal_lut\[122\] _0292_ _0298_ _0311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1494_ _0270_ _0962_ _0271_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2115_ _0133_ clknet_leaf_4_clk cal_lut\[152\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2046_ _0064_ clknet_leaf_5_clk ctr\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_36_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input67_I i_wb_we vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_1_1__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1256__A2 _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._070_ dec1._017_ dec1._020_ dec1._019_ dec1._021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_137_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1192__A1 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_18_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_4_Left_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_41_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1928__C _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0994_ ctr\[8\] ctr\[10\] ctr\[11\] ctr\[12\] _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_26_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1955__B1 _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1615_ net1 _0341_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1546_ _0247_ _0282_ _0302_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_5_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1477_ cal_lut\[55\] _0231_ _0977_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1238__A2 _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2029_ _0047_ clknet_leaf_4_clk cal_lut\[112\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1477__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._053_ dec1.i_bin\[3\] dec1._004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_70_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1400_ _0953_ _0954_ _0957_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__1165__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1331_ _0562_ _0846_ _0892_ _0893_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_36_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1262_ _0817_ _0821_ _0822_ _0828_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xinput6 i_wb_addr[14] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1468__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1193_ _0598_ _0585_ _0761_ dec1.i_bin\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_148_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_52_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1996__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1658__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1640__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_58_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1529_ _0230_ _0282_ _0293_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_109_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1459__A2 _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_67_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2001__CLK clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1849__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1631__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2151__CLK clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0979__I dec1.i_ones vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1147__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_85_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_56_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1870__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1622__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1880_ _0975_ _0496_ _0503_ _0430_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_113_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_wire4_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1314_ _0603_ _0585_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2024__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1245_ _0593_ cal_lut\[156\] _0595_ _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__1310__A1 _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1176_ cal_lut\[160\] _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_78_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2174__CLK clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1129__B2 cal_lut\[135\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1129__A1 cal_lut\[153\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1852__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1368__A1 _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2047__CLK clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1135__A4 _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1540__A1 _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_1_1__f__0889_ clknet_0__0889_ clknet_1_1__leaf__0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1030_ _0598_ _0595_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2197__CLK clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1843__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1932_ _0276_ _0497_ _0530_ _0963_ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_140_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1863_ _0383_ _0492_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_141_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput31 i_wb_addr[8] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput20 i_wb_addr[27] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1794_ cal_lut\[67\] _0451_ _0453_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput64 i_wb_data[8] net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput42 i_wb_data[17] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 i_wb_data[27] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1952__B _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1531__A1 _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1228_ cal_lut\[89\] _0795_ _0617_ cal_lut\[95\] _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1834__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1159_ _0585_ _0728_ _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1047__B1 _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xseg1._30_ dec1.o_dec\[0\] seg1._03_ seg1._04_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1522__A1 _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1825__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1589__A1 ctr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1756__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2200_ _0218_ clknet_leaf_7_clk en_dbg\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2131_ _0149_ clknet_leaf_17_clk cal_lut\[72\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2062_ _0080_ clknet_leaf_14_clk cal_lut\[163\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1013_ cal_ena _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XANTENNA__1816__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_32_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1029__B1 _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_14_clk clknet_1_0__leaf_clk clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1915_ cal_lut\[23\] _0506_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1044__A3 _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1666__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1846_ _0270_ _0451_ _0481_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_71_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1777_ _0443_ _0386_ _0444_ _0430_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1201__B1 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input12_I i_wb_addr[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1807__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1701__I cal_lut\[132\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_40_Left_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[1\].vdac_batch._8_ temp1.dac.parallel_cells\[1\].vdac_batch._0_
+ temp1.dac.parallel_cells\[1\].vdac_batch._1_ temp1.dac.parallel_cells\[1\].vdac_batch.en_vref
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1259__B1 _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1700_ _0391_ _0385_ _0392_ _0388_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1631_ cal_lut\[166\] _0346_ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_53_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1562_ _0263_ _0283_ _0310_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1493_ cal_lut\[60\] _0231_ _0266_ _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_3_clk clknet_1_1__leaf_clk clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input4_I i_wb_addr[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2114_ _0132_ clknet_leaf_4_clk cal_lut\[151\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_146_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2045_ _0063_ clknet_leaf_11_clk cal_lut\[128\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_146_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1973__A1 ctr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1829_ cal_lut\[84\] _0461_ _0453_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2108__CLK clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1964__A1 _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1247__A3 _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0993_ ctr\[0\] ctr\[1\] _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1614_ net12 _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1545_ cal_lut\[113\] _0292_ _0298_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1476_ net48 _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_66_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_105_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2028_ _0046_ clknet_leaf_4_clk cal_lut\[111\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_114_Left_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_119_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_17_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_123_Left_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_130_Right_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2080__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_132_Left_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xdec1._052_ dec1.i_bin\[4\] dec1._003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_140_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_141_Left_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1330_ seg1.o_segments\[3\] _0849_ _0846_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1261_ _0824_ _0825_ _0826_ _0827_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_127_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 i_wb_addr[15] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1192_ _0585_ _0760_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_36_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1928__A1 _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1674__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1528_ cal_lut\[105\] _0292_ _0266_ _0293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1459_ cal_lut\[49\] _0231_ _0977_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1092__A1 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1759__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1083__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_1_0__f__0553_ clknet_0__0553_ clknet_1_0__leaf__0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_138_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1313_ _0877_ io_out[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_138_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1244_ _0598_ cal_lut\[36\] _0612_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_47_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1175_ cal_lut\[82\] _0679_ _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_129_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1074__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_12_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1377__A2 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input42_I i_wb_data[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1704__I cal_lut\[133\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_112_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1986__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1540__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1056__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1931_ cal_lut\[31\] _0495_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1862_ _0963_ _0491_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xinput10 i_wb_addr[18] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 i_wb_addr[28] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput32 i_wb_addr[9] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput43 i_wb_data[18] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1793_ _0967_ _0450_ _0454_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput54 i_wb_data[28] net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput65 i_wb_data[9] net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1531__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1227_ _0587_ _0584_ _0580_ _0609_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__2141__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1158_ _0698_ _0592_ _0705_ _0727_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_TAPCELL_ROW_82_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1089_ _0651_ _0654_ _0657_ _0660_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_74_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1770__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1522__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1434__I _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_140_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2014__CLK clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1210__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1761__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1513__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2164__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2130_ _0148_ clknet_leaf_17_clk cal_lut\[71\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2061_ _0079_ clknet_leaf_17_clk cal_lut\[162\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1012_ _0583_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XANTENNA__1029__B2 cal_lut\[133\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1914_ _0257_ _0497_ _0521_ _0508_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_60_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1845_ cal_lut\[92\] _0461_ _0976_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1776_ net53 _0404_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1682__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1752__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2037__CLK clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2187__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1743__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[1\].vdac_batch._7_ temp1.dac.i_enable temp1.dac.parallel_cells\[1\].vdac_batch._0_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_0_temp1.i_precharge_n temp1.i_precharge_n clknet_0_temp1.i_precharge_n vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1630_ _0973_ _0345_ _0352_ _0348_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_53_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_144_Right_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1734__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1561_ cal_lut\[121\] _0292_ _0298_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1492_ net53 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_39_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2113_ _0131_ clknet_leaf_4_clk cal_lut\[150\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2044_ _0062_ clknet_leaf_12_clk cal_lut\[127\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1670__A1 _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1828_ _0251_ _0450_ _0472_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1725__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1186__B1 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1759_ _0431_ _0386_ _0432_ _0430_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_96_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1964__A2 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2202__CLK clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1652__A1 _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0992_ _0572_ temp1.dac.i_enable vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_26_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1955__A2 _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1613_ _0954_ _0339_ _0340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_67_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1544_ _0245_ _0282_ _0301_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1475_ _0257_ _0962_ _0258_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2027_ _0045_ clknet_leaf_3_clk cal_lut\[110\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1643__A1 _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1707__I cal_lut\[134\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1870__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1882__A1 _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1598__B _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1634__A1 _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._051_ dec1.i_bin\[5\] dec1.i_bin\[4\] dec1._002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_118_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1165__A3 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1260_ cal_lut\[192\] _0620_ _0659_ cal_lut\[120\] _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput8 i_wb_addr[16] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1191_ _0730_ _0592_ _0737_ _0759_ _0760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_36_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1625__A1 cal_lut\[163\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1301__B _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1928__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1527__I _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1527_ _0281_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1458_ net41 _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_1389_ net14 net13 net16 net15 _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_93_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1919__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1147__A3 _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1607__A1 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1312_ _0874_ _0876_ _0877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_47_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1243_ cal_lut\[78\] _0610_ _0810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1174_ _0739_ _0740_ _0741_ _0742_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1846__A1 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1074__A2 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2070__CLK clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input35_I i_wb_data[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1720__I cal_lut\[138\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_17_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1828__A1 _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1056__A2 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1930_ _0274_ _0497_ _0529_ _0963_ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1861_ net28 net27 _0490_ _0956_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_TAPCELL_ROW_12_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput11 i_wb_addr[19] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput22 i_wb_addr[29] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput33 i_wb_cyc net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput44 i_wb_data[19] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1792_ cal_lut\[66\] _0451_ _0453_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput55 i_wb_data[29] net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput66 i_wb_stb net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_58_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_0__f_clk clknet_0_clk clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1226_ _0791_ _0792_ _0793_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1157_ _0706_ _0711_ _0721_ _0726_ _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_TAPCELL_ROW_82_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1088_ cal_lut\[175\] _0658_ _0659_ cal_lut\[115\] _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1047__A2 _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1210__A2 cal_lut\[131\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2060_ _0078_ clknet_leaf_14_clk cal_lut\[161\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1011_ dbg3\[1\] _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_60_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1913_ cal_lut\[22\] _0506_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1844_ _0268_ _0451_ _0480_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1775_ cal_lut\[156\] _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1201__A2 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1209_ _0593_ cal_lut\[161\] _0772_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_0_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2189_ _0207_ clknet_leaf_11_clk cal_lut\[32\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0__0889_ _0889_ clknet_0__0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_105_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[1\].vdac_batch._6_ temp1.dac.parallel_cells\[1\].vdac_batch._2_
+ temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1259__A2 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1431__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2131__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1560_ _0261_ _0283_ _0309_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1783__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1491_ _0268_ _0962_ _0269_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2112_ _0130_ clknet_leaf_4_clk cal_lut\[149\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2043_ _0061_ clknet_leaf_13_clk cal_lut\[126\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1999__CLK clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.vdac_single._4__80 net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1670__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1827_ cal_lut\[83\] _0461_ _0453_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1974__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1186__A1 cal_lut\[100\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1758_ net47 _0404_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1689_ _0336_ _0383_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__2004__CLK clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1661__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2154__CLK clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1177__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1652__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0991_ dec1.i_ones ctr\[11\] ctr\[12\] _0571_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_26_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1794__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1612_ _0949_ _0951_ _0952_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_41_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1543_ cal_lut\[112\] _0292_ _0298_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1474_ cal_lut\[54\] _0231_ _0977_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2027__CLK clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XPHY_EDGE_ROW_19_Left_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1891__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2026_ _0044_ clknet_leaf_3_clk cal_lut\[109\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2177__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1643__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Left_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_32_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input65_I i_wb_data[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1159__A1 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._5__A1 temp1.dac.i_enable vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Left_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1331__A1 _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1882__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1095__B1 _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1634__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._050_ dec1.i_bin\[1\] dec1._001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_46_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1119__B _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1570__A1 _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1190_ _0738_ _0743_ _0753_ _0758_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1322__A1 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput9 i_wb_addr[17] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_118_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1789__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1873__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1625__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1526_ _0228_ _0282_ _0291_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1457_ _0245_ _0961_ _0246_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1388_ net26 _0941_ _0945_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1864__A2 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2009_ _0027_ clknet_leaf_11_clk cal_lut\[60\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1552__A1 _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_1_0__f__0551_ clknet_0__0551_ clknet_1_0__leaf__0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_54_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1083__A3 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_138_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1311_ ctr\[0\] _0564_ _0875_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1242_ cal_lut\[96\] _0617_ _0602_ cal_lut\[60\] _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_146_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_139_Right_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1173_ cal_lut\[184\] _0630_ _0631_ cal_lut\[52\] _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1846__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_72_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_144_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1074__A3 _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1538__I _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1782__A1 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_81_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1509_ _0281_ _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_input28_I i_wb_addr[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1837__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_120_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1876__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1828__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1056__A3 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1860_ _0944_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_83_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput12 i_wb_addr[1] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1791_ _0964_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xinput23 i_wb_addr[2] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput34 i_wb_data[0] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput45 i_wb_data[1] net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput56 i_wb_data[2] net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput67 i_wb_we net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1516__A1 _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1225_ cal_lut\[185\] _0630_ _0623_ cal_lut\[47\] _0793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1819__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1156_ _0722_ _0723_ _0724_ _0725_ _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
Xclkbuf_leaf_17_clk clknet_1_0__leaf_clk clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1087_ _0598_ _0591_ _0607_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_90_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1989_ _0007_ clknet_leaf_3_clk cal_lut\[40\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA_clkbuf_leaf_19_clk_I clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1210__A3 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2060__CLK clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1010_ _0582_ dec1.i_bin\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1912_ _0255_ _0497_ _0520_ _0508_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_60_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1843_ cal_lut\[91\] _0461_ _0976_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1774_ _0441_ _0386_ _0442_ _0430_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_114_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_6_clk clknet_1_1__leaf_clk clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_0_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1208_ _0773_ _0774_ _0775_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_79_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2188_ _0206_ clknet_leaf_12_clk cal_lut\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1139_ cal_lut\[165\] _0626_ _0628_ cal_lut\[123\] _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1976__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[1\].vdac_batch._5_ temp1.dac.i_enable temp1.dac.parallel_cells\[1\].vdac_batch._1_
+ temp1.dac.parallel_cells\[1\].vdac_batch._2_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2083__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1900__A1 _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1195__A2 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1490_ cal_lut\[59\] _0231_ _0266_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2111_ _0129_ clknet_leaf_1_clk cal_lut\[148\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_146_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2042_ _0060_ clknet_leaf_13_clk cal_lut\[125\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_71_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1958__A1 _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1826_ _0249_ _0450_ _0471_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1186__A2 _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1757_ cal_lut\[150\] _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1688_ _0338_ net23 _0340_ _0342_ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input10_I i_wb_addr[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_67_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1884__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_73_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0990_ ctr\[10\] _0570_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_26_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1611_ net26 _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_41_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1542_ _0243_ _0282_ _0300_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1473_ net47 _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_5_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I i_wb_addr[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2025_ _0043_ clknet_leaf_17_clk cal_lut\[108\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1809_ cal_lut\[74\] _0461_ _0453_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input58_I i_wb_data[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2121__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1095__B2 cal_lut\[134\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XPHY_EDGE_ROW_101_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1989__CLK clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1570__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1322__A2 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1525_ cal_lut\[104\] _0283_ _0266_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1561__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1456_ cal_lut\[48\] _0231_ _0977_ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1387_ net1 net12 _0944_ _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__2144__CLK clknet_leaf_8_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2008_ _0026_ clknet_leaf_12_clk cal_lut\[59\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_65_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1001__A1 _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1552__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1068__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._101_ dec1._048_ dec1.o_dec\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_123_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2017__CLK clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2167__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1543__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1310_ _0575_ _0837_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_47_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1241_ cal_lut\[150\] _0653_ _0605_ cal_lut\[66\] _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_146_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1172_ cal_lut\[166\] _0626_ _0628_ cal_lut\[124\] _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_2_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1059__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_62_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1782__A2 _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1534__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1508_ net26 net23 _0280_ _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1439_ _0233_ _0961_ _0234_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_85_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1222__A1 _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1892__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1773__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1525__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_temp1.dac._5__A2 temp1.dac.i_data\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput13 i_wb_addr[20] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1790_ _0940_ _0450_ _0452_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_83_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput24 i_wb_addr[30] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 i_wb_data[10] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput46 i_wb_data[20] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput68 reset net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1764__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput57 i_wb_data[30] net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1516__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1323__B _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1224_ _0593_ cal_lut\[155\] _0595_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_74_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1155_ cal_lut\[177\] _0658_ _0659_ cal_lut\[117\] _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1086_ _0597_ _0583_ _0581_ _0609_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_90_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1204__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1988_ _0006_ clknet_leaf_11_clk cal_lut\[39\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1217__C _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input40_I i_wb_data[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1140__B1 _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1746__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1408__B _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2205__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1131__B1 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1682__A1 _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1911_ cal_lut\[21\] _0506_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_60_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1842_ _0265_ _0451_ _0479_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1737__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1773_ net52 _0404_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_100_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_139_Left_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_85_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1207_ cal_lut\[173\] _0655_ _0650_ cal_lut\[143\] _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__1122__B1 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2187_ _0205_ clknet_leaf_11_clk cal_lut\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1138_ cal_lut\[45\] _0623_ _0624_ cal_lut\[21\] _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_148_Left_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_47_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1069_ cal_lut\[85\] _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1728__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[1\].vdac_batch._4_ temp1.dac.i_data\[1\] temp1.dac.i_data\[5\]
+ temp1.dac.parallel_cells\[1\].vdac_batch._1_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1900__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1664__A1 _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1719__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2110_ _0128_ clknet_leaf_1_clk cal_lut\[147\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2041_ _0059_ clknet_leaf_13_clk cal_lut\[124\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1104__B1 _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_18_clk_I clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1825_ cal_lut\[82\] _0461_ _0453_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1756_ _0428_ _0386_ _0429_ _0430_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_111_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1687_ cal_lut\[129\] _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_96_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1894__A1 _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1511__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1949__A2 _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2050__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1101__A3 _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_4
XFILLER_0_26_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1647__I _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1610_ _0336_ _0337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_41_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1168__A3 _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1541_ cal_lut\[111\] _0292_ _0298_ _0300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1472_ _0255_ _0962_ _0256_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1876__A1 _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2024_ _0042_ clknet_leaf_17_clk cal_lut\[107\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1628__A1 _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2073__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1808_ _0230_ _0450_ _0462_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1739_ net40 _0404_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_1_0__f__0902_ clknet_0__0902_ clknet_1_0__leaf__0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_126_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1086__A2 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1524_ _0226_ _0282_ _0290_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_77_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1455_ net40 _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1386_ _0942_ _0943_ _0944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2007_ _0025_ clknet_leaf_11_clk cal_lut\[58\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1068__A2 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._100_ dec1._029_ dec1._044_ dec1._046_ dec1._047_ dec1._000_ dec1._048_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_TAPCELL_ROW_123_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1240_ _0803_ _0804_ _0805_ _0806_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_TAPCELL_ROW_146_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1171_ cal_lut\[46\] _0623_ _0624_ cal_lut\[22\] _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_47_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1059__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_12_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2111__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_120_Left_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1507_ _0945_ _0958_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1438_ cal_lut\[42\] _0231_ _0977_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1369_ _0927_ _0928_ _0919_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_44_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2134__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput14 i_wb_addr[21] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput25 i_wb_addr[31] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput36 i_wb_data[11] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput47 i_wb_data[21] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput58 i_wb_data[31] net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1223_ cal_lut\[77\] _0610_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_67_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1154_ cal_lut\[171\] _0655_ _0656_ cal_lut\[15\] _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1085_ cal_lut\[169\] _0655_ _0656_ cal_lut\[13\] _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_74_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1987_ _0005_ clknet_leaf_3_clk cal_lut\[38\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1204__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input33_I i_wb_cyc vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2007__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2157__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1682__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1910_ _0253_ _0496_ _0519_ _0508_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_60_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1841_ cal_lut\[90\] _0461_ _0976_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1198__A1 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1772_ cal_lut\[155\] _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1370__A1 ctr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1206_ _0598_ cal_lut\[35\] _0612_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_0_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2186_ _0204_ clknet_leaf_11_clk cal_lut\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1137_ cal_lut\[189\] _0620_ _0621_ cal_lut\[105\] _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1673__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1068_ _0598_ _0583_ _0581_ _0635_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__1425__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[1\].vdac_batch._3_ temp1.dac.i_data\[1\] temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1898__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1664__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2040_ _0058_ clknet_leaf_13_clk cal_lut\[123\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1655__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1824_ _0247_ _0450_ _0470_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_4_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1755_ _0963_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_111_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1591__A1 ctr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1686_ _0278_ _0346_ _0381_ _0362_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1343__A1 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1894__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1646__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2169_ _0187_ clknet_leaf_1_clk cal_lut\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1582__A1 ctr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1753__I cal_lut\[149\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1168__A4 _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1540_ _0241_ _0282_ _0299_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1471_ cal_lut\[53\] _0231_ _0977_ _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1876__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2023_ _0041_ clknet_leaf_15_clk cal_lut\[106\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1628__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1800__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1807_ cal_lut\[73\] _0461_ _0453_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1564__A1 _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1738_ cal_lut\[144\] _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_40_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1669_ cal_lut\[184\] _0356_ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_134_Right_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1252__B1 _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_15_Left_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_17_clk_I clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1858__A2 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_24_Left_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_126_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1086__A3 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_33_Left_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1546__A1 _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1523_ cal_lut\[103\] _0283_ _0266_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1454_ _0243_ _0961_ _0244_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_58_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1385_ net32 net31 net3 net2 _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__1849__A2 _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Left_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2040__CLK clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2006_ _0024_ clknet_leaf_12_clk cal_lut\[57\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2190__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input63_I i_wb_data[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1537__A1 _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1517__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_96_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1068__A3 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_123_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2063__CLK clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1170_ cal_lut\[190\] _0620_ _0621_ cal_lut\[106\] _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_63_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1216__B1 _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1519__A1 cal_lut\[101\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1506_ _0278_ _0962_ _0279_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1437_ net65 _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_1368_ _0575_ _0846_ _0844_ _0928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1299_ ctr\[3\] _0846_ _0862_ _0863_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_93_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1800__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1207__B1 _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2086__CLK clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1930__A1 _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput26 i_wb_addr[3] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput15 i_wb_addr[22] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput37 i_wb_data[12] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput59 i_wb_data[3] net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput48 i_wb_data[22] net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1222_ _0786_ _0787_ _0788_ _0789_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_1153_ cal_lut\[99\] _0652_ _0653_ cal_lut\[147\] _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1084_ _0587_ _0584_ _0580_ _0591_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_TAPCELL_ROW_102_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1986_ _0004_ clknet_leaf_7_clk cal_lut\[37\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1204__A3 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_9_clk clknet_1_1__leaf_clk clknet_leaf_9_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_30_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1912__A1 _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input26_I i_wb_addr[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1140__A2 _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1530__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1979__A1 ctr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1131__A2 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2101__CLK clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1840_ _0263_ _0451_ _0478_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_114_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_7_Left_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1198__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1771_ _0439_ _0386_ _0440_ _0430_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_122_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_0__f_temp1.i_precharge_n clknet_0_temp1.i_precharge_n clknet_1_0__leaf_temp1.i_precharge_n
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1205_ _0598_ cal_lut\[65\] _0772_ _0773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2185_ _0203_ clknet_leaf_4_clk cal_lut\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_0_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1122__A2 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1136_ cal_lut\[93\] _0617_ _0618_ cal_lut\[9\] _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1350__B _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1067_ cal_lut\[37\] _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1969_ ctr\[2\] clknet_1_0__leaf__0553_ _0554_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1525__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2124__CLK clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1486__I _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_148_Right_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1435__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1823_ cal_lut\[81\] _0461_ _0453_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1754_ net46 _0404_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_88_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1040__A1 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._7__I temp1.dac.i_enable vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1685_ cal_lut\[192\] _0344_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2147__CLK clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2168_ _0186_ clknet_leaf_2_clk cal_lut\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2099_ _0117_ clknet_leaf_0_clk cal_lut\[136\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1119_ cal_lut\[140\] _0650_ _0592_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_35_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1582__A2 _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1255__B _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1098__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1573__A2 _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_97_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1470_ net46 _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_129_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2022_ _0040_ clknet_leaf_14_clk cal_lut\[105\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1806_ _0449_ _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_31_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1737_ _0416_ _0385_ _0417_ _0388_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1564__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1668_ _0259_ _0346_ _0372_ _0362_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1599_ ctr\[11\] _0571_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1555__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_126_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1491__A1 _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1794__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1522_ _0975_ _0282_ _0289_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1546__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1453_ cal_lut\[47\] _0231_ _0977_ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1384_ net5 net4 net7 net6 _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_26_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2005_ _0023_ clknet_leaf_10_clk cal_lut\[56\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1785__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1537__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input56_I i_wb_data[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1170__B1 _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1068__A4 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1776__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1528__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1700__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1767__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._089_ dec1._001_ dec1._027_ dec1._025_ dec1._039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_42_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1519__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1505_ cal_lut\[64\] _0960_ _0266_ _0279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1436_ _0230_ _0961_ _0232_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_128_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1367_ _0830_ _0831_ _0849_ _0926_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1298_ seg1.o_segments\[1\] _0849_ _0846_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_16_clk_I clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1758__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1528__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1930__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
Xinput27 i_wb_addr[4] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput16 i_wb_addr[23] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1749__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput38 i_wb_data[13] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1438__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput49 i_wb_data[23] net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2030__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1921__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2180__CLK clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1221_ _0594_ _0590_ cal_lut\[29\] _0646_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_1152_ cal_lut\[141\] _0650_ _0592_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1083_ _0587_ _0627_ _0635_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_0_142_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1985_ _0003_ clknet_leaf_15_clk cal_lut\[36\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1204__A4 _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1912__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1419_ net60 _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1125__B1 _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1676__A1 _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1811__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input19_I i_wb_addr[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2053__CLK clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_129_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1600__A1 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_60_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1772__I cal_lut\[155\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1903__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1012__I _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1770_ net51 _0404_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1198__A3 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1658__A1 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1204_ _0594_ _0590_ _0584_ _0580_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_79_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2184_ _0202_ clknet_leaf_4_clk cal_lut\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_108_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1135_ _0699_ _0700_ _0701_ _0704_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1066_ _0598_ _0634_ _0604_ _0636_ _0637_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_34_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2076__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1830__A1 _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1968_ _0580_ clknet_1_0__leaf__0553_ _0976_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_117_Left_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1899_ cal_lut\[15\] _0506_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_126_Left_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1541__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_135_Left_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_53_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_144_Left_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1888__A1 _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2099__CLK clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1812__A1 _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1822_ _0245_ _0450_ _0469_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1753_ cal_lut\[149\] _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1684_ _0276_ _0346_ _0380_ _0362_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1040__A2 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2167_ _0185_ clknet_leaf_11_clk cal_lut\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2098_ _0116_ clknet_leaf_0_clk cal_lut\[135\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1118_ _0680_ _0682_ _0685_ _0688_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_137_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1049_ _0597_ _0583_ _0581_ _0591_ _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_75_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1803__A1 _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1536__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1255__C _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xseg1._49_ dec1.o_dec\[2\] seg1._13_ seg1._12_ seg1._19_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1325__A3 clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2021_ _0039_ clknet_leaf_14_clk cal_lut\[104\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1805_ _0228_ _0450_ _0460_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2114__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1736_ net39 _0404_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1667_ cal_lut\[183\] _0356_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1598_ _0571_ _0328_ _0965_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1252__A2 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1491__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2137__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1243__A2 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1521_ cal_lut\[102\] _0283_ _0266_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1452_ net39 _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__1690__I _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1383_ net23 _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_93_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2004_ _0022_ clknet_leaf_10_clk cal_lut\[55\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1719_ _0403_ _0385_ _0405_ _0388_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_13_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input49_I i_wb_data[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch._8_ temp1.dac.parallel_cells\[4\].vdac_batch._0_
+ temp1.dac.parallel_cells\[4\].vdac_batch._1_ temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__1170__B2 cal_lut\[106\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1225__A2 _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1775__I cal_lut\[156\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1216__A2 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._088_ dec1.i_bin\[1\] dec1._028_ dec1._038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_12_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.inv1_1 temp1.dcdel_capnode_notouch_ net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_88_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1504_ net58 _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_0_10_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1435_ cal_lut\[41\] _0231_ _0977_ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1366_ seg1.o_segments\[6\] _0849_ _0846_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1297_ _0585_ _0663_ _0847_ _0861_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_77_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1207__A2 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1809__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1694__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput28 i_wb_addr[5] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xinput17 i_wb_addr[24] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput39 i_wb_data[14] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1220_ cal_lut\[11\] _0618_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1151_ _0712_ _0714_ _0717_ _0720_ _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_TAPCELL_ROW_134_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1685__A2 _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1082_ cal_lut\[97\] _0652_ _0653_ cal_lut\[145\] _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_23_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1984_ _0002_ clknet_leaf_14_clk cal_lut\[35\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1373__A1 temp1.dac.i_enable vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1364__B _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1418_ _0971_ _0961_ _0972_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1676__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1349_ _0593_ _0842_ _0840_ _0911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_3_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1428__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1992__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1539__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1364__A1 temp1.dac.i_data\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1116__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1667__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._4__A2 temp1.dac.i_data\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1198__A4 _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_15_clk_I clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1203_ _0769_ _0770_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1107__A1 _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1658__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2183_ _0201_ clknet_leaf_4_clk cal_lut\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1134_ _0702_ _0703_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1065_ cal_lut\[79\] _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1830__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ _0552_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1594__A1 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1898_ _0241_ _0496_ _0513_ _0508_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_113_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1897__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input31_I i_wb_addr[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1649__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2020__CLK clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1821__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dcdc temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ clknet_1_0__leaf_temp1.i_precharge_n
+ temp1.dcdel_capnode_notouch_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_1
XANTENNA__2170__CLK clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1034__B1 _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1888__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1812__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1821_ cal_lut\[80\] _0461_ _0453_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_4_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1576__A1 _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1752_ _0426_ _0385_ _0427_ _0388_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xclkbuf_leaf_10_clk clknet_1_1__leaf_clk clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1693__I _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1683_ cal_lut\[191\] _0344_ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1040__A3 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1626__C _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1328__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1879__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2043__CLK clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2166_ _0184_ clknet_leaf_11_clk cal_lut\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1500__A1 _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1117_ _0686_ _0645_ _0687_ _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2097_ _0115_ clknet_leaf_0_clk cal_lut\[134\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__2193__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1048_ _0597_ _0609_ _0607_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__1868__I _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1803__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1817__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1319__A1 ctr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_1_1__f_clk clknet_0_clk clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1098__A3 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1558__A1 _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._48_ seg1._18_ seg1.o_segments\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2066__CLK clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1462__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2020_ _0038_ clknet_leaf_14_clk cal_lut\[103\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1797__A1 _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1261__A3 _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1804_ cal_lut\[72\] _0451_ _0453_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1735_ cal_lut\[143\] _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_79_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1666_ _0257_ _0346_ _0371_ _0362_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1597_ ctr\[10\] _0570_ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2149_ _0167_ clknet_leaf_7_clk cal_lut\[90\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1547__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1004__A3 clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2089__CLK clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1960__A1 _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1228__B1 _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp_sensor_70 io_oeb[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_109_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1520_ _0973_ _0282_ _0288_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1451_ _0241_ _0961_ _0242_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1382_ net34 _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XANTENNA__1904__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_1_1__f_net81 clknet_0_net81 clknet_1_1__leaf_net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_109_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2003_ _0021_ clknet_leaf_12_clk cal_lut\[54\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_11_Left_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_132_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_1_0__f__0889_ clknet_0__0889_ clknet_1_0__leaf__0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1718_ net64 _0404_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1649_ cal_lut\[174\] _0356_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xwire4 clk net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch._7_ temp1.dac.i_enable temp1.dac.parallel_cells\[4\].vdac_batch._0_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1170__A2 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2104__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1031__I _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xdec1._087_ dec1._009_ dec1._031_ dec1._036_ dec1._037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_42_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1503_ _0276_ _0962_ _0277_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1924__A1 _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1634__C _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1434_ _0960_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_137_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1365_ ctr\[0\] ctr\[1\] _0875_ _0924_ _0925_ io_out[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__1152__A2 _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1296_ _0584_ _0585_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input61_I i_wb_data[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1825__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2127__CLK clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XTAP_TAPCELL_ROW_111_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1719__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 i_wb_addr[25] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput29 i_wb_addr[6] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1906__A1 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1150_ _0718_ _0645_ _0719_ _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_134_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._5__A1 temp1.dac.i_enable vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1081_ _0587_ _0589_ _0603_ _0627_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_0_90_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1983_ _0001_ clknet_leaf_17_clk cal_lut\[34\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1070__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1373__A2 _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_143_Right_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1417_ cal_lut\[36\] _0962_ _0965_ _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1125__A2 _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1348_ _0856_ _0908_ _0909_ _0884_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1279_ _0833_ en_dbg\[1\] _0838_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_TAPCELL_ROW_81_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1061__A1 _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1555__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1364__A2 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1116__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1052__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1465__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1202_ cal_lut\[101\] _0652_ _0653_ cal_lut\[149\] _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1912__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2182_ _0200_ clknet_leaf_4_clk cal_lut\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1133_ _0593_ cal_lut\[129\] _0612_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_125_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1064_ _0598_ _0584_ _0580_ _0635_ _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1966_ temp_delay_last clknet_1_0__leaf__0551_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1897_ cal_lut\[14\] _0506_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input24_I i_wb_addr[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_3_Left_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_91_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_49_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1820_ _0243_ _0450_ _0468_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1576__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1751_ net44 _0404_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1682_ _0274_ _0346_ _0379_ _0362_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1040__A4 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1328__A2 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1982__CLK clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2165_ _0183_ clknet_leaf_11_clk cal_lut\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1500__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1116_ _0594_ _0590_ cal_lut\[26\] _0646_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_2096_ _0114_ clknet_leaf_19_clk cal_lut\[133\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1047_ cal_lut\[91\] _0617_ _0618_ cal_lut\[7\] _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1016__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1949_ _0541_ _0542_ _0348_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1567__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1833__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1255__A1 _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_14_clk_I clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_57_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1558__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._47_ seg1._16_ seg1._17_ seg1._18_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_66_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_66_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1730__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xtemp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1494__A1 _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1246__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1797__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_75_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_142_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1803_ _0226_ _0450_ _0459_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_31_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1549__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1734_ _0414_ _0385_ _0415_ _0388_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_40_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1665_ cal_lut\[182\] _0356_ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1596_ _0570_ _0327_ _0965_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2010__CLK clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1372__C _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1721__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2160__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2148_ _0166_ clknet_leaf_10_clk cal_lut\[89\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2079_ _0097_ clknet_leaf_16_clk cal_lut\[180\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_93_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1960__A2 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1563__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1712__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1173__B1 _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1779__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp_sensor_71 io_oeb[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_109_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2033__CLK clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1450_ cal_lut\[46\] _0231_ _0977_ _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1381_ _0872_ _0938_ _0939_ io_out[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2183__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1164__B1 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1703__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2002_ _0020_ clknet_leaf_13_clk cal_lut\[53\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1920__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1219__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1717_ _0384_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_6_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1648_ _0239_ _0345_ _0361_ _0362_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch._6_ temp1.dac.parallel_cells\[4\].vdac_batch._2_
+ temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__1155__B1 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1579_ ctr\[2\] _0565_ _0318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_138_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1630__A1 _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1933__A2 _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1740__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_114_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1468__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._086_ dec1._017_ dec1._020_ dec1._035_ dec1._036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_42_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1502_ cal_lut\[63\] _0960_ _0266_ _0277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1924__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1433_ net64 _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_10_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1137__B1 _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1364_ temp1.dac.i_data\[5\] _0870_ _0872_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1295_ _0837_ _0859_ _0860_ io_out[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_37_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1650__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2079__CLK clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1915__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input54_I i_wb_data[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1841__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1603__A1 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Left_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput19 i_wb_addr[26] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1906__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1080_ _0587_ _0627_ _0644_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XTAP_TAPCELL_ROW_35_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_23_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1842__A1 _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1982_ _0000_ clknet_leaf_14_clk cal_lut\[33\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xdec1._069_ dec1._011_ dec1._014_ dec1._018_ dec1._019_ dec1._020_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_15_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1645__C _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1416_ net59 _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_48_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1347_ ctr\[4\] _0853_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_3_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1278_ _0843_ _0844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_81_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1887__I _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1571__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1824__A1 _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_107_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_1_0__f_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1201_ cal_lut\[191\] _0620_ _0659_ cal_lut\[119\] _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2181_ _0199_ clknet_leaf_11_clk cal_lut\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1132_ _0598_ cal_lut\[33\] _0612_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1063_ _0589_ _0590_ _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_87_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_140_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1965_ net82 _0565_ _0575_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_7_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2117__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1896_ _0239_ _0496_ _0512_ _0508_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_113_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input17_I i_wb_addr[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_104_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_113_Left_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_29_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1750_ cal_lut\[148\] _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_122_Left_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1681_ cal_lut\[190\] _0344_ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input9_I i_wb_addr[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_131_Left_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2164_ _0182_ clknet_leaf_11_clk cal_lut\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1115_ cal_lut\[110\] _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2095_ _0113_ clknet_leaf_18_clk cal_lut\[132\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1046_ _0587_ _0583_ _0581_ _0591_ _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_75_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1264__A2 _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1016__A2 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1948_ _0900_ clknet_1_0__leaf__0902_ _0535_ _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1879_ cal_lut\[6\] _0497_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_101_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._46_ dec1.o_dec\[1\] dec1.o_dec\[0\] dec1.o_dec\[2\] seg1._11_ seg1._17_ vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__1743__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1494__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1802_ cal_lut\[71\] _0451_ _0453_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1918__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1733_ net38 _0404_ _0415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1664_ _0255_ _0346_ _0370_ _0362_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1595_ ctr\[8\] _0569_ ctr\[9\] _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1182__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2147_ _0165_ clknet_leaf_10_clk cal_lut\[88\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2078_ _0096_ clknet_leaf_15_clk cal_lut\[179\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_138_Right_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1237__A2 _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1029_ cal_lut\[151\] _0596_ _0600_ cal_lut\[133\] _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_72_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref temp1.dac.parallel_cells\[0\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_63_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xtemp_sensor_72 io_oeb[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0987__A1 _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._29_ dec1.o_dec\[2\] seg1._03_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1380_ net83 _0872_ _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_93_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2001_ _0019_ clknet_leaf_16_clk cal_lut\[52\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1648__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1716_ cal_lut\[137\] _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1647_ _0963_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_6_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch._5_ temp1.dac.i_enable temp1.dac.parallel_cells\[4\].vdac_batch._1_
+ temp1.dac.parallel_cells\[4\].vdac_batch._2_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1578_ _0565_ _0573_ _0965_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_13_clk_I clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1995__CLK clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1839__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1630__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1091__B1 _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_temp1.dac._4__I temp1.dac.i_enable vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1697__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2000__CLK clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1082__B1 _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._085_ dec1._032_ dec1._034_ dec1._035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_103_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2150__CLK clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1501_ net57 _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_1432_ _0228_ _0961_ _0229_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_128_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1363_ _0870_ _0923_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_37_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1294_ _0565_ _0575_ _0837_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_38_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1378__C _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1376__A1 ctr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input47_I i_wb_data[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1679__A2 _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2023__CLK clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1851__A2 _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1569__B _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2173__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1367__A1 _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1842__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1981_ _0965_ clknet_1_1__leaf__0551_ _0560_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xdec1._068_ dec1.i_bin\[2\] dec1._019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1070__A3 _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1926__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1358__A1 dec1.i_ones vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1415_ _0969_ _0961_ _0970_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_47_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1942__B _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2046__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1346_ ctr\[12\] _0907_ _0843_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1530__A1 cal_lut\[106\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1277_ _0833_ _0834_ _0835_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__2196__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1833__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1349__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1116__A4 _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1521__A1 cal_lut\[102\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1824__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1588__A1 _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1746__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2069__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1200_ _0763_ _0764_ _0765_ _0767_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2180_ _0198_ clknet_leaf_3_clk cal_lut\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1512__A1 _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1131_ cal_lut\[69\] _0608_ _0610_ cal_lut\[75\] _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1062_ cal_lut\[157\] _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1815__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_13_clk clknet_1_0__leaf_clk clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1964_ _0969_ _0493_ _0550_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1579__A1 ctr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1895_ cal_lut\[13\] _0506_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1656__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1503__A1 _0276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1329_ _0585_ _0728_ _0847_ _0891_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_91_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1847__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1582__B ctr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1981__A1 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1680_ _0272_ _0346_ _0378_ _0362_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_111_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2_clk clknet_1_0__leaf_clk clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2163_ _0181_ clknet_leaf_7_clk cal_lut\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1114_ _0593_ _0683_ _0599_ _0640_ _0684_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2094_ _0112_ clknet_leaf_19_clk cal_lut\[131\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1045_ _0587_ _0609_ _0607_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_90_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1947_ o_wb_data[3] _0533_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1016__A3 _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1878_ _0973_ _0496_ _0502_ _0430_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1972__A1 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._7__I temp1.dac.i_enable vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._45_ dec1.o_dec\[2\] seg1._12_ seg1._09_ seg1._00_ seg1._13_ seg1._16_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1191__A2 _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2107__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1246__A3 _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1801_ _0975_ _0450_ _0458_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1487__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1732_ cal_lut\[142\] _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1954__A1 _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1663_ cal_lut\[181\] _0356_ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1934__C _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1594_ _0965_ _0326_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1182__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2146_ _0164_ clknet_leaf_10_clk cal_lut\[87\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2077_ _0095_ clknet_leaf_2_clk cal_lut\[178\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1028_ _0598_ _0599_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_72_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1173__A2 _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0987__A2 ctr\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp_sensor_73 io_oeb[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_109_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._28_ dec1.o_dec\[1\] seg1._01_ dec1.o_dec\[2\] seg1._02_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_22_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1164__A2 _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2000_ _0018_ clknet_leaf_16_clk cal_lut\[51\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_117_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1219__A3 _0766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1945__B _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1715_ _0401_ _0385_ _0402_ _0388_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_115_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1646_ cal_lut\[173\] _0356_ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1664__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1577_ ctr\[0\] _0965_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xtemp1.dac.parallel_cells\[4\].vdac_batch._4_ temp1.dac.i_data\[4\] temp1.dac.i_data\[5\]
+ temp1.dac.parallel_cells\[4\].vdac_batch._1_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1155__A2 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2129_ _0147_ clknet_leaf_17_clk cal_lut\[70\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1918__A1 _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_114_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1749__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1082__A1 cal_lut\[97\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._084_ dec1._033_ dec1._015_ dec1._031_ dec1._034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1500_ _0274_ _0962_ _0275_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1431_ cal_lut\[40\] _0962_ _0977_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1137__A2 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1362_ dbg3\[5\] _0884_ _0920_ _0922_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1293_ temp1.dac.i_data\[0\] _0840_ _0858_ _0859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1073__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1629_ cal_lut\[165\] _0346_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1064__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1585__B _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1119__A2 _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1980_ _0563_ _0564_ _0576_ temp_delay_last _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_23_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1055__A1 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._067_ dec1.i_bin\[3\] dec1._008_ dec1._018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_clkbuf_leaf_12_clk_I clknet_1_0__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1414_ cal_lut\[35\] _0962_ _0965_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1985__CLK clknet_leaf_15_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1345_ ctr\[6\] _0846_ _0905_ _0906_ _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1530__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1276_ _0833_ _0841_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_3_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1294__A1 _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1046__A1 _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1349__A2 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1424__I _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1521__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2140__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1285__A1 ctr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1037__A1 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1762__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1512__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1130_ cal_lut\[57\] _0602_ _0605_ cal_lut\[63\] _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1061_ _0622_ _0625_ _0629_ _0632_ _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_34_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1028__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1963_ _0833_ _0493_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1894_ _0237_ _0496_ _0511_ _0508_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1579__A2 _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1509__I _0281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2013__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1672__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1751__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2163__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1503__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1328_ _0594_ _0585_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1259_ cal_lut\[72\] _0608_ _0621_ cal_lut\[108\] _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_148_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1019__A1 _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_18_Left_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1742__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1258__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_27_Left_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xtemp1.dac.vdac_single._4__79 net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2036__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_36_Left_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2186__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1733__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1497__A1 _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2162_ _0180_ clknet_leaf_8_clk cal_lut\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2093_ _0111_ clknet_leaf_19_clk cal_lut\[130\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1113_ cal_lut\[86\] _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_45_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1044_ _0601_ _0606_ _0611_ _0615_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1249__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1948__B _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1946_ _0539_ _0540_ _0348_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1421__A1 _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1877_ cal_lut\[5\] _0497_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_3_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1724__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input22_I i_wb_addr[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1488__A1 _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1660__A1 _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1412__A1 _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1963__A2 _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._44_ seg1._03_ seg1._00_ seg1._08_ seg1.o_segments\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1715__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1800_ cal_lut\[70\] _0451_ _0453_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1731_ _0412_ _0385_ _0413_ _0388_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_40_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1662_ _0253_ _0345_ _0369_ _0362_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1593_ ctr\[8\] _0569_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1706__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_53_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2145_ _0163_ clknet_leaf_7_clk cal_lut\[86\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2201__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2076_ _0094_ clknet_leaf_2_clk cal_lut\[177\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1890__A1 _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1027_ _0594_ _0590_ _0583_ _0581_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XPHY_EDGE_ROW_62_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1929_ cal_lut\[30\] _0495_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_71_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp_sensor_74 io_oeb[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_109_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._27_ dec1.o_dec\[0\] seg1._01_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_22_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1872__A1 _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_18_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1624__A1 _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1714_ net63 _0386_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1927__A2 _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1645_ _0237_ _0345_ _0360_ _0348_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_13_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1576_ _0278_ _0283_ _0317_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.parallel_cells\[4\].vdac_batch._3_ temp1.dac.i_data\[4\] temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XANTENNA__1680__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2128_ _0146_ clknet_leaf_17_clk cal_lut\[69\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2059_ _0077_ clknet_leaf_9_clk dec1.i_ones vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_64_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1091__A2 _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1918__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_87_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1854__A1 _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA__1606__A1 temp1.dac.i_enable vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xdec1._083_ dec1.i_bin\[4\] dec1._009_ dec1.i_bin\[3\] dec1._033_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1082__A2 _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1909__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1765__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1430_ net63 _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_128_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1361_ _0884_ _0921_ _0922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1292_ _0581_ _0842_ _0854_ _0857_ _0840_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_37_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1073__A2 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1628_ _0971_ _0345_ _0351_ _0348_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_78_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1559_ cal_lut\[120\] _0292_ _0298_ _0309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_69_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1836__A1 _0259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1710__I cal_lut\[135\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1064__A2 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0996__I _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1055__A2 _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xdec1._066_ dec1._011_ dec1._014_ dec1._016_ dec1._017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1413_ net56 _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_48_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1344_ seg1.o_segments\[4\] _0849_ _0846_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_66_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1275_ en_dbg\[1\] _0835_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__1818__A1 _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1294__A2 _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1046__A2 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2092__CLK clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input52_I i_wb_data[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1037__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1596__B _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1060_ cal_lut\[181\] _0630_ _0631_ cal_lut\[49\] _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1028__A2 _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1962_ _0967_ _0493_ _0549_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1893_ cal_lut\[12\] _0506_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_50_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._049_ dec1.i_tens dec1._000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_0_119_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1327_ _0890_ io_out[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_75_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1258_ _0593_ cal_lut\[132\] _0612_ _0825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1189_ _0754_ _0755_ _0756_ _0757_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1019__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_11_clk_I clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1258__A2 cal_lut\[132\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_133_Right_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_139_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1497__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2161_ _0179_ clknet_leaf_7_clk cal_lut\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2092_ _0110_ clknet_leaf_18_clk cal_lut\[129\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1112_ cal_lut\[38\] _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1043_ _0613_ _0614_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1249__A2 _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
X_1945_ _0888_ clknet_1_0__leaf__0889_ _0535_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1957__B1 _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1421__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1876_ _0971_ _0496_ _0501_ _0430_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2130__CLK clknet_leaf_17_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1488__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input15_I i_wb_addr[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1998__CLK clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0999__A1 ctr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1660__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1412__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._43_ seg1._10_ seg1._15_ seg1.o_segments\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2003__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1651__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1768__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2153__CLK clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1939__B1 _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1730_ net37 _0404_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1661_ cal_lut\[180\] _0356_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1592_ _0965_ _0325_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1182__A4 _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input7_I i_wb_addr[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_0_Left_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2144_ _0162_ clknet_leaf_8_clk cal_lut\[85\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2075_ _0093_ clknet_leaf_2_clk cal_lut\[176\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1890__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1026_ _0597_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1642__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1678__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1928_ _0272_ _0497_ _0528_ _0963_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_31_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1859_ _0489_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1713__I cal_lut\[136\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2026__CLK clknet_leaf_3_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1881__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2176__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1633__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp_sensor_75 io_oeb[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_109_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._26_ dec1.o_dec\[3\] seg1._00_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_132_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1149__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1872__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1085__B1 _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1624__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_115_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1713_ cal_lut\[136\] _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_13_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1644_ cal_lut\[172\] _0356_ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_6_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1575_ cal_lut\[128\] _0281_ _0298_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2049__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1560__A1 _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2199__CLK clknet_leaf_7_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2127_ _0145_ clknet_leaf_15_clk cal_lut\[68\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2058_ _0076_ clknet_leaf_9_clk ctr\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1009_ _0581_ cal_ena _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_64_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1379__A1 temp1.dac.i_enable vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1303__A1 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1854__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_122_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_15_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._082_ dec1._009_ dec1._032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_23_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1618__I _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1790__A1 _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1781__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1360_ _0562_ _0856_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1542__A1 _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1291_ ctr\[0\] _0856_ _0842_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1845__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_90_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1073__A3 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
X_1627_ cal_lut\[164\] _0346_ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_111_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1972__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1533__A1 _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1558_ _0259_ _0283_ _0308_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_69_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1489_ net52 _0268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XPHY_EDGE_ROW_129_Left_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1836__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1064__A3 _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_138_Left_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_20_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1524__A1 _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_147_Left_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1827__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xdec1._065_ dec1._005_ dec1._015_ dec1._012_ dec1._016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1792__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1412_ _0967_ _0961_ _0968_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1515__A1 cal_lut\[99\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1343_ _0585_ _0760_ _0847_ _0904_ _0905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1274_ _0833_ _0839_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_147_Right_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1818__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_16_clk clknet_1_0__leaf_clk clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_80_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1686__C _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1046__A3 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0989_ ctr\[9\] ctr\[8\] _0569_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_input45_I i_wb_data[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1506__A1 _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1809__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1961_ en_dbg\[1\] _0493_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1892_ _0235_ _0496_ _0510_ _0508_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1806__I _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_5_clk clknet_1_1__leaf_clk clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1326_ _0888_ clknet_1_1__leaf__0889_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_75_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1257_ _0593_ cal_lut\[114\] _0644_ _0823_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_1188_ cal_lut\[178\] _0658_ _0659_ cal_lut\[118\] _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_78_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1975__A1 _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1716__I cal_lut\[137\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1258__A3 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2082__CLK clknet_leaf_13_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2160_ _0178_ clknet_leaf_11_clk cal_lut\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2091_ _0109_ clknet_leaf_12_clk cal_lut\[192\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1111_ _0598_ _0681_ _0604_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1042_ _0593_ cal_lut\[127\] _0612_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1944_ o_wb_data[2] _0533_ _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1875_ cal_lut\[4\] _0497_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_101_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1185__A2 _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1309_ _0867_ _0868_ _0873_ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._42_ seg1._11_ seg1._14_ seg1._15_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1874__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1660_ _0251_ _0345_ _0368_ _0362_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_103_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1591_ ctr\[7\] _0568_ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_56_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2143_ _0161_ clknet_leaf_2_clk cal_lut\[84\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2074_ _0092_ clknet_leaf_17_clk cal_lut\[175\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1025_ _0587_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_8
XFILLER_0_72_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1927_ cal_lut\[29\] _0495_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1694__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1858_ net66 _0965_ _0946_ _0488_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XANTENNA_clkbuf_leaf_10_clk_I clknet_1_1__leaf_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._4__A2 temp1.dac.i_data\[5\] vdd
+ vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1789_ cal_lut\[65\] _0451_ _0298_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1158__A2 _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_110_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_109_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp_sensor_76 io_oeb[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_117_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1149__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1779__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2120__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1712_ _0399_ _0385_ _0400_ _0388_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1643_ _0235_ _0345_ _0359_ _0348_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_6_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1574_ _0276_ _0283_ _0316_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1988__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1560__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2126_ _0144_ clknet_leaf_14_clk cal_lut\[67\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2057_ _0075_ clknet_leaf_9_clk ctr\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtemp1.dac.parallel_cells\[2\].vdac_batch._8_ temp1.dac.parallel_cells\[2\].vdac_batch._0_
+ temp1.dac.parallel_cells\[2\].vdac_batch._1_ temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1008_ _0580_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_8
XFILLER_0_8_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1379__A2 _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1000__A1 ctr\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1551__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2143__CLK clknet_leaf_2_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1303__A2 _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].pupd temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
Xdec1._081_ dec1._017_ dec1._020_ dec1._031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_128_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1790__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1542__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1290_ _0835_ _0855_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XTAP_TAPCELL_ROW_46_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.vdac_single._8_ temp1.dac.vdac_single._0_ temp1.dac.vdac_single._1_ temp1.dac.vdac_single.en_vref
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2016__CLK clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1626_ _0969_ _0345_ _0350_ _0348_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1781__A2 _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1557_ cal_lut\[119\] _0292_ _0298_ _0308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2166__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1533__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1488_ _0265_ _0962_ _0267_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_94_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1297__A1 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2109_ _0127_ clknet_leaf_1_clk cal_lut\[146\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1064__A4 _0635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1221__A1 _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1882__C _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1524__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2039__CLK clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1460__A1 _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._064_ dec1.i_bin\[4\] dec1._009_ dec1.i_bin\[5\] dec1._015_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2189__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1411_ cal_lut\[34\] _0962_ _0965_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1515__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1342_ _0598_ _0585_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1273_ en_dbg\[1\] _0838_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1451__A1 _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0988_ _0561_ _0568_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1754__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1609_ net28 _0944_ _0335_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__1506__A2 _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input38_I i_wb_data[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1442__A1 _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1745__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1130__B1 _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1960_ _0940_ _0493_ _0548_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1891_ cal_lut\[11\] _0506_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1736__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1308__B _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1325_ _0563_ ctr\[1\] clknet_leaf_6_clk _0875_ _0889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__2204__CLK clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1256_ _0584_ _0580_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1121__B1 _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1187_ cal_lut\[172\] _0655_ _0656_ cal_lut\[16\] _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1672__A1 _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1978__B _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1697__C _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1727__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1188__B1 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1415__A1 _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1718__A2 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1110_ cal_lut\[158\] _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_136_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2090_ _0108_ clknet_leaf_13_clk cal_lut\[191\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1103__B1 _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1041_ _0598_ cal_lut\[31\] _0612_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1798__B _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1654__A1 _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_14_Left_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1943_ _0537_ _0538_ _0348_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1957__A2 _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1874_ _0969_ _0496_ _0500_ _0430_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1709__A2 _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_23_Left_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1308_ temp1.dac.i_data\[1\] _0870_ _0872_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1239_ cal_lut\[90\] _0795_ _0624_ cal_lut\[24\] _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__1645__A1 _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_32_Left_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._5__A1 temp1.dac.i_enable vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xseg1._41_ dec1.o_dec\[2\] seg1._12_ seg1._13_ seg1._14_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_EDGE_ROW_41_Left_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1890__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1884__A1 _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1636__A1 _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1411__B _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1939__A2 _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1637__I _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1590_ _0965_ _0324_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2142_ _0160_ clknet_leaf_2_clk cal_lut\[83\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2073_ _0091_ clknet_leaf_17_clk cal_lut\[174\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1024_ _0593_ _0595_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_16_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1926_ _0270_ _0497_ _0527_ _0508_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1857_ _0953_ _0487_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_112_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1788_ _0449_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_97_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input20_I i_wb_addr[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp_sensor_77 o_wb_stall vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__2072__CLK clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1085__A2 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1711_ net62 _0386_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_108_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1642_ cal_lut\[171\] _0356_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_123_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1573_ cal_lut\[127\] _0281_ _0298_ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1848__A1 _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2125_ _0143_ clknet_leaf_2_clk cal_lut\[66\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2056_ _0074_ clknet_leaf_9_clk ctr\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtemp1.dac.parallel_cells\[2\].vdac_batch._7_ temp1.dac.i_enable temp1.dac.parallel_cells\[2\].vdac_batch._0_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1007_ dbg3\[0\] _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2095__CLK clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1909_ cal_lut\[20\] _0506_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input68_I reset vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xdec1._080_ dec1._000_ dec1._028_ dec1._029_ dec1._030_ dec1.o_dec\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XTAP_TAPCELL_ROW_23_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_105_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1058__A2 _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtemp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
Xtemp1.dac.vdac_single._7_ temp1.dac._0_ temp1.dac.vdac_single._0_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1625_ cal_lut\[163\] _0346_ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1556_ _0257_ _0283_ _0307_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1487_ cal_lut\[58\] _0231_ _0266_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Left_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2108_ _0126_ clknet_leaf_0_clk cal_lut\[145\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2039_ _0057_ clknet_leaf_16_clk cal_lut\[122\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1049__A2 _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1221__A2 _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2110__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1460__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xdec1._063_ dec1._013_ dec1._014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_125_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1410_ net45 _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_3
X_1341_ _0903_ io_out[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1272_ _0835_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1451__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2133__CLK clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0987_ _0562_ ctr\[6\] _0567_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_131_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1608_ net27 _0956_ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1539_ cal_lut\[110\] _0292_ _0298_ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_72_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1442__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1414__B _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_69_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2006__CLK clknet_leaf_12_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1681__A2 _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2156__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_78_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1890_ _0233_ _0496_ _0509_ _0508_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].pupd temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_70_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1197__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1324_ _0885_ _0886_ _0887_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_EDGE_ROW_87_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].pupd temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
+ temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1255_ _0603_ cal_lut\[30\] _0646_ _0594_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1186_ cal_lut\[100\] _0652_ _0653_ cal_lut\[148\] _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_91_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1672__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_96_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input50_I i_wb_data[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2029__CLK clknet_leaf_4_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1360__A1 _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2179__CLK clknet_leaf_11_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1663__A2 _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1888__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1415__A2 _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_45_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1040_ _0589_ _0603_ _0583_ _0581_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__1654__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1942_ _0874_ _0876_ _0535_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1873_ cal_lut\[3\] _0497_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1590__A1 _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1342__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1893__A2 _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1307_ _0871_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1238_ cal_lut\[138\] _0600_ _0652_ cal_lut\[102\] _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__1645__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1169_ cal_lut\[94\] _0617_ _0618_ cal_lut\[10\] _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xseg1._40_ dec1.o_dec\[1\] dec1.o_dec\[0\] seg1._13_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1333__A1 ctr\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1884__A2 _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1097__B1 _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1636__A2 _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1572__A1 _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2141_ _0159_ clknet_leaf_7_clk cal_lut\[82\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1875__A2 _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2072_ _0090_ clknet_leaf_18_clk cal_lut\[173\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1088__B1 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1023_ _0594_ _0590_ _0583_ _0581_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_72_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1627__A2 _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._7__I temp1.dac.i_enable vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1925_ cal_lut\[28\] _0506_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_16_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1856_ _0956_ _0486_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1260__B1 _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1787_ _0449_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__1315__A1 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input13_I i_wb_addr[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1251__B1 _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1149__A4 _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1554__A1 _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1710_ cal_lut\[135\] _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_108_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1641_ _0233_ _0345_ _0358_ _0348_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_13_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1793__A1 _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1572_ _0274_ _0283_ _0315_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_67_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I i_wb_addr[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2124_ _0142_ clknet_leaf_15_clk cal_lut\[65\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1848__A2 _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2055_ _0073_ clknet_leaf_9_clk ctr\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtemp1.dac.parallel_cells\[2\].vdac_batch._6_ temp1.dac.parallel_cells\[2\].vdac_batch._2_
+ temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1006_ _0579_ temp1.i_precharge_n vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_131_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1908_ _0251_ _0496_ _0518_ _0508_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1839_ cal_lut\[89\] _0461_ _0976_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1784__A1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1839__A2 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_142_Right_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_79_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1896__C _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1417__B _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref_I temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1152__B _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1058__A3 _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtemp1.dac.vdac_single._6_ temp1.dac.vdac_single._2_ temp1.dac.vdac_single.en_pupd
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1624_ _0967_ _0345_ _0349_ _0348_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1518__A1 _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1555_ cal_lut\[118\] _0292_ _0298_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1486_ _0976_ _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_136_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2062__CLK clknet_leaf_14_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_19_clk clknet_1_0__leaf_clk clknet_leaf_19_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2107_ _0125_ clknet_leaf_1_clk cal_lut\[144\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2038_ _0056_ clknet_leaf_12_clk cal_lut\[121\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1049__A3 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_107_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_99_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_116_Left_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xdec1._062_ dec1.i_bin\[3\] dec1._012_ dec1._013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_125_Left_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1340_ _0900_ clknet_1_1__leaf__0902_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2085__CLK clknet_leaf_16_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1920__A1 _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1271_ _0833_ _0836_ _0837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_134_Left_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_133_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_80_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_143_Left_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0986_ ctr\[4\] _0566_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_89_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_8_clk clknet_1_1__leaf_clk clknet_leaf_8_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1607_ _0965_ _0334_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1538_ _0976_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1469_ _0253_ _0961_ _0254_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_80_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1902__A1 _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1969__A1 ctr\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1323_ temp1.dac.i_data\[2\] _0870_ _0872_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1254_ _0818_ _0819_ _0820_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1121__A2 _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1185_ cal_lut\[142\] _0650_ _0592_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2100__CLK clknet_leaf_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1188__A2 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XANTENNA_input43_I i_wb_data[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1515__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtemp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
+ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_ temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__invz_3
XFILLER_0_37_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1425__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2123__CLK clknet_leaf_5_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1103__A2 _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1941_ o_wb_data[1] _0533_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1872_ _0967_ _0496_ _0499_ _0430_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_50_7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1342__A2 _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1306_ _0833_ _0836_ _0871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1237_ cal_lut\[54\] _0631_ _0623_ cal_lut\[48\] _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1168_ _0731_ _0732_ _0733_ _0736_ _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_35_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1099_ _0593_ cal_lut\[128\] _0612_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_19_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1030__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2146__CLK clknet_leaf_10_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1572__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ _0158_ clknet_leaf_11_clk cal_lut\[81\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2071_ _0089_ clknet_leaf_18_clk cal_lut\[172\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1022_ _0589_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_8
XTAP_TAPCELL_ROW_29_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2019__CLK clknet_leaf_18_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1924_ _0268_ _0497_ _0526_ _0508_ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_112_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1855_ net28 net27 _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1786_ net26 _0941_ _0280_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__2169__CLK clknet_leaf_1_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1563__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1003__A1 ctr\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1554__A2 _0283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1640_ cal_lut\[170\] _0356_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1793__A2 _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1571_ cal_lut\[126\] _0281_ _0298_ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1545__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_148_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2123_ _0141_ clknet_leaf_5_clk cal_lut\[160\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_108_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2054_ _0072_ clknet_leaf_8_clk ctr\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtemp1.dac.parallel_cells\[2\].vdac_batch._5_ temp1.dac.i_enable temp1.dac.parallel_cells\[2\].vdac_batch._1_
+ temp1.dac.parallel_cells\[2\].vdac_batch._2_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1005_ _0577_ _0578_ _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_29_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1481__A1 _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1907_ cal_lut\[19\] _0506_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1838_ _0261_ _0451_ _0477_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1784__A2 _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1536__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1769_ cal_lut\[154\] _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1523__B _0266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1472__A1 _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1224__A1 _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_105_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1463__A1 _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtemp1.dac.vdac_single._5_ temp1.dac._0_ temp1.dac.vdac_single._1_ temp1.dac.vdac_single._2_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_41_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1623_ cal_lut\[162\] _0346_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1518__A2 _0282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1554_ _0255_ _0283_ _0306_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1485_ net51 _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__2207__CLK clknet_leaf_6_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
.ends

