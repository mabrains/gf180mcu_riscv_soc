magic
tech gf180mcuD
magscale 1 5
timestamp 1702289190
<< obsm1 >>
rect 672 754 14360 59401
<< metal2 >>
rect 672 59800 728 60000
rect 1568 59800 1624 60000
rect 2464 59800 2520 60000
rect 3360 59800 3416 60000
rect 4256 59800 4312 60000
rect 5152 59800 5208 60000
rect 6048 59800 6104 60000
rect 6944 59800 7000 60000
rect 7840 59800 7896 60000
rect 8736 59800 8792 60000
rect 9632 59800 9688 60000
rect 10528 59800 10584 60000
rect 11424 59800 11480 60000
rect 12320 59800 12376 60000
rect 13216 59800 13272 60000
rect 14112 59800 14168 60000
rect 1344 0 1400 200
rect 1680 0 1736 200
rect 2016 0 2072 200
rect 2352 0 2408 200
rect 2688 0 2744 200
rect 3024 0 3080 200
rect 3360 0 3416 200
rect 3696 0 3752 200
rect 4032 0 4088 200
rect 4368 0 4424 200
rect 4704 0 4760 200
rect 5040 0 5096 200
rect 5376 0 5432 200
rect 5712 0 5768 200
rect 6048 0 6104 200
rect 6384 0 6440 200
rect 6720 0 6776 200
rect 7056 0 7112 200
rect 7392 0 7448 200
rect 7728 0 7784 200
rect 8064 0 8120 200
rect 8400 0 8456 200
rect 8736 0 8792 200
rect 9072 0 9128 200
rect 9408 0 9464 200
rect 9744 0 9800 200
rect 10080 0 10136 200
rect 10416 0 10472 200
rect 10752 0 10808 200
rect 11088 0 11144 200
rect 11424 0 11480 200
rect 11760 0 11816 200
rect 12096 0 12152 200
rect 12432 0 12488 200
rect 12768 0 12824 200
rect 13104 0 13160 200
rect 13440 0 13496 200
<< obsm2 >>
rect 758 59770 1538 59850
rect 1654 59770 2434 59850
rect 2550 59770 3330 59850
rect 3446 59770 4226 59850
rect 4342 59770 5122 59850
rect 5238 59770 6018 59850
rect 6134 59770 6914 59850
rect 7030 59770 7810 59850
rect 7926 59770 8706 59850
rect 8822 59770 9602 59850
rect 9718 59770 10498 59850
rect 10614 59770 11394 59850
rect 11510 59770 12290 59850
rect 12406 59770 13186 59850
rect 13302 59770 14082 59850
rect 14198 59770 14346 59850
rect 686 230 14346 59770
rect 686 200 1314 230
rect 1430 200 1650 230
rect 1766 200 1986 230
rect 2102 200 2322 230
rect 2438 200 2658 230
rect 2774 200 2994 230
rect 3110 200 3330 230
rect 3446 200 3666 230
rect 3782 200 4002 230
rect 4118 200 4338 230
rect 4454 200 4674 230
rect 4790 200 5010 230
rect 5126 200 5346 230
rect 5462 200 5682 230
rect 5798 200 6018 230
rect 6134 200 6354 230
rect 6470 200 6690 230
rect 6806 200 7026 230
rect 7142 200 7362 230
rect 7478 200 7698 230
rect 7814 200 8034 230
rect 8150 200 8370 230
rect 8486 200 8706 230
rect 8822 200 9042 230
rect 9158 200 9378 230
rect 9494 200 9714 230
rect 9830 200 10050 230
rect 10166 200 10386 230
rect 10502 200 10722 230
rect 10838 200 11058 230
rect 11174 200 11394 230
rect 11510 200 11730 230
rect 11846 200 12066 230
rect 12182 200 12402 230
rect 12518 200 12738 230
rect 12854 200 13074 230
rect 13190 200 13410 230
rect 13526 200 14346 230
<< metal3 >>
rect 0 57456 200 57512
rect 0 56112 200 56168
rect 0 54768 200 54824
rect 0 53424 200 53480
rect 0 52080 200 52136
rect 0 50736 200 50792
rect 0 49392 200 49448
rect 0 48048 200 48104
rect 0 46704 200 46760
rect 0 45360 200 45416
rect 0 44016 200 44072
rect 0 42672 200 42728
rect 0 41328 200 41384
rect 0 39984 200 40040
rect 0 38640 200 38696
rect 0 37296 200 37352
rect 0 35952 200 36008
rect 0 34608 200 34664
rect 0 33264 200 33320
rect 0 31920 200 31976
rect 0 30576 200 30632
rect 0 29232 200 29288
rect 0 27888 200 27944
rect 0 26544 200 26600
rect 0 25200 200 25256
rect 0 23856 200 23912
rect 0 22512 200 22568
rect 0 21168 200 21224
rect 0 19824 200 19880
rect 0 18480 200 18536
rect 0 17136 200 17192
rect 0 15792 200 15848
rect 0 14448 200 14504
rect 0 13104 200 13160
rect 0 11760 200 11816
rect 0 10416 200 10472
rect 0 9072 200 9128
rect 0 7728 200 7784
rect 0 6384 200 6440
rect 0 5040 200 5096
rect 0 3696 200 3752
rect 0 2352 200 2408
<< obsm3 >>
rect 200 57542 14351 59206
rect 230 57426 14351 57542
rect 200 56198 14351 57426
rect 230 56082 14351 56198
rect 200 54854 14351 56082
rect 230 54738 14351 54854
rect 200 53510 14351 54738
rect 230 53394 14351 53510
rect 200 52166 14351 53394
rect 230 52050 14351 52166
rect 200 50822 14351 52050
rect 230 50706 14351 50822
rect 200 49478 14351 50706
rect 230 49362 14351 49478
rect 200 48134 14351 49362
rect 230 48018 14351 48134
rect 200 46790 14351 48018
rect 230 46674 14351 46790
rect 200 45446 14351 46674
rect 230 45330 14351 45446
rect 200 44102 14351 45330
rect 230 43986 14351 44102
rect 200 42758 14351 43986
rect 230 42642 14351 42758
rect 200 41414 14351 42642
rect 230 41298 14351 41414
rect 200 40070 14351 41298
rect 230 39954 14351 40070
rect 200 38726 14351 39954
rect 230 38610 14351 38726
rect 200 37382 14351 38610
rect 230 37266 14351 37382
rect 200 36038 14351 37266
rect 230 35922 14351 36038
rect 200 34694 14351 35922
rect 230 34578 14351 34694
rect 200 33350 14351 34578
rect 230 33234 14351 33350
rect 200 32006 14351 33234
rect 230 31890 14351 32006
rect 200 30662 14351 31890
rect 230 30546 14351 30662
rect 200 29318 14351 30546
rect 230 29202 14351 29318
rect 200 27974 14351 29202
rect 230 27858 14351 27974
rect 200 26630 14351 27858
rect 230 26514 14351 26630
rect 200 25286 14351 26514
rect 230 25170 14351 25286
rect 200 23942 14351 25170
rect 230 23826 14351 23942
rect 200 22598 14351 23826
rect 230 22482 14351 22598
rect 200 21254 14351 22482
rect 230 21138 14351 21254
rect 200 19910 14351 21138
rect 230 19794 14351 19910
rect 200 18566 14351 19794
rect 230 18450 14351 18566
rect 200 17222 14351 18450
rect 230 17106 14351 17222
rect 200 15878 14351 17106
rect 230 15762 14351 15878
rect 200 14534 14351 15762
rect 230 14418 14351 14534
rect 200 13190 14351 14418
rect 230 13074 14351 13190
rect 200 11846 14351 13074
rect 230 11730 14351 11846
rect 200 10502 14351 11730
rect 230 10386 14351 10502
rect 200 9158 14351 10386
rect 230 9042 14351 9158
rect 200 7814 14351 9042
rect 230 7698 14351 7814
rect 200 6470 14351 7698
rect 230 6354 14351 6470
rect 200 5126 14351 6354
rect 230 5010 14351 5126
rect 200 3782 14351 5010
rect 230 3666 14351 3782
rect 200 2438 14351 3666
rect 230 2322 14351 2438
rect 200 238 14351 2322
<< metal4 >>
rect 2293 754 2453 59222
rect 3994 754 4154 59222
rect 5695 754 5855 59222
rect 7396 754 7556 59222
rect 9097 754 9257 59222
rect 10798 754 10958 59222
rect 12499 754 12659 59222
rect 14200 754 14360 59222
<< obsm4 >>
rect 1190 1073 2263 52855
rect 2483 1073 3964 52855
rect 4184 1073 5665 52855
rect 5885 1073 7366 52855
rect 7586 1073 9067 52855
rect 9287 1073 10768 52855
rect 10988 1073 12469 52855
rect 12689 1073 14042 52855
<< labels >>
rlabel metal2 s 1680 0 1736 200 6 clk
port 1 nsew signal input
rlabel metal2 s 12432 0 12488 200 6 i_wb_addr[0]
port 2 nsew signal input
rlabel metal2 s 9072 0 9128 200 6 i_wb_addr[10]
port 3 nsew signal input
rlabel metal2 s 8736 0 8792 200 6 i_wb_addr[11]
port 4 nsew signal input
rlabel metal2 s 8400 0 8456 200 6 i_wb_addr[12]
port 5 nsew signal input
rlabel metal2 s 8064 0 8120 200 6 i_wb_addr[13]
port 6 nsew signal input
rlabel metal2 s 7728 0 7784 200 6 i_wb_addr[14]
port 7 nsew signal input
rlabel metal2 s 7392 0 7448 200 6 i_wb_addr[15]
port 8 nsew signal input
rlabel metal2 s 7056 0 7112 200 6 i_wb_addr[16]
port 9 nsew signal input
rlabel metal2 s 6720 0 6776 200 6 i_wb_addr[17]
port 10 nsew signal input
rlabel metal2 s 6384 0 6440 200 6 i_wb_addr[18]
port 11 nsew signal input
rlabel metal2 s 6048 0 6104 200 6 i_wb_addr[19]
port 12 nsew signal input
rlabel metal2 s 12096 0 12152 200 6 i_wb_addr[1]
port 13 nsew signal input
rlabel metal2 s 5712 0 5768 200 6 i_wb_addr[20]
port 14 nsew signal input
rlabel metal2 s 5376 0 5432 200 6 i_wb_addr[21]
port 15 nsew signal input
rlabel metal2 s 5040 0 5096 200 6 i_wb_addr[22]
port 16 nsew signal input
rlabel metal2 s 4704 0 4760 200 6 i_wb_addr[23]
port 17 nsew signal input
rlabel metal2 s 4368 0 4424 200 6 i_wb_addr[24]
port 18 nsew signal input
rlabel metal2 s 4032 0 4088 200 6 i_wb_addr[25]
port 19 nsew signal input
rlabel metal2 s 3696 0 3752 200 6 i_wb_addr[26]
port 20 nsew signal input
rlabel metal2 s 3360 0 3416 200 6 i_wb_addr[27]
port 21 nsew signal input
rlabel metal2 s 3024 0 3080 200 6 i_wb_addr[28]
port 22 nsew signal input
rlabel metal2 s 2688 0 2744 200 6 i_wb_addr[29]
port 23 nsew signal input
rlabel metal2 s 11760 0 11816 200 6 i_wb_addr[2]
port 24 nsew signal input
rlabel metal2 s 2352 0 2408 200 6 i_wb_addr[30]
port 25 nsew signal input
rlabel metal2 s 2016 0 2072 200 6 i_wb_addr[31]
port 26 nsew signal input
rlabel metal2 s 11424 0 11480 200 6 i_wb_addr[3]
port 27 nsew signal input
rlabel metal2 s 11088 0 11144 200 6 i_wb_addr[4]
port 28 nsew signal input
rlabel metal2 s 10752 0 10808 200 6 i_wb_addr[5]
port 29 nsew signal input
rlabel metal2 s 10416 0 10472 200 6 i_wb_addr[6]
port 30 nsew signal input
rlabel metal2 s 10080 0 10136 200 6 i_wb_addr[7]
port 31 nsew signal input
rlabel metal2 s 9744 0 9800 200 6 i_wb_addr[8]
port 32 nsew signal input
rlabel metal2 s 9408 0 9464 200 6 i_wb_addr[9]
port 33 nsew signal input
rlabel metal2 s 13440 0 13496 200 6 i_wb_cyc
port 34 nsew signal input
rlabel metal3 s 0 2352 200 2408 6 i_wb_data[0]
port 35 nsew signal input
rlabel metal3 s 0 15792 200 15848 6 i_wb_data[10]
port 36 nsew signal input
rlabel metal3 s 0 17136 200 17192 6 i_wb_data[11]
port 37 nsew signal input
rlabel metal3 s 0 18480 200 18536 6 i_wb_data[12]
port 38 nsew signal input
rlabel metal3 s 0 19824 200 19880 6 i_wb_data[13]
port 39 nsew signal input
rlabel metal3 s 0 21168 200 21224 6 i_wb_data[14]
port 40 nsew signal input
rlabel metal3 s 0 22512 200 22568 6 i_wb_data[15]
port 41 nsew signal input
rlabel metal3 s 0 23856 200 23912 6 i_wb_data[16]
port 42 nsew signal input
rlabel metal3 s 0 25200 200 25256 6 i_wb_data[17]
port 43 nsew signal input
rlabel metal3 s 0 26544 200 26600 6 i_wb_data[18]
port 44 nsew signal input
rlabel metal3 s 0 27888 200 27944 6 i_wb_data[19]
port 45 nsew signal input
rlabel metal3 s 0 3696 200 3752 6 i_wb_data[1]
port 46 nsew signal input
rlabel metal3 s 0 29232 200 29288 6 i_wb_data[20]
port 47 nsew signal input
rlabel metal3 s 0 30576 200 30632 6 i_wb_data[21]
port 48 nsew signal input
rlabel metal3 s 0 31920 200 31976 6 i_wb_data[22]
port 49 nsew signal input
rlabel metal3 s 0 33264 200 33320 6 i_wb_data[23]
port 50 nsew signal input
rlabel metal3 s 0 34608 200 34664 6 i_wb_data[24]
port 51 nsew signal input
rlabel metal3 s 0 35952 200 36008 6 i_wb_data[25]
port 52 nsew signal input
rlabel metal3 s 0 37296 200 37352 6 i_wb_data[26]
port 53 nsew signal input
rlabel metal3 s 0 38640 200 38696 6 i_wb_data[27]
port 54 nsew signal input
rlabel metal3 s 0 39984 200 40040 6 i_wb_data[28]
port 55 nsew signal input
rlabel metal3 s 0 41328 200 41384 6 i_wb_data[29]
port 56 nsew signal input
rlabel metal3 s 0 5040 200 5096 6 i_wb_data[2]
port 57 nsew signal input
rlabel metal3 s 0 42672 200 42728 6 i_wb_data[30]
port 58 nsew signal input
rlabel metal3 s 0 44016 200 44072 6 i_wb_data[31]
port 59 nsew signal input
rlabel metal3 s 0 6384 200 6440 6 i_wb_data[3]
port 60 nsew signal input
rlabel metal3 s 0 7728 200 7784 6 i_wb_data[4]
port 61 nsew signal input
rlabel metal3 s 0 9072 200 9128 6 i_wb_data[5]
port 62 nsew signal input
rlabel metal3 s 0 10416 200 10472 6 i_wb_data[6]
port 63 nsew signal input
rlabel metal3 s 0 11760 200 11816 6 i_wb_data[7]
port 64 nsew signal input
rlabel metal3 s 0 13104 200 13160 6 i_wb_data[8]
port 65 nsew signal input
rlabel metal3 s 0 14448 200 14504 6 i_wb_data[9]
port 66 nsew signal input
rlabel metal2 s 13104 0 13160 200 6 i_wb_stb
port 67 nsew signal input
rlabel metal2 s 12768 0 12824 200 6 i_wb_we
port 68 nsew signal input
rlabel metal2 s 6944 59800 7000 60000 6 io_oeb[0]
port 69 nsew signal output
rlabel metal2 s 6048 59800 6104 60000 6 io_oeb[1]
port 70 nsew signal output
rlabel metal2 s 5152 59800 5208 60000 6 io_oeb[2]
port 71 nsew signal output
rlabel metal2 s 4256 59800 4312 60000 6 io_oeb[3]
port 72 nsew signal output
rlabel metal2 s 3360 59800 3416 60000 6 io_oeb[4]
port 73 nsew signal output
rlabel metal2 s 2464 59800 2520 60000 6 io_oeb[5]
port 74 nsew signal output
rlabel metal2 s 1568 59800 1624 60000 6 io_oeb[6]
port 75 nsew signal output
rlabel metal2 s 672 59800 728 60000 6 io_oeb[7]
port 76 nsew signal output
rlabel metal2 s 14112 59800 14168 60000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 13216 59800 13272 60000 6 io_out[1]
port 78 nsew signal output
rlabel metal2 s 12320 59800 12376 60000 6 io_out[2]
port 79 nsew signal output
rlabel metal2 s 11424 59800 11480 60000 6 io_out[3]
port 80 nsew signal output
rlabel metal2 s 10528 59800 10584 60000 6 io_out[4]
port 81 nsew signal output
rlabel metal2 s 9632 59800 9688 60000 6 io_out[5]
port 82 nsew signal output
rlabel metal2 s 8736 59800 8792 60000 6 io_out[6]
port 83 nsew signal output
rlabel metal2 s 7840 59800 7896 60000 6 io_out[7]
port 84 nsew signal output
rlabel metal3 s 0 45360 200 45416 6 o_wb_ack
port 85 nsew signal output
rlabel metal3 s 0 46704 200 46760 6 o_wb_data[0]
port 86 nsew signal output
rlabel metal3 s 0 48048 200 48104 6 o_wb_data[1]
port 87 nsew signal output
rlabel metal3 s 0 49392 200 49448 6 o_wb_data[2]
port 88 nsew signal output
rlabel metal3 s 0 50736 200 50792 6 o_wb_data[3]
port 89 nsew signal output
rlabel metal3 s 0 52080 200 52136 6 o_wb_data[4]
port 90 nsew signal output
rlabel metal3 s 0 53424 200 53480 6 o_wb_data[5]
port 91 nsew signal output
rlabel metal3 s 0 54768 200 54824 6 o_wb_data[6]
port 92 nsew signal output
rlabel metal3 s 0 56112 200 56168 6 o_wb_data[7]
port 93 nsew signal output
rlabel metal3 s 0 57456 200 57512 6 o_wb_stall
port 94 nsew signal output
rlabel metal2 s 1344 0 1400 200 6 reset
port 95 nsew signal input
rlabel metal4 s 2293 754 2453 59222 6 vdd
port 96 nsew power bidirectional
rlabel metal4 s 5695 754 5855 59222 6 vdd
port 96 nsew power bidirectional
rlabel metal4 s 9097 754 9257 59222 6 vdd
port 96 nsew power bidirectional
rlabel metal4 s 12499 754 12659 59222 6 vdd
port 96 nsew power bidirectional
rlabel metal4 s 3994 754 4154 59222 6 vss
port 97 nsew ground bidirectional
rlabel metal4 s 7396 754 7556 59222 6 vss
port 97 nsew ground bidirectional
rlabel metal4 s 10798 754 10958 59222 6 vss
port 97 nsew ground bidirectional
rlabel metal4 s 14200 754 14360 59222 6 vss
port 97 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 15000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4219490
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/temp_sensor/runs/23_12_11_12_00/results/signoff/temp_sensor.magic.gds
string GDS_START 425314
<< end >>

