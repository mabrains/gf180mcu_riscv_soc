VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO temp_sensor
  CLASS BLOCK ;
  FOREIGN temp_sensor ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 400.000 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 7.540 23.840 392.300 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 7.540 177.440 392.300 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 7.540 100.640 392.300 ;
    END
  END VSS
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 14.560 2.000 15.120 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.200 2.000 39.760 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 63.840 2.000 64.400 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 88.480 2.000 89.040 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 113.120 2.000 113.680 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 2.000 138.320 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 162.400 2.000 162.960 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.040 2.000 187.600 ;
    END
  END io_in[7]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.680 2.000 212.240 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.304800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 236.320 2.000 236.880 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 260.960 2.000 261.520 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 285.600 2.000 286.160 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.276000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.240 2.000 310.800 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.304800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.880 2.000 335.440 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.182800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 359.520 2.000 360.080 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.145600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 384.160 2.000 384.720 ;
    END
  END io_out[7]
  OBS
      LAYER Metal1 ;
        RECT 6.720 7.540 243.040 392.300 ;
      LAYER Metal2 ;
        RECT 7.980 7.650 240.660 392.190 ;
      LAYER Metal3 ;
        RECT 1.260 385.020 240.710 392.140 ;
        RECT 2.300 383.860 240.710 385.020 ;
        RECT 1.260 360.380 240.710 383.860 ;
        RECT 2.300 359.220 240.710 360.380 ;
        RECT 1.260 335.740 240.710 359.220 ;
        RECT 2.300 334.580 240.710 335.740 ;
        RECT 1.260 311.100 240.710 334.580 ;
        RECT 2.300 309.940 240.710 311.100 ;
        RECT 1.260 286.460 240.710 309.940 ;
        RECT 2.300 285.300 240.710 286.460 ;
        RECT 1.260 261.820 240.710 285.300 ;
        RECT 2.300 260.660 240.710 261.820 ;
        RECT 1.260 237.180 240.710 260.660 ;
        RECT 2.300 236.020 240.710 237.180 ;
        RECT 1.260 212.540 240.710 236.020 ;
        RECT 2.300 211.380 240.710 212.540 ;
        RECT 1.260 187.900 240.710 211.380 ;
        RECT 2.300 186.740 240.710 187.900 ;
        RECT 1.260 163.260 240.710 186.740 ;
        RECT 2.300 162.100 240.710 163.260 ;
        RECT 1.260 138.620 240.710 162.100 ;
        RECT 2.300 137.460 240.710 138.620 ;
        RECT 1.260 113.980 240.710 137.460 ;
        RECT 2.300 112.820 240.710 113.980 ;
        RECT 1.260 89.340 240.710 112.820 ;
        RECT 2.300 88.180 240.710 89.340 ;
        RECT 1.260 64.700 240.710 88.180 ;
        RECT 2.300 63.540 240.710 64.700 ;
        RECT 1.260 40.060 240.710 63.540 ;
        RECT 2.300 38.900 240.710 40.060 ;
        RECT 1.260 15.420 240.710 38.900 ;
        RECT 2.300 14.260 240.710 15.420 ;
        RECT 1.260 7.700 240.710 14.260 ;
      LAYER Metal4 ;
        RECT 11.340 18.570 21.940 338.150 ;
        RECT 24.140 18.570 98.740 338.150 ;
        RECT 100.940 18.570 175.540 338.150 ;
        RECT 177.740 18.570 199.780 338.150 ;
  END
END temp_sensor
END LIBRARY

