magic
tech gf180mcuD
magscale 1 10
timestamp 1700411247
<< metal1 >>
rect 1344 78426 48608 78460
rect 1344 78374 19838 78426
rect 19890 78374 19942 78426
rect 19994 78374 20046 78426
rect 20098 78374 48608 78426
rect 1344 78340 48608 78374
rect 1810 77982 1822 78034
rect 1874 77982 1886 78034
rect 3154 77982 3166 78034
rect 3218 77982 3230 78034
rect 2942 77922 2994 77934
rect 2942 77858 2994 77870
rect 1344 77642 48608 77676
rect 1344 77590 4478 77642
rect 4530 77590 4582 77642
rect 4634 77590 4686 77642
rect 4738 77590 35198 77642
rect 35250 77590 35302 77642
rect 35354 77590 35406 77642
rect 35458 77590 48608 77642
rect 1344 77556 48608 77590
rect 2942 77362 2994 77374
rect 33282 77310 33294 77362
rect 33346 77310 33358 77362
rect 2942 77298 2994 77310
rect 9886 77250 9938 77262
rect 1810 77198 1822 77250
rect 1874 77198 1886 77250
rect 3154 77198 3166 77250
rect 3218 77198 3230 77250
rect 8866 77198 8878 77250
rect 8930 77198 8942 77250
rect 30482 77198 30494 77250
rect 30546 77198 30558 77250
rect 9886 77186 9938 77198
rect 27806 77138 27858 77150
rect 31154 77086 31166 77138
rect 31218 77086 31230 77138
rect 27806 77074 27858 77086
rect 6190 77026 6242 77038
rect 6190 76962 6242 76974
rect 6638 77026 6690 77038
rect 6638 76962 6690 76974
rect 7310 77026 7362 77038
rect 7310 76962 7362 76974
rect 7534 77026 7586 77038
rect 7534 76962 7586 76974
rect 21534 77026 21586 77038
rect 21534 76962 21586 76974
rect 28142 77026 28194 77038
rect 28142 76962 28194 76974
rect 33742 77026 33794 77038
rect 33742 76962 33794 76974
rect 1344 76858 48608 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 48608 76858
rect 1344 76772 48608 76806
rect 3054 76690 3106 76702
rect 3054 76626 3106 76638
rect 3614 76690 3666 76702
rect 3614 76626 3666 76638
rect 10110 76690 10162 76702
rect 10110 76626 10162 76638
rect 30942 76690 30994 76702
rect 30942 76626 30994 76638
rect 33518 76578 33570 76590
rect 27906 76526 27918 76578
rect 27970 76526 27982 76578
rect 33518 76514 33570 76526
rect 5966 76466 6018 76478
rect 10446 76466 10498 76478
rect 13022 76466 13074 76478
rect 30606 76466 30658 76478
rect 1810 76414 1822 76466
rect 1874 76414 1886 76466
rect 3266 76414 3278 76466
rect 3330 76414 3342 76466
rect 4946 76414 4958 76466
rect 5010 76414 5022 76466
rect 6290 76414 6302 76466
rect 6354 76414 6366 76466
rect 7074 76414 7086 76466
rect 7138 76414 7150 76466
rect 11218 76414 11230 76466
rect 11282 76414 11294 76466
rect 13794 76414 13806 76466
rect 13858 76414 13870 76466
rect 18498 76414 18510 76466
rect 18562 76414 18574 76466
rect 21746 76414 21758 76466
rect 21810 76414 21822 76466
rect 27122 76414 27134 76466
rect 27186 76414 27198 76466
rect 33954 76414 33966 76466
rect 34018 76414 34030 76466
rect 5966 76402 6018 76414
rect 10446 76402 10498 76414
rect 13022 76402 13074 76414
rect 30606 76402 30658 76414
rect 8206 76354 8258 76366
rect 8206 76290 8258 76302
rect 18174 76354 18226 76366
rect 26798 76354 26850 76366
rect 33182 76354 33234 76366
rect 19282 76302 19294 76354
rect 19346 76302 19358 76354
rect 21410 76302 21422 76354
rect 21474 76302 21486 76354
rect 22530 76302 22542 76354
rect 22594 76302 22606 76354
rect 24658 76302 24670 76354
rect 24722 76302 24734 76354
rect 30034 76302 30046 76354
rect 30098 76302 30110 76354
rect 34738 76302 34750 76354
rect 34802 76302 34814 76354
rect 36866 76302 36878 76354
rect 36930 76302 36942 76354
rect 18174 76290 18226 76302
rect 26798 76290 26850 76302
rect 33182 76290 33234 76302
rect 12574 76242 12626 76254
rect 12574 76178 12626 76190
rect 15150 76242 15202 76254
rect 15150 76178 15202 76190
rect 33630 76242 33682 76254
rect 33630 76178 33682 76190
rect 1344 76074 48608 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 48608 76074
rect 1344 75988 48608 76022
rect 8318 75906 8370 75918
rect 8318 75842 8370 75854
rect 12014 75906 12066 75918
rect 12014 75842 12066 75854
rect 21310 75906 21362 75918
rect 21310 75842 21362 75854
rect 27806 75906 27858 75918
rect 27806 75842 27858 75854
rect 30494 75906 30546 75918
rect 30494 75842 30546 75854
rect 4286 75794 4338 75806
rect 4286 75730 4338 75742
rect 12686 75794 12738 75806
rect 12686 75730 12738 75742
rect 22878 75794 22930 75806
rect 22878 75730 22930 75742
rect 23550 75794 23602 75806
rect 23550 75730 23602 75742
rect 24110 75794 24162 75806
rect 28142 75794 28194 75806
rect 27458 75742 27470 75794
rect 27522 75742 27534 75794
rect 24110 75730 24162 75742
rect 28142 75730 28194 75742
rect 30158 75794 30210 75806
rect 30158 75730 30210 75742
rect 30942 75794 30994 75806
rect 36430 75794 36482 75806
rect 34178 75742 34190 75794
rect 34242 75742 34254 75794
rect 34738 75742 34750 75794
rect 34802 75742 34814 75794
rect 30942 75730 30994 75742
rect 36430 75730 36482 75742
rect 6190 75682 6242 75694
rect 9886 75682 9938 75694
rect 20750 75682 20802 75694
rect 3042 75630 3054 75682
rect 3106 75630 3118 75682
rect 6962 75630 6974 75682
rect 7026 75630 7038 75682
rect 10882 75630 10894 75682
rect 10946 75630 10958 75682
rect 6190 75618 6242 75630
rect 9886 75618 9938 75630
rect 20750 75618 20802 75630
rect 21646 75682 21698 75694
rect 21646 75618 21698 75630
rect 22430 75682 22482 75694
rect 22430 75618 22482 75630
rect 22766 75682 22818 75694
rect 23438 75682 23490 75694
rect 23090 75630 23102 75682
rect 23154 75630 23166 75682
rect 22766 75618 22818 75630
rect 23438 75618 23490 75630
rect 24222 75682 24274 75694
rect 29262 75682 29314 75694
rect 24546 75630 24558 75682
rect 24610 75630 24622 75682
rect 24222 75618 24274 75630
rect 29262 75618 29314 75630
rect 29934 75682 29986 75694
rect 35310 75682 35362 75694
rect 31266 75630 31278 75682
rect 31330 75630 31342 75682
rect 32050 75630 32062 75682
rect 32114 75630 32126 75682
rect 29934 75618 29986 75630
rect 35310 75618 35362 75630
rect 4398 75570 4450 75582
rect 28366 75570 28418 75582
rect 25330 75518 25342 75570
rect 25394 75518 25406 75570
rect 4398 75506 4450 75518
rect 28366 75506 28418 75518
rect 34526 75570 34578 75582
rect 34526 75506 34578 75518
rect 34750 75570 34802 75582
rect 34750 75506 34802 75518
rect 5854 75458 5906 75470
rect 5854 75394 5906 75406
rect 9550 75458 9602 75470
rect 9550 75394 9602 75406
rect 21422 75458 21474 75470
rect 21422 75394 21474 75406
rect 36318 75458 36370 75470
rect 36318 75394 36370 75406
rect 1344 75290 48608 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 48608 75290
rect 1344 75204 48608 75238
rect 4286 75122 4338 75134
rect 4286 75058 4338 75070
rect 5742 75122 5794 75134
rect 5742 75058 5794 75070
rect 8430 75122 8482 75134
rect 8430 75058 8482 75070
rect 8990 75122 9042 75134
rect 8990 75058 9042 75070
rect 25566 75122 25618 75134
rect 25566 75058 25618 75070
rect 25342 75010 25394 75022
rect 25342 74946 25394 74958
rect 33630 75010 33682 75022
rect 33630 74946 33682 74958
rect 4398 74898 4450 74910
rect 3042 74846 3054 74898
rect 3106 74846 3118 74898
rect 4398 74834 4450 74846
rect 6078 74898 6130 74910
rect 25230 74898 25282 74910
rect 6962 74846 6974 74898
rect 7026 74846 7038 74898
rect 9650 74846 9662 74898
rect 9714 74846 9726 74898
rect 10546 74846 10558 74898
rect 10610 74846 10622 74898
rect 6078 74834 6130 74846
rect 25230 74834 25282 74846
rect 25902 74898 25954 74910
rect 34962 74846 34974 74898
rect 35026 74846 35038 74898
rect 25902 74834 25954 74846
rect 24222 74786 24274 74798
rect 24222 74722 24274 74734
rect 27582 74786 27634 74798
rect 27582 74722 27634 74734
rect 30942 74786 30994 74798
rect 30942 74722 30994 74734
rect 32510 74786 32562 74798
rect 32510 74722 32562 74734
rect 33406 74786 33458 74798
rect 34190 74786 34242 74798
rect 33730 74734 33742 74786
rect 33794 74734 33806 74786
rect 33406 74722 33458 74734
rect 34190 74722 34242 74734
rect 34638 74786 34690 74798
rect 35746 74734 35758 74786
rect 35810 74734 35822 74786
rect 37874 74734 37886 74786
rect 37938 74734 37950 74786
rect 34638 74722 34690 74734
rect 11678 74674 11730 74686
rect 33954 74622 33966 74674
rect 34018 74671 34030 74674
rect 34626 74671 34638 74674
rect 34018 74625 34638 74671
rect 34018 74622 34030 74625
rect 34626 74622 34638 74625
rect 34690 74622 34702 74674
rect 11678 74610 11730 74622
rect 1344 74506 48608 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 48608 74506
rect 1344 74420 48608 74454
rect 12798 74338 12850 74350
rect 12798 74274 12850 74286
rect 36990 74338 37042 74350
rect 36990 74274 37042 74286
rect 10334 74226 10386 74238
rect 21310 74226 21362 74238
rect 20738 74174 20750 74226
rect 20802 74174 20814 74226
rect 10334 74162 10386 74174
rect 21310 74162 21362 74174
rect 33518 74226 33570 74238
rect 37102 74226 37154 74238
rect 35746 74174 35758 74226
rect 35810 74174 35822 74226
rect 33518 74162 33570 74174
rect 37102 74162 37154 74174
rect 10670 74114 10722 74126
rect 11442 74062 11454 74114
rect 11506 74062 11518 74114
rect 17826 74062 17838 74114
rect 17890 74062 17902 74114
rect 35634 74062 35646 74114
rect 35698 74062 35710 74114
rect 10670 74050 10722 74062
rect 17502 74002 17554 74014
rect 21422 74002 21474 74014
rect 18610 73950 18622 74002
rect 18674 73950 18686 74002
rect 17502 73938 17554 73950
rect 21422 73938 21474 73950
rect 30270 74002 30322 74014
rect 30270 73938 30322 73950
rect 30382 74002 30434 74014
rect 30382 73938 30434 73950
rect 33406 74002 33458 74014
rect 33406 73938 33458 73950
rect 35310 74002 35362 74014
rect 35310 73938 35362 73950
rect 35982 74002 36034 74014
rect 35982 73938 36034 73950
rect 29934 73890 29986 73902
rect 29934 73826 29986 73838
rect 30606 73890 30658 73902
rect 30606 73826 30658 73838
rect 1344 73722 48608 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 48608 73722
rect 1344 73636 48608 73670
rect 19406 73554 19458 73566
rect 19406 73490 19458 73502
rect 31266 73390 31278 73442
rect 31330 73390 31342 73442
rect 9650 73278 9662 73330
rect 9714 73278 9726 73330
rect 10322 73278 10334 73330
rect 10386 73278 10398 73330
rect 12226 73278 12238 73330
rect 12290 73278 12302 73330
rect 13010 73278 13022 73330
rect 13074 73278 13086 73330
rect 19618 73278 19630 73330
rect 19682 73278 19694 73330
rect 25890 73278 25902 73330
rect 25954 73278 25966 73330
rect 31938 73278 31950 73330
rect 32002 73278 32014 73330
rect 8990 73218 9042 73230
rect 8990 73154 9042 73166
rect 18958 73218 19010 73230
rect 18958 73154 19010 73166
rect 25566 73218 25618 73230
rect 33182 73218 33234 73230
rect 26674 73166 26686 73218
rect 26738 73166 26750 73218
rect 28802 73166 28814 73218
rect 28866 73166 28878 73218
rect 29138 73166 29150 73218
rect 29202 73166 29214 73218
rect 25566 73154 25618 73166
rect 33182 73154 33234 73166
rect 33854 73218 33906 73230
rect 33854 73154 33906 73166
rect 11678 73106 11730 73118
rect 11678 73042 11730 73054
rect 14254 73106 14306 73118
rect 14254 73042 14306 73054
rect 19294 73106 19346 73118
rect 19294 73042 19346 73054
rect 33070 73106 33122 73118
rect 33070 73042 33122 73054
rect 1344 72938 48608 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 48608 72938
rect 1344 72852 48608 72886
rect 34850 72718 34862 72770
rect 34914 72767 34926 72770
rect 35186 72767 35198 72770
rect 34914 72721 35198 72767
rect 34914 72718 34926 72721
rect 35186 72718 35198 72721
rect 35250 72718 35262 72770
rect 5070 72658 5122 72670
rect 35198 72658 35250 72670
rect 33618 72606 33630 72658
rect 33682 72606 33694 72658
rect 5070 72594 5122 72606
rect 35198 72594 35250 72606
rect 30046 72546 30098 72558
rect 1810 72494 1822 72546
rect 1874 72494 1886 72546
rect 3154 72494 3166 72546
rect 3218 72494 3230 72546
rect 6066 72494 6078 72546
rect 6130 72494 6142 72546
rect 6962 72494 6974 72546
rect 7026 72494 7038 72546
rect 9202 72494 9214 72546
rect 9266 72494 9278 72546
rect 10098 72494 10110 72546
rect 10162 72494 10174 72546
rect 30046 72482 30098 72494
rect 30382 72546 30434 72558
rect 30818 72494 30830 72546
rect 30882 72494 30894 72546
rect 30382 72482 30434 72494
rect 31490 72382 31502 72434
rect 31554 72382 31566 72434
rect 2942 72322 2994 72334
rect 2942 72258 2994 72270
rect 8318 72322 8370 72334
rect 8318 72258 8370 72270
rect 8766 72322 8818 72334
rect 8766 72258 8818 72270
rect 11454 72322 11506 72334
rect 11454 72258 11506 72270
rect 11790 72322 11842 72334
rect 11790 72258 11842 72270
rect 23550 72322 23602 72334
rect 23550 72258 23602 72270
rect 29262 72322 29314 72334
rect 29262 72258 29314 72270
rect 29822 72322 29874 72334
rect 29822 72258 29874 72270
rect 30270 72322 30322 72334
rect 30270 72258 30322 72270
rect 34302 72322 34354 72334
rect 34302 72258 34354 72270
rect 34750 72322 34802 72334
rect 34750 72258 34802 72270
rect 37102 72322 37154 72334
rect 37102 72258 37154 72270
rect 37550 72322 37602 72334
rect 37550 72258 37602 72270
rect 1344 72154 48608 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 48608 72154
rect 1344 72068 48608 72102
rect 5070 71986 5122 71998
rect 5070 71922 5122 71934
rect 5518 71986 5570 71998
rect 5518 71922 5570 71934
rect 33182 71986 33234 71998
rect 33182 71922 33234 71934
rect 3838 71874 3890 71886
rect 3838 71810 3890 71822
rect 23998 71874 24050 71886
rect 23998 71810 24050 71822
rect 24110 71874 24162 71886
rect 24110 71810 24162 71822
rect 6302 71762 6354 71774
rect 20302 71762 20354 71774
rect 23774 71762 23826 71774
rect 34862 71762 34914 71774
rect 36542 71762 36594 71774
rect 2706 71710 2718 71762
rect 2770 71710 2782 71762
rect 4050 71710 4062 71762
rect 4114 71710 4126 71762
rect 7074 71710 7086 71762
rect 7138 71710 7150 71762
rect 9650 71710 9662 71762
rect 9714 71710 9726 71762
rect 10322 71710 10334 71762
rect 10386 71710 10398 71762
rect 20738 71710 20750 71762
rect 20802 71710 20814 71762
rect 33394 71710 33406 71762
rect 33458 71710 33470 71762
rect 35074 71710 35086 71762
rect 35138 71710 35150 71762
rect 36082 71710 36094 71762
rect 36146 71710 36158 71762
rect 37538 71710 37550 71762
rect 37602 71710 37614 71762
rect 6302 71698 6354 71710
rect 20302 71698 20354 71710
rect 23774 71698 23826 71710
rect 34862 71698 34914 71710
rect 36542 71698 36594 71710
rect 6078 71650 6130 71662
rect 6078 71586 6130 71598
rect 8654 71650 8706 71662
rect 8654 71586 8706 71598
rect 8990 71650 9042 71662
rect 24558 71650 24610 71662
rect 21410 71598 21422 71650
rect 21474 71598 21486 71650
rect 8990 71586 9042 71598
rect 23538 71571 23550 71623
rect 23602 71571 23614 71623
rect 24558 71586 24610 71598
rect 25566 71650 25618 71662
rect 25566 71586 25618 71598
rect 26126 71650 26178 71662
rect 26126 71586 26178 71598
rect 32510 71650 32562 71662
rect 32510 71586 32562 71598
rect 33070 71650 33122 71662
rect 33070 71586 33122 71598
rect 33854 71650 33906 71662
rect 33854 71586 33906 71598
rect 34302 71650 34354 71662
rect 34302 71586 34354 71598
rect 37998 71650 38050 71662
rect 37998 71586 38050 71598
rect 11678 71538 11730 71550
rect 11678 71474 11730 71486
rect 24446 71538 24498 71550
rect 24446 71474 24498 71486
rect 25678 71538 25730 71550
rect 37214 71538 37266 71550
rect 36194 71486 36206 71538
rect 36258 71486 36270 71538
rect 25678 71474 25730 71486
rect 37214 71474 37266 71486
rect 37550 71538 37602 71550
rect 37550 71474 37602 71486
rect 1344 71370 48608 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 48608 71370
rect 1344 71284 48608 71318
rect 21646 71202 21698 71214
rect 21646 71138 21698 71150
rect 26350 71202 26402 71214
rect 36082 71150 36094 71202
rect 36146 71150 36158 71202
rect 26350 71138 26402 71150
rect 3502 71090 3554 71102
rect 3502 71026 3554 71038
rect 10334 71090 10386 71102
rect 10334 71026 10386 71038
rect 20750 71090 20802 71102
rect 29486 71090 29538 71102
rect 21410 71038 21422 71090
rect 21474 71038 21486 71090
rect 23538 71038 23550 71090
rect 23602 71038 23614 71090
rect 25666 71038 25678 71090
rect 25730 71038 25742 71090
rect 26002 71038 26014 71090
rect 26066 71038 26078 71090
rect 32946 71038 32958 71090
rect 33010 71038 33022 71090
rect 33842 71038 33854 71090
rect 33906 71038 33918 71090
rect 34850 71038 34862 71090
rect 34914 71038 34926 71090
rect 37762 71038 37774 71090
rect 37826 71038 37838 71090
rect 39890 71038 39902 71090
rect 39954 71038 39966 71090
rect 20750 71026 20802 71038
rect 29486 71026 29538 71038
rect 4174 70978 4226 70990
rect 6414 70978 6466 70990
rect 10670 70978 10722 70990
rect 36430 70978 36482 70990
rect 2370 70926 2382 70978
rect 2434 70926 2446 70978
rect 4610 70926 4622 70978
rect 4674 70926 4686 70978
rect 7186 70926 7198 70978
rect 7250 70926 7262 70978
rect 11666 70926 11678 70978
rect 11730 70926 11742 70978
rect 22866 70926 22878 70978
rect 22930 70926 22942 70978
rect 32834 70926 32846 70978
rect 32898 70926 32910 70978
rect 33618 70926 33630 70978
rect 33682 70926 33694 70978
rect 34962 70926 34974 70978
rect 35026 70926 35038 70978
rect 35970 70926 35982 70978
rect 36034 70926 36046 70978
rect 36978 70926 36990 70978
rect 37042 70926 37054 70978
rect 4174 70914 4226 70926
rect 6414 70914 6466 70926
rect 10670 70914 10722 70926
rect 36430 70914 36482 70926
rect 3614 70866 3666 70878
rect 5966 70866 6018 70878
rect 5618 70814 5630 70866
rect 5682 70814 5694 70866
rect 33282 70814 33294 70866
rect 33346 70814 33358 70866
rect 3614 70802 3666 70814
rect 5966 70802 6018 70814
rect 8766 70754 8818 70766
rect 8766 70690 8818 70702
rect 13022 70754 13074 70766
rect 13022 70690 13074 70702
rect 21422 70754 21474 70766
rect 21422 70690 21474 70702
rect 22430 70754 22482 70766
rect 22430 70690 22482 70702
rect 26126 70754 26178 70766
rect 26126 70690 26178 70702
rect 26910 70754 26962 70766
rect 26910 70690 26962 70702
rect 1344 70586 48608 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 48608 70586
rect 1344 70500 48608 70534
rect 16830 70418 16882 70430
rect 4386 70366 4398 70418
rect 4450 70366 4462 70418
rect 6290 70366 6302 70418
rect 6354 70366 6366 70418
rect 16830 70354 16882 70366
rect 34078 70418 34130 70430
rect 34078 70354 34130 70366
rect 38334 70418 38386 70430
rect 38334 70354 38386 70366
rect 38782 70418 38834 70430
rect 38782 70354 38834 70366
rect 34414 70306 34466 70318
rect 4946 70254 4958 70306
rect 5010 70254 5022 70306
rect 34414 70242 34466 70254
rect 34638 70306 34690 70318
rect 34638 70242 34690 70254
rect 38894 70306 38946 70318
rect 38894 70242 38946 70254
rect 6750 70194 6802 70206
rect 12350 70194 12402 70206
rect 14702 70194 14754 70206
rect 26574 70194 26626 70206
rect 28030 70194 28082 70206
rect 5618 70142 5630 70194
rect 5682 70142 5694 70194
rect 7522 70142 7534 70194
rect 7586 70142 7598 70194
rect 9874 70142 9886 70194
rect 9938 70142 9950 70194
rect 10770 70142 10782 70194
rect 10834 70142 10846 70194
rect 13346 70142 13358 70194
rect 13410 70142 13422 70194
rect 17714 70142 17726 70194
rect 17778 70142 17790 70194
rect 23090 70142 23102 70194
rect 23154 70142 23166 70194
rect 23426 70142 23438 70194
rect 23490 70142 23502 70194
rect 23986 70142 23998 70194
rect 24050 70142 24062 70194
rect 25442 70142 25454 70194
rect 25506 70142 25518 70194
rect 25778 70142 25790 70194
rect 25842 70142 25854 70194
rect 26898 70142 26910 70194
rect 26962 70142 26974 70194
rect 6750 70130 6802 70142
rect 12350 70130 12402 70142
rect 14702 70130 14754 70142
rect 26574 70130 26626 70142
rect 28030 70130 28082 70142
rect 29038 70194 29090 70206
rect 29038 70130 29090 70142
rect 29934 70194 29986 70206
rect 29934 70130 29986 70142
rect 31166 70194 31218 70206
rect 38446 70194 38498 70206
rect 35074 70142 35086 70194
rect 35138 70142 35150 70194
rect 31166 70130 31218 70142
rect 38446 70130 38498 70142
rect 3838 70082 3890 70094
rect 3838 70018 3890 70030
rect 9102 70082 9154 70094
rect 20862 70082 20914 70094
rect 28366 70082 28418 70094
rect 18386 70030 18398 70082
rect 18450 70030 18462 70082
rect 20514 70030 20526 70082
rect 20578 70030 20590 70082
rect 23314 70030 23326 70082
rect 23378 70030 23390 70082
rect 24434 70030 24446 70082
rect 24498 70030 24510 70082
rect 26002 70030 26014 70082
rect 26066 70030 26078 70082
rect 9102 70018 9154 70030
rect 20862 70018 20914 70030
rect 28366 70018 28418 70030
rect 29262 70082 29314 70094
rect 29262 70018 29314 70030
rect 29710 70082 29762 70094
rect 29710 70018 29762 70030
rect 30718 70082 30770 70094
rect 30718 70018 30770 70030
rect 31614 70082 31666 70094
rect 31614 70018 31666 70030
rect 33630 70082 33682 70094
rect 34738 70030 34750 70082
rect 34802 70030 34814 70082
rect 35858 70030 35870 70082
rect 35922 70030 35934 70082
rect 37986 70030 37998 70082
rect 38050 70030 38062 70082
rect 33630 70018 33682 70030
rect 4062 69970 4114 69982
rect 4062 69906 4114 69918
rect 11902 69970 11954 69982
rect 11902 69906 11954 69918
rect 20974 69970 21026 69982
rect 28702 69970 28754 69982
rect 24210 69918 24222 69970
rect 24274 69918 24286 69970
rect 26786 69918 26798 69970
rect 26850 69918 26862 69970
rect 20974 69906 21026 69918
rect 28702 69906 28754 69918
rect 30270 69970 30322 69982
rect 30270 69906 30322 69918
rect 1344 69802 48608 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 48608 69802
rect 1344 69716 48608 69750
rect 5630 69634 5682 69646
rect 35970 69582 35982 69634
rect 36034 69582 36046 69634
rect 5630 69570 5682 69582
rect 4622 69522 4674 69534
rect 4622 69458 4674 69470
rect 5742 69522 5794 69534
rect 5742 69458 5794 69470
rect 6190 69522 6242 69534
rect 6190 69458 6242 69470
rect 6638 69522 6690 69534
rect 6638 69458 6690 69470
rect 13022 69522 13074 69534
rect 23426 69470 23438 69522
rect 23490 69470 23502 69522
rect 25666 69470 25678 69522
rect 25730 69470 25742 69522
rect 27794 69470 27806 69522
rect 27858 69470 27870 69522
rect 32498 69470 32510 69522
rect 32562 69470 32574 69522
rect 34962 69470 34974 69522
rect 35026 69470 35038 69522
rect 13022 69458 13074 69470
rect 10670 69410 10722 69422
rect 18734 69410 18786 69422
rect 11442 69358 11454 69410
rect 11506 69358 11518 69410
rect 10670 69346 10722 69358
rect 18734 69346 18786 69358
rect 21422 69410 21474 69422
rect 28590 69410 28642 69422
rect 37102 69410 37154 69422
rect 21858 69358 21870 69410
rect 21922 69358 21934 69410
rect 22530 69358 22542 69410
rect 22594 69358 22606 69410
rect 23090 69358 23102 69410
rect 23154 69358 23166 69410
rect 24994 69358 25006 69410
rect 25058 69358 25070 69410
rect 29586 69358 29598 69410
rect 29650 69358 29662 69410
rect 34850 69358 34862 69410
rect 34914 69358 34926 69410
rect 35634 69358 35646 69410
rect 35698 69358 35710 69410
rect 35858 69358 35870 69410
rect 35922 69358 35934 69410
rect 21422 69346 21474 69358
rect 28590 69346 28642 69358
rect 37102 69346 37154 69358
rect 18510 69298 18562 69310
rect 18510 69234 18562 69246
rect 19070 69298 19122 69310
rect 19070 69234 19122 69246
rect 22318 69298 22370 69310
rect 30370 69246 30382 69298
rect 30434 69246 30446 69298
rect 22318 69234 22370 69246
rect 9438 69186 9490 69198
rect 9438 69122 9490 69134
rect 10334 69186 10386 69198
rect 10334 69122 10386 69134
rect 18958 69186 19010 69198
rect 18958 69122 19010 69134
rect 24110 69186 24162 69198
rect 24110 69122 24162 69134
rect 24558 69186 24610 69198
rect 24558 69122 24610 69134
rect 28254 69186 28306 69198
rect 28254 69122 28306 69134
rect 32958 69186 33010 69198
rect 32958 69122 33010 69134
rect 34190 69186 34242 69198
rect 34190 69122 34242 69134
rect 1344 69018 48608 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 48608 69018
rect 1344 68932 48608 68966
rect 12014 68850 12066 68862
rect 12014 68786 12066 68798
rect 19742 68850 19794 68862
rect 19742 68786 19794 68798
rect 23774 68850 23826 68862
rect 23774 68786 23826 68798
rect 25342 68850 25394 68862
rect 25342 68786 25394 68798
rect 30494 68850 30546 68862
rect 30494 68786 30546 68798
rect 35534 68850 35586 68862
rect 35534 68786 35586 68798
rect 2494 68738 2546 68750
rect 2494 68674 2546 68686
rect 2942 68738 2994 68750
rect 2942 68674 2994 68686
rect 3390 68738 3442 68750
rect 3390 68674 3442 68686
rect 24670 68738 24722 68750
rect 33070 68738 33122 68750
rect 28018 68686 28030 68738
rect 28082 68686 28094 68738
rect 24670 68674 24722 68686
rect 33070 68674 33122 68686
rect 20302 68626 20354 68638
rect 22430 68626 22482 68638
rect 20850 68574 20862 68626
rect 20914 68574 20926 68626
rect 21410 68574 21422 68626
rect 21474 68574 21486 68626
rect 21970 68574 21982 68626
rect 22034 68574 22046 68626
rect 20302 68562 20354 68574
rect 22430 68562 22482 68574
rect 23102 68626 23154 68638
rect 33406 68626 33458 68638
rect 27346 68574 27358 68626
rect 27410 68574 27422 68626
rect 30706 68574 30718 68626
rect 30770 68574 30782 68626
rect 23102 68562 23154 68574
rect 33406 68562 33458 68574
rect 19630 68514 19682 68526
rect 19630 68450 19682 68462
rect 24222 68514 24274 68526
rect 24222 68450 24274 68462
rect 25790 68514 25842 68526
rect 25790 68450 25842 68462
rect 26910 68514 26962 68526
rect 35646 68514 35698 68526
rect 30146 68462 30158 68514
rect 30210 68462 30222 68514
rect 26910 68450 26962 68462
rect 35646 68450 35698 68462
rect 21858 68350 21870 68402
rect 21922 68350 21934 68402
rect 24210 68350 24222 68402
rect 24274 68399 24286 68402
rect 24546 68399 24558 68402
rect 24274 68353 24558 68399
rect 24274 68350 24286 68353
rect 24546 68350 24558 68353
rect 24610 68399 24622 68402
rect 24770 68399 24782 68402
rect 24610 68353 24782 68399
rect 24610 68350 24622 68353
rect 24770 68350 24782 68353
rect 24834 68350 24846 68402
rect 1344 68234 48608 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 48608 68234
rect 1344 68148 48608 68182
rect 3838 68066 3890 68078
rect 10782 68066 10834 68078
rect 5730 68014 5742 68066
rect 5794 68014 5806 68066
rect 3838 68002 3890 68014
rect 10782 68002 10834 68014
rect 20302 68066 20354 68078
rect 20302 68002 20354 68014
rect 8318 67954 8370 67966
rect 6402 67902 6414 67954
rect 6466 67902 6478 67954
rect 8318 67890 8370 67902
rect 16382 67954 16434 67966
rect 23326 67954 23378 67966
rect 19618 67902 19630 67954
rect 19682 67902 19694 67954
rect 32610 67902 32622 67954
rect 32674 67902 32686 67954
rect 34738 67902 34750 67954
rect 34802 67902 34814 67954
rect 16382 67890 16434 67902
rect 23326 67890 23378 67902
rect 2942 67842 2994 67854
rect 2942 67778 2994 67790
rect 3166 67842 3218 67854
rect 3166 67778 3218 67790
rect 3502 67842 3554 67854
rect 7646 67842 7698 67854
rect 6066 67790 6078 67842
rect 6130 67790 6142 67842
rect 8754 67790 8766 67842
rect 8818 67790 8830 67842
rect 9650 67790 9662 67842
rect 9714 67790 9726 67842
rect 16818 67790 16830 67842
rect 16882 67790 16894 67842
rect 31826 67790 31838 67842
rect 31890 67790 31902 67842
rect 3502 67778 3554 67790
rect 7646 67778 7698 67790
rect 2270 67730 2322 67742
rect 20414 67730 20466 67742
rect 2594 67678 2606 67730
rect 2658 67678 2670 67730
rect 17490 67678 17502 67730
rect 17554 67678 17566 67730
rect 2270 67666 2322 67678
rect 20414 67666 20466 67678
rect 21422 67730 21474 67742
rect 21422 67666 21474 67678
rect 1934 67618 1986 67630
rect 1934 67554 1986 67566
rect 3726 67618 3778 67630
rect 3726 67554 3778 67566
rect 7198 67618 7250 67630
rect 7198 67554 7250 67566
rect 22878 67618 22930 67630
rect 22878 67554 22930 67566
rect 31502 67618 31554 67630
rect 31502 67554 31554 67566
rect 1344 67450 48608 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 48608 67450
rect 1344 67364 48608 67398
rect 3726 67282 3778 67294
rect 3726 67218 3778 67230
rect 17950 67282 18002 67294
rect 17950 67218 18002 67230
rect 3614 67170 3666 67182
rect 3614 67106 3666 67118
rect 6526 67170 6578 67182
rect 33618 67118 33630 67170
rect 33682 67118 33694 67170
rect 35074 67118 35086 67170
rect 35138 67118 35150 67170
rect 37202 67118 37214 67170
rect 37266 67118 37278 67170
rect 39218 67118 39230 67170
rect 39282 67118 39294 67170
rect 6526 67106 6578 67118
rect 3054 67058 3106 67070
rect 6862 67058 6914 67070
rect 1810 67006 1822 67058
rect 1874 67006 1886 67058
rect 4050 67006 4062 67058
rect 4114 67006 4126 67058
rect 5506 67006 5518 67058
rect 5570 67006 5582 67058
rect 3054 66994 3106 67006
rect 6862 66994 6914 67006
rect 7310 67058 7362 67070
rect 18286 67058 18338 67070
rect 7522 67006 7534 67058
rect 7586 67006 7598 67058
rect 10770 67006 10782 67058
rect 10834 67006 10846 67058
rect 11666 67006 11678 67058
rect 11730 67006 11742 67058
rect 27458 67006 27470 67058
rect 27522 67006 27534 67058
rect 35298 67006 35310 67058
rect 35362 67006 35374 67058
rect 36978 67006 36990 67058
rect 37042 67006 37054 67058
rect 38546 67006 38558 67058
rect 38610 67006 38622 67058
rect 7310 66994 7362 67006
rect 18286 66994 18338 67006
rect 2942 66946 2994 66958
rect 2942 66882 2994 66894
rect 4846 66946 4898 66958
rect 4846 66882 4898 66894
rect 6078 66946 6130 66958
rect 25342 66946 25394 66958
rect 8754 66894 8766 66946
rect 8818 66894 8830 66946
rect 6078 66882 6130 66894
rect 25342 66882 25394 66894
rect 27246 66946 27298 66958
rect 27246 66882 27298 66894
rect 28030 66946 28082 66958
rect 28030 66882 28082 66894
rect 28590 66946 28642 66958
rect 28590 66882 28642 66894
rect 32622 66946 32674 66958
rect 32622 66882 32674 66894
rect 33070 66946 33122 66958
rect 33070 66882 33122 66894
rect 34190 66946 34242 66958
rect 34190 66882 34242 66894
rect 34526 66946 34578 66958
rect 34526 66882 34578 66894
rect 6974 66834 7026 66846
rect 6974 66770 7026 66782
rect 9662 66834 9714 66846
rect 9662 66770 9714 66782
rect 27806 66834 27858 66846
rect 27806 66770 27858 66782
rect 33294 66834 33346 66846
rect 33294 66770 33346 66782
rect 1344 66666 48608 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 48608 66666
rect 1344 66580 48608 66614
rect 7870 66498 7922 66510
rect 2594 66446 2606 66498
rect 2658 66446 2670 66498
rect 7186 66446 7198 66498
rect 7250 66446 7262 66498
rect 33618 66446 33630 66498
rect 33682 66495 33694 66498
rect 34178 66495 34190 66498
rect 33682 66449 34190 66495
rect 33682 66446 33694 66449
rect 34178 66446 34190 66449
rect 34242 66446 34254 66498
rect 7870 66434 7922 66446
rect 3614 66386 3666 66398
rect 2930 66334 2942 66386
rect 2994 66334 3006 66386
rect 3614 66322 3666 66334
rect 4286 66386 4338 66398
rect 4286 66322 4338 66334
rect 4734 66386 4786 66398
rect 14702 66386 14754 66398
rect 33630 66386 33682 66398
rect 6738 66334 6750 66386
rect 6802 66334 6814 66386
rect 9426 66334 9438 66386
rect 9490 66334 9502 66386
rect 25218 66334 25230 66386
rect 25282 66334 25294 66386
rect 28466 66334 28478 66386
rect 28530 66334 28542 66386
rect 39890 66334 39902 66386
rect 39954 66334 39966 66386
rect 4734 66322 4786 66334
rect 14702 66322 14754 66334
rect 33630 66322 33682 66334
rect 7646 66274 7698 66286
rect 21758 66274 21810 66286
rect 2706 66222 2718 66274
rect 2770 66222 2782 66274
rect 6626 66222 6638 66274
rect 6690 66222 6702 66274
rect 11106 66222 11118 66274
rect 11170 66222 11182 66274
rect 12450 66222 12462 66274
rect 12514 66222 12526 66274
rect 13458 66222 13470 66274
rect 13522 66222 13534 66274
rect 22306 66222 22318 66274
rect 22370 66222 22382 66274
rect 25666 66222 25678 66274
rect 25730 66222 25742 66274
rect 36194 66222 36206 66274
rect 36258 66222 36270 66274
rect 36978 66222 36990 66274
rect 37042 66222 37054 66274
rect 7646 66210 7698 66222
rect 21758 66210 21810 66222
rect 3502 66162 3554 66174
rect 14814 66162 14866 66174
rect 36430 66162 36482 66174
rect 8194 66110 8206 66162
rect 8258 66110 8270 66162
rect 8530 66110 8542 66162
rect 8594 66110 8606 66162
rect 23090 66110 23102 66162
rect 23154 66110 23166 66162
rect 26338 66110 26350 66162
rect 26402 66110 26414 66162
rect 37762 66110 37774 66162
rect 37826 66110 37838 66162
rect 3502 66098 3554 66110
rect 14814 66098 14866 66110
rect 36430 66098 36482 66110
rect 3726 66050 3778 66062
rect 3726 65986 3778 65998
rect 4174 66050 4226 66062
rect 4174 65986 4226 65998
rect 10222 66050 10274 66062
rect 10222 65986 10274 65998
rect 11342 66050 11394 66062
rect 11342 65986 11394 65998
rect 21422 66050 21474 66062
rect 21422 65986 21474 65998
rect 21870 66050 21922 66062
rect 21870 65986 21922 65998
rect 34078 66050 34130 66062
rect 34078 65986 34130 65998
rect 35758 66050 35810 66062
rect 35758 65986 35810 65998
rect 1344 65882 48608 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 48608 65882
rect 1344 65796 48608 65830
rect 7310 65714 7362 65726
rect 7310 65650 7362 65662
rect 14366 65714 14418 65726
rect 14366 65650 14418 65662
rect 26462 65714 26514 65726
rect 38098 65662 38110 65714
rect 38162 65662 38174 65714
rect 26462 65650 26514 65662
rect 25342 65602 25394 65614
rect 25342 65538 25394 65550
rect 30494 65602 30546 65614
rect 34738 65550 34750 65602
rect 34802 65550 34814 65602
rect 37426 65550 37438 65602
rect 37490 65550 37502 65602
rect 30494 65538 30546 65550
rect 2718 65490 2770 65502
rect 2718 65426 2770 65438
rect 7758 65490 7810 65502
rect 12126 65490 12178 65502
rect 14478 65490 14530 65502
rect 30830 65490 30882 65502
rect 9538 65438 9550 65490
rect 9602 65438 9614 65490
rect 10770 65438 10782 65490
rect 10834 65438 10846 65490
rect 13122 65438 13134 65490
rect 13186 65438 13198 65490
rect 17938 65438 17950 65490
rect 18002 65438 18014 65490
rect 21186 65438 21198 65490
rect 21250 65438 21262 65490
rect 26674 65438 26686 65490
rect 26738 65438 26750 65490
rect 7758 65426 7810 65438
rect 12126 65426 12178 65438
rect 14478 65426 14530 65438
rect 30830 65426 30882 65438
rect 32062 65490 32114 65502
rect 32062 65426 32114 65438
rect 33742 65490 33794 65502
rect 39230 65490 39282 65502
rect 34178 65438 34190 65490
rect 34242 65438 34254 65490
rect 35970 65438 35982 65490
rect 36034 65438 36046 65490
rect 38322 65438 38334 65490
rect 38386 65438 38398 65490
rect 33742 65426 33794 65438
rect 39230 65426 39282 65438
rect 4062 65378 4114 65390
rect 4062 65314 4114 65326
rect 8206 65378 8258 65390
rect 8206 65314 8258 65326
rect 8990 65378 9042 65390
rect 8990 65314 9042 65326
rect 12014 65378 12066 65390
rect 12014 65314 12066 65326
rect 17614 65378 17666 65390
rect 24446 65378 24498 65390
rect 18722 65326 18734 65378
rect 18786 65326 18798 65378
rect 20850 65326 20862 65378
rect 20914 65326 20926 65378
rect 21970 65326 21982 65378
rect 22034 65326 22046 65378
rect 24098 65326 24110 65378
rect 24162 65326 24174 65378
rect 17614 65314 17666 65326
rect 24446 65314 24498 65326
rect 32510 65378 32562 65390
rect 32510 65314 32562 65326
rect 39006 65378 39058 65390
rect 39006 65314 39058 65326
rect 39678 65378 39730 65390
rect 39678 65314 39730 65326
rect 2830 65266 2882 65278
rect 24558 65266 24610 65278
rect 10098 65214 10110 65266
rect 10162 65214 10174 65266
rect 2830 65202 2882 65214
rect 24558 65202 24610 65214
rect 25454 65266 25506 65278
rect 33518 65266 33570 65278
rect 33170 65214 33182 65266
rect 33234 65214 33246 65266
rect 38658 65214 38670 65266
rect 38722 65214 38734 65266
rect 25454 65202 25506 65214
rect 33518 65202 33570 65214
rect 1344 65098 48608 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 48608 65098
rect 1344 65012 48608 65046
rect 21422 64930 21474 64942
rect 21422 64866 21474 64878
rect 22094 64930 22146 64942
rect 36978 64878 36990 64930
rect 37042 64878 37054 64930
rect 22094 64866 22146 64878
rect 23538 64766 23550 64818
rect 23602 64766 23614 64818
rect 25666 64766 25678 64818
rect 25730 64766 25742 64818
rect 30146 64766 30158 64818
rect 30210 64766 30222 64818
rect 32274 64766 32286 64818
rect 32338 64766 32350 64818
rect 35746 64766 35758 64818
rect 35810 64766 35822 64818
rect 37986 64766 37998 64818
rect 38050 64766 38062 64818
rect 10782 64706 10834 64718
rect 37326 64706 37378 64718
rect 9426 64654 9438 64706
rect 9490 64654 9502 64706
rect 28578 64654 28590 64706
rect 28642 64654 28654 64706
rect 29362 64654 29374 64706
rect 29426 64654 29438 64706
rect 32834 64654 32846 64706
rect 32898 64654 32910 64706
rect 10782 64642 10834 64654
rect 37326 64642 37378 64654
rect 37550 64706 37602 64718
rect 40786 64654 40798 64706
rect 40850 64654 40862 64706
rect 37550 64642 37602 64654
rect 18510 64594 18562 64606
rect 18510 64530 18562 64542
rect 21758 64594 21810 64606
rect 21758 64530 21810 64542
rect 22430 64594 22482 64606
rect 22430 64530 22482 64542
rect 23326 64594 23378 64606
rect 27794 64542 27806 64594
rect 27858 64542 27870 64594
rect 33618 64542 33630 64594
rect 33682 64542 33694 64594
rect 40114 64542 40126 64594
rect 40178 64542 40190 64594
rect 23326 64530 23378 64542
rect 10670 64482 10722 64494
rect 10670 64418 10722 64430
rect 18622 64482 18674 64494
rect 18622 64418 18674 64430
rect 20750 64482 20802 64494
rect 20750 64418 20802 64430
rect 21534 64482 21586 64494
rect 21534 64418 21586 64430
rect 22206 64482 22258 64494
rect 22206 64418 22258 64430
rect 22878 64482 22930 64494
rect 22878 64418 22930 64430
rect 23550 64482 23602 64494
rect 23550 64418 23602 64430
rect 24110 64482 24162 64494
rect 24110 64418 24162 64430
rect 25342 64482 25394 64494
rect 25342 64418 25394 64430
rect 36430 64482 36482 64494
rect 36430 64418 36482 64430
rect 1344 64314 48608 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 48608 64314
rect 1344 64228 48608 64262
rect 5294 64146 5346 64158
rect 5294 64082 5346 64094
rect 21982 64146 22034 64158
rect 21982 64082 22034 64094
rect 27918 64146 27970 64158
rect 27918 64082 27970 64094
rect 30606 64146 30658 64158
rect 33854 64146 33906 64158
rect 30930 64094 30942 64146
rect 30994 64094 31006 64146
rect 30606 64082 30658 64094
rect 33854 64082 33906 64094
rect 34526 64146 34578 64158
rect 34526 64082 34578 64094
rect 39678 64146 39730 64158
rect 39678 64082 39730 64094
rect 22878 64034 22930 64046
rect 22878 63970 22930 63982
rect 33518 64034 33570 64046
rect 35186 63982 35198 64034
rect 35250 63982 35262 64034
rect 33518 63970 33570 63982
rect 16830 63922 16882 63934
rect 22766 63922 22818 63934
rect 10770 63870 10782 63922
rect 10834 63870 10846 63922
rect 12114 63870 12126 63922
rect 12178 63870 12190 63922
rect 17378 63870 17390 63922
rect 17442 63870 17454 63922
rect 16830 63858 16882 63870
rect 22766 63858 22818 63870
rect 28254 63922 28306 63934
rect 28254 63858 28306 63870
rect 28702 63922 28754 63934
rect 28702 63858 28754 63870
rect 31278 63922 31330 63934
rect 31278 63858 31330 63870
rect 31502 63922 31554 63934
rect 31502 63858 31554 63870
rect 32510 63922 32562 63934
rect 32510 63858 32562 63870
rect 33182 63922 33234 63934
rect 37774 63922 37826 63934
rect 35298 63870 35310 63922
rect 35362 63870 35374 63922
rect 37090 63870 37102 63922
rect 37154 63870 37166 63922
rect 38546 63870 38558 63922
rect 38610 63870 38622 63922
rect 33182 63858 33234 63870
rect 37774 63858 37826 63870
rect 11902 63810 11954 63822
rect 37662 63810 37714 63822
rect 18162 63758 18174 63810
rect 18226 63758 18238 63810
rect 20290 63758 20302 63810
rect 20354 63758 20366 63810
rect 11902 63746 11954 63758
rect 37662 63746 37714 63758
rect 1344 63530 48608 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 48608 63530
rect 1344 63444 48608 63478
rect 7758 63362 7810 63374
rect 4050 63310 4062 63362
rect 4114 63359 4126 63362
rect 4946 63359 4958 63362
rect 4114 63313 4958 63359
rect 4114 63310 4126 63313
rect 4946 63310 4958 63313
rect 5010 63310 5022 63362
rect 7758 63298 7810 63310
rect 19182 63362 19234 63374
rect 19182 63298 19234 63310
rect 30382 63362 30434 63374
rect 30382 63298 30434 63310
rect 4062 63250 4114 63262
rect 4062 63186 4114 63198
rect 4510 63250 4562 63262
rect 4510 63186 4562 63198
rect 4958 63250 5010 63262
rect 30606 63250 30658 63262
rect 16370 63198 16382 63250
rect 16434 63198 16446 63250
rect 18498 63198 18510 63250
rect 18562 63198 18574 63250
rect 18946 63198 18958 63250
rect 19010 63198 19022 63250
rect 4958 63186 5010 63198
rect 30606 63186 30658 63198
rect 31054 63250 31106 63262
rect 31054 63186 31106 63198
rect 31950 63250 32002 63262
rect 31950 63186 32002 63198
rect 37550 63250 37602 63262
rect 37550 63186 37602 63198
rect 37998 63250 38050 63262
rect 37998 63186 38050 63198
rect 39230 63250 39282 63262
rect 39230 63186 39282 63198
rect 5630 63138 5682 63150
rect 14814 63138 14866 63150
rect 19630 63138 19682 63150
rect 37326 63138 37378 63150
rect 6402 63086 6414 63138
rect 6466 63086 6478 63138
rect 8306 63086 8318 63138
rect 8370 63086 8382 63138
rect 13458 63086 13470 63138
rect 13522 63086 13534 63138
rect 15586 63086 15598 63138
rect 15650 63086 15662 63138
rect 18834 63086 18846 63138
rect 18898 63086 18910 63138
rect 32386 63086 32398 63138
rect 32450 63086 32462 63138
rect 33954 63086 33966 63138
rect 34018 63086 34030 63138
rect 36418 63086 36430 63138
rect 36482 63086 36494 63138
rect 38546 63086 38558 63138
rect 38610 63086 38622 63138
rect 5630 63074 5682 63086
rect 14814 63074 14866 63086
rect 19630 63074 19682 63086
rect 37326 63074 37378 63086
rect 2718 63026 2770 63038
rect 2718 62962 2770 62974
rect 9550 63026 9602 63038
rect 38782 63026 38834 63038
rect 32946 62974 32958 63026
rect 33010 62974 33022 63026
rect 35634 62974 35646 63026
rect 35698 62974 35710 63026
rect 9550 62962 9602 62974
rect 38782 62962 38834 62974
rect 2382 62914 2434 62926
rect 2382 62850 2434 62862
rect 9438 62914 9490 62926
rect 9438 62850 9490 62862
rect 14702 62914 14754 62926
rect 34862 62914 34914 62926
rect 30034 62862 30046 62914
rect 30098 62862 30110 62914
rect 36978 62862 36990 62914
rect 37042 62862 37054 62914
rect 14702 62850 14754 62862
rect 34862 62850 34914 62862
rect 1344 62746 48608 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 48608 62746
rect 1344 62660 48608 62694
rect 3054 62578 3106 62590
rect 7422 62578 7474 62590
rect 3714 62526 3726 62578
rect 3778 62526 3790 62578
rect 3054 62514 3106 62526
rect 7422 62514 7474 62526
rect 14254 62578 14306 62590
rect 14254 62514 14306 62526
rect 35982 62578 36034 62590
rect 35982 62514 36034 62526
rect 17726 62466 17778 62478
rect 17726 62402 17778 62414
rect 17950 62466 18002 62478
rect 17950 62402 18002 62414
rect 18510 62466 18562 62478
rect 18510 62402 18562 62414
rect 18958 62466 19010 62478
rect 18958 62402 19010 62414
rect 19630 62466 19682 62478
rect 19630 62402 19682 62414
rect 23326 62466 23378 62478
rect 23326 62402 23378 62414
rect 23662 62466 23714 62478
rect 23662 62402 23714 62414
rect 23774 62466 23826 62478
rect 23774 62402 23826 62414
rect 4286 62354 4338 62366
rect 1922 62302 1934 62354
rect 1986 62302 1998 62354
rect 3266 62302 3278 62354
rect 3330 62302 3342 62354
rect 4286 62290 4338 62302
rect 4622 62354 4674 62366
rect 31726 62354 31778 62366
rect 5170 62302 5182 62354
rect 5234 62302 5246 62354
rect 6066 62302 6078 62354
rect 6130 62302 6142 62354
rect 10322 62302 10334 62354
rect 10386 62302 10398 62354
rect 11666 62302 11678 62354
rect 11730 62302 11742 62354
rect 13010 62302 13022 62354
rect 13074 62302 13086 62354
rect 14466 62302 14478 62354
rect 14530 62302 14542 62354
rect 28354 62302 28366 62354
rect 28418 62302 28430 62354
rect 39106 62302 39118 62354
rect 39170 62302 39182 62354
rect 4622 62290 4674 62302
rect 31726 62290 31778 62302
rect 11454 62242 11506 62254
rect 18050 62190 18062 62242
rect 18114 62190 18126 62242
rect 29138 62190 29150 62242
rect 29202 62190 29214 62242
rect 31266 62190 31278 62242
rect 31330 62190 31342 62242
rect 36306 62190 36318 62242
rect 36370 62190 36382 62242
rect 38434 62190 38446 62242
rect 38498 62190 38510 62242
rect 11454 62178 11506 62190
rect 4062 62130 4114 62142
rect 4062 62066 4114 62078
rect 4734 62130 4786 62142
rect 4734 62066 4786 62078
rect 19742 62130 19794 62142
rect 19742 62066 19794 62078
rect 23774 62130 23826 62142
rect 23774 62066 23826 62078
rect 1344 61962 48608 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 48608 61962
rect 1344 61876 48608 61910
rect 32958 61794 33010 61806
rect 4274 61742 4286 61794
rect 4338 61742 4350 61794
rect 32958 61730 33010 61742
rect 3054 61682 3106 61694
rect 3054 61618 3106 61630
rect 5742 61682 5794 61694
rect 5742 61618 5794 61630
rect 14702 61682 14754 61694
rect 21646 61682 21698 61694
rect 26238 61682 26290 61694
rect 20738 61630 20750 61682
rect 20802 61630 20814 61682
rect 23762 61630 23774 61682
rect 23826 61630 23838 61682
rect 25890 61630 25902 61682
rect 25954 61630 25966 61682
rect 14702 61618 14754 61630
rect 21646 61618 21698 61630
rect 26238 61618 26290 61630
rect 33182 61682 33234 61694
rect 33182 61618 33234 61630
rect 33630 61682 33682 61694
rect 33630 61618 33682 61630
rect 39566 61682 39618 61694
rect 42802 61630 42814 61682
rect 42866 61630 42878 61682
rect 39566 61618 39618 61630
rect 4622 61570 4674 61582
rect 14814 61570 14866 61582
rect 30046 61570 30098 61582
rect 1922 61518 1934 61570
rect 1986 61518 1998 61570
rect 3266 61518 3278 61570
rect 3330 61518 3342 61570
rect 3938 61518 3950 61570
rect 4002 61518 4014 61570
rect 7634 61518 7646 61570
rect 7698 61518 7710 61570
rect 9426 61518 9438 61570
rect 9490 61518 9502 61570
rect 13458 61518 13470 61570
rect 13522 61518 13534 61570
rect 17826 61518 17838 61570
rect 17890 61518 17902 61570
rect 22978 61518 22990 61570
rect 23042 61518 23054 61570
rect 4622 61506 4674 61518
rect 14814 61506 14866 61518
rect 30046 61506 30098 61518
rect 37102 61570 37154 61582
rect 39890 61518 39902 61570
rect 39954 61518 39966 61570
rect 37102 61506 37154 61518
rect 5630 61458 5682 61470
rect 5630 61394 5682 61406
rect 5854 61458 5906 61470
rect 5854 61394 5906 61406
rect 8878 61458 8930 61470
rect 8878 61394 8930 61406
rect 10782 61458 10834 61470
rect 29710 61458 29762 61470
rect 18610 61406 18622 61458
rect 18674 61406 18686 61458
rect 40674 61406 40686 61458
rect 40738 61406 40750 61458
rect 10782 61394 10834 61406
rect 29710 61394 29762 61406
rect 8766 61346 8818 61358
rect 8766 61282 8818 61294
rect 10670 61346 10722 61358
rect 10670 61282 10722 61294
rect 17502 61346 17554 61358
rect 17502 61282 17554 61294
rect 21758 61346 21810 61358
rect 21758 61282 21810 61294
rect 22654 61346 22706 61358
rect 22654 61282 22706 61294
rect 26350 61346 26402 61358
rect 37438 61346 37490 61358
rect 32610 61294 32622 61346
rect 32674 61294 32686 61346
rect 26350 61282 26402 61294
rect 37438 61282 37490 61294
rect 1344 61178 48608 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 48608 61178
rect 1344 61092 48608 61126
rect 19854 61010 19906 61022
rect 19854 60946 19906 60958
rect 20638 61010 20690 61022
rect 20638 60946 20690 60958
rect 24558 61010 24610 61022
rect 24558 60946 24610 60958
rect 19966 60898 20018 60910
rect 16482 60846 16494 60898
rect 16546 60846 16558 60898
rect 19966 60834 20018 60846
rect 32174 60898 32226 60910
rect 32174 60834 32226 60846
rect 32510 60898 32562 60910
rect 32510 60834 32562 60846
rect 40238 60898 40290 60910
rect 40238 60834 40290 60846
rect 8766 60786 8818 60798
rect 7522 60734 7534 60786
rect 7586 60734 7598 60786
rect 15362 60734 15374 60786
rect 15426 60734 15438 60786
rect 20962 60734 20974 60786
rect 21026 60734 21038 60786
rect 25218 60734 25230 60786
rect 25282 60734 25294 60786
rect 33170 60734 33182 60786
rect 33234 60734 33246 60786
rect 40898 60734 40910 60786
rect 40962 60734 40974 60786
rect 8766 60722 8818 60734
rect 3726 60674 3778 60686
rect 3726 60610 3778 60622
rect 3838 60674 3890 60686
rect 3838 60610 3890 60622
rect 5070 60674 5122 60686
rect 5070 60610 5122 60622
rect 8654 60674 8706 60686
rect 8654 60610 8706 60622
rect 15150 60674 15202 60686
rect 15150 60610 15202 60622
rect 19406 60674 19458 60686
rect 39678 60674 39730 60686
rect 21746 60622 21758 60674
rect 21810 60622 21822 60674
rect 23874 60622 23886 60674
rect 23938 60622 23950 60674
rect 24658 60622 24670 60674
rect 24722 60622 24734 60674
rect 26002 60622 26014 60674
rect 26066 60622 26078 60674
rect 28130 60622 28142 60674
rect 28194 60622 28206 60674
rect 33842 60622 33854 60674
rect 33906 60622 33918 60674
rect 35970 60622 35982 60674
rect 36034 60622 36046 60674
rect 40338 60622 40350 60674
rect 40402 60622 40414 60674
rect 41682 60622 41694 60674
rect 41746 60622 41758 60674
rect 43810 60622 43822 60674
rect 43874 60622 43886 60674
rect 19406 60610 19458 60622
rect 39678 60610 39730 60622
rect 19742 60562 19794 60574
rect 19742 60498 19794 60510
rect 24334 60562 24386 60574
rect 24334 60498 24386 60510
rect 40014 60562 40066 60574
rect 40014 60498 40066 60510
rect 1344 60394 48608 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 48608 60394
rect 1344 60308 48608 60342
rect 7646 60226 7698 60238
rect 7646 60162 7698 60174
rect 23774 60226 23826 60238
rect 23774 60162 23826 60174
rect 26462 60226 26514 60238
rect 26462 60162 26514 60174
rect 41246 60226 41298 60238
rect 41246 60162 41298 60174
rect 18286 60114 18338 60126
rect 17826 60062 17838 60114
rect 17890 60062 17902 60114
rect 18286 60050 18338 60062
rect 23886 60114 23938 60126
rect 23886 60050 23938 60062
rect 24894 60114 24946 60126
rect 24894 60050 24946 60062
rect 30718 60114 30770 60126
rect 30718 60050 30770 60062
rect 40126 60114 40178 60126
rect 40126 60050 40178 60062
rect 42366 60114 42418 60126
rect 42366 60050 42418 60062
rect 42814 60114 42866 60126
rect 42814 60050 42866 60062
rect 21982 60002 22034 60014
rect 15026 59950 15038 60002
rect 15090 59950 15102 60002
rect 21982 59938 22034 59950
rect 24334 60002 24386 60014
rect 24334 59938 24386 59950
rect 26798 60002 26850 60014
rect 27570 59950 27582 60002
rect 27634 59950 27646 60002
rect 31266 59950 31278 60002
rect 31330 59950 31342 60002
rect 41234 59950 41246 60002
rect 41298 59950 41310 60002
rect 26798 59938 26850 59950
rect 7534 59890 7586 59902
rect 21646 59890 21698 59902
rect 7074 59838 7086 59890
rect 7138 59838 7150 59890
rect 15698 59838 15710 59890
rect 15762 59838 15774 59890
rect 7534 59826 7586 59838
rect 21646 59826 21698 59838
rect 27022 59890 27074 59902
rect 40910 59890 40962 59902
rect 31826 59838 31838 59890
rect 31890 59838 31902 59890
rect 27022 59826 27074 59838
rect 40910 59826 40962 59838
rect 6750 59778 6802 59790
rect 6750 59714 6802 59726
rect 21758 59778 21810 59790
rect 21758 59714 21810 59726
rect 22318 59778 22370 59790
rect 22318 59714 22370 59726
rect 26126 59778 26178 59790
rect 26126 59714 26178 59726
rect 27358 59778 27410 59790
rect 27358 59714 27410 59726
rect 32734 59778 32786 59790
rect 32734 59714 32786 59726
rect 40574 59778 40626 59790
rect 40574 59714 40626 59726
rect 42254 59778 42306 59790
rect 42254 59714 42306 59726
rect 42702 59778 42754 59790
rect 42702 59714 42754 59726
rect 1344 59610 48608 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 48608 59610
rect 1344 59524 48608 59558
rect 5854 59442 5906 59454
rect 16942 59442 16994 59454
rect 6738 59390 6750 59442
rect 6802 59390 6814 59442
rect 5854 59378 5906 59390
rect 16942 59378 16994 59390
rect 18062 59442 18114 59454
rect 18062 59378 18114 59390
rect 26014 59442 26066 59454
rect 26014 59378 26066 59390
rect 33406 59442 33458 59454
rect 33406 59378 33458 59390
rect 2382 59330 2434 59342
rect 2382 59266 2434 59278
rect 12014 59330 12066 59342
rect 17390 59330 17442 59342
rect 30606 59330 30658 59342
rect 15586 59278 15598 59330
rect 15650 59278 15662 59330
rect 16370 59278 16382 59330
rect 16434 59278 16446 59330
rect 27122 59278 27134 59330
rect 27186 59278 27198 59330
rect 12014 59266 12066 59278
rect 17390 59266 17442 59278
rect 30606 59266 30658 59278
rect 6190 59218 6242 59230
rect 18398 59218 18450 59230
rect 22878 59218 22930 59230
rect 33070 59218 33122 59230
rect 10658 59166 10670 59218
rect 10722 59166 10734 59218
rect 12786 59166 12798 59218
rect 12850 59166 12862 59218
rect 14242 59166 14254 59218
rect 14306 59166 14318 59218
rect 17602 59166 17614 59218
rect 17666 59166 17678 59218
rect 21970 59166 21982 59218
rect 22034 59166 22046 59218
rect 22418 59166 22430 59218
rect 22482 59166 22494 59218
rect 23426 59166 23438 59218
rect 23490 59166 23502 59218
rect 26338 59166 26350 59218
rect 26402 59166 26414 59218
rect 6190 59154 6242 59166
rect 18398 59154 18450 59166
rect 22878 59154 22930 59166
rect 33070 59154 33122 59166
rect 34638 59218 34690 59230
rect 35074 59166 35086 59218
rect 35138 59166 35150 59218
rect 34638 59154 34690 59166
rect 4174 59106 4226 59118
rect 4174 59042 4226 59054
rect 4622 59106 4674 59118
rect 4622 59042 4674 59054
rect 5406 59106 5458 59118
rect 5406 59042 5458 59054
rect 11902 59106 11954 59118
rect 11902 59042 11954 59054
rect 14030 59106 14082 59118
rect 14030 59042 14082 59054
rect 18846 59106 18898 59118
rect 18846 59042 18898 59054
rect 19630 59106 19682 59118
rect 22766 59106 22818 59118
rect 22082 59054 22094 59106
rect 22146 59054 22158 59106
rect 19630 59042 19682 59054
rect 22766 59042 22818 59054
rect 24334 59106 24386 59118
rect 24334 59042 24386 59054
rect 24782 59106 24834 59118
rect 24782 59042 24834 59054
rect 25454 59106 25506 59118
rect 31054 59106 31106 59118
rect 29250 59054 29262 59106
rect 29314 59054 29326 59106
rect 35746 59054 35758 59106
rect 35810 59054 35822 59106
rect 37874 59054 37886 59106
rect 37938 59054 37950 59106
rect 25454 59042 25506 59054
rect 31054 59042 31106 59054
rect 2270 58994 2322 59006
rect 2270 58930 2322 58942
rect 2606 58994 2658 59006
rect 2606 58930 2658 58942
rect 6414 58994 6466 59006
rect 6414 58930 6466 58942
rect 30046 58994 30098 59006
rect 30046 58930 30098 58942
rect 30382 58994 30434 59006
rect 30382 58930 30434 58942
rect 1344 58826 48608 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 48608 58826
rect 1344 58740 48608 58774
rect 27470 58658 27522 58670
rect 24658 58606 24670 58658
rect 24722 58606 24734 58658
rect 29138 58606 29150 58658
rect 29202 58606 29214 58658
rect 27470 58594 27522 58606
rect 5070 58546 5122 58558
rect 5070 58482 5122 58494
rect 6638 58546 6690 58558
rect 25678 58546 25730 58558
rect 41134 58546 41186 58558
rect 16258 58494 16270 58546
rect 16322 58494 16334 58546
rect 18386 58494 18398 58546
rect 18450 58494 18462 58546
rect 23762 58494 23774 58546
rect 23826 58494 23838 58546
rect 24770 58494 24782 58546
rect 24834 58494 24846 58546
rect 31602 58494 31614 58546
rect 31666 58494 31678 58546
rect 33730 58494 33742 58546
rect 33794 58494 33806 58546
rect 40674 58494 40686 58546
rect 40738 58494 40750 58546
rect 6638 58482 6690 58494
rect 25678 58482 25730 58494
rect 41134 58482 41186 58494
rect 4062 58434 4114 58446
rect 6526 58434 6578 58446
rect 12014 58434 12066 58446
rect 14814 58434 14866 58446
rect 26126 58434 26178 58446
rect 1810 58382 1822 58434
rect 1874 58382 1886 58434
rect 2706 58382 2718 58434
rect 2770 58382 2782 58434
rect 4498 58382 4510 58434
rect 4562 58382 4574 58434
rect 6290 58382 6302 58434
rect 6354 58382 6366 58434
rect 10658 58382 10670 58434
rect 10722 58382 10734 58434
rect 13458 58382 13470 58434
rect 13522 58382 13534 58434
rect 15586 58382 15598 58434
rect 15650 58382 15662 58434
rect 23538 58382 23550 58434
rect 23602 58382 23614 58434
rect 24210 58382 24222 58434
rect 24274 58382 24286 58434
rect 24546 58382 24558 58434
rect 24610 58382 24622 58434
rect 4062 58370 4114 58382
rect 6526 58370 6578 58382
rect 12014 58370 12066 58382
rect 14814 58370 14866 58382
rect 26126 58370 26178 58382
rect 27134 58434 27186 58446
rect 27134 58370 27186 58382
rect 27806 58434 27858 58446
rect 27806 58370 27858 58382
rect 29486 58434 29538 58446
rect 29486 58370 29538 58382
rect 29710 58434 29762 58446
rect 34302 58434 34354 58446
rect 37550 58434 37602 58446
rect 30930 58382 30942 58434
rect 30994 58382 31006 58434
rect 35634 58382 35646 58434
rect 35698 58382 35710 58434
rect 37874 58382 37886 58434
rect 37938 58382 37950 58434
rect 29710 58370 29762 58382
rect 34302 58370 34354 58382
rect 37550 58370 37602 58382
rect 18846 58322 18898 58334
rect 18846 58258 18898 58270
rect 19294 58322 19346 58334
rect 19294 58258 19346 58270
rect 19854 58322 19906 58334
rect 19854 58258 19906 58270
rect 20302 58322 20354 58334
rect 20302 58258 20354 58270
rect 28030 58322 28082 58334
rect 28030 58258 28082 58270
rect 35870 58322 35922 58334
rect 41022 58322 41074 58334
rect 38546 58270 38558 58322
rect 38610 58270 38622 58322
rect 35870 58258 35922 58270
rect 41022 58258 41074 58270
rect 4286 58210 4338 58222
rect 4286 58146 4338 58158
rect 7198 58210 7250 58222
rect 7198 58146 7250 58158
rect 11902 58210 11954 58222
rect 11902 58146 11954 58158
rect 14702 58210 14754 58222
rect 14702 58146 14754 58158
rect 19070 58210 19122 58222
rect 19070 58146 19122 58158
rect 19406 58210 19458 58222
rect 19406 58146 19458 58158
rect 28478 58210 28530 58222
rect 28478 58146 28530 58158
rect 30158 58210 30210 58222
rect 30158 58146 30210 58158
rect 1344 58042 48608 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 48608 58042
rect 1344 57956 48608 57990
rect 2270 57874 2322 57886
rect 2270 57810 2322 57822
rect 5294 57874 5346 57886
rect 5294 57810 5346 57822
rect 6414 57874 6466 57886
rect 6414 57810 6466 57822
rect 14030 57874 14082 57886
rect 32286 57874 32338 57886
rect 17378 57822 17390 57874
rect 17442 57822 17454 57874
rect 14030 57810 14082 57822
rect 32286 57810 32338 57822
rect 32398 57874 32450 57886
rect 32398 57810 32450 57822
rect 34078 57874 34130 57886
rect 36094 57874 36146 57886
rect 35634 57822 35646 57874
rect 35698 57822 35710 57874
rect 34078 57810 34130 57822
rect 36094 57810 36146 57822
rect 2606 57762 2658 57774
rect 2606 57698 2658 57710
rect 10894 57762 10946 57774
rect 10894 57698 10946 57710
rect 17950 57762 18002 57774
rect 17950 57698 18002 57710
rect 18734 57762 18786 57774
rect 23326 57762 23378 57774
rect 20850 57710 20862 57762
rect 20914 57710 20926 57762
rect 18734 57698 18786 57710
rect 23326 57698 23378 57710
rect 31838 57762 31890 57774
rect 31838 57698 31890 57710
rect 38558 57762 38610 57774
rect 38558 57698 38610 57710
rect 38782 57762 38834 57774
rect 38782 57698 38834 57710
rect 1934 57650 1986 57662
rect 5406 57650 5458 57662
rect 8990 57650 9042 57662
rect 22430 57650 22482 57662
rect 27918 57650 27970 57662
rect 32062 57650 32114 57662
rect 3266 57598 3278 57650
rect 3330 57598 3342 57650
rect 4162 57598 4174 57650
rect 4226 57598 4238 57650
rect 7970 57598 7982 57650
rect 8034 57598 8046 57650
rect 12114 57598 12126 57650
rect 12178 57598 12190 57650
rect 12786 57598 12798 57650
rect 12850 57598 12862 57650
rect 14242 57598 14254 57650
rect 14306 57598 14318 57650
rect 18274 57598 18286 57650
rect 18338 57598 18350 57650
rect 18498 57598 18510 57650
rect 18562 57598 18574 57650
rect 18946 57598 18958 57650
rect 19010 57598 19022 57650
rect 19954 57598 19966 57650
rect 20018 57598 20030 57650
rect 20290 57598 20302 57650
rect 20354 57598 20366 57650
rect 22754 57598 22766 57650
rect 22818 57598 22830 57650
rect 25442 57598 25454 57650
rect 25506 57598 25518 57650
rect 25666 57598 25678 57650
rect 25730 57598 25742 57650
rect 26786 57598 26798 57650
rect 26850 57598 26862 57650
rect 31490 57598 31502 57650
rect 31554 57598 31566 57650
rect 1934 57586 1986 57598
rect 5406 57586 5458 57598
rect 8990 57586 9042 57598
rect 22430 57586 22482 57598
rect 27918 57586 27970 57598
rect 32062 57586 32114 57598
rect 35310 57650 35362 57662
rect 35310 57586 35362 57598
rect 2158 57538 2210 57550
rect 11006 57538 11058 57550
rect 3042 57486 3054 57538
rect 3106 57486 3118 57538
rect 2158 57474 2210 57486
rect 11006 57474 11058 57486
rect 18846 57538 18898 57550
rect 18846 57474 18898 57486
rect 22542 57538 22594 57550
rect 32174 57538 32226 57550
rect 25330 57486 25342 57538
rect 25394 57486 25406 57538
rect 26898 57486 26910 57538
rect 26962 57486 26974 57538
rect 28578 57486 28590 57538
rect 28642 57486 28654 57538
rect 30706 57486 30718 57538
rect 30770 57486 30782 57538
rect 22542 57474 22594 57486
rect 32174 57474 32226 57486
rect 33182 57538 33234 57550
rect 33182 57474 33234 57486
rect 33742 57538 33794 57550
rect 33742 57474 33794 57486
rect 35086 57538 35138 57550
rect 35086 57474 35138 57486
rect 38110 57538 38162 57550
rect 38434 57486 38446 57538
rect 38498 57486 38510 57538
rect 38110 57474 38162 57486
rect 6862 57426 6914 57438
rect 6862 57362 6914 57374
rect 17726 57426 17778 57438
rect 20066 57374 20078 57426
rect 20130 57374 20142 57426
rect 26338 57374 26350 57426
rect 26402 57374 26414 57426
rect 17726 57362 17778 57374
rect 1344 57258 48608 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 48608 57258
rect 1344 57172 48608 57206
rect 3166 57090 3218 57102
rect 5070 57090 5122 57102
rect 3490 57038 3502 57090
rect 3554 57038 3566 57090
rect 3166 57026 3218 57038
rect 5070 57026 5122 57038
rect 9550 57090 9602 57102
rect 9550 57026 9602 57038
rect 12126 57090 12178 57102
rect 25454 57090 25506 57102
rect 19842 57038 19854 57090
rect 19906 57038 19918 57090
rect 12126 57026 12178 57038
rect 25454 57026 25506 57038
rect 32062 57090 32114 57102
rect 32062 57026 32114 57038
rect 4958 56978 5010 56990
rect 26238 56978 26290 56990
rect 6626 56926 6638 56978
rect 6690 56926 6702 56978
rect 25778 56926 25790 56978
rect 25842 56926 25854 56978
rect 4958 56914 5010 56926
rect 26238 56914 26290 56926
rect 30718 56978 30770 56990
rect 30718 56914 30770 56926
rect 34302 56978 34354 56990
rect 34302 56914 34354 56926
rect 34526 56978 34578 56990
rect 34526 56914 34578 56926
rect 34974 56978 35026 56990
rect 41346 56926 41358 56978
rect 41410 56926 41422 56978
rect 34974 56914 35026 56926
rect 2158 56866 2210 56878
rect 2158 56802 2210 56814
rect 2606 56866 2658 56878
rect 2606 56802 2658 56814
rect 2942 56866 2994 56878
rect 2942 56802 2994 56814
rect 5854 56866 5906 56878
rect 7086 56866 7138 56878
rect 9998 56866 10050 56878
rect 22990 56866 23042 56878
rect 6514 56814 6526 56866
rect 6578 56814 6590 56866
rect 7522 56814 7534 56866
rect 7586 56814 7598 56866
rect 8306 56814 8318 56866
rect 8370 56814 8382 56866
rect 10770 56814 10782 56866
rect 10834 56814 10846 56866
rect 19394 56814 19406 56866
rect 19458 56814 19470 56866
rect 19730 56814 19742 56866
rect 19794 56814 19806 56866
rect 20290 56814 20302 56866
rect 20354 56814 20366 56866
rect 23314 56814 23326 56866
rect 23378 56814 23390 56866
rect 31042 56814 31054 56866
rect 31106 56814 31118 56866
rect 44146 56814 44158 56866
rect 44210 56814 44222 56866
rect 5854 56802 5906 56814
rect 7086 56802 7138 56814
rect 9998 56802 10050 56814
rect 22990 56802 23042 56814
rect 5966 56754 6018 56766
rect 23886 56754 23938 56766
rect 21298 56702 21310 56754
rect 21362 56702 21374 56754
rect 5966 56690 6018 56702
rect 23886 56690 23938 56702
rect 25678 56754 25730 56766
rect 25678 56690 25730 56702
rect 29822 56754 29874 56766
rect 29822 56690 29874 56702
rect 30158 56754 30210 56766
rect 30158 56690 30210 56702
rect 38446 56754 38498 56766
rect 43474 56702 43486 56754
rect 43538 56702 43550 56754
rect 38446 56690 38498 56702
rect 4286 56642 4338 56654
rect 4286 56578 4338 56590
rect 4734 56642 4786 56654
rect 4734 56578 4786 56590
rect 18174 56642 18226 56654
rect 18174 56578 18226 56590
rect 18734 56642 18786 56654
rect 38558 56642 38610 56654
rect 22306 56590 22318 56642
rect 22370 56590 22382 56642
rect 33954 56590 33966 56642
rect 34018 56590 34030 56642
rect 18734 56578 18786 56590
rect 38558 56578 38610 56590
rect 41022 56642 41074 56654
rect 41022 56578 41074 56590
rect 1344 56474 48608 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 48608 56474
rect 1344 56388 48608 56422
rect 7982 56306 8034 56318
rect 7982 56242 8034 56254
rect 9662 56306 9714 56318
rect 9662 56242 9714 56254
rect 38670 56306 38722 56318
rect 38670 56242 38722 56254
rect 41918 56306 41970 56318
rect 41918 56242 41970 56254
rect 42142 56306 42194 56318
rect 42142 56242 42194 56254
rect 33406 56194 33458 56206
rect 26002 56142 26014 56194
rect 26066 56142 26078 56194
rect 33406 56130 33458 56142
rect 33742 56194 33794 56206
rect 33742 56130 33794 56142
rect 22766 56082 22818 56094
rect 41806 56082 41858 56094
rect 6290 56030 6302 56082
rect 6354 56030 6366 56082
rect 21858 56030 21870 56082
rect 21922 56030 21934 56082
rect 22306 56030 22318 56082
rect 22370 56030 22382 56082
rect 23426 56030 23438 56082
rect 23490 56030 23502 56082
rect 25218 56030 25230 56082
rect 25282 56030 25294 56082
rect 35410 56030 35422 56082
rect 35474 56030 35486 56082
rect 22766 56018 22818 56030
rect 41806 56018 41858 56030
rect 42478 56082 42530 56094
rect 42478 56018 42530 56030
rect 20974 55970 21026 55982
rect 24782 55970 24834 55982
rect 41246 55970 41298 55982
rect 3154 55918 3166 55970
rect 3218 55918 3230 55970
rect 23090 55918 23102 55970
rect 23154 55918 23166 55970
rect 28130 55918 28142 55970
rect 28194 55918 28206 55970
rect 36082 55918 36094 55970
rect 36146 55918 36158 55970
rect 38210 55918 38222 55970
rect 38274 55918 38286 55970
rect 20974 55906 21026 55918
rect 24782 55906 24834 55918
rect 41246 55906 41298 55918
rect 20962 55806 20974 55858
rect 21026 55855 21038 55858
rect 21410 55855 21422 55858
rect 21026 55809 21422 55855
rect 21026 55806 21038 55809
rect 21410 55806 21422 55809
rect 21474 55806 21486 55858
rect 23314 55806 23326 55858
rect 23378 55806 23390 55858
rect 41234 55806 41246 55858
rect 41298 55855 41310 55858
rect 41570 55855 41582 55858
rect 41298 55809 41582 55855
rect 41298 55806 41310 55809
rect 41570 55806 41582 55809
rect 41634 55806 41646 55858
rect 1344 55690 48608 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 48608 55690
rect 1344 55604 48608 55638
rect 17054 55522 17106 55534
rect 2706 55470 2718 55522
rect 2770 55519 2782 55522
rect 3266 55519 3278 55522
rect 2770 55473 3278 55519
rect 2770 55470 2782 55473
rect 3266 55470 3278 55473
rect 3330 55470 3342 55522
rect 17054 55458 17106 55470
rect 18062 55410 18114 55422
rect 22430 55410 22482 55422
rect 42366 55410 42418 55422
rect 21298 55358 21310 55410
rect 21362 55358 21374 55410
rect 33506 55358 33518 55410
rect 33570 55358 33582 55410
rect 35634 55358 35646 55410
rect 35698 55358 35710 55410
rect 41234 55358 41246 55410
rect 41298 55358 41310 55410
rect 41906 55358 41918 55410
rect 41970 55358 41982 55410
rect 18062 55346 18114 55358
rect 22430 55346 22482 55358
rect 42366 55346 42418 55358
rect 42814 55410 42866 55422
rect 42814 55346 42866 55358
rect 1934 55298 1986 55310
rect 1934 55234 1986 55246
rect 3278 55298 3330 55310
rect 3278 55234 3330 55246
rect 4622 55298 4674 55310
rect 4622 55234 4674 55246
rect 6638 55298 6690 55310
rect 17838 55298 17890 55310
rect 7970 55246 7982 55298
rect 8034 55246 8046 55298
rect 8866 55246 8878 55298
rect 8930 55246 8942 55298
rect 19506 55246 19518 55298
rect 19570 55246 19582 55298
rect 20178 55246 20190 55298
rect 20242 55246 20254 55298
rect 20626 55246 20638 55298
rect 20690 55246 20702 55298
rect 24322 55246 24334 55298
rect 24386 55246 24398 55298
rect 24770 55246 24782 55298
rect 24834 55246 24846 55298
rect 32834 55246 32846 55298
rect 32898 55246 32910 55298
rect 38434 55246 38446 55298
rect 38498 55246 38510 55298
rect 6638 55234 6690 55246
rect 17838 55234 17890 55246
rect 3726 55186 3778 55198
rect 3726 55122 3778 55134
rect 6190 55186 6242 55198
rect 6190 55122 6242 55134
rect 16942 55186 16994 55198
rect 21422 55186 21474 55198
rect 20738 55134 20750 55186
rect 20802 55134 20814 55186
rect 16942 55122 16994 55134
rect 21422 55122 21474 55134
rect 21646 55186 21698 55198
rect 25342 55186 25394 55198
rect 41582 55186 41634 55198
rect 22754 55134 22766 55186
rect 22818 55134 22830 55186
rect 39106 55134 39118 55186
rect 39170 55134 39182 55186
rect 21646 55122 21698 55134
rect 25342 55122 25394 55134
rect 41582 55122 41634 55134
rect 41806 55186 41858 55198
rect 41806 55122 41858 55134
rect 2382 55074 2434 55086
rect 2382 55010 2434 55022
rect 2942 55074 2994 55086
rect 2942 55010 2994 55022
rect 4174 55074 4226 55086
rect 4174 55010 4226 55022
rect 5182 55074 5234 55086
rect 5182 55010 5234 55022
rect 5742 55074 5794 55086
rect 5742 55010 5794 55022
rect 5966 55074 6018 55086
rect 5966 55010 6018 55022
rect 6078 55074 6130 55086
rect 18510 55074 18562 55086
rect 32398 55074 32450 55086
rect 17490 55022 17502 55074
rect 17554 55022 17566 55074
rect 24210 55022 24222 55074
rect 24274 55022 24286 55074
rect 6078 55010 6130 55022
rect 18510 55010 18562 55022
rect 32398 55010 32450 55022
rect 42254 55074 42306 55086
rect 42254 55010 42306 55022
rect 1344 54906 48608 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 48608 54906
rect 1344 54820 48608 54854
rect 13134 54738 13186 54750
rect 13134 54674 13186 54686
rect 19518 54738 19570 54750
rect 19518 54674 19570 54686
rect 19630 54738 19682 54750
rect 19630 54674 19682 54686
rect 29710 54738 29762 54750
rect 29710 54674 29762 54686
rect 35198 54738 35250 54750
rect 35198 54674 35250 54686
rect 41022 54738 41074 54750
rect 41022 54674 41074 54686
rect 17390 54626 17442 54638
rect 24110 54626 24162 54638
rect 21298 54574 21310 54626
rect 21362 54574 21374 54626
rect 17390 54562 17442 54574
rect 24110 54562 24162 54574
rect 25342 54626 25394 54638
rect 25342 54562 25394 54574
rect 28030 54626 28082 54638
rect 28030 54562 28082 54574
rect 29262 54626 29314 54638
rect 29262 54562 29314 54574
rect 30494 54626 30546 54638
rect 30494 54562 30546 54574
rect 38334 54626 38386 54638
rect 38334 54562 38386 54574
rect 38894 54626 38946 54638
rect 42130 54574 42142 54626
rect 42194 54574 42206 54626
rect 38894 54562 38946 54574
rect 25230 54514 25282 54526
rect 1810 54462 1822 54514
rect 1874 54462 1886 54514
rect 3154 54462 3166 54514
rect 3218 54462 3230 54514
rect 3602 54462 3614 54514
rect 3666 54462 3678 54514
rect 13794 54462 13806 54514
rect 13858 54462 13870 54514
rect 17602 54462 17614 54514
rect 17666 54462 17678 54514
rect 19842 54462 19854 54514
rect 19906 54462 19918 54514
rect 20066 54462 20078 54514
rect 20130 54462 20142 54514
rect 20514 54462 20526 54514
rect 20578 54462 20590 54514
rect 25230 54450 25282 54462
rect 25566 54514 25618 54526
rect 25566 54450 25618 54462
rect 25902 54514 25954 54526
rect 25902 54450 25954 54462
rect 28926 54514 28978 54526
rect 28926 54450 28978 54462
rect 30158 54514 30210 54526
rect 30158 54450 30210 54462
rect 34862 54514 34914 54526
rect 41346 54462 41358 54514
rect 41410 54462 41422 54514
rect 34862 54450 34914 54462
rect 2494 54402 2546 54414
rect 18174 54402 18226 54414
rect 6290 54350 6302 54402
rect 6354 54350 6366 54402
rect 14466 54350 14478 54402
rect 14530 54350 14542 54402
rect 16594 54350 16606 54402
rect 16658 54350 16670 54402
rect 2494 54338 2546 54350
rect 18174 54338 18226 54350
rect 18846 54402 18898 54414
rect 18846 54338 18898 54350
rect 19294 54402 19346 54414
rect 23998 54402 24050 54414
rect 23426 54350 23438 54402
rect 23490 54350 23502 54402
rect 19294 54338 19346 54350
rect 23998 54338 24050 54350
rect 24558 54402 24610 54414
rect 24558 54338 24610 54350
rect 27806 54402 27858 54414
rect 27806 54338 27858 54350
rect 28590 54402 28642 54414
rect 28590 54338 28642 54350
rect 33294 54402 33346 54414
rect 33294 54338 33346 54350
rect 33742 54402 33794 54414
rect 33742 54338 33794 54350
rect 38670 54402 38722 54414
rect 38994 54350 39006 54402
rect 39058 54350 39070 54402
rect 44258 54350 44270 54402
rect 44322 54350 44334 54402
rect 38670 54338 38722 54350
rect 28254 54290 28306 54302
rect 28254 54226 28306 54238
rect 1344 54122 48608 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 48608 54122
rect 1344 54036 48608 54070
rect 7198 53954 7250 53966
rect 7198 53890 7250 53902
rect 29710 53954 29762 53966
rect 29710 53890 29762 53902
rect 34190 53954 34242 53966
rect 40898 53902 40910 53954
rect 40962 53902 40974 53954
rect 34190 53890 34242 53902
rect 2606 53842 2658 53854
rect 2606 53778 2658 53790
rect 2942 53842 2994 53854
rect 2942 53778 2994 53790
rect 3726 53842 3778 53854
rect 3726 53778 3778 53790
rect 6638 53842 6690 53854
rect 6638 53778 6690 53790
rect 7646 53842 7698 53854
rect 7646 53778 7698 53790
rect 9438 53842 9490 53854
rect 33854 53842 33906 53854
rect 44046 53842 44098 53854
rect 17042 53790 17054 53842
rect 17106 53790 17118 53842
rect 19170 53790 19182 53842
rect 19234 53790 19246 53842
rect 23426 53790 23438 53842
rect 23490 53790 23502 53842
rect 30930 53790 30942 53842
rect 30994 53790 31006 53842
rect 33058 53790 33070 53842
rect 33122 53790 33134 53842
rect 41122 53790 41134 53842
rect 41186 53790 41198 53842
rect 42130 53790 42142 53842
rect 42194 53790 42206 53842
rect 9438 53778 9490 53790
rect 33854 53778 33906 53790
rect 44046 53778 44098 53790
rect 1934 53730 1986 53742
rect 1934 53666 1986 53678
rect 3166 53730 3218 53742
rect 3166 53666 3218 53678
rect 3614 53730 3666 53742
rect 3614 53666 3666 53678
rect 4286 53730 4338 53742
rect 6974 53730 7026 53742
rect 4498 53678 4510 53730
rect 4562 53678 4574 53730
rect 4286 53666 4338 53678
rect 6974 53666 7026 53678
rect 12686 53730 12738 53742
rect 15934 53730 15986 53742
rect 26014 53730 26066 53742
rect 28590 53730 28642 53742
rect 14466 53678 14478 53730
rect 14530 53678 14542 53730
rect 16370 53678 16382 53730
rect 16434 53678 16446 53730
rect 23314 53678 23326 53730
rect 23378 53678 23390 53730
rect 24098 53678 24110 53730
rect 24162 53678 24174 53730
rect 26338 53678 26350 53730
rect 26402 53678 26414 53730
rect 12686 53666 12738 53678
rect 15934 53666 15986 53678
rect 26014 53666 26066 53678
rect 28590 53666 28642 53678
rect 29374 53730 29426 53742
rect 33630 53730 33682 53742
rect 30146 53678 30158 53730
rect 30210 53678 30222 53730
rect 41010 53678 41022 53730
rect 41074 53678 41086 53730
rect 41682 53678 41694 53730
rect 41746 53678 41758 53730
rect 42242 53678 42254 53730
rect 42306 53678 42318 53730
rect 29374 53666 29426 53678
rect 33630 53666 33682 53678
rect 5630 53618 5682 53630
rect 5630 53554 5682 53566
rect 6526 53618 6578 53630
rect 6526 53554 6578 53566
rect 7982 53618 8034 53630
rect 7982 53554 8034 53566
rect 8542 53618 8594 53630
rect 15038 53618 15090 53630
rect 13570 53566 13582 53618
rect 13634 53566 13646 53618
rect 8542 53554 8594 53566
rect 15038 53554 15090 53566
rect 15374 53618 15426 53630
rect 26910 53618 26962 53630
rect 23202 53566 23214 53618
rect 23266 53566 23278 53618
rect 24434 53566 24446 53618
rect 24498 53566 24510 53618
rect 15374 53554 15426 53566
rect 26910 53554 26962 53566
rect 29150 53618 29202 53630
rect 29150 53554 29202 53566
rect 35982 53618 36034 53630
rect 35982 53554 36034 53566
rect 38558 53618 38610 53630
rect 38558 53554 38610 53566
rect 2046 53506 2098 53518
rect 2046 53442 2098 53454
rect 2494 53506 2546 53518
rect 2494 53442 2546 53454
rect 2718 53506 2770 53518
rect 2718 53442 2770 53454
rect 3838 53506 3890 53518
rect 3838 53442 3890 53454
rect 4846 53506 4898 53518
rect 4846 53442 4898 53454
rect 4958 53506 5010 53518
rect 4958 53442 5010 53454
rect 5070 53506 5122 53518
rect 5070 53442 5122 53454
rect 5742 53506 5794 53518
rect 5742 53442 5794 53454
rect 5966 53506 6018 53518
rect 5966 53442 6018 53454
rect 6750 53506 6802 53518
rect 6750 53442 6802 53454
rect 7534 53506 7586 53518
rect 7534 53442 7586 53454
rect 7758 53506 7810 53518
rect 7758 53442 7810 53454
rect 8430 53506 8482 53518
rect 8430 53442 8482 53454
rect 8990 53506 9042 53518
rect 8990 53442 9042 53454
rect 12126 53506 12178 53518
rect 12126 53442 12178 53454
rect 12350 53506 12402 53518
rect 12350 53442 12402 53454
rect 12574 53506 12626 53518
rect 12574 53442 12626 53454
rect 20302 53506 20354 53518
rect 34638 53506 34690 53518
rect 25330 53454 25342 53506
rect 25394 53454 25406 53506
rect 20302 53442 20354 53454
rect 34638 53442 34690 53454
rect 36318 53506 36370 53518
rect 36318 53442 36370 53454
rect 38670 53506 38722 53518
rect 38670 53442 38722 53454
rect 40238 53506 40290 53518
rect 40238 53442 40290 53454
rect 43150 53506 43202 53518
rect 43150 53442 43202 53454
rect 43934 53506 43986 53518
rect 43934 53442 43986 53454
rect 1344 53338 48608 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 48608 53338
rect 1344 53252 48608 53286
rect 4174 53170 4226 53182
rect 3266 53118 3278 53170
rect 3330 53118 3342 53170
rect 4174 53106 4226 53118
rect 5182 53170 5234 53182
rect 5182 53106 5234 53118
rect 8430 53170 8482 53182
rect 8430 53106 8482 53118
rect 8878 53170 8930 53182
rect 8878 53106 8930 53118
rect 22766 53170 22818 53182
rect 22766 53106 22818 53118
rect 23998 53170 24050 53182
rect 23998 53106 24050 53118
rect 24110 53170 24162 53182
rect 38894 53170 38946 53182
rect 32386 53118 32398 53170
rect 32450 53118 32462 53170
rect 24110 53106 24162 53118
rect 38894 53106 38946 53118
rect 42366 53170 42418 53182
rect 42366 53106 42418 53118
rect 42814 53170 42866 53182
rect 42814 53106 42866 53118
rect 3726 53058 3778 53070
rect 3726 52994 3778 53006
rect 4286 53058 4338 53070
rect 4286 52994 4338 53006
rect 4510 53058 4562 53070
rect 20638 53058 20690 53070
rect 6178 53006 6190 53058
rect 6242 53006 6254 53058
rect 11890 53006 11902 53058
rect 11954 53006 11966 53058
rect 4510 52994 4562 53006
rect 20638 52994 20690 53006
rect 23214 53058 23266 53070
rect 26002 53006 26014 53058
rect 26066 53006 26078 53058
rect 29250 53006 29262 53058
rect 29314 53006 29326 53058
rect 36306 53006 36318 53058
rect 36370 53006 36382 53058
rect 23214 52994 23266 53006
rect 4062 52946 4114 52958
rect 2930 52894 2942 52946
rect 2994 52894 3006 52946
rect 3490 52894 3502 52946
rect 3554 52894 3566 52946
rect 4062 52882 4114 52894
rect 5406 52946 5458 52958
rect 19406 52946 19458 52958
rect 20302 52946 20354 52958
rect 5506 52894 5518 52946
rect 5570 52894 5582 52946
rect 6738 52894 6750 52946
rect 6802 52894 6814 52946
rect 7522 52894 7534 52946
rect 7586 52894 7598 52946
rect 11106 52894 11118 52946
rect 11170 52894 11182 52946
rect 19954 52894 19966 52946
rect 20018 52894 20030 52946
rect 5406 52882 5458 52894
rect 19406 52882 19458 52894
rect 20302 52882 20354 52894
rect 23438 52946 23490 52958
rect 33630 52946 33682 52958
rect 23762 52894 23774 52946
rect 23826 52894 23838 52946
rect 25218 52894 25230 52946
rect 25282 52894 25294 52946
rect 28578 52894 28590 52946
rect 28642 52894 28654 52946
rect 35522 52894 35534 52946
rect 35586 52894 35598 52946
rect 43138 52894 43150 52946
rect 43202 52894 43214 52946
rect 23438 52882 23490 52894
rect 33630 52882 33682 52894
rect 2270 52834 2322 52846
rect 2270 52770 2322 52782
rect 2606 52834 2658 52846
rect 2606 52770 2658 52782
rect 3278 52834 3330 52846
rect 3278 52770 3330 52782
rect 5294 52834 5346 52846
rect 5294 52770 5346 52782
rect 6414 52834 6466 52846
rect 6414 52770 6466 52782
rect 8094 52834 8146 52846
rect 14478 52834 14530 52846
rect 14018 52782 14030 52834
rect 14082 52782 14094 52834
rect 8094 52770 8146 52782
rect 14478 52770 14530 52782
rect 14926 52834 14978 52846
rect 14926 52770 14978 52782
rect 19070 52834 19122 52846
rect 19070 52770 19122 52782
rect 24670 52834 24722 52846
rect 31838 52834 31890 52846
rect 28130 52782 28142 52834
rect 28194 52782 28206 52834
rect 31378 52782 31390 52834
rect 31442 52782 31454 52834
rect 24670 52770 24722 52782
rect 31838 52770 31890 52782
rect 33182 52834 33234 52846
rect 41022 52834 41074 52846
rect 38434 52782 38446 52834
rect 38498 52782 38510 52834
rect 33182 52770 33234 52782
rect 41022 52770 41074 52782
rect 41470 52834 41522 52846
rect 43922 52782 43934 52834
rect 43986 52782 43998 52834
rect 46050 52782 46062 52834
rect 46114 52782 46126 52834
rect 41470 52770 41522 52782
rect 5854 52722 5906 52734
rect 2146 52670 2158 52722
rect 2210 52719 2222 52722
rect 2706 52719 2718 52722
rect 2210 52673 2718 52719
rect 2210 52670 2222 52673
rect 2706 52670 2718 52673
rect 2770 52670 2782 52722
rect 5854 52658 5906 52670
rect 19630 52722 19682 52734
rect 32062 52722 32114 52734
rect 22642 52670 22654 52722
rect 22706 52719 22718 52722
rect 23090 52719 23102 52722
rect 22706 52673 23102 52719
rect 22706 52670 22718 52673
rect 23090 52670 23102 52673
rect 23154 52670 23166 52722
rect 19630 52658 19682 52670
rect 32062 52658 32114 52670
rect 1344 52554 48608 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 48608 52554
rect 1344 52468 48608 52502
rect 4734 52386 4786 52398
rect 4050 52334 4062 52386
rect 4114 52334 4126 52386
rect 4734 52322 4786 52334
rect 22654 52386 22706 52398
rect 22654 52322 22706 52334
rect 35646 52386 35698 52398
rect 37326 52386 37378 52398
rect 43598 52386 43650 52398
rect 35970 52334 35982 52386
rect 36034 52334 36046 52386
rect 39666 52334 39678 52386
rect 39730 52334 39742 52386
rect 42466 52334 42478 52386
rect 42530 52334 42542 52386
rect 35646 52322 35698 52334
rect 37326 52322 37378 52334
rect 43598 52322 43650 52334
rect 43934 52386 43986 52398
rect 43934 52322 43986 52334
rect 3166 52274 3218 52286
rect 23214 52274 23266 52286
rect 7634 52222 7646 52274
rect 7698 52222 7710 52274
rect 3166 52210 3218 52222
rect 23214 52210 23266 52222
rect 30718 52274 30770 52286
rect 30718 52210 30770 52222
rect 36430 52274 36482 52286
rect 45054 52274 45106 52286
rect 38210 52222 38222 52274
rect 38274 52222 38286 52274
rect 42130 52222 42142 52274
rect 42194 52222 42206 52274
rect 36430 52210 36482 52222
rect 45054 52210 45106 52222
rect 45166 52274 45218 52286
rect 45166 52210 45218 52222
rect 2270 52162 2322 52174
rect 2270 52098 2322 52110
rect 3502 52162 3554 52174
rect 3502 52098 3554 52110
rect 3726 52162 3778 52174
rect 12014 52162 12066 52174
rect 6290 52110 6302 52162
rect 6354 52110 6366 52162
rect 3726 52098 3778 52110
rect 12014 52098 12066 52110
rect 33518 52162 33570 52174
rect 33518 52098 33570 52110
rect 35086 52162 35138 52174
rect 35086 52098 35138 52110
rect 35422 52162 35474 52174
rect 40238 52162 40290 52174
rect 41694 52162 41746 52174
rect 37650 52110 37662 52162
rect 37714 52110 37726 52162
rect 38322 52110 38334 52162
rect 38386 52110 38398 52162
rect 39218 52110 39230 52162
rect 39282 52110 39294 52162
rect 39554 52110 39566 52162
rect 39618 52110 39630 52162
rect 41122 52110 41134 52162
rect 41186 52110 41198 52162
rect 42018 52110 42030 52162
rect 42082 52110 42094 52162
rect 42354 52110 42366 52162
rect 42418 52110 42430 52162
rect 43922 52110 43934 52162
rect 43986 52110 43998 52162
rect 35422 52098 35474 52110
rect 40238 52098 40290 52110
rect 41694 52098 41746 52110
rect 4398 52050 4450 52062
rect 4398 51986 4450 51998
rect 11230 52050 11282 52062
rect 11230 51986 11282 51998
rect 22766 52050 22818 52062
rect 22766 51986 22818 51998
rect 32734 52050 32786 52062
rect 32734 51986 32786 51998
rect 2718 51938 2770 51950
rect 2718 51874 2770 51886
rect 4622 51938 4674 51950
rect 4622 51874 4674 51886
rect 11342 51938 11394 51950
rect 11342 51874 11394 51886
rect 11566 51938 11618 51950
rect 11566 51874 11618 51886
rect 31166 51938 31218 51950
rect 31166 51874 31218 51886
rect 31838 51938 31890 51950
rect 31838 51874 31890 51886
rect 32286 51938 32338 51950
rect 32286 51874 32338 51886
rect 34526 51938 34578 51950
rect 34526 51874 34578 51886
rect 37438 51938 37490 51950
rect 37438 51874 37490 51886
rect 1344 51770 48608 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 48608 51770
rect 1344 51684 48608 51718
rect 29822 51602 29874 51614
rect 29822 51538 29874 51550
rect 30718 51602 30770 51614
rect 30718 51538 30770 51550
rect 39902 51602 39954 51614
rect 39902 51538 39954 51550
rect 40350 51602 40402 51614
rect 40350 51538 40402 51550
rect 43710 51602 43762 51614
rect 43710 51538 43762 51550
rect 44158 51602 44210 51614
rect 44158 51538 44210 51550
rect 14702 51490 14754 51502
rect 26574 51490 26626 51502
rect 6962 51438 6974 51490
rect 7026 51438 7038 51490
rect 10322 51438 10334 51490
rect 10386 51438 10398 51490
rect 20626 51438 20638 51490
rect 20690 51438 20702 51490
rect 38658 51438 38670 51490
rect 38722 51438 38734 51490
rect 14702 51426 14754 51438
rect 26574 51426 26626 51438
rect 4510 51378 4562 51390
rect 6302 51378 6354 51390
rect 14366 51378 14418 51390
rect 4834 51326 4846 51378
rect 4898 51326 4910 51378
rect 6738 51326 6750 51378
rect 6802 51326 6814 51378
rect 7298 51326 7310 51378
rect 7362 51326 7374 51378
rect 7634 51326 7646 51378
rect 7698 51326 7710 51378
rect 9650 51326 9662 51378
rect 9714 51326 9726 51378
rect 12786 51326 12798 51378
rect 12850 51326 12862 51378
rect 4510 51314 4562 51326
rect 6302 51314 6354 51326
rect 14366 51314 14418 51326
rect 19518 51378 19570 51390
rect 23438 51378 23490 51390
rect 19842 51326 19854 51378
rect 19906 51326 19918 51378
rect 19518 51314 19570 51326
rect 23438 51314 23490 51326
rect 23662 51378 23714 51390
rect 41134 51378 41186 51390
rect 42142 51378 42194 51390
rect 26786 51326 26798 51378
rect 26850 51326 26862 51378
rect 33058 51326 33070 51378
rect 33122 51326 33134 51378
rect 39442 51326 39454 51378
rect 39506 51326 39518 51378
rect 41346 51326 41358 51378
rect 41410 51326 41422 51378
rect 42242 51326 42254 51378
rect 42306 51326 42318 51378
rect 42802 51326 42814 51378
rect 42866 51326 42878 51378
rect 23662 51314 23714 51326
rect 41134 51314 41186 51326
rect 42142 51314 42194 51326
rect 3278 51266 3330 51278
rect 3278 51202 3330 51214
rect 3726 51266 3778 51278
rect 3726 51202 3778 51214
rect 4174 51266 4226 51278
rect 4174 51202 4226 51214
rect 8542 51266 8594 51278
rect 30270 51266 30322 51278
rect 12450 51214 12462 51266
rect 12514 51214 12526 51266
rect 13458 51214 13470 51266
rect 13522 51214 13534 51266
rect 22754 51214 22766 51266
rect 22818 51214 22830 51266
rect 8542 51202 8594 51214
rect 30270 51202 30322 51214
rect 31390 51266 31442 51278
rect 31390 51202 31442 51214
rect 31838 51266 31890 51278
rect 31838 51202 31890 51214
rect 32286 51266 32338 51278
rect 33842 51214 33854 51266
rect 33906 51214 33918 51266
rect 35970 51214 35982 51266
rect 36034 51214 36046 51266
rect 36530 51214 36542 51266
rect 36594 51214 36606 51266
rect 32286 51202 32338 51214
rect 23090 51102 23102 51154
rect 23154 51102 23166 51154
rect 30594 51102 30606 51154
rect 30658 51151 30670 51154
rect 31378 51151 31390 51154
rect 30658 51105 31390 51151
rect 30658 51102 30670 51105
rect 31378 51102 31390 51105
rect 31442 51102 31454 51154
rect 42690 51102 42702 51154
rect 42754 51102 42766 51154
rect 1344 50986 48608 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 48608 50986
rect 1344 50900 48608 50934
rect 27582 50818 27634 50830
rect 3714 50766 3726 50818
rect 3778 50766 3790 50818
rect 13906 50766 13918 50818
rect 13970 50766 13982 50818
rect 27582 50754 27634 50766
rect 33854 50818 33906 50830
rect 33854 50754 33906 50766
rect 34190 50818 34242 50830
rect 37090 50766 37102 50818
rect 37154 50815 37166 50818
rect 37314 50815 37326 50818
rect 37154 50769 37326 50815
rect 37154 50766 37166 50769
rect 37314 50766 37326 50769
rect 37378 50766 37390 50818
rect 34190 50754 34242 50766
rect 10782 50706 10834 50718
rect 10782 50642 10834 50654
rect 11454 50706 11506 50718
rect 11454 50642 11506 50654
rect 12686 50706 12738 50718
rect 12686 50642 12738 50654
rect 14478 50706 14530 50718
rect 27246 50706 27298 50718
rect 15810 50654 15822 50706
rect 15874 50654 15886 50706
rect 17938 50654 17950 50706
rect 18002 50654 18014 50706
rect 25778 50654 25790 50706
rect 25842 50654 25854 50706
rect 14478 50642 14530 50654
rect 27246 50642 27298 50654
rect 27806 50706 27858 50718
rect 27806 50642 27858 50654
rect 28254 50706 28306 50718
rect 32734 50706 32786 50718
rect 29474 50654 29486 50706
rect 29538 50654 29550 50706
rect 28254 50642 28306 50654
rect 32734 50642 32786 50654
rect 33294 50706 33346 50718
rect 33294 50642 33346 50654
rect 35758 50706 35810 50718
rect 35758 50642 35810 50654
rect 37102 50706 37154 50718
rect 37102 50642 37154 50654
rect 37662 50706 37714 50718
rect 37662 50642 37714 50654
rect 42030 50706 42082 50718
rect 42030 50642 42082 50654
rect 3950 50594 4002 50606
rect 3950 50530 4002 50542
rect 4398 50594 4450 50606
rect 4398 50530 4450 50542
rect 4846 50594 4898 50606
rect 4846 50530 4898 50542
rect 7310 50594 7362 50606
rect 14254 50594 14306 50606
rect 22542 50594 22594 50606
rect 32398 50594 32450 50606
rect 7858 50542 7870 50594
rect 7922 50542 7934 50594
rect 18722 50542 18734 50594
rect 18786 50542 18798 50594
rect 22978 50542 22990 50594
rect 23042 50542 23054 50594
rect 29698 50542 29710 50594
rect 29762 50542 29774 50594
rect 30482 50542 30494 50594
rect 30546 50542 30558 50594
rect 7310 50530 7362 50542
rect 14254 50530 14306 50542
rect 22542 50530 22594 50542
rect 32398 50530 32450 50542
rect 34750 50594 34802 50606
rect 34750 50530 34802 50542
rect 34862 50594 34914 50606
rect 34862 50530 34914 50542
rect 35086 50594 35138 50606
rect 36206 50594 36258 50606
rect 35298 50542 35310 50594
rect 35362 50542 35374 50594
rect 35086 50530 35138 50542
rect 36206 50530 36258 50542
rect 26238 50482 26290 50494
rect 8642 50430 8654 50482
rect 8706 50430 8718 50482
rect 23650 50430 23662 50482
rect 23714 50430 23726 50482
rect 26238 50418 26290 50430
rect 26910 50482 26962 50494
rect 31502 50482 31554 50494
rect 29362 50430 29374 50482
rect 29426 50430 29438 50482
rect 26910 50418 26962 50430
rect 31502 50418 31554 50430
rect 33966 50482 34018 50494
rect 33966 50418 34018 50430
rect 41358 50482 41410 50494
rect 41358 50418 41410 50430
rect 6078 50370 6130 50382
rect 6078 50306 6130 50318
rect 14926 50370 14978 50382
rect 14926 50306 14978 50318
rect 15486 50370 15538 50382
rect 15486 50306 15538 50318
rect 26574 50370 26626 50382
rect 26574 50306 26626 50318
rect 30382 50370 30434 50382
rect 30382 50306 30434 50318
rect 34974 50370 35026 50382
rect 34974 50306 35026 50318
rect 1344 50202 48608 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 48608 50202
rect 1344 50116 48608 50150
rect 23662 50034 23714 50046
rect 23662 49970 23714 49982
rect 24110 50034 24162 50046
rect 24110 49970 24162 49982
rect 25342 50034 25394 50046
rect 31054 50034 31106 50046
rect 29698 49982 29710 50034
rect 29762 49982 29774 50034
rect 25342 49970 25394 49982
rect 31054 49970 31106 49982
rect 31166 50034 31218 50046
rect 31166 49970 31218 49982
rect 10670 49922 10722 49934
rect 23326 49922 23378 49934
rect 31278 49922 31330 49934
rect 42030 49922 42082 49934
rect 14914 49870 14926 49922
rect 14978 49870 14990 49922
rect 19282 49870 19294 49922
rect 19346 49870 19358 49922
rect 26450 49870 26462 49922
rect 26514 49870 26526 49922
rect 33954 49870 33966 49922
rect 34018 49870 34030 49922
rect 10670 49858 10722 49870
rect 23326 49858 23378 49870
rect 31278 49858 31330 49870
rect 42030 49858 42082 49870
rect 5294 49810 5346 49822
rect 29710 49810 29762 49822
rect 31390 49810 31442 49822
rect 1810 49758 1822 49810
rect 1874 49758 1886 49810
rect 6850 49758 6862 49810
rect 6914 49758 6926 49810
rect 7298 49758 7310 49810
rect 7362 49758 7374 49810
rect 8418 49758 8430 49810
rect 8482 49758 8494 49810
rect 9762 49758 9774 49810
rect 9826 49758 9838 49810
rect 15586 49758 15598 49810
rect 15650 49758 15662 49810
rect 19618 49758 19630 49810
rect 19682 49758 19694 49810
rect 20626 49758 20638 49810
rect 20690 49758 20702 49810
rect 25666 49758 25678 49810
rect 25730 49758 25742 49810
rect 29810 49758 29822 49810
rect 29874 49758 29886 49810
rect 30818 49758 30830 49810
rect 30882 49758 30894 49810
rect 33058 49758 33070 49810
rect 33122 49758 33134 49810
rect 34738 49758 34750 49810
rect 34802 49758 34814 49810
rect 41682 49758 41694 49810
rect 41746 49758 41758 49810
rect 42354 49758 42366 49810
rect 42418 49758 42430 49810
rect 5294 49746 5346 49758
rect 29710 49746 29762 49758
rect 31390 49746 31442 49758
rect 4622 49698 4674 49710
rect 11118 49698 11170 49710
rect 16158 49698 16210 49710
rect 21086 49698 21138 49710
rect 2482 49646 2494 49698
rect 2546 49646 2558 49698
rect 9986 49646 9998 49698
rect 10050 49646 10062 49698
rect 12786 49646 12798 49698
rect 12850 49646 12862 49698
rect 20066 49646 20078 49698
rect 20130 49646 20142 49698
rect 20626 49646 20638 49698
rect 20690 49695 20702 49698
rect 20690 49649 20911 49695
rect 20690 49646 20702 49649
rect 4622 49634 4674 49646
rect 11118 49634 11170 49646
rect 16158 49634 16210 49646
rect 7746 49534 7758 49586
rect 7810 49534 7822 49586
rect 20865 49583 20911 49649
rect 21086 49634 21138 49646
rect 21534 49698 21586 49710
rect 21534 49634 21586 49646
rect 23102 49698 23154 49710
rect 31950 49698 32002 49710
rect 28578 49646 28590 49698
rect 28642 49646 28654 49698
rect 30146 49646 30158 49698
rect 30210 49646 30222 49698
rect 23102 49634 23154 49646
rect 31950 49634 32002 49646
rect 32398 49698 32450 49710
rect 36206 49698 36258 49710
rect 34066 49646 34078 49698
rect 34130 49646 34142 49698
rect 32398 49634 32450 49646
rect 36206 49634 36258 49646
rect 36542 49698 36594 49710
rect 36542 49634 36594 49646
rect 41134 49698 41186 49710
rect 41134 49634 41186 49646
rect 41918 49698 41970 49710
rect 43138 49646 43150 49698
rect 43202 49646 43214 49698
rect 45266 49646 45278 49698
rect 45330 49646 45342 49698
rect 41918 49634 41970 49646
rect 21186 49583 21198 49586
rect 20865 49537 21198 49583
rect 21186 49534 21198 49537
rect 21250 49534 21262 49586
rect 1344 49418 48608 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 48608 49418
rect 1344 49332 48608 49366
rect 21198 49250 21250 49262
rect 5954 49198 5966 49250
rect 6018 49198 6030 49250
rect 21198 49186 21250 49198
rect 27694 49250 27746 49262
rect 27694 49186 27746 49198
rect 28030 49250 28082 49262
rect 34414 49250 34466 49262
rect 29810 49198 29822 49250
rect 29874 49198 29886 49250
rect 28030 49186 28082 49198
rect 34414 49186 34466 49198
rect 35758 49250 35810 49262
rect 42242 49198 42254 49250
rect 42306 49247 42318 49250
rect 43026 49247 43038 49250
rect 42306 49201 43038 49247
rect 42306 49198 42318 49201
rect 43026 49198 43038 49201
rect 43090 49198 43102 49250
rect 35758 49186 35810 49198
rect 2606 49138 2658 49150
rect 7982 49138 8034 49150
rect 4498 49086 4510 49138
rect 4562 49086 4574 49138
rect 6402 49086 6414 49138
rect 6466 49086 6478 49138
rect 2606 49074 2658 49086
rect 7982 49074 8034 49086
rect 8990 49138 9042 49150
rect 8990 49074 9042 49086
rect 14926 49138 14978 49150
rect 18734 49138 18786 49150
rect 28254 49138 28306 49150
rect 18386 49086 18398 49138
rect 18450 49086 18462 49138
rect 20178 49086 20190 49138
rect 20242 49086 20254 49138
rect 25778 49086 25790 49138
rect 25842 49086 25854 49138
rect 14926 49074 14978 49086
rect 18734 49074 18786 49086
rect 28254 49074 28306 49086
rect 29262 49138 29314 49150
rect 29262 49074 29314 49086
rect 31054 49138 31106 49150
rect 41582 49138 41634 49150
rect 41122 49086 41134 49138
rect 41186 49086 41198 49138
rect 31054 49074 31106 49086
rect 41582 49074 41634 49086
rect 42590 49138 42642 49150
rect 42590 49074 42642 49086
rect 43038 49138 43090 49150
rect 43038 49074 43090 49086
rect 44942 49138 44994 49150
rect 44942 49074 44994 49086
rect 2718 49026 2770 49038
rect 2718 48962 2770 48974
rect 3278 49026 3330 49038
rect 8206 49026 8258 49038
rect 3938 48974 3950 49026
rect 4002 48974 4014 49026
rect 6290 48974 6302 49026
rect 6354 48974 6366 49026
rect 6850 48974 6862 49026
rect 6914 48974 6926 49026
rect 3278 48962 3330 48974
rect 8206 48962 8258 48974
rect 14702 49026 14754 49038
rect 21310 49026 21362 49038
rect 15474 48974 15486 49026
rect 15538 48974 15550 49026
rect 19506 48974 19518 49026
rect 19570 48974 19582 49026
rect 20066 48974 20078 49026
rect 20130 48974 20142 49026
rect 21858 48974 21870 49026
rect 21922 48974 21934 49026
rect 22530 48974 22542 49026
rect 22594 48974 22606 49026
rect 24434 48974 24446 49026
rect 24498 48974 24510 49026
rect 27346 48974 27358 49026
rect 27410 48974 27422 49026
rect 32386 48974 32398 49026
rect 32450 48974 32462 49026
rect 33730 48974 33742 49026
rect 33794 48974 33806 49026
rect 38322 48974 38334 49026
rect 38386 48974 38398 49026
rect 14702 48962 14754 48974
rect 21310 48962 21362 48974
rect 1934 48914 1986 48926
rect 1934 48850 1986 48862
rect 2270 48914 2322 48926
rect 2270 48850 2322 48862
rect 7422 48914 7474 48926
rect 7422 48850 7474 48862
rect 7646 48914 7698 48926
rect 30270 48914 30322 48926
rect 8530 48862 8542 48914
rect 8594 48862 8606 48914
rect 16258 48862 16270 48914
rect 16322 48862 16334 48914
rect 20738 48862 20750 48914
rect 20802 48862 20814 48914
rect 22642 48862 22654 48914
rect 22706 48862 22718 48914
rect 24994 48862 25006 48914
rect 25058 48862 25070 48914
rect 25666 48862 25678 48914
rect 25730 48862 25742 48914
rect 7646 48850 7698 48862
rect 30270 48850 30322 48862
rect 30382 48914 30434 48926
rect 30382 48850 30434 48862
rect 30494 48914 30546 48926
rect 35870 48914 35922 48926
rect 32946 48862 32958 48914
rect 33010 48862 33022 48914
rect 33842 48862 33854 48914
rect 33906 48862 33918 48914
rect 38994 48862 39006 48914
rect 39058 48862 39070 48914
rect 30494 48850 30546 48862
rect 35870 48850 35922 48862
rect 2494 48802 2546 48814
rect 2494 48738 2546 48750
rect 3054 48802 3106 48814
rect 3054 48738 3106 48750
rect 3166 48802 3218 48814
rect 3166 48738 3218 48750
rect 3502 48802 3554 48814
rect 3502 48738 3554 48750
rect 7534 48802 7586 48814
rect 7534 48738 7586 48750
rect 8878 48802 8930 48814
rect 8878 48738 8930 48750
rect 9102 48802 9154 48814
rect 9102 48738 9154 48750
rect 9326 48802 9378 48814
rect 9326 48738 9378 48750
rect 9886 48802 9938 48814
rect 9886 48738 9938 48750
rect 10334 48802 10386 48814
rect 10334 48738 10386 48750
rect 14030 48802 14082 48814
rect 18846 48802 18898 48814
rect 14354 48750 14366 48802
rect 14418 48750 14430 48802
rect 14030 48738 14082 48750
rect 18846 48738 18898 48750
rect 23326 48802 23378 48814
rect 23326 48738 23378 48750
rect 23886 48802 23938 48814
rect 23886 48738 23938 48750
rect 31502 48802 31554 48814
rect 31502 48738 31554 48750
rect 36318 48802 36370 48814
rect 36318 48738 36370 48750
rect 37102 48802 37154 48814
rect 37102 48738 37154 48750
rect 41694 48802 41746 48814
rect 41694 48738 41746 48750
rect 42142 48802 42194 48814
rect 42142 48738 42194 48750
rect 44830 48802 44882 48814
rect 44830 48738 44882 48750
rect 1344 48634 48608 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 48608 48634
rect 1344 48548 48608 48582
rect 2830 48466 2882 48478
rect 2830 48402 2882 48414
rect 15150 48466 15202 48478
rect 15150 48402 15202 48414
rect 16158 48466 16210 48478
rect 16158 48402 16210 48414
rect 16382 48466 16434 48478
rect 16382 48402 16434 48414
rect 24222 48466 24274 48478
rect 24222 48402 24274 48414
rect 37662 48466 37714 48478
rect 37662 48402 37714 48414
rect 40126 48466 40178 48478
rect 40126 48402 40178 48414
rect 42926 48466 42978 48478
rect 42926 48402 42978 48414
rect 9662 48354 9714 48366
rect 3042 48351 3054 48354
rect 2945 48305 3054 48351
rect 1934 48130 1986 48142
rect 1934 48066 1986 48078
rect 2382 48130 2434 48142
rect 2382 48066 2434 48078
rect 1922 47966 1934 48018
rect 1986 48015 1998 48018
rect 2945 48015 2991 48305
rect 3042 48302 3054 48305
rect 3106 48302 3118 48354
rect 9662 48290 9714 48302
rect 14142 48354 14194 48366
rect 14142 48290 14194 48302
rect 16606 48354 16658 48366
rect 16606 48290 16658 48302
rect 16718 48354 16770 48366
rect 36766 48354 36818 48366
rect 18834 48302 18846 48354
rect 18898 48302 18910 48354
rect 26786 48302 26798 48354
rect 26850 48302 26862 48354
rect 27570 48302 27582 48354
rect 27634 48302 27646 48354
rect 16718 48290 16770 48302
rect 36766 48290 36818 48302
rect 38782 48354 38834 48366
rect 41234 48302 41246 48354
rect 41298 48302 41310 48354
rect 38782 48290 38834 48302
rect 13806 48242 13858 48254
rect 18622 48242 18674 48254
rect 20302 48242 20354 48254
rect 36430 48242 36482 48254
rect 7858 48190 7870 48242
rect 7922 48190 7934 48242
rect 13234 48190 13246 48242
rect 13298 48190 13310 48242
rect 14354 48190 14366 48242
rect 14418 48190 14430 48242
rect 18946 48190 18958 48242
rect 19010 48190 19022 48242
rect 19730 48190 19742 48242
rect 19794 48190 19806 48242
rect 20626 48190 20638 48242
rect 20690 48190 20702 48242
rect 25218 48190 25230 48242
rect 25282 48190 25294 48242
rect 28354 48190 28366 48242
rect 28418 48190 28430 48242
rect 32498 48190 32510 48242
rect 32562 48190 32574 48242
rect 33058 48190 33070 48242
rect 33122 48190 33134 48242
rect 13806 48178 13858 48190
rect 18622 48178 18674 48190
rect 20302 48178 20354 48190
rect 36430 48178 36482 48190
rect 41022 48242 41074 48254
rect 41570 48190 41582 48242
rect 41634 48190 41646 48242
rect 42242 48190 42254 48242
rect 42306 48190 42318 48242
rect 41022 48178 41074 48190
rect 8990 48130 9042 48142
rect 3826 48078 3838 48130
rect 3890 48078 3902 48130
rect 8990 48066 9042 48078
rect 10446 48130 10498 48142
rect 18062 48130 18114 48142
rect 24670 48130 24722 48142
rect 28926 48130 28978 48142
rect 12562 48078 12574 48130
rect 12626 48078 12638 48130
rect 21410 48078 21422 48130
rect 21474 48078 21486 48130
rect 23538 48078 23550 48130
rect 23602 48078 23614 48130
rect 26114 48078 26126 48130
rect 26178 48078 26190 48130
rect 10446 48066 10498 48078
rect 18062 48066 18114 48078
rect 24670 48066 24722 48078
rect 28926 48066 28978 48078
rect 29598 48130 29650 48142
rect 37214 48130 37266 48142
rect 31378 48078 31390 48130
rect 31442 48078 31454 48130
rect 33842 48078 33854 48130
rect 33906 48078 33918 48130
rect 35970 48078 35982 48130
rect 36034 48078 36046 48130
rect 29598 48066 29650 48078
rect 37214 48066 37266 48078
rect 38222 48130 38274 48142
rect 39342 48130 39394 48142
rect 38882 48078 38894 48130
rect 38946 48078 38958 48130
rect 38222 48066 38274 48078
rect 39342 48066 39394 48078
rect 43374 48130 43426 48142
rect 43374 48066 43426 48078
rect 38558 48018 38610 48030
rect 1986 47969 2991 48015
rect 1986 47966 1998 47969
rect 13570 47966 13582 48018
rect 13634 48015 13646 48018
rect 13906 48015 13918 48018
rect 13634 47969 13918 48015
rect 13634 47966 13646 47969
rect 13906 47966 13918 47969
rect 13970 47966 13982 48018
rect 19506 47966 19518 48018
rect 19570 47966 19582 48018
rect 36978 47966 36990 48018
rect 37042 48015 37054 48018
rect 38210 48015 38222 48018
rect 37042 47969 38222 48015
rect 37042 47966 37054 47969
rect 38210 47966 38222 47969
rect 38274 47966 38286 48018
rect 38558 47954 38610 47966
rect 40910 48018 40962 48030
rect 40910 47954 40962 47966
rect 1344 47850 48608 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 48608 47850
rect 1344 47764 48608 47798
rect 2942 47682 2994 47694
rect 6738 47630 6750 47682
rect 6802 47630 6814 47682
rect 36418 47630 36430 47682
rect 36482 47630 36494 47682
rect 2942 47618 2994 47630
rect 2718 47570 2770 47582
rect 23998 47570 24050 47582
rect 29598 47570 29650 47582
rect 4162 47518 4174 47570
rect 4226 47518 4238 47570
rect 6178 47518 6190 47570
rect 6242 47518 6254 47570
rect 14242 47518 14254 47570
rect 14306 47518 14318 47570
rect 16370 47518 16382 47570
rect 16434 47518 16446 47570
rect 26674 47518 26686 47570
rect 26738 47518 26750 47570
rect 2718 47506 2770 47518
rect 23998 47506 24050 47518
rect 29598 47506 29650 47518
rect 29822 47570 29874 47582
rect 40350 47570 40402 47582
rect 42702 47570 42754 47582
rect 33170 47518 33182 47570
rect 33234 47518 33246 47570
rect 37762 47518 37774 47570
rect 37826 47518 37838 47570
rect 39890 47518 39902 47570
rect 39954 47518 39966 47570
rect 41122 47518 41134 47570
rect 41186 47518 41198 47570
rect 41458 47518 41470 47570
rect 41522 47518 41534 47570
rect 29822 47506 29874 47518
rect 40350 47506 40402 47518
rect 42702 47506 42754 47518
rect 42926 47570 42978 47582
rect 42926 47506 42978 47518
rect 2494 47458 2546 47470
rect 2494 47394 2546 47406
rect 3166 47458 3218 47470
rect 3166 47394 3218 47406
rect 3502 47458 3554 47470
rect 3502 47394 3554 47406
rect 3726 47458 3778 47470
rect 9998 47458 10050 47470
rect 4050 47406 4062 47458
rect 4114 47406 4126 47458
rect 5842 47406 5854 47458
rect 5906 47406 5918 47458
rect 7522 47406 7534 47458
rect 7586 47406 7598 47458
rect 3726 47394 3778 47406
rect 9998 47394 10050 47406
rect 10334 47458 10386 47470
rect 11902 47458 11954 47470
rect 24446 47458 24498 47470
rect 27918 47458 27970 47470
rect 10546 47406 10558 47458
rect 10610 47406 10622 47458
rect 13570 47406 13582 47458
rect 13634 47406 13646 47458
rect 26114 47406 26126 47458
rect 26178 47406 26190 47458
rect 10334 47394 10386 47406
rect 11902 47394 11954 47406
rect 24446 47394 24498 47406
rect 27918 47394 27970 47406
rect 28590 47458 28642 47470
rect 34414 47458 34466 47470
rect 31490 47406 31502 47458
rect 31554 47406 31566 47458
rect 32162 47406 32174 47458
rect 32226 47406 32238 47458
rect 28590 47394 28642 47406
rect 34414 47394 34466 47406
rect 34638 47458 34690 47470
rect 34638 47394 34690 47406
rect 35870 47458 35922 47470
rect 35870 47394 35922 47406
rect 36094 47458 36146 47470
rect 37090 47406 37102 47458
rect 37154 47406 37166 47458
rect 40898 47406 40910 47458
rect 40962 47406 40974 47458
rect 41682 47406 41694 47458
rect 41746 47406 41758 47458
rect 36094 47394 36146 47406
rect 2270 47346 2322 47358
rect 2270 47282 2322 47294
rect 2382 47346 2434 47358
rect 2382 47282 2434 47294
rect 9662 47346 9714 47358
rect 9662 47282 9714 47294
rect 11230 47346 11282 47358
rect 11230 47282 11282 47294
rect 11566 47346 11618 47358
rect 11566 47282 11618 47294
rect 11678 47346 11730 47358
rect 11678 47282 11730 47294
rect 12238 47346 12290 47358
rect 12238 47282 12290 47294
rect 22094 47346 22146 47358
rect 22094 47282 22146 47294
rect 22430 47346 22482 47358
rect 43822 47346 43874 47358
rect 25666 47294 25678 47346
rect 25730 47294 25742 47346
rect 26562 47294 26574 47346
rect 26626 47294 26638 47346
rect 31378 47294 31390 47346
rect 31442 47294 31454 47346
rect 32050 47294 32062 47346
rect 32114 47294 32126 47346
rect 22430 47282 22482 47294
rect 43822 47282 43874 47294
rect 4174 47234 4226 47246
rect 4174 47170 4226 47182
rect 4398 47234 4450 47246
rect 4398 47170 4450 47182
rect 4958 47234 5010 47246
rect 4958 47170 5010 47182
rect 8878 47234 8930 47246
rect 8878 47170 8930 47182
rect 9326 47234 9378 47246
rect 9326 47170 9378 47182
rect 9774 47234 9826 47246
rect 9774 47170 9826 47182
rect 16830 47234 16882 47246
rect 16830 47170 16882 47182
rect 18510 47234 18562 47246
rect 18510 47170 18562 47182
rect 19518 47234 19570 47246
rect 19518 47170 19570 47182
rect 19966 47234 20018 47246
rect 19966 47170 20018 47182
rect 20414 47234 20466 47246
rect 20414 47170 20466 47182
rect 21422 47234 21474 47246
rect 21422 47170 21474 47182
rect 29262 47234 29314 47246
rect 35086 47234 35138 47246
rect 30146 47182 30158 47234
rect 30210 47182 30222 47234
rect 34066 47182 34078 47234
rect 34130 47182 34142 47234
rect 29262 47170 29314 47182
rect 35086 47170 35138 47182
rect 35534 47234 35586 47246
rect 44158 47234 44210 47246
rect 43250 47182 43262 47234
rect 43314 47182 43326 47234
rect 35534 47170 35586 47182
rect 44158 47170 44210 47182
rect 1344 47066 48608 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 48608 47066
rect 1344 46980 48608 47014
rect 4174 46898 4226 46910
rect 3154 46846 3166 46898
rect 3218 46846 3230 46898
rect 4174 46834 4226 46846
rect 4510 46898 4562 46910
rect 4510 46834 4562 46846
rect 4622 46898 4674 46910
rect 8542 46898 8594 46910
rect 7970 46846 7982 46898
rect 8034 46846 8046 46898
rect 4622 46834 4674 46846
rect 8542 46834 8594 46846
rect 17614 46898 17666 46910
rect 17614 46834 17666 46846
rect 25902 46898 25954 46910
rect 25902 46834 25954 46846
rect 28590 46898 28642 46910
rect 33854 46898 33906 46910
rect 31826 46846 31838 46898
rect 31890 46846 31902 46898
rect 28590 46834 28642 46846
rect 33854 46834 33906 46846
rect 38894 46898 38946 46910
rect 41234 46846 41246 46898
rect 41298 46846 41310 46898
rect 38894 46834 38946 46846
rect 4846 46786 4898 46798
rect 8766 46786 8818 46798
rect 28142 46786 28194 46798
rect 34638 46786 34690 46798
rect 39006 46786 39058 46798
rect 5506 46734 5518 46786
rect 5570 46734 5582 46786
rect 10098 46734 10110 46786
rect 10162 46734 10174 46786
rect 10434 46734 10446 46786
rect 10498 46734 10510 46786
rect 21522 46734 21534 46786
rect 21586 46734 21598 46786
rect 22306 46734 22318 46786
rect 22370 46734 22382 46786
rect 26562 46734 26574 46786
rect 26626 46734 26638 46786
rect 32386 46734 32398 46786
rect 32450 46734 32462 46786
rect 36194 46734 36206 46786
rect 36258 46734 36270 46786
rect 37090 46734 37102 46786
rect 37154 46734 37166 46786
rect 4846 46722 4898 46734
rect 8766 46722 8818 46734
rect 28142 46722 28194 46734
rect 34638 46722 34690 46734
rect 39006 46722 39058 46734
rect 39902 46786 39954 46798
rect 43598 46786 43650 46798
rect 41122 46734 41134 46786
rect 41186 46734 41198 46786
rect 45938 46734 45950 46786
rect 46002 46734 46014 46786
rect 39902 46722 39954 46734
rect 43598 46722 43650 46734
rect 4398 46674 4450 46686
rect 7422 46674 7474 46686
rect 6178 46622 6190 46674
rect 6242 46622 6254 46674
rect 6850 46622 6862 46674
rect 6914 46622 6926 46674
rect 7186 46622 7198 46674
rect 7250 46622 7262 46674
rect 4398 46610 4450 46622
rect 7422 46610 7474 46622
rect 7534 46674 7586 46686
rect 7534 46610 7586 46622
rect 8318 46674 8370 46686
rect 8318 46610 8370 46622
rect 9662 46674 9714 46686
rect 44718 46674 44770 46686
rect 19394 46622 19406 46674
rect 19458 46622 19470 46674
rect 20402 46622 20414 46674
rect 20466 46622 20478 46674
rect 21634 46622 21646 46674
rect 21698 46622 21710 46674
rect 23986 46622 23998 46674
rect 24050 46622 24062 46674
rect 26226 46622 26238 46674
rect 26290 46622 26302 46674
rect 32274 46622 32286 46674
rect 32338 46622 32350 46674
rect 34066 46622 34078 46674
rect 34130 46622 34142 46674
rect 35522 46622 35534 46674
rect 35586 46622 35598 46674
rect 38546 46622 38558 46674
rect 38610 46622 38622 46674
rect 39666 46622 39678 46674
rect 39730 46622 39742 46674
rect 41010 46622 41022 46674
rect 41074 46622 41086 46674
rect 45154 46622 45166 46674
rect 45218 46622 45230 46674
rect 9662 46610 9714 46622
rect 44718 46610 44770 46622
rect 2270 46562 2322 46574
rect 2270 46498 2322 46510
rect 2606 46562 2658 46574
rect 2606 46498 2658 46510
rect 3614 46562 3666 46574
rect 8430 46562 8482 46574
rect 5954 46510 5966 46562
rect 6018 46510 6030 46562
rect 3614 46498 3666 46510
rect 8430 46498 8482 46510
rect 9438 46562 9490 46574
rect 9438 46498 9490 46510
rect 11118 46562 11170 46574
rect 11118 46498 11170 46510
rect 15374 46562 15426 46574
rect 15374 46498 15426 46510
rect 18286 46562 18338 46574
rect 18286 46498 18338 46510
rect 18846 46562 18898 46574
rect 29038 46562 29090 46574
rect 19842 46510 19854 46562
rect 19906 46510 19918 46562
rect 20066 46510 20078 46562
rect 20130 46510 20142 46562
rect 23426 46510 23438 46562
rect 23490 46510 23502 46562
rect 18846 46498 18898 46510
rect 29038 46498 29090 46510
rect 29822 46562 29874 46574
rect 29822 46498 29874 46510
rect 30382 46562 30434 46574
rect 30382 46498 30434 46510
rect 33294 46562 33346 46574
rect 40350 46562 40402 46574
rect 37874 46510 37886 46562
rect 37938 46510 37950 46562
rect 48066 46510 48078 46562
rect 48130 46510 48142 46562
rect 33294 46498 33346 46510
rect 40350 46498 40402 46510
rect 2830 46450 2882 46462
rect 2830 46386 2882 46398
rect 17502 46450 17554 46462
rect 17502 46386 17554 46398
rect 17838 46450 17890 46462
rect 29810 46398 29822 46450
rect 29874 46447 29886 46450
rect 30594 46447 30606 46450
rect 29874 46401 30606 46447
rect 29874 46398 29886 46401
rect 30594 46398 30606 46401
rect 30658 46398 30670 46450
rect 17838 46386 17890 46398
rect 1344 46282 48608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48608 46282
rect 1344 46196 48608 46230
rect 2942 46114 2994 46126
rect 22654 46114 22706 46126
rect 20402 46062 20414 46114
rect 20466 46062 20478 46114
rect 42466 46062 42478 46114
rect 42530 46111 42542 46114
rect 43138 46111 43150 46114
rect 42530 46065 43150 46111
rect 42530 46062 42542 46065
rect 43138 46062 43150 46065
rect 43202 46062 43214 46114
rect 2942 46050 2994 46062
rect 22654 46050 22706 46062
rect 2158 46002 2210 46014
rect 2158 45938 2210 45950
rect 3054 46002 3106 46014
rect 3054 45938 3106 45950
rect 4174 46002 4226 46014
rect 29150 46002 29202 46014
rect 37774 46002 37826 46014
rect 43150 46002 43202 46014
rect 9090 45950 9102 46002
rect 9154 45950 9166 46002
rect 16818 45950 16830 46002
rect 16882 45950 16894 46002
rect 18946 45950 18958 46002
rect 19010 45950 19022 46002
rect 33506 45950 33518 46002
rect 33570 45950 33582 46002
rect 40114 45950 40126 46002
rect 40178 45950 40190 46002
rect 42242 45950 42254 46002
rect 42306 45950 42318 46002
rect 4174 45938 4226 45950
rect 29150 45938 29202 45950
rect 37774 45938 37826 45950
rect 43150 45938 43202 45950
rect 1934 45890 1986 45902
rect 1934 45826 1986 45838
rect 2606 45890 2658 45902
rect 3614 45890 3666 45902
rect 3266 45838 3278 45890
rect 3330 45838 3342 45890
rect 2606 45826 2658 45838
rect 3614 45826 3666 45838
rect 3726 45890 3778 45902
rect 20750 45890 20802 45902
rect 9874 45838 9886 45890
rect 9938 45838 9950 45890
rect 14466 45838 14478 45890
rect 14530 45838 14542 45890
rect 16146 45838 16158 45890
rect 16210 45838 16222 45890
rect 19282 45838 19294 45890
rect 19346 45838 19358 45890
rect 20178 45838 20190 45890
rect 20242 45838 20254 45890
rect 3726 45826 3778 45838
rect 20750 45826 20802 45838
rect 22318 45890 22370 45902
rect 22318 45826 22370 45838
rect 22990 45890 23042 45902
rect 22990 45826 23042 45838
rect 23662 45890 23714 45902
rect 23662 45826 23714 45838
rect 29934 45890 29986 45902
rect 36094 45890 36146 45902
rect 30370 45838 30382 45890
rect 30434 45838 30446 45890
rect 31266 45838 31278 45890
rect 31330 45838 31342 45890
rect 35186 45838 35198 45890
rect 35250 45838 35262 45890
rect 39442 45838 39454 45890
rect 39506 45838 39518 45890
rect 29934 45826 29986 45838
rect 36094 45826 36146 45838
rect 2382 45778 2434 45790
rect 19518 45778 19570 45790
rect 14914 45726 14926 45778
rect 14978 45726 14990 45778
rect 2382 45714 2434 45726
rect 19518 45714 19570 45726
rect 23214 45778 23266 45790
rect 23214 45714 23266 45726
rect 29374 45778 29426 45790
rect 30718 45778 30770 45790
rect 29586 45726 29598 45778
rect 29650 45726 29662 45778
rect 34626 45726 34638 45778
rect 34690 45726 34702 45778
rect 29374 45714 29426 45726
rect 30718 45714 30770 45726
rect 4622 45666 4674 45678
rect 4622 45602 4674 45614
rect 5070 45666 5122 45678
rect 5070 45602 5122 45614
rect 6078 45666 6130 45678
rect 6078 45602 6130 45614
rect 6414 45666 6466 45678
rect 10334 45666 10386 45678
rect 6850 45614 6862 45666
rect 6914 45614 6926 45666
rect 6414 45602 6466 45614
rect 10334 45602 10386 45614
rect 15710 45666 15762 45678
rect 15710 45602 15762 45614
rect 21422 45666 21474 45678
rect 21422 45602 21474 45614
rect 21870 45666 21922 45678
rect 21870 45602 21922 45614
rect 26462 45666 26514 45678
rect 26462 45602 26514 45614
rect 28142 45666 28194 45678
rect 28142 45602 28194 45614
rect 28590 45666 28642 45678
rect 28590 45602 28642 45614
rect 30158 45666 30210 45678
rect 30158 45602 30210 45614
rect 30606 45666 30658 45678
rect 37326 45666 37378 45678
rect 34290 45614 34302 45666
rect 34354 45614 34366 45666
rect 30606 45602 30658 45614
rect 37326 45602 37378 45614
rect 38222 45666 38274 45678
rect 38222 45602 38274 45614
rect 38670 45666 38722 45678
rect 38670 45602 38722 45614
rect 42702 45666 42754 45678
rect 42702 45602 42754 45614
rect 43598 45666 43650 45678
rect 43598 45602 43650 45614
rect 44046 45666 44098 45678
rect 44046 45602 44098 45614
rect 44942 45666 44994 45678
rect 44942 45602 44994 45614
rect 1344 45498 48608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48608 45498
rect 1344 45412 48608 45446
rect 2830 45330 2882 45342
rect 2830 45266 2882 45278
rect 19182 45330 19234 45342
rect 19182 45266 19234 45278
rect 26910 45330 26962 45342
rect 26910 45266 26962 45278
rect 27134 45330 27186 45342
rect 27134 45266 27186 45278
rect 31166 45330 31218 45342
rect 31166 45266 31218 45278
rect 32510 45330 32562 45342
rect 32510 45266 32562 45278
rect 34302 45330 34354 45342
rect 34302 45266 34354 45278
rect 35086 45330 35138 45342
rect 35086 45266 35138 45278
rect 35534 45330 35586 45342
rect 39666 45278 39678 45330
rect 39730 45278 39742 45330
rect 35534 45266 35586 45278
rect 19070 45218 19122 45230
rect 23326 45218 23378 45230
rect 8082 45166 8094 45218
rect 8146 45166 8158 45218
rect 22194 45166 22206 45218
rect 22258 45166 22270 45218
rect 19070 45154 19122 45166
rect 23326 45154 23378 45166
rect 28030 45218 28082 45230
rect 31614 45218 31666 45230
rect 29026 45166 29038 45218
rect 29090 45166 29102 45218
rect 30482 45166 30494 45218
rect 30546 45166 30558 45218
rect 28030 45154 28082 45166
rect 31614 45154 31666 45166
rect 33070 45218 33122 45230
rect 41906 45166 41918 45218
rect 41970 45166 41982 45218
rect 33070 45154 33122 45166
rect 22990 45106 23042 45118
rect 3490 45054 3502 45106
rect 3554 45054 3566 45106
rect 12898 45054 12910 45106
rect 12962 45054 12974 45106
rect 20962 45054 20974 45106
rect 21026 45054 21038 45106
rect 22082 45054 22094 45106
rect 22146 45054 22158 45106
rect 22990 45042 23042 45054
rect 25454 45106 25506 45118
rect 25454 45042 25506 45054
rect 25678 45106 25730 45118
rect 27918 45106 27970 45118
rect 31390 45106 31442 45118
rect 26674 45054 26686 45106
rect 26738 45054 26750 45106
rect 27346 45054 27358 45106
rect 27410 45054 27422 45106
rect 28242 45054 28254 45106
rect 28306 45054 28318 45106
rect 28914 45054 28926 45106
rect 28978 45054 28990 45106
rect 29922 45054 29934 45106
rect 29986 45054 29998 45106
rect 30930 45054 30942 45106
rect 30994 45054 31006 45106
rect 25678 45042 25730 45054
rect 27918 45042 27970 45054
rect 31390 45042 31442 45054
rect 33294 45106 33346 45118
rect 41694 45106 41746 45118
rect 33618 45054 33630 45106
rect 33682 45054 33694 45106
rect 37538 45054 37550 45106
rect 37602 45054 37614 45106
rect 38098 45054 38110 45106
rect 38162 45054 38174 45106
rect 38770 45054 38782 45106
rect 38834 45054 38846 45106
rect 42354 45054 42366 45106
rect 42418 45054 42430 45106
rect 42914 45054 42926 45106
rect 42978 45054 42990 45106
rect 43474 45054 43486 45106
rect 43538 45054 43550 45106
rect 33294 45042 33346 45054
rect 41694 45042 41746 45054
rect 2382 44994 2434 45006
rect 19630 44994 19682 45006
rect 23662 44994 23714 45006
rect 16482 44942 16494 44994
rect 16546 44942 16558 44994
rect 21746 44942 21758 44994
rect 21810 44942 21822 44994
rect 2382 44930 2434 44942
rect 19630 44930 19682 44942
rect 23662 44930 23714 44942
rect 24222 44994 24274 45006
rect 24222 44930 24274 44942
rect 24670 44994 24722 45006
rect 27694 44994 27746 45006
rect 31278 44994 31330 45006
rect 27234 44942 27246 44994
rect 27298 44942 27310 44994
rect 29362 44942 29374 44994
rect 29426 44942 29438 44994
rect 24670 44930 24722 44942
rect 27694 44930 27746 44942
rect 31278 44930 31330 44942
rect 32062 44994 32114 45006
rect 32062 44930 32114 44942
rect 34638 44994 34690 45006
rect 34638 44930 34690 44942
rect 35982 44994 36034 45006
rect 35982 44930 36034 44942
rect 36766 44994 36818 45006
rect 36766 44930 36818 44942
rect 37102 44994 37154 45006
rect 39118 44994 39170 45006
rect 38546 44942 38558 44994
rect 38610 44942 38622 44994
rect 37102 44930 37154 44942
rect 39118 44930 39170 44942
rect 39342 44994 39394 45006
rect 39342 44930 39394 44942
rect 40126 44994 40178 45006
rect 40126 44930 40178 44942
rect 41246 44994 41298 45006
rect 44258 44942 44270 44994
rect 44322 44942 44334 44994
rect 46386 44942 46398 44994
rect 46450 44942 46462 44994
rect 41246 44930 41298 44942
rect 23998 44882 24050 44894
rect 28702 44882 28754 44894
rect 41582 44882 41634 44894
rect 26002 44830 26014 44882
rect 26066 44830 26078 44882
rect 35522 44830 35534 44882
rect 35586 44879 35598 44882
rect 35858 44879 35870 44882
rect 35586 44833 35870 44879
rect 35586 44830 35598 44833
rect 35858 44830 35870 44833
rect 35922 44830 35934 44882
rect 23998 44818 24050 44830
rect 28702 44818 28754 44830
rect 41582 44818 41634 44830
rect 1344 44714 48608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48608 44714
rect 1344 44628 48608 44662
rect 38782 44546 38834 44558
rect 21970 44494 21982 44546
rect 22034 44543 22046 44546
rect 22530 44543 22542 44546
rect 22034 44497 22542 44543
rect 22034 44494 22046 44497
rect 22530 44494 22542 44497
rect 22594 44494 22606 44546
rect 38782 44482 38834 44494
rect 44046 44546 44098 44558
rect 44046 44482 44098 44494
rect 6302 44434 6354 44446
rect 13582 44434 13634 44446
rect 6738 44382 6750 44434
rect 6802 44382 6814 44434
rect 12898 44382 12910 44434
rect 12962 44382 12974 44434
rect 6302 44370 6354 44382
rect 13582 44370 13634 44382
rect 16606 44434 16658 44446
rect 16606 44370 16658 44382
rect 18622 44434 18674 44446
rect 18622 44370 18674 44382
rect 21422 44434 21474 44446
rect 21422 44370 21474 44382
rect 21982 44434 22034 44446
rect 27358 44434 27410 44446
rect 23538 44382 23550 44434
rect 23602 44382 23614 44434
rect 25666 44382 25678 44434
rect 25730 44382 25742 44434
rect 21982 44370 22034 44382
rect 27358 44370 27410 44382
rect 28030 44434 28082 44446
rect 39902 44434 39954 44446
rect 33394 44382 33406 44434
rect 33458 44382 33470 44434
rect 28030 44370 28082 44382
rect 39902 44370 39954 44382
rect 40350 44434 40402 44446
rect 40350 44370 40402 44382
rect 42702 44434 42754 44446
rect 42702 44370 42754 44382
rect 43374 44434 43426 44446
rect 43374 44370 43426 44382
rect 43710 44434 43762 44446
rect 43710 44370 43762 44382
rect 2494 44322 2546 44334
rect 2494 44258 2546 44270
rect 2942 44322 2994 44334
rect 2942 44258 2994 44270
rect 3502 44322 3554 44334
rect 3502 44258 3554 44270
rect 4398 44322 4450 44334
rect 5966 44322 6018 44334
rect 4722 44270 4734 44322
rect 4786 44270 4798 44322
rect 4398 44258 4450 44270
rect 5966 44258 6018 44270
rect 6190 44322 6242 44334
rect 6190 44258 6242 44270
rect 6526 44322 6578 44334
rect 16382 44322 16434 44334
rect 9650 44270 9662 44322
rect 9714 44270 9726 44322
rect 10098 44270 10110 44322
rect 10162 44270 10174 44322
rect 6526 44258 6578 44270
rect 16382 44258 16434 44270
rect 19182 44322 19234 44334
rect 28366 44322 28418 44334
rect 35422 44322 35474 44334
rect 39006 44322 39058 44334
rect 22754 44270 22766 44322
rect 22818 44270 22830 44322
rect 29138 44270 29150 44322
rect 29202 44270 29214 44322
rect 30594 44270 30606 44322
rect 30658 44270 30670 44322
rect 32162 44270 32174 44322
rect 32226 44270 32238 44322
rect 33058 44270 33070 44322
rect 33122 44270 33134 44322
rect 34962 44270 34974 44322
rect 35026 44270 35038 44322
rect 37650 44270 37662 44322
rect 37714 44270 37726 44322
rect 38322 44270 38334 44322
rect 38386 44270 38398 44322
rect 41570 44270 41582 44322
rect 41634 44270 41646 44322
rect 42578 44270 42590 44322
rect 42642 44270 42654 44322
rect 44034 44270 44046 44322
rect 44098 44270 44110 44322
rect 19182 44258 19234 44270
rect 28366 44258 28418 44270
rect 35422 44258 35474 44270
rect 39006 44258 39058 44270
rect 2830 44210 2882 44222
rect 2830 44146 2882 44158
rect 4174 44210 4226 44222
rect 15486 44210 15538 44222
rect 19070 44210 19122 44222
rect 8866 44158 8878 44210
rect 8930 44158 8942 44210
rect 10770 44158 10782 44210
rect 10834 44158 10846 44210
rect 16034 44158 16046 44210
rect 16098 44158 16110 44210
rect 4174 44146 4226 44158
rect 15486 44146 15538 44158
rect 19070 44146 19122 44158
rect 26126 44210 26178 44222
rect 26126 44146 26178 44158
rect 26238 44210 26290 44222
rect 26238 44146 26290 44158
rect 28478 44210 28530 44222
rect 35982 44210 36034 44222
rect 30370 44158 30382 44210
rect 30434 44158 30446 44210
rect 31938 44158 31950 44210
rect 32002 44158 32014 44210
rect 32946 44158 32958 44210
rect 33010 44158 33022 44210
rect 28478 44146 28530 44158
rect 35982 44146 36034 44158
rect 37774 44210 37826 44222
rect 37774 44146 37826 44158
rect 39454 44210 39506 44222
rect 39454 44146 39506 44158
rect 40798 44210 40850 44222
rect 42802 44158 42814 44210
rect 42866 44158 42878 44210
rect 40798 44146 40850 44158
rect 2606 44098 2658 44110
rect 2606 44034 2658 44046
rect 3838 44098 3890 44110
rect 3838 44034 3890 44046
rect 15150 44098 15202 44110
rect 15150 44034 15202 44046
rect 17054 44098 17106 44110
rect 17054 44034 17106 44046
rect 17502 44098 17554 44110
rect 17502 44034 17554 44046
rect 18846 44098 18898 44110
rect 18846 44034 18898 44046
rect 20638 44098 20690 44110
rect 20638 44034 20690 44046
rect 22430 44098 22482 44110
rect 22430 44034 22482 44046
rect 26462 44098 26514 44110
rect 26462 44034 26514 44046
rect 26798 44098 26850 44110
rect 26798 44034 26850 44046
rect 28702 44098 28754 44110
rect 31166 44098 31218 44110
rect 29250 44046 29262 44098
rect 29314 44046 29326 44098
rect 29474 44046 29486 44098
rect 29538 44046 29550 44098
rect 28702 44034 28754 44046
rect 31166 44034 31218 44046
rect 35198 44098 35250 44110
rect 35198 44034 35250 44046
rect 35310 44098 35362 44110
rect 35310 44034 35362 44046
rect 35534 44098 35586 44110
rect 35534 44034 35586 44046
rect 36318 44098 36370 44110
rect 36318 44034 36370 44046
rect 37214 44098 37266 44110
rect 37214 44034 37266 44046
rect 41246 44098 41298 44110
rect 41246 44034 41298 44046
rect 1344 43930 48608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48608 43930
rect 1344 43844 48608 43878
rect 8654 43762 8706 43774
rect 8654 43698 8706 43710
rect 8878 43762 8930 43774
rect 8878 43698 8930 43710
rect 9886 43762 9938 43774
rect 9886 43698 9938 43710
rect 10334 43762 10386 43774
rect 10334 43698 10386 43710
rect 11342 43762 11394 43774
rect 11342 43698 11394 43710
rect 17838 43762 17890 43774
rect 41794 43710 41806 43762
rect 41858 43710 41870 43762
rect 17838 43698 17890 43710
rect 28814 43650 28866 43662
rect 8194 43598 8206 43650
rect 8258 43598 8270 43650
rect 14690 43598 14702 43650
rect 14754 43598 14766 43650
rect 18946 43598 18958 43650
rect 19010 43598 19022 43650
rect 22866 43598 22878 43650
rect 22930 43598 22942 43650
rect 23986 43598 23998 43650
rect 24050 43598 24062 43650
rect 28814 43586 28866 43598
rect 30942 43650 30994 43662
rect 41022 43650 41074 43662
rect 34738 43598 34750 43650
rect 34802 43598 34814 43650
rect 35522 43598 35534 43650
rect 35586 43598 35598 43650
rect 38210 43598 38222 43650
rect 38274 43598 38286 43650
rect 30942 43586 30994 43598
rect 41022 43586 41074 43598
rect 42814 43650 42866 43662
rect 42814 43586 42866 43598
rect 44270 43650 44322 43662
rect 44270 43586 44322 43598
rect 45950 43650 46002 43662
rect 45950 43586 46002 43598
rect 7534 43538 7586 43550
rect 6626 43486 6638 43538
rect 6690 43486 6702 43538
rect 7534 43474 7586 43486
rect 7870 43538 7922 43550
rect 7870 43474 7922 43486
rect 8542 43538 8594 43550
rect 30382 43538 30434 43550
rect 13906 43486 13918 43538
rect 13970 43486 13982 43538
rect 18274 43486 18286 43538
rect 18338 43486 18350 43538
rect 21410 43486 21422 43538
rect 21474 43486 21486 43538
rect 23538 43486 23550 43538
rect 23602 43486 23614 43538
rect 8542 43474 8594 43486
rect 30382 43474 30434 43486
rect 32286 43538 32338 43550
rect 34626 43486 34638 43538
rect 34690 43486 34702 43538
rect 37090 43486 37102 43538
rect 37154 43486 37166 43538
rect 37426 43486 37438 43538
rect 37490 43486 37502 43538
rect 43250 43486 43262 43538
rect 43314 43486 43326 43538
rect 43698 43486 43710 43538
rect 43762 43486 43774 43538
rect 32286 43474 32338 43486
rect 10894 43426 10946 43438
rect 2706 43374 2718 43426
rect 2770 43374 2782 43426
rect 10894 43362 10946 43374
rect 11790 43426 11842 43438
rect 25342 43426 25394 43438
rect 16818 43374 16830 43426
rect 16882 43374 16894 43426
rect 21074 43374 21086 43426
rect 21138 43374 21150 43426
rect 21746 43374 21758 43426
rect 21810 43374 21822 43426
rect 11790 43362 11842 43374
rect 25342 43362 25394 43374
rect 29262 43426 29314 43438
rect 29262 43362 29314 43374
rect 30046 43426 30098 43438
rect 30046 43362 30098 43374
rect 31502 43426 31554 43438
rect 31502 43362 31554 43374
rect 31838 43426 31890 43438
rect 31838 43362 31890 43374
rect 33182 43426 33234 43438
rect 40338 43374 40350 43426
rect 40402 43374 40414 43426
rect 33182 43362 33234 43374
rect 7422 43314 7474 43326
rect 33966 43314 34018 43326
rect 10770 43262 10782 43314
rect 10834 43311 10846 43314
rect 11442 43311 11454 43314
rect 10834 43265 11454 43311
rect 10834 43262 10846 43265
rect 11442 43262 11454 43265
rect 11506 43262 11518 43314
rect 32946 43262 32958 43314
rect 33010 43311 33022 43314
rect 33506 43311 33518 43314
rect 33010 43265 33518 43311
rect 33010 43262 33022 43265
rect 33506 43262 33518 43265
rect 33570 43262 33582 43314
rect 7422 43250 7474 43262
rect 33966 43250 34018 43262
rect 45838 43314 45890 43326
rect 45838 43250 45890 43262
rect 1344 43146 48608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48608 43146
rect 1344 43060 48608 43094
rect 20862 42978 20914 42990
rect 25666 42926 25678 42978
rect 25730 42975 25742 42978
rect 26562 42975 26574 42978
rect 25730 42929 26574 42975
rect 25730 42926 25742 42929
rect 26562 42926 26574 42929
rect 26626 42926 26638 42978
rect 27794 42926 27806 42978
rect 27858 42926 27870 42978
rect 20862 42914 20914 42926
rect 2606 42866 2658 42878
rect 2606 42802 2658 42814
rect 4062 42866 4114 42878
rect 4062 42802 4114 42814
rect 6750 42866 6802 42878
rect 6750 42802 6802 42814
rect 7198 42866 7250 42878
rect 7198 42802 7250 42814
rect 7758 42866 7810 42878
rect 7758 42802 7810 42814
rect 11454 42866 11506 42878
rect 11454 42802 11506 42814
rect 16158 42866 16210 42878
rect 16158 42802 16210 42814
rect 17614 42866 17666 42878
rect 17614 42802 17666 42814
rect 18958 42866 19010 42878
rect 18958 42802 19010 42814
rect 21310 42866 21362 42878
rect 21310 42802 21362 42814
rect 26574 42866 26626 42878
rect 26574 42802 26626 42814
rect 29262 42866 29314 42878
rect 29262 42802 29314 42814
rect 29822 42866 29874 42878
rect 29822 42802 29874 42814
rect 30718 42866 30770 42878
rect 30718 42802 30770 42814
rect 31166 42866 31218 42878
rect 35198 42866 35250 42878
rect 32946 42814 32958 42866
rect 33010 42814 33022 42866
rect 31166 42802 31218 42814
rect 35198 42802 35250 42814
rect 1934 42754 1986 42766
rect 1934 42690 1986 42702
rect 2270 42754 2322 42766
rect 4398 42754 4450 42766
rect 20750 42754 20802 42766
rect 2482 42702 2494 42754
rect 2546 42702 2558 42754
rect 2706 42702 2718 42754
rect 2770 42702 2782 42754
rect 3490 42702 3502 42754
rect 3554 42702 3566 42754
rect 6178 42702 6190 42754
rect 6242 42702 6254 42754
rect 6514 42702 6526 42754
rect 6578 42702 6590 42754
rect 10546 42702 10558 42754
rect 10610 42702 10622 42754
rect 13906 42702 13918 42754
rect 13970 42702 13982 42754
rect 19282 42702 19294 42754
rect 19346 42702 19358 42754
rect 20066 42702 20078 42754
rect 20130 42702 20142 42754
rect 2270 42690 2322 42702
rect 4398 42690 4450 42702
rect 20750 42690 20802 42702
rect 27246 42754 27298 42766
rect 35534 42754 35586 42766
rect 37550 42754 37602 42766
rect 33282 42702 33294 42754
rect 33346 42702 33358 42754
rect 33506 42702 33518 42754
rect 33570 42702 33582 42754
rect 35746 42702 35758 42754
rect 35810 42702 35822 42754
rect 27246 42690 27298 42702
rect 35534 42690 35586 42702
rect 37550 42690 37602 42702
rect 37662 42754 37714 42766
rect 37662 42690 37714 42702
rect 39790 42754 39842 42766
rect 39790 42690 39842 42702
rect 40238 42754 40290 42766
rect 40238 42690 40290 42702
rect 2942 42642 2994 42654
rect 2942 42578 2994 42590
rect 3278 42642 3330 42654
rect 3278 42578 3330 42590
rect 3726 42642 3778 42654
rect 3726 42578 3778 42590
rect 4174 42642 4226 42654
rect 11006 42642 11058 42654
rect 9874 42590 9886 42642
rect 9938 42590 9950 42642
rect 4174 42578 4226 42590
rect 11006 42578 11058 42590
rect 11230 42642 11282 42654
rect 11230 42578 11282 42590
rect 11566 42642 11618 42654
rect 27134 42642 27186 42654
rect 19394 42590 19406 42642
rect 19458 42590 19470 42642
rect 11566 42578 11618 42590
rect 27134 42578 27186 42590
rect 27358 42642 27410 42654
rect 35422 42642 35474 42654
rect 33170 42590 33182 42642
rect 33234 42590 33246 42642
rect 33954 42590 33966 42642
rect 34018 42590 34030 42642
rect 27358 42578 27410 42590
rect 35422 42578 35474 42590
rect 37438 42642 37490 42654
rect 37438 42578 37490 42590
rect 38670 42642 38722 42654
rect 38670 42578 38722 42590
rect 40686 42642 40738 42654
rect 40686 42578 40738 42590
rect 2046 42530 2098 42542
rect 2046 42466 2098 42478
rect 3838 42530 3890 42542
rect 3838 42466 3890 42478
rect 4846 42530 4898 42542
rect 4846 42466 4898 42478
rect 4958 42530 5010 42542
rect 4958 42466 5010 42478
rect 5070 42530 5122 42542
rect 5070 42466 5122 42478
rect 12126 42530 12178 42542
rect 12126 42466 12178 42478
rect 12574 42530 12626 42542
rect 12574 42466 12626 42478
rect 12910 42530 12962 42542
rect 12910 42466 12962 42478
rect 17166 42530 17218 42542
rect 17166 42466 17218 42478
rect 18062 42530 18114 42542
rect 18062 42466 18114 42478
rect 18510 42530 18562 42542
rect 18510 42466 18562 42478
rect 21422 42530 21474 42542
rect 21422 42466 21474 42478
rect 21870 42530 21922 42542
rect 21870 42466 21922 42478
rect 22318 42530 22370 42542
rect 22318 42466 22370 42478
rect 26014 42530 26066 42542
rect 26014 42466 26066 42478
rect 28254 42530 28306 42542
rect 28254 42466 28306 42478
rect 30270 42530 30322 42542
rect 30270 42466 30322 42478
rect 36206 42530 36258 42542
rect 42478 42530 42530 42542
rect 36978 42478 36990 42530
rect 37042 42478 37054 42530
rect 38210 42478 38222 42530
rect 38274 42478 38286 42530
rect 36206 42466 36258 42478
rect 42478 42466 42530 42478
rect 42926 42530 42978 42542
rect 42926 42466 42978 42478
rect 1344 42362 48608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48608 42362
rect 1344 42276 48608 42310
rect 2270 42194 2322 42206
rect 2270 42130 2322 42142
rect 8990 42194 9042 42206
rect 8990 42130 9042 42142
rect 9438 42194 9490 42206
rect 9438 42130 9490 42142
rect 9662 42194 9714 42206
rect 9662 42130 9714 42142
rect 10558 42194 10610 42206
rect 10558 42130 10610 42142
rect 14814 42194 14866 42206
rect 14814 42130 14866 42142
rect 16606 42194 16658 42206
rect 16606 42130 16658 42142
rect 23326 42194 23378 42206
rect 23326 42130 23378 42142
rect 28814 42194 28866 42206
rect 28814 42130 28866 42142
rect 34974 42194 35026 42206
rect 34974 42130 35026 42142
rect 2718 42082 2770 42094
rect 2718 42018 2770 42030
rect 10446 42082 10498 42094
rect 10446 42018 10498 42030
rect 17502 42082 17554 42094
rect 17502 42018 17554 42030
rect 18622 42082 18674 42094
rect 18622 42018 18674 42030
rect 23438 42082 23490 42094
rect 23438 42018 23490 42030
rect 29262 42082 29314 42094
rect 40126 42082 40178 42094
rect 30258 42030 30270 42082
rect 30322 42030 30334 42082
rect 32274 42030 32286 42082
rect 32338 42030 32350 42082
rect 33058 42030 33070 42082
rect 33122 42030 33134 42082
rect 36082 42030 36094 42082
rect 36146 42030 36158 42082
rect 37314 42030 37326 42082
rect 37378 42030 37390 42082
rect 29262 42018 29314 42030
rect 40126 42018 40178 42030
rect 40238 42082 40290 42094
rect 40238 42018 40290 42030
rect 2830 41970 2882 41982
rect 9774 41970 9826 41982
rect 10670 41970 10722 41982
rect 16158 41970 16210 41982
rect 3826 41918 3838 41970
rect 3890 41918 3902 41970
rect 10098 41918 10110 41970
rect 10162 41918 10174 41970
rect 10994 41918 11006 41970
rect 11058 41918 11070 41970
rect 14466 41918 14478 41970
rect 14530 41918 14542 41970
rect 2830 41906 2882 41918
rect 9774 41906 9826 41918
rect 10670 41906 10722 41918
rect 16158 41906 16210 41918
rect 17726 41970 17778 41982
rect 17726 41906 17778 41918
rect 18398 41970 18450 41982
rect 18398 41906 18450 41918
rect 18734 41970 18786 41982
rect 23102 41970 23154 41982
rect 19058 41918 19070 41970
rect 19122 41918 19134 41970
rect 19394 41918 19406 41970
rect 19458 41918 19470 41970
rect 21970 41918 21982 41970
rect 22034 41918 22046 41970
rect 18734 41906 18786 41918
rect 23102 41906 23154 41918
rect 24670 41970 24722 41982
rect 38670 41970 38722 41982
rect 25218 41918 25230 41970
rect 25282 41918 25294 41970
rect 29362 41918 29374 41970
rect 29426 41918 29438 41970
rect 30034 41918 30046 41970
rect 30098 41918 30110 41970
rect 31490 41918 31502 41970
rect 31554 41918 31566 41970
rect 33842 41918 33854 41970
rect 33906 41918 33918 41970
rect 35522 41918 35534 41970
rect 35586 41918 35598 41970
rect 24670 41906 24722 41918
rect 38670 41906 38722 41918
rect 39118 41970 39170 41982
rect 41234 41918 41246 41970
rect 41298 41918 41310 41970
rect 41458 41918 41470 41970
rect 41522 41918 41534 41970
rect 42242 41918 42254 41970
rect 42306 41918 42318 41970
rect 42802 41918 42814 41970
rect 42866 41918 42878 41970
rect 43810 41918 43822 41970
rect 43874 41918 43886 41970
rect 39118 41906 39170 41918
rect 16494 41858 16546 41870
rect 7522 41806 7534 41858
rect 7586 41806 7598 41858
rect 11778 41806 11790 41858
rect 11842 41806 11854 41858
rect 13906 41806 13918 41858
rect 13970 41806 13982 41858
rect 16494 41794 16546 41806
rect 19966 41858 20018 41870
rect 19966 41794 20018 41806
rect 23886 41858 23938 41870
rect 44606 41858 44658 41870
rect 26002 41806 26014 41858
rect 26066 41806 26078 41858
rect 28130 41806 28142 41858
rect 28194 41806 28206 41858
rect 30258 41806 30270 41858
rect 30322 41806 30334 41858
rect 31826 41806 31838 41858
rect 31890 41806 31902 41858
rect 33954 41806 33966 41858
rect 34018 41806 34030 41858
rect 35970 41806 35982 41858
rect 36034 41806 36046 41858
rect 43362 41806 43374 41858
rect 43426 41806 43438 41858
rect 23886 41794 23938 41806
rect 44606 41794 44658 41806
rect 2942 41746 2994 41758
rect 2942 41682 2994 41694
rect 18062 41746 18114 41758
rect 18062 41682 18114 41694
rect 22654 41746 22706 41758
rect 39342 41746 39394 41758
rect 40238 41746 40290 41758
rect 23650 41694 23662 41746
rect 23714 41743 23726 41746
rect 23874 41743 23886 41746
rect 23714 41697 23886 41743
rect 23714 41694 23726 41697
rect 23874 41694 23886 41697
rect 23938 41694 23950 41746
rect 39666 41694 39678 41746
rect 39730 41694 39742 41746
rect 41906 41694 41918 41746
rect 41970 41694 41982 41746
rect 43586 41694 43598 41746
rect 43650 41694 43662 41746
rect 22654 41682 22706 41694
rect 39342 41682 39394 41694
rect 40238 41682 40290 41694
rect 1344 41578 48608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48608 41578
rect 1344 41492 48608 41526
rect 25566 41410 25618 41422
rect 25566 41346 25618 41358
rect 27470 41410 27522 41422
rect 27470 41346 27522 41358
rect 27806 41410 27858 41422
rect 27806 41346 27858 41358
rect 36094 41410 36146 41422
rect 36094 41346 36146 41358
rect 44270 41410 44322 41422
rect 44270 41346 44322 41358
rect 45166 41410 45218 41422
rect 45166 41346 45218 41358
rect 11454 41298 11506 41310
rect 2482 41246 2494 41298
rect 2546 41246 2558 41298
rect 4610 41246 4622 41298
rect 4674 41246 4686 41298
rect 8418 41246 8430 41298
rect 8482 41246 8494 41298
rect 11454 41234 11506 41246
rect 13694 41298 13746 41310
rect 19966 41298 20018 41310
rect 15922 41246 15934 41298
rect 15986 41246 15998 41298
rect 17938 41246 17950 41298
rect 18002 41246 18014 41298
rect 13694 41234 13746 41246
rect 19966 41234 20018 41246
rect 20750 41298 20802 41310
rect 25790 41298 25842 41310
rect 22082 41246 22094 41298
rect 22146 41246 22158 41298
rect 24210 41246 24222 41298
rect 24274 41246 24286 41298
rect 20750 41234 20802 41246
rect 25790 41234 25842 41246
rect 28254 41298 28306 41310
rect 28254 41234 28306 41246
rect 29934 41298 29986 41310
rect 37102 41298 37154 41310
rect 44158 41298 44210 41310
rect 32386 41246 32398 41298
rect 32450 41246 32462 41298
rect 36306 41246 36318 41298
rect 36370 41246 36382 41298
rect 40450 41246 40462 41298
rect 40514 41246 40526 41298
rect 41682 41246 41694 41298
rect 41746 41246 41758 41298
rect 43810 41246 43822 41298
rect 43874 41246 43886 41298
rect 44818 41246 44830 41298
rect 44882 41246 44894 41298
rect 29934 41234 29986 41246
rect 37102 41234 37154 41246
rect 44158 41234 44210 41246
rect 11566 41186 11618 41198
rect 1810 41134 1822 41186
rect 1874 41134 1886 41186
rect 6514 41134 6526 41186
rect 6578 41134 6590 41186
rect 11566 41122 11618 41134
rect 11902 41186 11954 41198
rect 11902 41122 11954 41134
rect 12350 41186 12402 41198
rect 12350 41122 12402 41134
rect 12462 41186 12514 41198
rect 26798 41186 26850 41198
rect 14018 41134 14030 41186
rect 14082 41134 14094 41186
rect 19058 41134 19070 41186
rect 19122 41134 19134 41186
rect 21410 41134 21422 41186
rect 21474 41134 21486 41186
rect 24658 41134 24670 41186
rect 24722 41134 24734 41186
rect 25218 41134 25230 41186
rect 25282 41134 25294 41186
rect 12462 41122 12514 41134
rect 26798 41122 26850 41134
rect 26910 41186 26962 41198
rect 26910 41122 26962 41134
rect 29710 41186 29762 41198
rect 29710 41122 29762 41134
rect 30046 41186 30098 41198
rect 30706 41134 30718 41186
rect 30770 41134 30782 41186
rect 33282 41134 33294 41186
rect 33346 41134 33358 41186
rect 34402 41134 34414 41186
rect 34466 41134 34478 41186
rect 35634 41134 35646 41186
rect 35698 41134 35710 41186
rect 37538 41134 37550 41186
rect 37602 41134 37614 41186
rect 38322 41134 38334 41186
rect 38386 41134 38398 41186
rect 40898 41134 40910 41186
rect 40962 41134 40974 41186
rect 30046 41122 30098 41134
rect 11342 41074 11394 41086
rect 11342 41010 11394 41022
rect 12686 41074 12738 41086
rect 12686 41010 12738 41022
rect 27022 41074 27074 41086
rect 27022 41010 27074 41022
rect 27582 41074 27634 41086
rect 32162 41022 32174 41074
rect 32226 41022 32238 41074
rect 33058 41022 33070 41074
rect 33122 41022 33134 41074
rect 35522 41022 35534 41074
rect 35586 41022 35598 41074
rect 27582 41010 27634 41022
rect 5070 40962 5122 40974
rect 5070 40898 5122 40910
rect 12238 40962 12290 40974
rect 12238 40898 12290 40910
rect 24894 40962 24946 40974
rect 29262 40962 29314 40974
rect 26338 40910 26350 40962
rect 26402 40910 26414 40962
rect 24894 40898 24946 40910
rect 29262 40898 29314 40910
rect 29822 40962 29874 40974
rect 29822 40898 29874 40910
rect 30158 40962 30210 40974
rect 30158 40898 30210 40910
rect 34526 40962 34578 40974
rect 36318 40962 36370 40974
rect 34626 40910 34638 40962
rect 34690 40910 34702 40962
rect 34526 40898 34578 40910
rect 36318 40898 36370 40910
rect 44942 40962 44994 40974
rect 44942 40898 44994 40910
rect 1344 40794 48608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48608 40794
rect 1344 40708 48608 40742
rect 2494 40626 2546 40638
rect 2494 40562 2546 40574
rect 3614 40626 3666 40638
rect 3614 40562 3666 40574
rect 4398 40626 4450 40638
rect 4398 40562 4450 40574
rect 24670 40626 24722 40638
rect 40238 40626 40290 40638
rect 28914 40574 28926 40626
rect 28978 40574 28990 40626
rect 32498 40574 32510 40626
rect 32562 40574 32574 40626
rect 24670 40562 24722 40574
rect 40238 40562 40290 40574
rect 42814 40626 42866 40638
rect 42814 40562 42866 40574
rect 9550 40514 9602 40526
rect 17502 40514 17554 40526
rect 5618 40462 5630 40514
rect 5682 40462 5694 40514
rect 6290 40462 6302 40514
rect 6354 40462 6366 40514
rect 7970 40462 7982 40514
rect 8034 40462 8046 40514
rect 8306 40462 8318 40514
rect 8370 40462 8382 40514
rect 12226 40462 12238 40514
rect 12290 40462 12302 40514
rect 9550 40450 9602 40462
rect 17502 40450 17554 40462
rect 18734 40514 18786 40526
rect 18734 40450 18786 40462
rect 18958 40514 19010 40526
rect 18958 40450 19010 40462
rect 20526 40514 20578 40526
rect 20526 40450 20578 40462
rect 26462 40514 26514 40526
rect 26462 40450 26514 40462
rect 28478 40514 28530 40526
rect 31950 40514 32002 40526
rect 40350 40514 40402 40526
rect 29810 40462 29822 40514
rect 29874 40462 29886 40514
rect 33618 40462 33630 40514
rect 33682 40462 33694 40514
rect 34850 40462 34862 40514
rect 34914 40462 34926 40514
rect 40898 40462 40910 40514
rect 40962 40462 40974 40514
rect 44370 40462 44382 40514
rect 44434 40462 44446 40514
rect 28478 40450 28530 40462
rect 31950 40450 32002 40462
rect 40350 40450 40402 40462
rect 2718 40402 2770 40414
rect 2718 40338 2770 40350
rect 3166 40402 3218 40414
rect 11006 40402 11058 40414
rect 18174 40402 18226 40414
rect 21758 40402 21810 40414
rect 4834 40350 4846 40402
rect 4898 40350 4910 40402
rect 5506 40350 5518 40402
rect 5570 40350 5582 40402
rect 6402 40350 6414 40402
rect 6466 40350 6478 40402
rect 7074 40350 7086 40402
rect 7138 40350 7150 40402
rect 7634 40350 7646 40402
rect 7698 40350 7710 40402
rect 8418 40350 8430 40402
rect 8482 40350 8494 40402
rect 9986 40350 9998 40402
rect 10050 40350 10062 40402
rect 15362 40350 15374 40402
rect 15426 40350 15438 40402
rect 19170 40350 19182 40402
rect 19234 40350 19246 40402
rect 19954 40350 19966 40402
rect 20018 40350 20030 40402
rect 3166 40338 3218 40350
rect 11006 40338 11058 40350
rect 18174 40338 18226 40350
rect 21758 40338 21810 40350
rect 26910 40402 26962 40414
rect 26910 40338 26962 40350
rect 27358 40402 27410 40414
rect 27358 40338 27410 40350
rect 29486 40402 29538 40414
rect 30146 40350 30158 40402
rect 30210 40350 30222 40402
rect 33506 40350 33518 40402
rect 33570 40350 33582 40402
rect 34738 40350 34750 40402
rect 34802 40350 34814 40402
rect 36642 40350 36654 40402
rect 36706 40350 36718 40402
rect 37426 40350 37438 40402
rect 37490 40350 37502 40402
rect 38322 40350 38334 40402
rect 38386 40350 38398 40402
rect 38546 40350 38558 40402
rect 38610 40350 38622 40402
rect 39666 40350 39678 40402
rect 39730 40350 39742 40402
rect 41010 40350 41022 40402
rect 41074 40350 41086 40402
rect 43586 40350 43598 40402
rect 43650 40350 43662 40402
rect 29486 40338 29538 40350
rect 2158 40290 2210 40302
rect 2158 40226 2210 40238
rect 2606 40290 2658 40302
rect 2606 40226 2658 40238
rect 3726 40290 3778 40302
rect 21870 40290 21922 40302
rect 43262 40290 43314 40302
rect 9874 40238 9886 40290
rect 9938 40238 9950 40290
rect 35858 40238 35870 40290
rect 35922 40238 35934 40290
rect 39442 40238 39454 40290
rect 39506 40238 39518 40290
rect 41346 40238 41358 40290
rect 41410 40238 41422 40290
rect 46498 40238 46510 40290
rect 46562 40238 46574 40290
rect 3726 40226 3778 40238
rect 21870 40226 21922 40238
rect 43262 40226 43314 40238
rect 3838 40178 3890 40190
rect 3838 40114 3890 40126
rect 30718 40178 30770 40190
rect 30718 40114 30770 40126
rect 32174 40178 32226 40190
rect 32174 40114 32226 40126
rect 1344 40010 48608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48608 40010
rect 1344 39924 48608 39958
rect 30158 39842 30210 39854
rect 5058 39790 5070 39842
rect 5122 39790 5134 39842
rect 30158 39778 30210 39790
rect 38334 39842 38386 39854
rect 45054 39842 45106 39854
rect 39890 39839 39902 39842
rect 38334 39778 38386 39790
rect 39121 39793 39902 39839
rect 2830 39730 2882 39742
rect 2830 39666 2882 39678
rect 3838 39730 3890 39742
rect 3838 39666 3890 39678
rect 4510 39730 4562 39742
rect 13582 39730 13634 39742
rect 28142 39730 28194 39742
rect 5842 39678 5854 39730
rect 5906 39678 5918 39730
rect 10882 39678 10894 39730
rect 10946 39678 10958 39730
rect 16818 39678 16830 39730
rect 16882 39678 16894 39730
rect 17938 39678 17950 39730
rect 18002 39678 18014 39730
rect 20066 39678 20078 39730
rect 20130 39678 20142 39730
rect 4510 39666 4562 39678
rect 13582 39666 13634 39678
rect 28142 39666 28194 39678
rect 28590 39730 28642 39742
rect 28590 39666 28642 39678
rect 29374 39730 29426 39742
rect 29374 39666 29426 39678
rect 31278 39730 31330 39742
rect 31278 39666 31330 39678
rect 35198 39730 35250 39742
rect 35198 39666 35250 39678
rect 36430 39730 36482 39742
rect 36430 39666 36482 39678
rect 37102 39730 37154 39742
rect 37102 39666 37154 39678
rect 4734 39618 4786 39630
rect 21982 39618 22034 39630
rect 26126 39618 26178 39630
rect 1810 39566 1822 39618
rect 1874 39566 1886 39618
rect 5730 39566 5742 39618
rect 5794 39566 5806 39618
rect 6962 39566 6974 39618
rect 7026 39566 7038 39618
rect 7186 39566 7198 39618
rect 7250 39566 7262 39618
rect 12786 39566 12798 39618
rect 12850 39566 12862 39618
rect 13906 39566 13918 39618
rect 13970 39566 13982 39618
rect 17266 39566 17278 39618
rect 17330 39566 17342 39618
rect 23426 39566 23438 39618
rect 23490 39566 23502 39618
rect 25890 39566 25902 39618
rect 25954 39566 25966 39618
rect 4734 39554 4786 39566
rect 21982 39554 22034 39566
rect 26126 39554 26178 39566
rect 27246 39618 27298 39630
rect 33058 39566 33070 39618
rect 33122 39566 33134 39618
rect 33394 39566 33406 39618
rect 33458 39566 33470 39618
rect 37762 39566 37774 39618
rect 37826 39566 37838 39618
rect 27246 39554 27298 39566
rect 24222 39506 24274 39518
rect 5954 39454 5966 39506
rect 6018 39454 6030 39506
rect 14690 39454 14702 39506
rect 14754 39454 14766 39506
rect 23538 39454 23550 39506
rect 23602 39454 23614 39506
rect 24222 39442 24274 39454
rect 26238 39506 26290 39518
rect 26238 39442 26290 39454
rect 27358 39506 27410 39518
rect 27358 39442 27410 39454
rect 27582 39506 27634 39518
rect 27582 39442 27634 39454
rect 32510 39506 32562 39518
rect 32510 39442 32562 39454
rect 33966 39506 34018 39518
rect 39121 39506 39167 39793
rect 39890 39790 39902 39793
rect 39954 39790 39966 39842
rect 45054 39778 45106 39790
rect 39902 39730 39954 39742
rect 39902 39666 39954 39678
rect 40350 39730 40402 39742
rect 40350 39666 40402 39678
rect 40910 39730 40962 39742
rect 40910 39666 40962 39678
rect 41358 39730 41410 39742
rect 44270 39730 44322 39742
rect 42130 39678 42142 39730
rect 42194 39678 42206 39730
rect 41358 39666 41410 39678
rect 44270 39666 44322 39678
rect 46510 39730 46562 39742
rect 46510 39666 46562 39678
rect 44830 39618 44882 39630
rect 41458 39566 41470 39618
rect 41522 39566 41534 39618
rect 42578 39566 42590 39618
rect 42642 39566 42654 39618
rect 44830 39554 44882 39566
rect 46398 39618 46450 39630
rect 46398 39554 46450 39566
rect 45726 39506 45778 39518
rect 39106 39454 39118 39506
rect 39170 39454 39182 39506
rect 42914 39454 42926 39506
rect 42978 39454 42990 39506
rect 45378 39454 45390 39506
rect 45442 39454 45454 39506
rect 33966 39442 34018 39454
rect 45726 39442 45778 39454
rect 2046 39394 2098 39406
rect 2046 39330 2098 39342
rect 3278 39394 3330 39406
rect 3278 39330 3330 39342
rect 4286 39394 4338 39406
rect 4286 39330 4338 39342
rect 20526 39394 20578 39406
rect 20526 39330 20578 39342
rect 21422 39394 21474 39406
rect 26350 39394 26402 39406
rect 23650 39342 23662 39394
rect 23714 39342 23726 39394
rect 21422 39330 21474 39342
rect 26350 39330 26402 39342
rect 26462 39394 26514 39406
rect 26462 39330 26514 39342
rect 29934 39394 29986 39406
rect 29934 39330 29986 39342
rect 30046 39394 30098 39406
rect 30046 39330 30098 39342
rect 30718 39394 30770 39406
rect 30718 39330 30770 39342
rect 34974 39394 35026 39406
rect 34974 39330 35026 39342
rect 39454 39394 39506 39406
rect 39454 39330 39506 39342
rect 46062 39394 46114 39406
rect 46062 39330 46114 39342
rect 1344 39226 48608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48608 39226
rect 1344 39140 48608 39174
rect 2270 39058 2322 39070
rect 2270 38994 2322 39006
rect 2382 39058 2434 39070
rect 2382 38994 2434 39006
rect 2494 39058 2546 39070
rect 2494 38994 2546 39006
rect 3166 39058 3218 39070
rect 3166 38994 3218 39006
rect 10110 39058 10162 39070
rect 10110 38994 10162 39006
rect 10558 39058 10610 39070
rect 10558 38994 10610 39006
rect 11454 39058 11506 39070
rect 11454 38994 11506 39006
rect 15374 39058 15426 39070
rect 15374 38994 15426 39006
rect 16270 39058 16322 39070
rect 16270 38994 16322 39006
rect 20526 39058 20578 39070
rect 20526 38994 20578 39006
rect 21086 39058 21138 39070
rect 21086 38994 21138 39006
rect 21310 39058 21362 39070
rect 21310 38994 21362 39006
rect 21982 39058 22034 39070
rect 33182 39058 33234 39070
rect 31826 39006 31838 39058
rect 31890 39006 31902 39058
rect 21982 38994 22034 39006
rect 33182 38994 33234 39006
rect 33630 39058 33682 39070
rect 33630 38994 33682 39006
rect 34078 39058 34130 39070
rect 34078 38994 34130 39006
rect 38446 39058 38498 39070
rect 38446 38994 38498 39006
rect 38894 39058 38946 39070
rect 38894 38994 38946 39006
rect 41022 39058 41074 39070
rect 41022 38994 41074 39006
rect 41918 39058 41970 39070
rect 41918 38994 41970 39006
rect 42366 39058 42418 39070
rect 42366 38994 42418 39006
rect 43486 39058 43538 39070
rect 43486 38994 43538 39006
rect 3054 38946 3106 38958
rect 20862 38946 20914 38958
rect 39342 38946 39394 38958
rect 3938 38894 3950 38946
rect 4002 38894 4014 38946
rect 26450 38894 26462 38946
rect 26514 38894 26526 38946
rect 26786 38894 26798 38946
rect 26850 38894 26862 38946
rect 29586 38894 29598 38946
rect 29650 38894 29662 38946
rect 30482 38894 30494 38946
rect 30546 38894 30558 38946
rect 31938 38894 31950 38946
rect 32002 38894 32014 38946
rect 3054 38882 3106 38894
rect 20862 38882 20914 38894
rect 39342 38882 39394 38894
rect 1822 38834 1874 38846
rect 1822 38770 1874 38782
rect 2830 38834 2882 38846
rect 2830 38770 2882 38782
rect 3502 38834 3554 38846
rect 9662 38834 9714 38846
rect 15710 38834 15762 38846
rect 7522 38782 7534 38834
rect 7586 38782 7598 38834
rect 11778 38782 11790 38834
rect 11842 38782 11854 38834
rect 3502 38770 3554 38782
rect 9662 38770 9714 38782
rect 15710 38770 15762 38782
rect 16606 38834 16658 38846
rect 21534 38834 21586 38846
rect 17938 38782 17950 38834
rect 18002 38782 18014 38834
rect 16606 38770 16658 38782
rect 21534 38770 21586 38782
rect 21646 38834 21698 38846
rect 27358 38834 27410 38846
rect 39678 38834 39730 38846
rect 41470 38834 41522 38846
rect 26898 38782 26910 38834
rect 26962 38782 26974 38834
rect 28018 38782 28030 38834
rect 28082 38782 28094 38834
rect 30818 38782 30830 38834
rect 30882 38782 30894 38834
rect 32274 38782 32286 38834
rect 32338 38782 32350 38834
rect 37426 38782 37438 38834
rect 37490 38782 37502 38834
rect 40002 38782 40014 38834
rect 40066 38782 40078 38834
rect 21646 38770 21698 38782
rect 27358 38770 27410 38782
rect 39678 38770 39730 38782
rect 41470 38770 41522 38782
rect 11006 38722 11058 38734
rect 26350 38722 26402 38734
rect 38110 38722 38162 38734
rect 12562 38670 12574 38722
rect 12626 38670 12638 38722
rect 14690 38670 14702 38722
rect 14754 38670 14766 38722
rect 19170 38670 19182 38722
rect 19234 38670 19246 38722
rect 28690 38670 28702 38722
rect 28754 38670 28766 38722
rect 34626 38670 34638 38722
rect 34690 38670 34702 38722
rect 36754 38670 36766 38722
rect 36818 38670 36830 38722
rect 11006 38658 11058 38670
rect 26350 38658 26402 38670
rect 38110 38658 38162 38670
rect 42814 38722 42866 38734
rect 42814 38658 42866 38670
rect 9550 38610 9602 38622
rect 40014 38610 40066 38622
rect 10658 38558 10670 38610
rect 10722 38607 10734 38610
rect 11330 38607 11342 38610
rect 10722 38561 11342 38607
rect 10722 38558 10734 38561
rect 11330 38558 11342 38561
rect 11394 38558 11406 38610
rect 15922 38558 15934 38610
rect 15986 38607 15998 38610
rect 16146 38607 16158 38610
rect 15986 38561 16158 38607
rect 15986 38558 15998 38561
rect 16146 38558 16158 38561
rect 16210 38558 16222 38610
rect 41122 38558 41134 38610
rect 41186 38607 41198 38610
rect 41682 38607 41694 38610
rect 41186 38561 41694 38607
rect 41186 38558 41198 38561
rect 41682 38558 41694 38561
rect 41746 38607 41758 38610
rect 42466 38607 42478 38610
rect 41746 38561 42478 38607
rect 41746 38558 41758 38561
rect 42466 38558 42478 38561
rect 42530 38558 42542 38610
rect 9550 38546 9602 38558
rect 40014 38546 40066 38558
rect 1344 38442 48608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48608 38442
rect 1344 38356 48608 38390
rect 19966 38274 20018 38286
rect 43822 38274 43874 38286
rect 29250 38222 29262 38274
rect 29314 38271 29326 38274
rect 29922 38271 29934 38274
rect 29314 38225 29934 38271
rect 29314 38222 29326 38225
rect 29922 38222 29934 38225
rect 29986 38222 29998 38274
rect 19966 38210 20018 38222
rect 43822 38210 43874 38222
rect 10670 38162 10722 38174
rect 1698 38110 1710 38162
rect 1762 38110 1774 38162
rect 4050 38110 4062 38162
rect 4114 38110 4126 38162
rect 10670 38098 10722 38110
rect 12350 38162 12402 38174
rect 20190 38162 20242 38174
rect 28254 38162 28306 38174
rect 18386 38110 18398 38162
rect 18450 38110 18462 38162
rect 24210 38110 24222 38162
rect 24274 38110 24286 38162
rect 27234 38110 27246 38162
rect 27298 38110 27310 38162
rect 12350 38098 12402 38110
rect 20190 38098 20242 38110
rect 28254 38098 28306 38110
rect 29262 38162 29314 38174
rect 29262 38098 29314 38110
rect 29710 38162 29762 38174
rect 29710 38098 29762 38110
rect 30718 38162 30770 38174
rect 30718 38098 30770 38110
rect 35870 38162 35922 38174
rect 41358 38162 41410 38174
rect 37986 38110 37998 38162
rect 38050 38110 38062 38162
rect 40114 38110 40126 38162
rect 40178 38110 40190 38162
rect 35870 38098 35922 38110
rect 41358 38098 41410 38110
rect 4958 38050 5010 38062
rect 11454 38050 11506 38062
rect 1810 37998 1822 38050
rect 1874 37998 1886 38050
rect 2818 37998 2830 38050
rect 2882 37998 2894 38050
rect 3266 37998 3278 38050
rect 3330 37998 3342 38050
rect 4386 37998 4398 38050
rect 4450 37998 4462 38050
rect 6290 37998 6302 38050
rect 6354 37998 6366 38050
rect 7634 37998 7646 38050
rect 7698 37998 7710 38050
rect 9426 37998 9438 38050
rect 9490 37998 9502 38050
rect 4958 37986 5010 37998
rect 11454 37986 11506 37998
rect 11902 38050 11954 38062
rect 11902 37986 11954 37998
rect 12126 38050 12178 38062
rect 27582 38050 27634 38062
rect 36094 38050 36146 38062
rect 41918 38050 41970 38062
rect 15362 37998 15374 38050
rect 15426 37998 15438 38050
rect 21298 37998 21310 38050
rect 21362 37998 21374 38050
rect 27794 37998 27806 38050
rect 27858 37998 27870 38050
rect 33282 37998 33294 38050
rect 33346 37998 33358 38050
rect 33730 37998 33742 38050
rect 33794 37998 33806 38050
rect 37202 37998 37214 38050
rect 37266 37998 37278 38050
rect 40898 37998 40910 38050
rect 40962 37998 40974 38050
rect 12126 37986 12178 37998
rect 27582 37986 27634 37998
rect 36094 37986 36146 37998
rect 41918 37986 41970 37998
rect 42142 38050 42194 38062
rect 42142 37986 42194 37998
rect 42926 38050 42978 38062
rect 42926 37986 42978 37998
rect 2158 37938 2210 37950
rect 4622 37938 4674 37950
rect 11118 37938 11170 37950
rect 4274 37886 4286 37938
rect 4338 37886 4350 37938
rect 6514 37886 6526 37938
rect 6578 37886 6590 37938
rect 9986 37886 9998 37938
rect 10050 37886 10062 37938
rect 2158 37874 2210 37886
rect 4622 37874 4674 37886
rect 11118 37874 11170 37886
rect 12462 37938 12514 37950
rect 27246 37938 27298 37950
rect 22082 37886 22094 37938
rect 22146 37886 22158 37938
rect 12462 37874 12514 37886
rect 27246 37874 27298 37886
rect 31278 37938 31330 37950
rect 31278 37874 31330 37886
rect 32286 37938 32338 37950
rect 32286 37874 32338 37886
rect 34302 37938 34354 37950
rect 36990 37938 37042 37950
rect 36418 37886 36430 37938
rect 36482 37886 36494 37938
rect 34302 37874 34354 37886
rect 36990 37874 37042 37886
rect 42590 37938 42642 37950
rect 42590 37874 42642 37886
rect 44046 37938 44098 37950
rect 44046 37874 44098 37886
rect 2270 37826 2322 37838
rect 2270 37762 2322 37774
rect 2494 37826 2546 37838
rect 2494 37762 2546 37774
rect 4846 37826 4898 37838
rect 4846 37762 4898 37774
rect 5854 37826 5906 37838
rect 5854 37762 5906 37774
rect 11342 37826 11394 37838
rect 11342 37762 11394 37774
rect 11566 37826 11618 37838
rect 11566 37762 11618 37774
rect 12910 37826 12962 37838
rect 12910 37762 12962 37774
rect 13582 37826 13634 37838
rect 20750 37826 20802 37838
rect 19618 37774 19630 37826
rect 19682 37774 19694 37826
rect 13582 37762 13634 37774
rect 20750 37762 20802 37774
rect 27358 37826 27410 37838
rect 27358 37762 27410 37774
rect 30158 37826 30210 37838
rect 30158 37762 30210 37774
rect 34974 37826 35026 37838
rect 34974 37762 35026 37774
rect 42366 37826 42418 37838
rect 42366 37762 42418 37774
rect 42702 37826 42754 37838
rect 42702 37762 42754 37774
rect 43038 37826 43090 37838
rect 43038 37762 43090 37774
rect 43150 37826 43202 37838
rect 43150 37762 43202 37774
rect 43374 37826 43426 37838
rect 43374 37762 43426 37774
rect 43934 37826 43986 37838
rect 43934 37762 43986 37774
rect 1344 37658 48608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48608 37658
rect 1344 37572 48608 37606
rect 5182 37490 5234 37502
rect 5182 37426 5234 37438
rect 5630 37490 5682 37502
rect 5630 37426 5682 37438
rect 9886 37490 9938 37502
rect 17950 37490 18002 37502
rect 26126 37490 26178 37502
rect 16146 37438 16158 37490
rect 16210 37438 16222 37490
rect 21186 37438 21198 37490
rect 21250 37438 21262 37490
rect 9886 37426 9938 37438
rect 17950 37426 18002 37438
rect 26126 37426 26178 37438
rect 27022 37490 27074 37502
rect 27022 37426 27074 37438
rect 28142 37490 28194 37502
rect 30606 37490 30658 37502
rect 29586 37438 29598 37490
rect 29650 37438 29662 37490
rect 28142 37426 28194 37438
rect 30606 37426 30658 37438
rect 30942 37490 30994 37502
rect 30942 37426 30994 37438
rect 32510 37490 32562 37502
rect 32510 37426 32562 37438
rect 36766 37490 36818 37502
rect 36766 37426 36818 37438
rect 41134 37490 41186 37502
rect 41570 37438 41582 37490
rect 41634 37438 41646 37490
rect 41134 37426 41186 37438
rect 8990 37378 9042 37390
rect 7186 37326 7198 37378
rect 7250 37326 7262 37378
rect 7522 37326 7534 37378
rect 7586 37326 7598 37378
rect 8990 37314 9042 37326
rect 9662 37378 9714 37390
rect 9662 37314 9714 37326
rect 9774 37378 9826 37390
rect 9774 37314 9826 37326
rect 19070 37378 19122 37390
rect 19070 37314 19122 37326
rect 19406 37378 19458 37390
rect 19406 37314 19458 37326
rect 26350 37378 26402 37390
rect 26350 37314 26402 37326
rect 27358 37378 27410 37390
rect 27358 37314 27410 37326
rect 29262 37378 29314 37390
rect 31838 37378 31890 37390
rect 42590 37378 42642 37390
rect 29474 37326 29486 37378
rect 29538 37326 29550 37378
rect 33954 37326 33966 37378
rect 34018 37326 34030 37378
rect 34738 37326 34750 37378
rect 34802 37326 34814 37378
rect 29262 37314 29314 37326
rect 31838 37314 31890 37326
rect 42590 37314 42642 37326
rect 44046 37378 44098 37390
rect 44046 37314 44098 37326
rect 8542 37266 8594 37278
rect 2146 37214 2158 37266
rect 2210 37214 2222 37266
rect 6066 37214 6078 37266
rect 6130 37214 6142 37266
rect 6738 37214 6750 37266
rect 6802 37214 6814 37266
rect 7858 37214 7870 37266
rect 7922 37214 7934 37266
rect 8542 37202 8594 37214
rect 8654 37266 8706 37278
rect 8654 37202 8706 37214
rect 10334 37266 10386 37278
rect 26462 37266 26514 37278
rect 10546 37214 10558 37266
rect 10610 37214 10622 37266
rect 19730 37214 19742 37266
rect 19794 37214 19806 37266
rect 24658 37214 24670 37266
rect 24722 37214 24734 37266
rect 10334 37202 10386 37214
rect 26462 37202 26514 37214
rect 27918 37266 27970 37278
rect 31390 37266 31442 37278
rect 36206 37266 36258 37278
rect 28354 37214 28366 37266
rect 28418 37214 28430 37266
rect 28578 37214 28590 37266
rect 28642 37214 28654 37266
rect 29810 37214 29822 37266
rect 29874 37214 29886 37266
rect 33058 37214 33070 37266
rect 33122 37214 33134 37266
rect 27918 37202 27970 37214
rect 31390 37202 31442 37214
rect 36206 37202 36258 37214
rect 37662 37266 37714 37278
rect 37662 37202 37714 37214
rect 43150 37266 43202 37278
rect 43150 37202 43202 37214
rect 45166 37266 45218 37278
rect 45166 37202 45218 37214
rect 45726 37266 45778 37278
rect 45726 37202 45778 37214
rect 1934 37154 1986 37166
rect 8878 37154 8930 37166
rect 16718 37154 16770 37166
rect 3602 37102 3614 37154
rect 3666 37102 3678 37154
rect 14354 37102 14366 37154
rect 14418 37102 14430 37154
rect 1934 37090 1986 37102
rect 8878 37090 8930 37102
rect 16718 37090 16770 37102
rect 17502 37154 17554 37166
rect 17502 37090 17554 37102
rect 18734 37154 18786 37166
rect 25342 37154 25394 37166
rect 21746 37102 21758 37154
rect 21810 37102 21822 37154
rect 23874 37102 23886 37154
rect 23938 37102 23950 37154
rect 18734 37090 18786 37102
rect 25342 37090 25394 37102
rect 25902 37154 25954 37166
rect 37214 37154 37266 37166
rect 28242 37102 28254 37154
rect 28306 37102 28318 37154
rect 25902 37090 25954 37102
rect 37214 37090 37266 37102
rect 38110 37154 38162 37166
rect 38110 37090 38162 37102
rect 16494 37042 16546 37054
rect 16494 36978 16546 36990
rect 29710 37042 29762 37054
rect 29710 36978 29762 36990
rect 34414 37042 34466 37054
rect 45614 37042 45666 37054
rect 37090 36990 37102 37042
rect 37154 37039 37166 37042
rect 37426 37039 37438 37042
rect 37154 36993 37438 37039
rect 37154 36990 37166 36993
rect 37426 36990 37438 36993
rect 37490 37039 37502 37042
rect 38098 37039 38110 37042
rect 37490 36993 38110 37039
rect 37490 36990 37502 36993
rect 38098 36990 38110 36993
rect 38162 36990 38174 37042
rect 34414 36978 34466 36990
rect 45614 36978 45666 36990
rect 1344 36874 48608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48608 36874
rect 1344 36788 48608 36822
rect 2046 36706 2098 36718
rect 24894 36706 24946 36718
rect 3378 36654 3390 36706
rect 3442 36654 3454 36706
rect 2046 36642 2098 36654
rect 24894 36642 24946 36654
rect 27582 36706 27634 36718
rect 27582 36642 27634 36654
rect 27806 36706 27858 36718
rect 27806 36642 27858 36654
rect 38110 36706 38162 36718
rect 38110 36642 38162 36654
rect 2382 36594 2434 36606
rect 2382 36530 2434 36542
rect 8094 36594 8146 36606
rect 32286 36594 32338 36606
rect 9202 36542 9214 36594
rect 9266 36542 9278 36594
rect 11330 36542 11342 36594
rect 11394 36542 11406 36594
rect 15698 36542 15710 36594
rect 15762 36542 15774 36594
rect 18610 36542 18622 36594
rect 18674 36542 18686 36594
rect 20738 36542 20750 36594
rect 20802 36542 20814 36594
rect 26114 36542 26126 36594
rect 26178 36542 26190 36594
rect 30818 36542 30830 36594
rect 30882 36542 30894 36594
rect 8094 36530 8146 36542
rect 32286 36530 32338 36542
rect 35422 36594 35474 36606
rect 35422 36530 35474 36542
rect 36990 36594 37042 36606
rect 36990 36530 37042 36542
rect 37998 36594 38050 36606
rect 37998 36530 38050 36542
rect 41358 36594 41410 36606
rect 43474 36542 43486 36594
rect 43538 36542 43550 36594
rect 45938 36542 45950 36594
rect 46002 36542 46014 36594
rect 48066 36542 48078 36594
rect 48130 36542 48142 36594
rect 41358 36530 41410 36542
rect 2942 36482 2994 36494
rect 25118 36482 25170 36494
rect 25790 36482 25842 36494
rect 3602 36430 3614 36482
rect 3666 36430 3678 36482
rect 6178 36430 6190 36482
rect 6242 36430 6254 36482
rect 6738 36430 6750 36482
rect 6802 36430 6814 36482
rect 8530 36430 8542 36482
rect 8594 36430 8606 36482
rect 14690 36430 14702 36482
rect 14754 36430 14766 36482
rect 17826 36430 17838 36482
rect 17890 36430 17902 36482
rect 25554 36430 25566 36482
rect 25618 36430 25630 36482
rect 2942 36418 2994 36430
rect 25118 36418 25170 36430
rect 25790 36418 25842 36430
rect 26910 36482 26962 36494
rect 29822 36482 29874 36494
rect 29586 36430 29598 36482
rect 29650 36430 29662 36482
rect 26910 36418 26962 36430
rect 29822 36418 29874 36430
rect 30158 36482 30210 36494
rect 35310 36482 35362 36494
rect 30930 36430 30942 36482
rect 30994 36430 31006 36482
rect 32610 36430 32622 36482
rect 32674 36430 32686 36482
rect 33618 36430 33630 36482
rect 33682 36430 33694 36482
rect 35074 36430 35086 36482
rect 35138 36430 35150 36482
rect 30158 36418 30210 36430
rect 35310 36418 35362 36430
rect 37214 36482 37266 36494
rect 37214 36418 37266 36430
rect 41134 36482 41186 36494
rect 41682 36430 41694 36482
rect 41746 36430 41758 36482
rect 45266 36430 45278 36482
rect 45330 36430 45342 36482
rect 41134 36418 41186 36430
rect 2606 36370 2658 36382
rect 17390 36370 17442 36382
rect 7186 36318 7198 36370
rect 7250 36318 7262 36370
rect 2606 36306 2658 36318
rect 17390 36306 17442 36318
rect 23774 36370 23826 36382
rect 23774 36306 23826 36318
rect 24110 36370 24162 36382
rect 26126 36370 26178 36382
rect 24546 36318 24558 36370
rect 24610 36318 24622 36370
rect 24110 36306 24162 36318
rect 26126 36306 26178 36318
rect 27246 36370 27298 36382
rect 27246 36306 27298 36318
rect 27470 36370 27522 36382
rect 27470 36306 27522 36318
rect 27918 36370 27970 36382
rect 27918 36306 27970 36318
rect 30270 36370 30322 36382
rect 35758 36370 35810 36382
rect 31602 36318 31614 36370
rect 31666 36318 31678 36370
rect 30270 36306 30322 36318
rect 35758 36306 35810 36318
rect 17054 36258 17106 36270
rect 6290 36206 6302 36258
rect 6354 36206 6366 36258
rect 17054 36194 17106 36206
rect 21422 36258 21474 36270
rect 21422 36194 21474 36206
rect 26014 36258 26066 36270
rect 26014 36194 26066 36206
rect 26686 36258 26738 36270
rect 26686 36194 26738 36206
rect 28366 36258 28418 36270
rect 35534 36258 35586 36270
rect 29250 36206 29262 36258
rect 29314 36206 29326 36258
rect 32946 36206 32958 36258
rect 33010 36206 33022 36258
rect 34626 36206 34638 36258
rect 34690 36206 34702 36258
rect 28366 36194 28418 36206
rect 35534 36194 35586 36206
rect 36206 36258 36258 36270
rect 40462 36258 40514 36270
rect 37538 36206 37550 36258
rect 37602 36206 37614 36258
rect 40786 36206 40798 36258
rect 40850 36206 40862 36258
rect 36206 36194 36258 36206
rect 40462 36194 40514 36206
rect 1344 36090 48608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48608 36090
rect 1344 36004 48608 36038
rect 2494 35922 2546 35934
rect 2494 35858 2546 35870
rect 2606 35922 2658 35934
rect 2606 35858 2658 35870
rect 3502 35922 3554 35934
rect 3502 35858 3554 35870
rect 6078 35922 6130 35934
rect 6078 35858 6130 35870
rect 10670 35922 10722 35934
rect 10670 35858 10722 35870
rect 12686 35922 12738 35934
rect 12686 35858 12738 35870
rect 28142 35922 28194 35934
rect 28142 35858 28194 35870
rect 31614 35922 31666 35934
rect 31614 35858 31666 35870
rect 32062 35922 32114 35934
rect 32062 35858 32114 35870
rect 41358 35922 41410 35934
rect 41358 35858 41410 35870
rect 2830 35810 2882 35822
rect 2830 35746 2882 35758
rect 5630 35810 5682 35822
rect 5630 35746 5682 35758
rect 6190 35810 6242 35822
rect 29598 35810 29650 35822
rect 18162 35758 18174 35810
rect 18226 35758 18238 35810
rect 6190 35746 6242 35758
rect 29598 35746 29650 35758
rect 30718 35810 30770 35822
rect 30718 35746 30770 35758
rect 37550 35810 37602 35822
rect 37550 35746 37602 35758
rect 37886 35810 37938 35822
rect 44034 35758 44046 35810
rect 44098 35758 44110 35810
rect 37886 35746 37938 35758
rect 2942 35698 2994 35710
rect 2942 35634 2994 35646
rect 5854 35698 5906 35710
rect 35198 35698 35250 35710
rect 11330 35646 11342 35698
rect 11394 35646 11406 35698
rect 19954 35646 19966 35698
rect 20018 35646 20030 35698
rect 30930 35646 30942 35698
rect 30994 35646 31006 35698
rect 31154 35646 31166 35698
rect 31218 35646 31230 35698
rect 43250 35646 43262 35698
rect 43314 35646 43326 35698
rect 5854 35634 5906 35646
rect 35198 35634 35250 35646
rect 8094 35586 8146 35598
rect 8094 35522 8146 35534
rect 8542 35586 8594 35598
rect 8542 35522 8594 35534
rect 15934 35586 15986 35598
rect 15934 35522 15986 35534
rect 16382 35586 16434 35598
rect 16382 35522 16434 35534
rect 16830 35586 16882 35598
rect 16830 35522 16882 35534
rect 20414 35586 20466 35598
rect 20414 35522 20466 35534
rect 25566 35586 25618 35598
rect 25566 35522 25618 35534
rect 30046 35586 30098 35598
rect 32510 35586 32562 35598
rect 30706 35534 30718 35586
rect 30770 35534 30782 35586
rect 30046 35522 30098 35534
rect 32510 35522 32562 35534
rect 34750 35586 34802 35598
rect 34750 35522 34802 35534
rect 35982 35586 36034 35598
rect 35982 35522 36034 35534
rect 36654 35586 36706 35598
rect 36654 35522 36706 35534
rect 42926 35586 42978 35598
rect 46162 35534 46174 35586
rect 46226 35534 46238 35586
rect 42926 35522 42978 35534
rect 34738 35422 34750 35474
rect 34802 35471 34814 35474
rect 34962 35471 34974 35474
rect 34802 35425 34974 35471
rect 34802 35422 34814 35425
rect 34962 35422 34974 35425
rect 35026 35422 35038 35474
rect 1344 35306 48608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48608 35306
rect 1344 35220 48608 35254
rect 2382 35138 2434 35150
rect 2382 35074 2434 35086
rect 4846 35138 4898 35150
rect 4846 35074 4898 35086
rect 18510 35138 18562 35150
rect 18510 35074 18562 35086
rect 12798 35026 12850 35038
rect 4162 34974 4174 35026
rect 4226 34974 4238 35026
rect 8754 34974 8766 35026
rect 8818 34974 8830 35026
rect 12798 34962 12850 34974
rect 17950 35026 18002 35038
rect 17950 34962 18002 34974
rect 19070 35026 19122 35038
rect 19070 34962 19122 34974
rect 19518 35026 19570 35038
rect 19518 34962 19570 34974
rect 25790 35026 25842 35038
rect 44942 35026 44994 35038
rect 37874 34974 37886 35026
rect 37938 34974 37950 35026
rect 40002 34974 40014 35026
rect 40066 34974 40078 35026
rect 25790 34962 25842 34974
rect 44942 34962 44994 34974
rect 8654 34914 8706 34926
rect 3042 34862 3054 34914
rect 3106 34862 3118 34914
rect 8654 34850 8706 34862
rect 10782 34914 10834 34926
rect 10782 34850 10834 34862
rect 11118 34914 11170 34926
rect 11118 34850 11170 34862
rect 11454 34914 11506 34926
rect 11454 34850 11506 34862
rect 11902 34914 11954 34926
rect 11902 34850 11954 34862
rect 12462 34914 12514 34926
rect 18846 34914 18898 34926
rect 14242 34862 14254 34914
rect 14306 34862 14318 34914
rect 12462 34850 12514 34862
rect 18846 34850 18898 34862
rect 30382 34914 30434 34926
rect 30382 34850 30434 34862
rect 32062 34914 32114 34926
rect 37202 34862 37214 34914
rect 37266 34862 37278 34914
rect 40786 34862 40798 34914
rect 40850 34862 40862 34914
rect 32062 34850 32114 34862
rect 3950 34802 4002 34814
rect 3950 34738 4002 34750
rect 4174 34802 4226 34814
rect 4174 34738 4226 34750
rect 4958 34802 5010 34814
rect 4958 34738 5010 34750
rect 6974 34802 7026 34814
rect 6974 34738 7026 34750
rect 21422 34802 21474 34814
rect 21422 34738 21474 34750
rect 21758 34802 21810 34814
rect 21758 34738 21810 34750
rect 31278 34802 31330 34814
rect 31278 34738 31330 34750
rect 34414 34802 34466 34814
rect 34414 34738 34466 34750
rect 4846 34690 4898 34702
rect 4846 34626 4898 34638
rect 6638 34690 6690 34702
rect 6638 34626 6690 34638
rect 7086 34690 7138 34702
rect 7086 34626 7138 34638
rect 7198 34690 7250 34702
rect 7198 34626 7250 34638
rect 7758 34690 7810 34702
rect 7758 34626 7810 34638
rect 8990 34690 9042 34702
rect 8990 34626 9042 34638
rect 10558 34690 10610 34702
rect 10558 34626 10610 34638
rect 11118 34690 11170 34702
rect 11118 34626 11170 34638
rect 11790 34690 11842 34702
rect 11790 34626 11842 34638
rect 12014 34690 12066 34702
rect 12014 34626 12066 34638
rect 13582 34690 13634 34702
rect 13582 34626 13634 34638
rect 27022 34690 27074 34702
rect 27022 34626 27074 34638
rect 27470 34690 27522 34702
rect 27470 34626 27522 34638
rect 27918 34690 27970 34702
rect 27918 34626 27970 34638
rect 29934 34690 29986 34702
rect 29934 34626 29986 34638
rect 31726 34690 31778 34702
rect 31726 34626 31778 34638
rect 34750 34690 34802 34702
rect 34750 34626 34802 34638
rect 36430 34690 36482 34702
rect 36430 34626 36482 34638
rect 40574 34690 40626 34702
rect 40574 34626 40626 34638
rect 1344 34522 48608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48608 34522
rect 1344 34436 48608 34470
rect 2830 34354 2882 34366
rect 2830 34290 2882 34302
rect 5854 34354 5906 34366
rect 5854 34290 5906 34302
rect 8766 34354 8818 34366
rect 39118 34354 39170 34366
rect 26114 34302 26126 34354
rect 26178 34302 26190 34354
rect 33618 34302 33630 34354
rect 33682 34302 33694 34354
rect 8766 34290 8818 34302
rect 39118 34290 39170 34302
rect 42702 34354 42754 34366
rect 42702 34290 42754 34302
rect 5630 34242 5682 34254
rect 4386 34190 4398 34242
rect 4450 34190 4462 34242
rect 4834 34190 4846 34242
rect 4898 34190 4910 34242
rect 5630 34178 5682 34190
rect 6302 34242 6354 34254
rect 25790 34242 25842 34254
rect 33070 34242 33122 34254
rect 39454 34242 39506 34254
rect 7634 34190 7646 34242
rect 7698 34190 7710 34242
rect 7970 34190 7982 34242
rect 8034 34190 8046 34242
rect 10770 34190 10782 34242
rect 10834 34190 10846 34242
rect 29250 34190 29262 34242
rect 29314 34190 29326 34242
rect 30146 34190 30158 34242
rect 30210 34190 30222 34242
rect 35410 34190 35422 34242
rect 35474 34190 35486 34242
rect 6302 34178 6354 34190
rect 25790 34178 25842 34190
rect 33070 34178 33122 34190
rect 39454 34178 39506 34190
rect 39678 34242 39730 34254
rect 39678 34178 39730 34190
rect 40238 34242 40290 34254
rect 40238 34178 40290 34190
rect 43038 34242 43090 34254
rect 43038 34178 43090 34190
rect 43262 34242 43314 34254
rect 43262 34178 43314 34190
rect 1934 34130 1986 34142
rect 1934 34066 1986 34078
rect 2158 34130 2210 34142
rect 5518 34130 5570 34142
rect 26462 34130 26514 34142
rect 40126 34130 40178 34142
rect 3938 34078 3950 34130
rect 4002 34078 4014 34130
rect 4722 34078 4734 34130
rect 4786 34078 4798 34130
rect 6850 34078 6862 34130
rect 6914 34078 6926 34130
rect 7074 34078 7086 34130
rect 7138 34078 7150 34130
rect 8306 34078 8318 34130
rect 8370 34078 8382 34130
rect 14354 34078 14366 34130
rect 14418 34078 14430 34130
rect 15922 34078 15934 34130
rect 15986 34078 15998 34130
rect 17602 34078 17614 34130
rect 17666 34078 17678 34130
rect 24546 34078 24558 34130
rect 24610 34078 24622 34130
rect 29362 34078 29374 34130
rect 29426 34078 29438 34130
rect 29698 34078 29710 34130
rect 29762 34078 29774 34130
rect 34626 34078 34638 34130
rect 34690 34078 34702 34130
rect 2158 34066 2210 34078
rect 5518 34066 5570 34078
rect 26462 34066 26514 34078
rect 40126 34066 40178 34078
rect 6078 34018 6130 34030
rect 4274 33966 4286 34018
rect 4338 33966 4350 34018
rect 6078 33954 6130 33966
rect 6190 34018 6242 34030
rect 19070 34018 19122 34030
rect 16370 33966 16382 34018
rect 16434 33966 16446 34018
rect 6190 33954 6242 33966
rect 19070 33954 19122 33966
rect 21422 34018 21474 34030
rect 26686 34018 26738 34030
rect 21746 33966 21758 34018
rect 21810 33966 21822 34018
rect 23874 33966 23886 34018
rect 23938 33966 23950 34018
rect 21422 33954 21474 33966
rect 26686 33954 26738 33966
rect 27134 34018 27186 34030
rect 32510 34018 32562 34030
rect 28802 33966 28814 34018
rect 28866 33966 28878 34018
rect 27134 33954 27186 33966
rect 32510 33954 32562 33966
rect 34302 34018 34354 34030
rect 37538 33966 37550 34018
rect 37602 33966 37614 34018
rect 34302 33954 34354 33966
rect 2382 33906 2434 33918
rect 2382 33842 2434 33854
rect 18398 33906 18450 33918
rect 18398 33842 18450 33854
rect 25230 33906 25282 33918
rect 25230 33842 25282 33854
rect 25566 33906 25618 33918
rect 25566 33842 25618 33854
rect 33294 33906 33346 33918
rect 33294 33842 33346 33854
rect 39790 33906 39842 33918
rect 39790 33842 39842 33854
rect 43374 33906 43426 33918
rect 43374 33842 43426 33854
rect 1344 33738 48608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48608 33738
rect 1344 33652 48608 33686
rect 8206 33570 8258 33582
rect 8206 33506 8258 33518
rect 14030 33570 14082 33582
rect 14030 33506 14082 33518
rect 14366 33570 14418 33582
rect 21646 33570 21698 33582
rect 44830 33570 44882 33582
rect 21298 33518 21310 33570
rect 21362 33518 21374 33570
rect 34178 33518 34190 33570
rect 34242 33518 34254 33570
rect 14366 33506 14418 33518
rect 21646 33506 21698 33518
rect 8094 33458 8146 33470
rect 20750 33458 20802 33470
rect 3602 33406 3614 33458
rect 3666 33406 3678 33458
rect 7410 33406 7422 33458
rect 7474 33406 7486 33458
rect 11442 33406 11454 33458
rect 11506 33406 11518 33458
rect 15810 33406 15822 33458
rect 15874 33406 15886 33458
rect 17938 33406 17950 33458
rect 18002 33406 18014 33458
rect 8094 33394 8146 33406
rect 20750 33394 20802 33406
rect 22542 33458 22594 33470
rect 22542 33394 22594 33406
rect 26574 33458 26626 33470
rect 26574 33394 26626 33406
rect 30270 33458 30322 33470
rect 33966 33458 34018 33470
rect 33506 33406 33518 33458
rect 33570 33406 33582 33458
rect 30270 33394 30322 33406
rect 33966 33394 34018 33406
rect 21870 33346 21922 33358
rect 2594 33294 2606 33346
rect 2658 33294 2670 33346
rect 4162 33294 4174 33346
rect 4226 33294 4238 33346
rect 6066 33294 6078 33346
rect 6130 33294 6142 33346
rect 6290 33294 6302 33346
rect 6354 33294 6366 33346
rect 7074 33294 7086 33346
rect 7138 33294 7150 33346
rect 8530 33294 8542 33346
rect 8594 33294 8606 33346
rect 15138 33294 15150 33346
rect 15202 33294 15214 33346
rect 21870 33282 21922 33294
rect 22766 33346 22818 33358
rect 22766 33282 22818 33294
rect 24222 33346 24274 33358
rect 24222 33282 24274 33294
rect 25230 33346 25282 33358
rect 28242 33294 28254 33346
rect 28306 33294 28318 33346
rect 30594 33294 30606 33346
rect 30658 33294 30670 33346
rect 25230 33282 25282 33294
rect 13806 33234 13858 33246
rect 3154 33182 3166 33234
rect 3218 33182 3230 33234
rect 7186 33182 7198 33234
rect 7250 33182 7262 33234
rect 9314 33182 9326 33234
rect 9378 33182 9390 33234
rect 13806 33170 13858 33182
rect 23438 33234 23490 33246
rect 23438 33170 23490 33182
rect 23774 33234 23826 33246
rect 27346 33182 27358 33234
rect 27410 33182 27422 33234
rect 31378 33182 31390 33234
rect 31442 33182 31454 33234
rect 23774 33170 23826 33182
rect 24894 33122 24946 33134
rect 23090 33070 23102 33122
rect 23154 33070 23166 33122
rect 24894 33058 24946 33070
rect 25566 33122 25618 33134
rect 25566 33058 25618 33070
rect 26126 33122 26178 33134
rect 27682 33070 27694 33122
rect 27746 33070 27758 33122
rect 34193 33119 34239 33518
rect 44830 33506 44882 33518
rect 44270 33458 44322 33470
rect 35746 33406 35758 33458
rect 35810 33406 35822 33458
rect 40002 33406 40014 33458
rect 40066 33406 40078 33458
rect 42130 33406 42142 33458
rect 42194 33406 42206 33458
rect 43362 33406 43374 33458
rect 43426 33406 43438 33458
rect 45154 33406 45166 33458
rect 45218 33406 45230 33458
rect 44270 33394 44322 33406
rect 34962 33294 34974 33346
rect 35026 33294 35038 33346
rect 39218 33294 39230 33346
rect 39282 33294 39294 33346
rect 42578 33294 42590 33346
rect 42642 33294 42654 33346
rect 43250 33294 43262 33346
rect 43314 33294 43326 33346
rect 43810 33182 43822 33234
rect 43874 33182 43886 33234
rect 34526 33122 34578 33134
rect 34402 33119 34414 33122
rect 34193 33073 34414 33119
rect 34402 33070 34414 33073
rect 34466 33070 34478 33122
rect 26126 33058 26178 33070
rect 34526 33058 34578 33070
rect 38894 33122 38946 33134
rect 38894 33058 38946 33070
rect 45054 33122 45106 33134
rect 45054 33058 45106 33070
rect 1344 32954 48608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48608 32954
rect 1344 32868 48608 32902
rect 7310 32786 7362 32798
rect 4498 32734 4510 32786
rect 4562 32734 4574 32786
rect 7310 32722 7362 32734
rect 7534 32786 7586 32798
rect 7534 32722 7586 32734
rect 8990 32786 9042 32798
rect 8990 32722 9042 32734
rect 9662 32786 9714 32798
rect 9662 32722 9714 32734
rect 10558 32786 10610 32798
rect 10558 32722 10610 32734
rect 10894 32786 10946 32798
rect 32510 32786 32562 32798
rect 29922 32734 29934 32786
rect 29986 32734 29998 32786
rect 10894 32722 10946 32734
rect 32510 32722 32562 32734
rect 34526 32786 34578 32798
rect 34526 32722 34578 32734
rect 42030 32786 42082 32798
rect 42030 32722 42082 32734
rect 42478 32786 42530 32798
rect 42478 32722 42530 32734
rect 2270 32674 2322 32686
rect 2270 32610 2322 32622
rect 3166 32674 3218 32686
rect 3166 32610 3218 32622
rect 6638 32674 6690 32686
rect 6638 32610 6690 32622
rect 10110 32674 10162 32686
rect 35870 32674 35922 32686
rect 42366 32674 42418 32686
rect 12226 32622 12238 32674
rect 12290 32622 12302 32674
rect 26002 32622 26014 32674
rect 26066 32622 26078 32674
rect 28578 32622 28590 32674
rect 28642 32622 28654 32674
rect 30034 32622 30046 32674
rect 30098 32622 30110 32674
rect 30594 32622 30606 32674
rect 30658 32622 30670 32674
rect 40114 32622 40126 32674
rect 40178 32622 40190 32674
rect 43810 32622 43822 32674
rect 43874 32622 43886 32674
rect 10110 32610 10162 32622
rect 35870 32610 35922 32622
rect 42366 32610 42418 32622
rect 1710 32562 1762 32574
rect 4398 32562 4450 32574
rect 2594 32510 2606 32562
rect 2658 32510 2670 32562
rect 1710 32498 1762 32510
rect 4398 32498 4450 32510
rect 6190 32562 6242 32574
rect 6190 32498 6242 32510
rect 6302 32562 6354 32574
rect 6302 32498 6354 32510
rect 6526 32562 6578 32574
rect 6526 32498 6578 32510
rect 7086 32562 7138 32574
rect 7086 32498 7138 32510
rect 7198 32562 7250 32574
rect 7198 32498 7250 32510
rect 7422 32562 7474 32574
rect 7422 32498 7474 32510
rect 9550 32562 9602 32574
rect 9550 32498 9602 32510
rect 9774 32562 9826 32574
rect 9774 32498 9826 32510
rect 10446 32562 10498 32574
rect 10446 32498 10498 32510
rect 10670 32562 10722 32574
rect 35534 32562 35586 32574
rect 46398 32562 46450 32574
rect 11442 32510 11454 32562
rect 11506 32510 11518 32562
rect 17938 32510 17950 32562
rect 18002 32510 18014 32562
rect 25218 32510 25230 32562
rect 25282 32510 25294 32562
rect 28466 32510 28478 32562
rect 28530 32510 28542 32562
rect 30146 32510 30158 32562
rect 30210 32510 30222 32562
rect 30706 32510 30718 32562
rect 30770 32510 30782 32562
rect 31490 32510 31502 32562
rect 31554 32510 31566 32562
rect 31826 32510 31838 32562
rect 31890 32510 31902 32562
rect 38882 32510 38894 32562
rect 38946 32510 38958 32562
rect 39666 32510 39678 32562
rect 39730 32510 39742 32562
rect 43026 32510 43038 32562
rect 43090 32510 43102 32562
rect 10670 32498 10722 32510
rect 35534 32498 35586 32510
rect 46398 32498 46450 32510
rect 8206 32450 8258 32462
rect 14814 32450 14866 32462
rect 14354 32398 14366 32450
rect 14418 32398 14430 32450
rect 8206 32386 8258 32398
rect 14814 32386 14866 32398
rect 15486 32450 15538 32462
rect 15486 32386 15538 32398
rect 17502 32450 17554 32462
rect 24670 32450 24722 32462
rect 33182 32450 33234 32462
rect 18610 32398 18622 32450
rect 18674 32398 18686 32450
rect 20738 32398 20750 32450
rect 20802 32398 20814 32450
rect 28130 32398 28142 32450
rect 28194 32398 28206 32450
rect 17502 32386 17554 32398
rect 24670 32386 24722 32398
rect 33182 32386 33234 32398
rect 33742 32450 33794 32462
rect 33742 32386 33794 32398
rect 34078 32450 34130 32462
rect 39330 32398 39342 32450
rect 39394 32398 39406 32450
rect 45938 32398 45950 32450
rect 46002 32398 46014 32450
rect 34078 32386 34130 32398
rect 30494 32338 30546 32350
rect 30494 32274 30546 32286
rect 46286 32338 46338 32350
rect 46286 32274 46338 32286
rect 1344 32170 48608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48608 32170
rect 1344 32084 48608 32118
rect 28254 32002 28306 32014
rect 11106 31950 11118 32002
rect 11170 31999 11182 32002
rect 11330 31999 11342 32002
rect 11170 31953 11342 31999
rect 11170 31950 11182 31953
rect 11330 31950 11342 31953
rect 11394 31950 11406 32002
rect 28254 31938 28306 31950
rect 28590 32002 28642 32014
rect 38894 32002 38946 32014
rect 31490 31950 31502 32002
rect 31554 31950 31566 32002
rect 28590 31938 28642 31950
rect 38894 31938 38946 31950
rect 42590 32002 42642 32014
rect 42590 31938 42642 31950
rect 1822 31890 1874 31902
rect 1822 31826 1874 31838
rect 4734 31890 4786 31902
rect 4734 31826 4786 31838
rect 11342 31890 11394 31902
rect 11342 31826 11394 31838
rect 11678 31890 11730 31902
rect 11678 31826 11730 31838
rect 14590 31890 14642 31902
rect 14590 31826 14642 31838
rect 18286 31890 18338 31902
rect 18286 31826 18338 31838
rect 18510 31890 18562 31902
rect 18510 31826 18562 31838
rect 19966 31890 20018 31902
rect 29262 31890 29314 31902
rect 26226 31838 26238 31890
rect 26290 31838 26302 31890
rect 19966 31826 20018 31838
rect 29262 31826 29314 31838
rect 30046 31890 30098 31902
rect 30046 31826 30098 31838
rect 32734 31890 32786 31902
rect 44270 31890 44322 31902
rect 36306 31838 36318 31890
rect 36370 31838 36382 31890
rect 45602 31838 45614 31890
rect 45666 31838 45678 31890
rect 47730 31838 47742 31890
rect 47794 31838 47806 31890
rect 32734 31826 32786 31838
rect 44270 31826 44322 31838
rect 2494 31778 2546 31790
rect 3950 31778 4002 31790
rect 3266 31726 3278 31778
rect 3330 31726 3342 31778
rect 2494 31714 2546 31726
rect 3950 31714 4002 31726
rect 4398 31778 4450 31790
rect 26126 31778 26178 31790
rect 29486 31778 29538 31790
rect 19394 31726 19406 31778
rect 19458 31726 19470 31778
rect 26786 31726 26798 31778
rect 26850 31726 26862 31778
rect 27458 31726 27470 31778
rect 27522 31726 27534 31778
rect 27906 31726 27918 31778
rect 27970 31726 27982 31778
rect 4398 31714 4450 31726
rect 26126 31714 26178 31726
rect 29486 31714 29538 31726
rect 30158 31778 30210 31790
rect 38670 31778 38722 31790
rect 31042 31726 31054 31778
rect 31106 31726 31118 31778
rect 31602 31726 31614 31778
rect 31666 31726 31678 31778
rect 32050 31726 32062 31778
rect 32114 31726 32126 31778
rect 33394 31726 33406 31778
rect 33458 31726 33470 31778
rect 39330 31726 39342 31778
rect 39394 31726 39406 31778
rect 40114 31726 40126 31778
rect 40178 31726 40190 31778
rect 41906 31726 41918 31778
rect 41970 31726 41982 31778
rect 42690 31726 42702 31778
rect 42754 31726 42766 31778
rect 43138 31726 43150 31778
rect 43202 31726 43214 31778
rect 44818 31726 44830 31778
rect 44882 31726 44894 31778
rect 30158 31714 30210 31726
rect 38670 31714 38722 31726
rect 2718 31666 2770 31678
rect 2718 31602 2770 31614
rect 2942 31666 2994 31678
rect 2942 31602 2994 31614
rect 3726 31666 3778 31678
rect 3726 31602 3778 31614
rect 13470 31666 13522 31678
rect 13470 31602 13522 31614
rect 17278 31666 17330 31678
rect 17278 31602 17330 31614
rect 19182 31666 19234 31678
rect 19182 31602 19234 31614
rect 25678 31666 25730 31678
rect 28478 31666 28530 31678
rect 37662 31666 37714 31678
rect 26674 31614 26686 31666
rect 26738 31614 26750 31666
rect 30930 31614 30942 31666
rect 30994 31614 31006 31666
rect 34178 31614 34190 31666
rect 34242 31614 34254 31666
rect 38882 31614 38894 31666
rect 38946 31614 38958 31666
rect 41794 31614 41806 31666
rect 41858 31614 41870 31666
rect 25678 31602 25730 31614
rect 28478 31602 28530 31614
rect 37662 31602 37714 31614
rect 4062 31554 4114 31566
rect 4062 31490 4114 31502
rect 6862 31554 6914 31566
rect 6862 31490 6914 31502
rect 13806 31554 13858 31566
rect 13806 31490 13858 31502
rect 16942 31554 16994 31566
rect 25902 31554 25954 31566
rect 17938 31502 17950 31554
rect 18002 31502 18014 31554
rect 16942 31490 16994 31502
rect 25902 31490 25954 31502
rect 26238 31554 26290 31566
rect 26238 31490 26290 31502
rect 29934 31554 29986 31566
rect 29934 31490 29986 31502
rect 38110 31554 38162 31566
rect 38110 31490 38162 31502
rect 40574 31554 40626 31566
rect 40574 31490 40626 31502
rect 41246 31554 41298 31566
rect 41246 31490 41298 31502
rect 43710 31554 43762 31566
rect 43710 31490 43762 31502
rect 1344 31386 48608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48608 31386
rect 1344 31300 48608 31334
rect 3166 31218 3218 31230
rect 3166 31154 3218 31166
rect 5518 31218 5570 31230
rect 5518 31154 5570 31166
rect 6190 31218 6242 31230
rect 26574 31218 26626 31230
rect 30494 31218 30546 31230
rect 19058 31166 19070 31218
rect 19122 31166 19134 31218
rect 29698 31166 29710 31218
rect 29762 31166 29774 31218
rect 6190 31154 6242 31166
rect 26574 31154 26626 31166
rect 30494 31154 30546 31166
rect 31278 31218 31330 31230
rect 31278 31154 31330 31166
rect 32286 31218 32338 31230
rect 32286 31154 32338 31166
rect 31838 31106 31890 31118
rect 2594 31054 2606 31106
rect 2658 31103 2670 31106
rect 2930 31103 2942 31106
rect 2658 31057 2942 31103
rect 2658 31054 2670 31057
rect 2930 31054 2942 31057
rect 2994 31054 3006 31106
rect 14130 31054 14142 31106
rect 14194 31054 14206 31106
rect 31838 31042 31890 31054
rect 32510 31106 32562 31118
rect 36430 31106 36482 31118
rect 46398 31106 46450 31118
rect 33618 31054 33630 31106
rect 33682 31054 33694 31106
rect 34626 31054 34638 31106
rect 34690 31054 34702 31106
rect 37426 31054 37438 31106
rect 37490 31054 37502 31106
rect 43922 31054 43934 31106
rect 43986 31054 43998 31106
rect 32510 31042 32562 31054
rect 36430 31042 36482 31054
rect 46398 31042 46450 31054
rect 4174 30994 4226 31006
rect 2258 30942 2270 30994
rect 2322 30942 2334 30994
rect 3154 30942 3166 30994
rect 3218 30942 3230 30994
rect 4174 30930 4226 30942
rect 4622 30994 4674 31006
rect 4622 30930 4674 30942
rect 4846 30994 4898 31006
rect 5742 30994 5794 31006
rect 5170 30942 5182 30994
rect 5234 30942 5246 30994
rect 4846 30930 4898 30942
rect 5742 30930 5794 30942
rect 10670 30994 10722 31006
rect 19406 30994 19458 31006
rect 29150 30994 29202 31006
rect 32062 30994 32114 31006
rect 46286 30994 46338 31006
rect 14802 30942 14814 30994
rect 14866 30942 14878 30994
rect 20066 30942 20078 30994
rect 20130 30942 20142 30994
rect 31490 30942 31502 30994
rect 31554 30942 31566 30994
rect 33058 30942 33070 30994
rect 33122 30942 33134 30994
rect 34738 30942 34750 30994
rect 34802 30942 34814 30994
rect 36642 30942 36654 30994
rect 36706 30942 36718 30994
rect 43026 30942 43038 30994
rect 43090 30942 43102 30994
rect 43586 30942 43598 30994
rect 43650 30942 43662 30994
rect 44370 30942 44382 30994
rect 44434 30942 44446 30994
rect 45490 30942 45502 30994
rect 45554 30942 45566 30994
rect 10670 30930 10722 30942
rect 19406 30930 19458 30942
rect 29150 30930 29202 30942
rect 32062 30930 32114 30942
rect 46286 30930 46338 30942
rect 4062 30882 4114 30894
rect 4062 30818 4114 30830
rect 4734 30882 4786 30894
rect 4734 30818 4786 30830
rect 5630 30882 5682 30894
rect 5630 30818 5682 30830
rect 11454 30882 11506 30894
rect 15374 30882 15426 30894
rect 12002 30830 12014 30882
rect 12066 30830 12078 30882
rect 11454 30818 11506 30830
rect 15374 30818 15426 30830
rect 18734 30882 18786 30894
rect 18734 30818 18786 30830
rect 19630 30882 19682 30894
rect 28814 30882 28866 30894
rect 41470 30882 41522 30894
rect 20738 30830 20750 30882
rect 20802 30830 20814 30882
rect 22866 30830 22878 30882
rect 22930 30830 22942 30882
rect 39554 30830 39566 30882
rect 39618 30830 39630 30882
rect 43362 30830 43374 30882
rect 43426 30830 43438 30882
rect 44706 30830 44718 30882
rect 44770 30830 44782 30882
rect 45042 30830 45054 30882
rect 45106 30830 45118 30882
rect 19630 30818 19682 30830
rect 28814 30818 28866 30830
rect 41470 30818 41522 30830
rect 2494 30770 2546 30782
rect 2494 30706 2546 30718
rect 10558 30770 10610 30782
rect 10558 30706 10610 30718
rect 29374 30770 29426 30782
rect 29374 30706 29426 30718
rect 31166 30770 31218 30782
rect 31166 30706 31218 30718
rect 32398 30770 32450 30782
rect 32398 30706 32450 30718
rect 1344 30602 48608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48608 30602
rect 1344 30516 48608 30550
rect 13470 30434 13522 30446
rect 6402 30382 6414 30434
rect 6466 30382 6478 30434
rect 13470 30370 13522 30382
rect 26238 30434 26290 30446
rect 33966 30434 34018 30446
rect 29474 30382 29486 30434
rect 29538 30382 29550 30434
rect 26238 30370 26290 30382
rect 33966 30370 34018 30382
rect 34190 30434 34242 30446
rect 34190 30370 34242 30382
rect 34526 30434 34578 30446
rect 34526 30370 34578 30382
rect 34862 30434 34914 30446
rect 34862 30370 34914 30382
rect 43150 30434 43202 30446
rect 43150 30370 43202 30382
rect 7534 30322 7586 30334
rect 3714 30270 3726 30322
rect 3778 30270 3790 30322
rect 6178 30270 6190 30322
rect 6242 30270 6254 30322
rect 7534 30258 7586 30270
rect 14478 30322 14530 30334
rect 14478 30258 14530 30270
rect 15150 30322 15202 30334
rect 19854 30322 19906 30334
rect 26574 30322 26626 30334
rect 18386 30270 18398 30322
rect 18450 30270 18462 30322
rect 25218 30270 25230 30322
rect 25282 30270 25294 30322
rect 15150 30258 15202 30270
rect 19854 30258 19906 30270
rect 26574 30258 26626 30270
rect 33742 30322 33794 30334
rect 33742 30258 33794 30270
rect 40798 30322 40850 30334
rect 40798 30258 40850 30270
rect 41246 30322 41298 30334
rect 41246 30258 41298 30270
rect 13806 30210 13858 30222
rect 31726 30210 31778 30222
rect 2930 30158 2942 30210
rect 2994 30158 3006 30210
rect 4050 30158 4062 30210
rect 4114 30158 4126 30210
rect 5954 30158 5966 30210
rect 6018 30158 6030 30210
rect 6290 30158 6302 30210
rect 6354 30158 6366 30210
rect 7970 30158 7982 30210
rect 8034 30158 8046 30210
rect 11778 30158 11790 30210
rect 11842 30158 11854 30210
rect 15586 30158 15598 30210
rect 15650 30158 15662 30210
rect 16258 30158 16270 30210
rect 16322 30158 16334 30210
rect 21522 30158 21534 30210
rect 21586 30158 21598 30210
rect 22306 30158 22318 30210
rect 22370 30158 22382 30210
rect 25890 30158 25902 30210
rect 25954 30158 25966 30210
rect 30034 30158 30046 30210
rect 30098 30158 30110 30210
rect 13806 30146 13858 30158
rect 31726 30146 31778 30158
rect 35758 30210 35810 30222
rect 35758 30146 35810 30158
rect 36206 30210 36258 30222
rect 36206 30146 36258 30158
rect 40350 30210 40402 30222
rect 44942 30210 44994 30222
rect 41570 30158 41582 30210
rect 41634 30158 41646 30210
rect 42466 30158 42478 30210
rect 42530 30158 42542 30210
rect 42802 30158 42814 30210
rect 42866 30158 42878 30210
rect 40350 30146 40402 30158
rect 44942 30146 44994 30158
rect 4958 30098 5010 30110
rect 2818 30046 2830 30098
rect 2882 30046 2894 30098
rect 4162 30046 4174 30098
rect 4226 30046 4238 30098
rect 4958 30034 5010 30046
rect 7422 30098 7474 30110
rect 7422 30034 7474 30046
rect 7646 30098 7698 30110
rect 7646 30034 7698 30046
rect 10222 30098 10274 30110
rect 10222 30034 10274 30046
rect 10670 30098 10722 30110
rect 10670 30034 10722 30046
rect 11118 30098 11170 30110
rect 11118 30034 11170 30046
rect 12126 30098 12178 30110
rect 12126 30034 12178 30046
rect 14030 30098 14082 30110
rect 14030 30034 14082 30046
rect 21310 30098 21362 30110
rect 25678 30098 25730 30110
rect 33518 30098 33570 30110
rect 23090 30046 23102 30098
rect 23154 30046 23166 30098
rect 30818 30046 30830 30098
rect 30882 30046 30894 30098
rect 21310 30034 21362 30046
rect 25678 30034 25730 30046
rect 33518 30034 33570 30046
rect 35310 30098 35362 30110
rect 41682 30046 41694 30098
rect 41746 30046 41758 30098
rect 35310 30034 35362 30046
rect 9886 29986 9938 29998
rect 9886 29922 9938 29934
rect 11006 29986 11058 29998
rect 11006 29922 11058 29934
rect 12238 29986 12290 29998
rect 12238 29922 12290 29934
rect 12350 29986 12402 29998
rect 12350 29922 12402 29934
rect 12798 29986 12850 29998
rect 12798 29922 12850 29934
rect 26126 29986 26178 29998
rect 26126 29922 26178 29934
rect 27134 29986 27186 29998
rect 27134 29922 27186 29934
rect 28590 29986 28642 29998
rect 33294 29986 33346 29998
rect 32610 29934 32622 29986
rect 32674 29934 32686 29986
rect 28590 29922 28642 29934
rect 33294 29922 33346 29934
rect 33406 29986 33458 29998
rect 33406 29922 33458 29934
rect 34638 29986 34690 29998
rect 34638 29922 34690 29934
rect 37102 29986 37154 29998
rect 37102 29922 37154 29934
rect 1344 29818 48608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48608 29818
rect 1344 29732 48608 29766
rect 5630 29650 5682 29662
rect 5630 29586 5682 29598
rect 5742 29650 5794 29662
rect 5742 29586 5794 29598
rect 6862 29650 6914 29662
rect 6862 29586 6914 29598
rect 6974 29650 7026 29662
rect 6974 29586 7026 29598
rect 8206 29650 8258 29662
rect 8206 29586 8258 29598
rect 9886 29650 9938 29662
rect 26462 29650 26514 29662
rect 32174 29650 32226 29662
rect 10658 29598 10670 29650
rect 10722 29598 10734 29650
rect 20962 29598 20974 29650
rect 21026 29598 21038 29650
rect 27122 29598 27134 29650
rect 27186 29598 27198 29650
rect 9886 29586 9938 29598
rect 26462 29586 26514 29598
rect 32174 29586 32226 29598
rect 33182 29650 33234 29662
rect 33182 29586 33234 29598
rect 33630 29650 33682 29662
rect 33630 29586 33682 29598
rect 34078 29650 34130 29662
rect 34078 29586 34130 29598
rect 34974 29650 35026 29662
rect 34974 29586 35026 29598
rect 35534 29650 35586 29662
rect 35534 29586 35586 29598
rect 36654 29650 36706 29662
rect 36654 29586 36706 29598
rect 38110 29650 38162 29662
rect 38110 29586 38162 29598
rect 40910 29650 40962 29662
rect 40910 29586 40962 29598
rect 41918 29650 41970 29662
rect 41918 29586 41970 29598
rect 42366 29650 42418 29662
rect 42366 29586 42418 29598
rect 43038 29650 43090 29662
rect 43038 29586 43090 29598
rect 7646 29538 7698 29550
rect 11230 29538 11282 29550
rect 3042 29486 3054 29538
rect 3106 29486 3118 29538
rect 10546 29486 10558 29538
rect 10610 29486 10622 29538
rect 7646 29474 7698 29486
rect 11230 29474 11282 29486
rect 13358 29538 13410 29550
rect 17390 29538 17442 29550
rect 16034 29486 16046 29538
rect 16098 29486 16110 29538
rect 13358 29474 13410 29486
rect 17390 29474 17442 29486
rect 21422 29538 21474 29550
rect 29710 29538 29762 29550
rect 27010 29486 27022 29538
rect 27074 29486 27086 29538
rect 21422 29474 21474 29486
rect 29710 29474 29762 29486
rect 32398 29538 32450 29550
rect 32398 29474 32450 29486
rect 39230 29538 39282 29550
rect 45166 29538 45218 29550
rect 43138 29486 43150 29538
rect 43202 29486 43214 29538
rect 39230 29474 39282 29486
rect 45166 29474 45218 29486
rect 5070 29426 5122 29438
rect 2258 29374 2270 29426
rect 2322 29374 2334 29426
rect 4162 29374 4174 29426
rect 4226 29374 4238 29426
rect 5070 29362 5122 29374
rect 5518 29426 5570 29438
rect 5518 29362 5570 29374
rect 6414 29426 6466 29438
rect 6414 29362 6466 29374
rect 7086 29426 7138 29438
rect 8542 29426 8594 29438
rect 8418 29374 8430 29426
rect 8482 29374 8494 29426
rect 7086 29362 7138 29374
rect 8542 29362 8594 29374
rect 8654 29426 8706 29438
rect 8654 29362 8706 29374
rect 8990 29426 9042 29438
rect 8990 29362 9042 29374
rect 9774 29426 9826 29438
rect 11006 29426 11058 29438
rect 13246 29426 13298 29438
rect 20638 29426 20690 29438
rect 10322 29374 10334 29426
rect 10386 29374 10398 29426
rect 11778 29374 11790 29426
rect 11842 29374 11854 29426
rect 12226 29374 12238 29426
rect 12290 29374 12302 29426
rect 12786 29374 12798 29426
rect 12850 29374 12862 29426
rect 16818 29374 16830 29426
rect 16882 29374 16894 29426
rect 17602 29374 17614 29426
rect 17666 29374 17678 29426
rect 9774 29362 9826 29374
rect 11006 29362 11058 29374
rect 13246 29362 13298 29374
rect 20638 29362 20690 29374
rect 26014 29426 26066 29438
rect 29150 29426 29202 29438
rect 28802 29374 28814 29426
rect 28866 29374 28878 29426
rect 26014 29362 26066 29374
rect 29150 29362 29202 29374
rect 31502 29426 31554 29438
rect 31502 29362 31554 29374
rect 31950 29426 32002 29438
rect 31950 29362 32002 29374
rect 34638 29426 34690 29438
rect 34638 29362 34690 29374
rect 41134 29426 41186 29438
rect 41134 29362 41186 29374
rect 41582 29426 41634 29438
rect 41582 29362 41634 29374
rect 42926 29426 42978 29438
rect 44830 29426 44882 29438
rect 43586 29374 43598 29426
rect 43650 29374 43662 29426
rect 44146 29374 44158 29426
rect 44210 29374 44222 29426
rect 45490 29374 45502 29426
rect 45554 29374 45566 29426
rect 42926 29362 42978 29374
rect 44830 29362 44882 29374
rect 1934 29314 1986 29326
rect 5294 29314 5346 29326
rect 20414 29314 20466 29326
rect 3826 29262 3838 29314
rect 3890 29262 3902 29314
rect 11890 29262 11902 29314
rect 11954 29262 11966 29314
rect 13906 29262 13918 29314
rect 13970 29262 13982 29314
rect 1934 29250 1986 29262
rect 5294 29250 5346 29262
rect 20414 29250 20466 29262
rect 21982 29314 22034 29326
rect 35870 29314 35922 29326
rect 32162 29262 32174 29314
rect 32226 29262 32238 29314
rect 21982 29250 22034 29262
rect 35870 29250 35922 29262
rect 38894 29314 38946 29326
rect 38894 29250 38946 29262
rect 41022 29314 41074 29326
rect 41022 29250 41074 29262
rect 9886 29202 9938 29214
rect 9886 29138 9938 29150
rect 10782 29202 10834 29214
rect 10782 29138 10834 29150
rect 31726 29202 31778 29214
rect 31726 29138 31778 29150
rect 39454 29202 39506 29214
rect 39454 29138 39506 29150
rect 39790 29202 39842 29214
rect 39790 29138 39842 29150
rect 45502 29202 45554 29214
rect 45502 29138 45554 29150
rect 1344 29034 48608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48608 29034
rect 1344 28948 48608 28982
rect 16270 28866 16322 28878
rect 16270 28802 16322 28814
rect 16606 28866 16658 28878
rect 16606 28802 16658 28814
rect 30158 28866 30210 28878
rect 33518 28866 33570 28878
rect 31378 28814 31390 28866
rect 31442 28863 31454 28866
rect 31714 28863 31726 28866
rect 31442 28817 31726 28863
rect 31442 28814 31454 28817
rect 31714 28814 31726 28817
rect 31778 28814 31790 28866
rect 30158 28802 30210 28814
rect 33518 28802 33570 28814
rect 33966 28866 34018 28878
rect 33966 28802 34018 28814
rect 36206 28866 36258 28878
rect 36206 28802 36258 28814
rect 6638 28754 6690 28766
rect 3378 28702 3390 28754
rect 3442 28702 3454 28754
rect 6638 28690 6690 28702
rect 12686 28754 12738 28766
rect 12686 28690 12738 28702
rect 17054 28754 17106 28766
rect 17054 28690 17106 28702
rect 17502 28754 17554 28766
rect 17502 28690 17554 28702
rect 24446 28754 24498 28766
rect 24446 28690 24498 28702
rect 25902 28754 25954 28766
rect 25902 28690 25954 28702
rect 26686 28754 26738 28766
rect 26686 28690 26738 28702
rect 27358 28754 27410 28766
rect 27358 28690 27410 28702
rect 27694 28754 27746 28766
rect 27694 28690 27746 28702
rect 28254 28754 28306 28766
rect 28254 28690 28306 28702
rect 29934 28754 29986 28766
rect 29934 28690 29986 28702
rect 31166 28754 31218 28766
rect 31166 28690 31218 28702
rect 31726 28754 31778 28766
rect 31726 28690 31778 28702
rect 32622 28754 32674 28766
rect 32622 28690 32674 28702
rect 33294 28754 33346 28766
rect 33294 28690 33346 28702
rect 33742 28754 33794 28766
rect 33742 28690 33794 28702
rect 38110 28754 38162 28766
rect 41694 28754 41746 28766
rect 38434 28702 38446 28754
rect 38498 28702 38510 28754
rect 40562 28702 40574 28754
rect 40626 28702 40638 28754
rect 38110 28690 38162 28702
rect 41694 28690 41746 28702
rect 42926 28754 42978 28766
rect 42926 28690 42978 28702
rect 43374 28754 43426 28766
rect 43374 28690 43426 28702
rect 43822 28754 43874 28766
rect 45714 28702 45726 28754
rect 45778 28702 45790 28754
rect 47842 28702 47854 28754
rect 47906 28702 47918 28754
rect 43822 28690 43874 28702
rect 6190 28642 6242 28654
rect 13582 28642 13634 28654
rect 34414 28642 34466 28654
rect 2930 28590 2942 28642
rect 2994 28590 3006 28642
rect 4162 28590 4174 28642
rect 4226 28590 4238 28642
rect 6962 28590 6974 28642
rect 7026 28590 7038 28642
rect 23538 28590 23550 28642
rect 23602 28590 23614 28642
rect 30594 28590 30606 28642
rect 30658 28590 30670 28642
rect 6190 28578 6242 28590
rect 13582 28578 13634 28590
rect 34414 28578 34466 28590
rect 34862 28642 34914 28654
rect 34862 28578 34914 28590
rect 35422 28642 35474 28654
rect 35422 28578 35474 28590
rect 35982 28642 36034 28654
rect 35982 28578 36034 28590
rect 36878 28642 36930 28654
rect 36878 28578 36930 28590
rect 36990 28642 37042 28654
rect 36990 28578 37042 28590
rect 37550 28642 37602 28654
rect 41806 28642 41858 28654
rect 41346 28590 41358 28642
rect 41410 28590 41422 28642
rect 37550 28578 37602 28590
rect 41806 28578 41858 28590
rect 42254 28642 42306 28654
rect 42254 28578 42306 28590
rect 42366 28642 42418 28654
rect 42366 28578 42418 28590
rect 44270 28642 44322 28654
rect 44930 28590 44942 28642
rect 44994 28590 45006 28642
rect 44270 28578 44322 28590
rect 1934 28530 1986 28542
rect 1934 28466 1986 28478
rect 2158 28530 2210 28542
rect 16046 28530 16098 28542
rect 3042 28478 3054 28530
rect 3106 28478 3118 28530
rect 10994 28478 11006 28530
rect 11058 28478 11070 28530
rect 2158 28466 2210 28478
rect 16046 28466 16098 28478
rect 23326 28530 23378 28542
rect 23326 28466 23378 28478
rect 30830 28530 30882 28542
rect 35310 28530 35362 28542
rect 31042 28478 31054 28530
rect 31106 28478 31118 28530
rect 30830 28466 30882 28478
rect 35310 28466 35362 28478
rect 35534 28530 35586 28542
rect 35534 28466 35586 28478
rect 36318 28530 36370 28542
rect 36318 28466 36370 28478
rect 2046 28418 2098 28430
rect 2046 28354 2098 28366
rect 27806 28418 27858 28430
rect 27806 28354 27858 28366
rect 32174 28418 32226 28430
rect 32174 28354 32226 28366
rect 37214 28418 37266 28430
rect 37214 28354 37266 28366
rect 37438 28418 37490 28430
rect 37438 28354 37490 28366
rect 42030 28418 42082 28430
rect 42030 28354 42082 28366
rect 1344 28250 48608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48608 28250
rect 1344 28164 48608 28198
rect 4398 28082 4450 28094
rect 10782 28082 10834 28094
rect 5170 28030 5182 28082
rect 5234 28030 5246 28082
rect 6290 28030 6302 28082
rect 6354 28030 6366 28082
rect 4398 28018 4450 28030
rect 10782 28018 10834 28030
rect 16270 28082 16322 28094
rect 16270 28018 16322 28030
rect 16830 28082 16882 28094
rect 16830 28018 16882 28030
rect 25678 28082 25730 28094
rect 25678 28018 25730 28030
rect 30158 28082 30210 28094
rect 30158 28018 30210 28030
rect 32286 28082 32338 28094
rect 32286 28018 32338 28030
rect 33182 28082 33234 28094
rect 33182 28018 33234 28030
rect 33630 28082 33682 28094
rect 33630 28018 33682 28030
rect 36878 28082 36930 28094
rect 36878 28018 36930 28030
rect 4734 27970 4786 27982
rect 8094 27970 8146 27982
rect 2818 27918 2830 27970
rect 2882 27918 2894 27970
rect 3714 27918 3726 27970
rect 3778 27918 3790 27970
rect 5954 27918 5966 27970
rect 6018 27918 6030 27970
rect 4734 27906 4786 27918
rect 8094 27906 8146 27918
rect 8878 27970 8930 27982
rect 25230 27970 25282 27982
rect 14130 27918 14142 27970
rect 14194 27918 14206 27970
rect 22754 27918 22766 27970
rect 22818 27918 22830 27970
rect 8878 27906 8930 27918
rect 25230 27906 25282 27918
rect 25790 27970 25842 27982
rect 29038 27970 29090 27982
rect 26562 27918 26574 27970
rect 26626 27918 26638 27970
rect 27010 27918 27022 27970
rect 27074 27918 27086 27970
rect 25790 27906 25842 27918
rect 29038 27906 29090 27918
rect 30494 27970 30546 27982
rect 30494 27906 30546 27918
rect 40014 27970 40066 27982
rect 40014 27906 40066 27918
rect 40350 27970 40402 27982
rect 40350 27906 40402 27918
rect 47294 27970 47346 27982
rect 47294 27906 47346 27918
rect 5070 27858 5122 27870
rect 8766 27858 8818 27870
rect 2146 27806 2158 27858
rect 2210 27806 2222 27858
rect 2706 27806 2718 27858
rect 2770 27806 2782 27858
rect 3826 27806 3838 27858
rect 3890 27806 3902 27858
rect 5282 27806 5294 27858
rect 5346 27806 5358 27858
rect 6290 27806 6302 27858
rect 6354 27806 6366 27858
rect 6850 27806 6862 27858
rect 6914 27806 6926 27858
rect 7410 27806 7422 27858
rect 7474 27806 7486 27858
rect 7746 27806 7758 27858
rect 7810 27806 7822 27858
rect 5070 27794 5122 27806
rect 8766 27794 8818 27806
rect 9102 27858 9154 27870
rect 24334 27858 24386 27870
rect 27470 27858 27522 27870
rect 9650 27806 9662 27858
rect 9714 27806 9726 27858
rect 10098 27806 10110 27858
rect 10162 27806 10174 27858
rect 11106 27806 11118 27858
rect 11170 27806 11182 27858
rect 13346 27806 13358 27858
rect 13410 27806 13422 27858
rect 15586 27806 15598 27858
rect 15650 27806 15662 27858
rect 17602 27806 17614 27858
rect 17666 27806 17678 27858
rect 23426 27806 23438 27858
rect 23490 27806 23502 27858
rect 25442 27806 25454 27858
rect 25506 27806 25518 27858
rect 9102 27794 9154 27806
rect 24334 27794 24386 27806
rect 27470 27794 27522 27806
rect 27694 27858 27746 27870
rect 37550 27858 37602 27870
rect 27906 27806 27918 27858
rect 27970 27806 27982 27858
rect 29922 27806 29934 27858
rect 29986 27806 29998 27858
rect 35074 27806 35086 27858
rect 35138 27806 35150 27858
rect 27694 27794 27746 27806
rect 37550 27794 37602 27806
rect 37774 27858 37826 27870
rect 41010 27806 41022 27858
rect 41074 27806 41086 27858
rect 37774 27794 37826 27806
rect 22206 27746 22258 27758
rect 3602 27694 3614 27746
rect 3666 27694 3678 27746
rect 12002 27694 12014 27746
rect 12066 27694 12078 27746
rect 13458 27694 13470 27746
rect 13522 27694 13534 27746
rect 15250 27694 15262 27746
rect 15314 27694 15326 27746
rect 18386 27694 18398 27746
rect 18450 27694 18462 27746
rect 20514 27694 20526 27746
rect 20578 27694 20590 27746
rect 22206 27682 22258 27694
rect 24670 27746 24722 27758
rect 24670 27682 24722 27694
rect 26126 27746 26178 27758
rect 26126 27682 26178 27694
rect 34414 27746 34466 27758
rect 34414 27682 34466 27694
rect 34750 27746 34802 27758
rect 34750 27682 34802 27694
rect 34862 27746 34914 27758
rect 34862 27682 34914 27694
rect 35534 27746 35586 27758
rect 35534 27682 35586 27694
rect 36430 27746 36482 27758
rect 36430 27682 36482 27694
rect 39678 27746 39730 27758
rect 41682 27694 41694 27746
rect 41746 27694 41758 27746
rect 43810 27694 43822 27746
rect 43874 27694 43886 27746
rect 39678 27682 39730 27694
rect 7758 27634 7810 27646
rect 47182 27634 47234 27646
rect 5282 27582 5294 27634
rect 5346 27582 5358 27634
rect 9650 27582 9662 27634
rect 9714 27582 9726 27634
rect 37202 27582 37214 27634
rect 37266 27582 37278 27634
rect 7758 27570 7810 27582
rect 47182 27570 47234 27582
rect 1344 27466 48608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48608 27466
rect 1344 27380 48608 27414
rect 5966 27298 6018 27310
rect 5966 27234 6018 27246
rect 6078 27298 6130 27310
rect 6078 27234 6130 27246
rect 6414 27298 6466 27310
rect 6414 27234 6466 27246
rect 10222 27298 10274 27310
rect 10222 27234 10274 27246
rect 10334 27298 10386 27310
rect 10334 27234 10386 27246
rect 10558 27298 10610 27310
rect 10558 27234 10610 27246
rect 10670 27298 10722 27310
rect 10670 27234 10722 27246
rect 23550 27298 23602 27310
rect 23550 27234 23602 27246
rect 23886 27298 23938 27310
rect 23886 27234 23938 27246
rect 26574 27298 26626 27310
rect 30606 27298 30658 27310
rect 27234 27246 27246 27298
rect 27298 27246 27310 27298
rect 30258 27246 30270 27298
rect 30322 27246 30334 27298
rect 26574 27234 26626 27246
rect 30606 27234 30658 27246
rect 3054 27186 3106 27198
rect 7422 27186 7474 27198
rect 4834 27134 4846 27186
rect 4898 27134 4910 27186
rect 3054 27122 3106 27134
rect 7422 27122 7474 27134
rect 11342 27186 11394 27198
rect 11342 27122 11394 27134
rect 14814 27186 14866 27198
rect 14814 27122 14866 27134
rect 23214 27186 23266 27198
rect 23214 27122 23266 27134
rect 24110 27186 24162 27198
rect 24110 27122 24162 27134
rect 25342 27186 25394 27198
rect 25342 27122 25394 27134
rect 25678 27186 25730 27198
rect 25678 27122 25730 27134
rect 26126 27186 26178 27198
rect 26126 27122 26178 27134
rect 28254 27186 28306 27198
rect 31838 27186 31890 27198
rect 29362 27134 29374 27186
rect 29426 27134 29438 27186
rect 28254 27122 28306 27134
rect 31838 27122 31890 27134
rect 32174 27186 32226 27198
rect 32174 27122 32226 27134
rect 32622 27186 32674 27198
rect 43038 27186 43090 27198
rect 34290 27134 34302 27186
rect 34354 27134 34366 27186
rect 36418 27134 36430 27186
rect 36482 27134 36494 27186
rect 36978 27134 36990 27186
rect 37042 27134 37054 27186
rect 40562 27134 40574 27186
rect 40626 27134 40638 27186
rect 32622 27122 32674 27134
rect 43038 27122 43090 27134
rect 43374 27186 43426 27198
rect 43374 27122 43426 27134
rect 2942 27074 2994 27086
rect 6302 27074 6354 27086
rect 3938 27022 3950 27074
rect 4002 27022 4014 27074
rect 2942 27010 2994 27022
rect 6302 27010 6354 27022
rect 7646 27074 7698 27086
rect 24558 27074 24610 27086
rect 7646 27010 7698 27022
rect 8206 27018 8258 27030
rect 21298 27022 21310 27074
rect 21362 27022 21374 27074
rect 22194 27022 22206 27074
rect 22258 27022 22270 27074
rect 3278 26962 3330 26974
rect 24558 27010 24610 27022
rect 25902 27074 25954 27086
rect 29486 27074 29538 27086
rect 27794 27022 27806 27074
rect 27858 27022 27870 27074
rect 28466 27022 28478 27074
rect 28530 27022 28542 27074
rect 29250 27022 29262 27074
rect 29314 27022 29326 27074
rect 25902 27010 25954 27022
rect 29486 27010 29538 27022
rect 30830 27074 30882 27086
rect 43598 27074 43650 27086
rect 33506 27022 33518 27074
rect 33570 27022 33582 27074
rect 39890 27022 39902 27074
rect 39954 27022 39966 27074
rect 30830 27010 30882 27022
rect 43598 27010 43650 27022
rect 3826 26910 3838 26962
rect 3890 26910 3902 26962
rect 8206 26954 8258 26966
rect 18062 26962 18114 26974
rect 3278 26898 3330 26910
rect 18062 26898 18114 26910
rect 18398 26962 18450 26974
rect 22542 26962 22594 26974
rect 29934 26962 29986 26974
rect 21410 26910 21422 26962
rect 21474 26910 21486 26962
rect 26898 26910 26910 26962
rect 26962 26910 26974 26962
rect 18398 26898 18450 26910
rect 22542 26898 22594 26910
rect 29934 26898 29986 26910
rect 31278 26962 31330 26974
rect 40238 26962 40290 26974
rect 39106 26910 39118 26962
rect 39170 26910 39182 26962
rect 31278 26898 31330 26910
rect 40238 26898 40290 26910
rect 40462 26962 40514 26974
rect 40462 26898 40514 26910
rect 7758 26850 7810 26862
rect 7758 26786 7810 26798
rect 7982 26850 8034 26862
rect 7982 26786 8034 26798
rect 8318 26850 8370 26862
rect 8318 26786 8370 26798
rect 8542 26850 8594 26862
rect 8542 26786 8594 26798
rect 9214 26850 9266 26862
rect 9214 26786 9266 26798
rect 9662 26850 9714 26862
rect 9662 26786 9714 26798
rect 11790 26850 11842 26862
rect 29710 26850 29762 26862
rect 22418 26798 22430 26850
rect 22482 26798 22494 26850
rect 11790 26786 11842 26798
rect 29710 26786 29762 26798
rect 33182 26850 33234 26862
rect 43922 26798 43934 26850
rect 43986 26798 43998 26850
rect 33182 26786 33234 26798
rect 1344 26682 48608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48608 26682
rect 1344 26596 48608 26630
rect 2158 26514 2210 26526
rect 2158 26450 2210 26462
rect 2606 26514 2658 26526
rect 6750 26514 6802 26526
rect 4050 26462 4062 26514
rect 4114 26462 4126 26514
rect 2606 26450 2658 26462
rect 6750 26450 6802 26462
rect 8206 26514 8258 26526
rect 8206 26450 8258 26462
rect 8878 26514 8930 26526
rect 25454 26514 25506 26526
rect 17714 26462 17726 26514
rect 17778 26462 17790 26514
rect 8878 26450 8930 26462
rect 25454 26450 25506 26462
rect 26014 26514 26066 26526
rect 26014 26450 26066 26462
rect 26686 26514 26738 26526
rect 26686 26450 26738 26462
rect 27806 26514 27858 26526
rect 27806 26450 27858 26462
rect 28478 26514 28530 26526
rect 28478 26450 28530 26462
rect 37662 26514 37714 26526
rect 37662 26450 37714 26462
rect 39902 26514 39954 26526
rect 39902 26450 39954 26462
rect 15150 26402 15202 26414
rect 7186 26350 7198 26402
rect 7250 26350 7262 26402
rect 14578 26350 14590 26402
rect 14642 26350 14654 26402
rect 15150 26338 15202 26350
rect 25566 26402 25618 26414
rect 25566 26338 25618 26350
rect 27582 26402 27634 26414
rect 27582 26338 27634 26350
rect 28814 26402 28866 26414
rect 28814 26338 28866 26350
rect 29038 26402 29090 26414
rect 29038 26338 29090 26350
rect 37326 26402 37378 26414
rect 37326 26338 37378 26350
rect 43822 26402 43874 26414
rect 43822 26338 43874 26350
rect 3502 26290 3554 26302
rect 2258 26238 2270 26290
rect 2322 26238 2334 26290
rect 3502 26226 3554 26238
rect 3726 26290 3778 26302
rect 7074 26238 7086 26290
rect 7138 26238 7150 26290
rect 15362 26238 15374 26290
rect 15426 26238 15438 26290
rect 21410 26238 21422 26290
rect 21474 26238 21486 26290
rect 32274 26238 32286 26290
rect 32338 26238 32350 26290
rect 33058 26238 33070 26290
rect 33122 26238 33134 26290
rect 44034 26238 44046 26290
rect 44098 26238 44110 26290
rect 3726 26226 3778 26238
rect 5630 26178 5682 26190
rect 3042 26126 3054 26178
rect 3106 26126 3118 26178
rect 5630 26114 5682 26126
rect 6190 26178 6242 26190
rect 6190 26114 6242 26126
rect 10894 26178 10946 26190
rect 10894 26114 10946 26126
rect 18286 26178 18338 26190
rect 18286 26114 18338 26126
rect 18734 26178 18786 26190
rect 18734 26114 18786 26126
rect 20974 26178 21026 26190
rect 36654 26178 36706 26190
rect 22082 26126 22094 26178
rect 22146 26126 22158 26178
rect 24210 26126 24222 26178
rect 24274 26126 24286 26178
rect 29138 26126 29150 26178
rect 29202 26126 29214 26178
rect 29474 26126 29486 26178
rect 29538 26126 29550 26178
rect 31602 26126 31614 26178
rect 31666 26126 31678 26178
rect 35186 26126 35198 26178
rect 35250 26126 35262 26178
rect 20974 26114 21026 26126
rect 36654 26114 36706 26126
rect 7870 26066 7922 26078
rect 7870 26002 7922 26014
rect 14030 26066 14082 26078
rect 14030 26002 14082 26014
rect 18062 26066 18114 26078
rect 18062 26002 18114 26014
rect 25454 26066 25506 26078
rect 25454 26002 25506 26014
rect 27918 26066 27970 26078
rect 27918 26002 27970 26014
rect 1344 25898 48608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48608 25898
rect 1344 25812 48608 25846
rect 10446 25730 10498 25742
rect 9202 25678 9214 25730
rect 9266 25727 9278 25730
rect 9426 25727 9438 25730
rect 9266 25681 9438 25727
rect 9266 25678 9278 25681
rect 9426 25678 9438 25681
rect 9490 25678 9502 25730
rect 10446 25666 10498 25678
rect 30494 25730 30546 25742
rect 30494 25666 30546 25678
rect 2382 25618 2434 25630
rect 2382 25554 2434 25566
rect 8990 25618 9042 25630
rect 8990 25554 9042 25566
rect 12574 25618 12626 25630
rect 28254 25618 28306 25630
rect 15138 25566 15150 25618
rect 15202 25566 15214 25618
rect 17266 25566 17278 25618
rect 17330 25566 17342 25618
rect 20626 25566 20638 25618
rect 20690 25566 20702 25618
rect 24546 25566 24558 25618
rect 24610 25566 24622 25618
rect 26674 25566 26686 25618
rect 26738 25566 26750 25618
rect 12574 25554 12626 25566
rect 28254 25554 28306 25566
rect 29262 25618 29314 25630
rect 29262 25554 29314 25566
rect 29710 25618 29762 25630
rect 29710 25554 29762 25566
rect 31950 25618 32002 25630
rect 31950 25554 32002 25566
rect 32398 25618 32450 25630
rect 32398 25554 32450 25566
rect 45390 25618 45442 25630
rect 45390 25554 45442 25566
rect 7982 25506 8034 25518
rect 7982 25442 8034 25454
rect 8542 25506 8594 25518
rect 23438 25506 23490 25518
rect 30270 25506 30322 25518
rect 10322 25454 10334 25506
rect 10386 25454 10398 25506
rect 11330 25454 11342 25506
rect 11394 25454 11406 25506
rect 11666 25454 11678 25506
rect 11730 25454 11742 25506
rect 14466 25454 14478 25506
rect 14530 25454 14542 25506
rect 17714 25454 17726 25506
rect 17778 25454 17790 25506
rect 23874 25454 23886 25506
rect 23938 25454 23950 25506
rect 8542 25442 8594 25454
rect 23438 25442 23490 25454
rect 30270 25442 30322 25454
rect 32622 25506 32674 25518
rect 32622 25442 32674 25454
rect 45166 25506 45218 25518
rect 45166 25442 45218 25454
rect 7870 25394 7922 25406
rect 10894 25394 10946 25406
rect 10658 25342 10670 25394
rect 10722 25342 10734 25394
rect 7870 25330 7922 25342
rect 10894 25330 10946 25342
rect 11230 25394 11282 25406
rect 21982 25394 22034 25406
rect 18498 25342 18510 25394
rect 18562 25342 18574 25394
rect 11230 25330 11282 25342
rect 21982 25330 22034 25342
rect 22318 25394 22370 25406
rect 31166 25394 31218 25406
rect 30818 25342 30830 25394
rect 30882 25342 30894 25394
rect 22318 25330 22370 25342
rect 31166 25330 31218 25342
rect 31502 25394 31554 25406
rect 31502 25330 31554 25342
rect 32958 25394 33010 25406
rect 32958 25330 33010 25342
rect 8094 25282 8146 25294
rect 8094 25218 8146 25230
rect 9326 25282 9378 25294
rect 9326 25218 9378 25230
rect 9774 25282 9826 25294
rect 9774 25218 9826 25230
rect 10110 25282 10162 25294
rect 10110 25218 10162 25230
rect 14030 25282 14082 25294
rect 14030 25218 14082 25230
rect 32846 25282 32898 25294
rect 32846 25218 32898 25230
rect 33406 25282 33458 25294
rect 33406 25218 33458 25230
rect 44270 25282 44322 25294
rect 44818 25230 44830 25282
rect 44882 25230 44894 25282
rect 44270 25218 44322 25230
rect 1344 25114 48608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48608 25114
rect 1344 25028 48608 25062
rect 2942 24946 2994 24958
rect 2942 24882 2994 24894
rect 4958 24946 5010 24958
rect 4958 24882 5010 24894
rect 6638 24946 6690 24958
rect 6638 24882 6690 24894
rect 7646 24946 7698 24958
rect 7646 24882 7698 24894
rect 16494 24946 16546 24958
rect 16494 24882 16546 24894
rect 17502 24946 17554 24958
rect 17502 24882 17554 24894
rect 18510 24946 18562 24958
rect 18510 24882 18562 24894
rect 29598 24946 29650 24958
rect 29598 24882 29650 24894
rect 37214 24946 37266 24958
rect 37214 24882 37266 24894
rect 42814 24946 42866 24958
rect 42814 24882 42866 24894
rect 8878 24834 8930 24846
rect 36654 24834 36706 24846
rect 3826 24782 3838 24834
rect 3890 24782 3902 24834
rect 4386 24782 4398 24834
rect 4450 24782 4462 24834
rect 5618 24782 5630 24834
rect 5682 24782 5694 24834
rect 5954 24782 5966 24834
rect 6018 24782 6030 24834
rect 10546 24782 10558 24834
rect 10610 24782 10622 24834
rect 12786 24782 12798 24834
rect 12850 24782 12862 24834
rect 8878 24770 8930 24782
rect 36654 24770 36706 24782
rect 42254 24834 42306 24846
rect 43922 24782 43934 24834
rect 43986 24782 43998 24834
rect 42254 24770 42306 24782
rect 7422 24722 7474 24734
rect 7422 24658 7474 24670
rect 7758 24722 7810 24734
rect 7758 24658 7810 24670
rect 8990 24722 9042 24734
rect 8990 24658 9042 24670
rect 9550 24722 9602 24734
rect 9550 24658 9602 24670
rect 9774 24722 9826 24734
rect 10098 24670 10110 24722
rect 10162 24670 10174 24722
rect 10770 24670 10782 24722
rect 10834 24670 10846 24722
rect 11890 24670 11902 24722
rect 11954 24670 11966 24722
rect 13234 24670 13246 24722
rect 13298 24670 13310 24722
rect 18274 24670 18286 24722
rect 18338 24670 18350 24722
rect 20962 24670 20974 24722
rect 21026 24670 21038 24722
rect 22306 24670 22318 24722
rect 22370 24670 22382 24722
rect 22978 24670 22990 24722
rect 23042 24670 23054 24722
rect 36418 24670 36430 24722
rect 36482 24670 36494 24722
rect 42018 24670 42030 24722
rect 42082 24670 42094 24722
rect 43250 24670 43262 24722
rect 43314 24670 43326 24722
rect 9774 24658 9826 24670
rect 7198 24610 7250 24622
rect 7198 24546 7250 24558
rect 8430 24610 8482 24622
rect 8430 24546 8482 24558
rect 9662 24610 9714 24622
rect 24670 24610 24722 24622
rect 13906 24558 13918 24610
rect 13970 24558 13982 24610
rect 16034 24558 16046 24610
rect 16098 24558 16110 24610
rect 19730 24558 19742 24610
rect 19794 24558 19806 24610
rect 23090 24558 23102 24610
rect 23154 24558 23166 24610
rect 9662 24546 9714 24558
rect 24670 24546 24722 24558
rect 25454 24610 25506 24622
rect 25454 24546 25506 24558
rect 30046 24610 30098 24622
rect 30046 24546 30098 24558
rect 32398 24610 32450 24622
rect 46050 24558 46062 24610
rect 46114 24558 46126 24610
rect 32398 24546 32450 24558
rect 4622 24498 4674 24510
rect 4622 24434 4674 24446
rect 6302 24498 6354 24510
rect 6302 24434 6354 24446
rect 8878 24498 8930 24510
rect 20178 24446 20190 24498
rect 20242 24446 20254 24498
rect 8878 24434 8930 24446
rect 1344 24330 48608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48608 24330
rect 1344 24244 48608 24278
rect 3950 24162 4002 24174
rect 3950 24098 4002 24110
rect 4286 24162 4338 24174
rect 21758 24162 21810 24174
rect 15138 24110 15150 24162
rect 15202 24110 15214 24162
rect 4286 24098 4338 24110
rect 21758 24098 21810 24110
rect 36990 24162 37042 24174
rect 42590 24162 42642 24174
rect 42242 24110 42254 24162
rect 42306 24110 42318 24162
rect 36990 24098 37042 24110
rect 42590 24098 42642 24110
rect 6750 24050 6802 24062
rect 13470 24050 13522 24062
rect 2370 23998 2382 24050
rect 2434 23998 2446 24050
rect 10770 23998 10782 24050
rect 10834 23998 10846 24050
rect 6750 23986 6802 23998
rect 13470 23986 13522 23998
rect 15710 24050 15762 24062
rect 15710 23986 15762 23998
rect 16830 24050 16882 24062
rect 16830 23986 16882 23998
rect 18510 24050 18562 24062
rect 18510 23986 18562 23998
rect 25342 24050 25394 24062
rect 25342 23986 25394 23998
rect 27022 24050 27074 24062
rect 27022 23986 27074 23998
rect 27694 24050 27746 24062
rect 27694 23986 27746 23998
rect 30942 24050 30994 24062
rect 30942 23986 30994 23998
rect 31950 24050 32002 24062
rect 31950 23986 32002 23998
rect 32510 24050 32562 24062
rect 41918 24050 41970 24062
rect 38546 23998 38558 24050
rect 38610 23998 38622 24050
rect 40674 23998 40686 24050
rect 40738 23998 40750 24050
rect 32510 23986 32562 23998
rect 41918 23986 41970 23998
rect 42814 24050 42866 24062
rect 47730 23998 47742 24050
rect 47794 23998 47806 24050
rect 42814 23986 42866 23998
rect 6190 23938 6242 23950
rect 7646 23938 7698 23950
rect 8766 23938 8818 23950
rect 13806 23938 13858 23950
rect 2258 23886 2270 23938
rect 2322 23886 2334 23938
rect 3378 23886 3390 23938
rect 3442 23886 3454 23938
rect 6514 23886 6526 23938
rect 6578 23886 6590 23938
rect 7410 23886 7422 23938
rect 7474 23886 7486 23938
rect 7858 23886 7870 23938
rect 7922 23886 7934 23938
rect 8530 23886 8542 23938
rect 8594 23886 8606 23938
rect 8978 23886 8990 23938
rect 9042 23886 9054 23938
rect 9874 23886 9886 23938
rect 9938 23886 9950 23938
rect 10882 23886 10894 23938
rect 10946 23886 10958 23938
rect 13570 23886 13582 23938
rect 13634 23886 13646 23938
rect 6190 23874 6242 23886
rect 7646 23874 7698 23886
rect 8766 23874 8818 23886
rect 13806 23874 13858 23886
rect 14814 23938 14866 23950
rect 14814 23874 14866 23886
rect 15486 23938 15538 23950
rect 15486 23874 15538 23886
rect 22094 23938 22146 23950
rect 22094 23874 22146 23886
rect 27582 23938 27634 23950
rect 27582 23874 27634 23886
rect 27806 23938 27858 23950
rect 27806 23874 27858 23886
rect 27918 23938 27970 23950
rect 27918 23874 27970 23886
rect 32174 23938 32226 23950
rect 44270 23938 44322 23950
rect 33058 23886 33070 23938
rect 33122 23886 33134 23938
rect 41458 23886 41470 23938
rect 41522 23886 41534 23938
rect 44818 23886 44830 23938
rect 44882 23886 44894 23938
rect 32174 23874 32226 23886
rect 44270 23874 44322 23886
rect 2718 23826 2770 23838
rect 5070 23826 5122 23838
rect 3154 23774 3166 23826
rect 3218 23774 3230 23826
rect 2718 23762 2770 23774
rect 5070 23762 5122 23774
rect 5854 23826 5906 23838
rect 5854 23762 5906 23774
rect 6638 23826 6690 23838
rect 6638 23762 6690 23774
rect 8094 23826 8146 23838
rect 8094 23762 8146 23774
rect 9214 23826 9266 23838
rect 16046 23826 16098 23838
rect 11666 23774 11678 23826
rect 11730 23774 11742 23826
rect 9214 23762 9266 23774
rect 16046 23762 16098 23774
rect 16382 23826 16434 23838
rect 16382 23762 16434 23774
rect 22318 23826 22370 23838
rect 22318 23762 22370 23774
rect 24334 23826 24386 23838
rect 24334 23762 24386 23774
rect 27358 23826 27410 23838
rect 27358 23762 27410 23774
rect 37102 23826 37154 23838
rect 45602 23774 45614 23826
rect 45666 23774 45678 23826
rect 37102 23762 37154 23774
rect 5518 23714 5570 23726
rect 5518 23650 5570 23662
rect 5742 23714 5794 23726
rect 5742 23650 5794 23662
rect 6862 23714 6914 23726
rect 6862 23650 6914 23662
rect 7310 23714 7362 23726
rect 7310 23650 7362 23662
rect 8430 23714 8482 23726
rect 8430 23650 8482 23662
rect 12910 23714 12962 23726
rect 12910 23650 12962 23662
rect 22766 23714 22818 23726
rect 22766 23650 22818 23662
rect 24894 23714 24946 23726
rect 24894 23650 24946 23662
rect 31614 23714 31666 23726
rect 31614 23650 31666 23662
rect 32846 23714 32898 23726
rect 32846 23650 32898 23662
rect 38222 23714 38274 23726
rect 38222 23650 38274 23662
rect 1344 23546 48608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48608 23546
rect 1344 23460 48608 23494
rect 5070 23378 5122 23390
rect 5070 23314 5122 23326
rect 5518 23378 5570 23390
rect 5518 23314 5570 23326
rect 6078 23378 6130 23390
rect 6078 23314 6130 23326
rect 6302 23378 6354 23390
rect 6302 23314 6354 23326
rect 6414 23378 6466 23390
rect 6414 23314 6466 23326
rect 8542 23378 8594 23390
rect 8542 23314 8594 23326
rect 10110 23378 10162 23390
rect 15486 23378 15538 23390
rect 25342 23378 25394 23390
rect 15026 23326 15038 23378
rect 15090 23326 15102 23378
rect 18274 23326 18286 23378
rect 18338 23326 18350 23378
rect 10110 23314 10162 23326
rect 15486 23314 15538 23326
rect 25342 23314 25394 23326
rect 25790 23378 25842 23390
rect 25790 23314 25842 23326
rect 33182 23378 33234 23390
rect 33182 23314 33234 23326
rect 40350 23378 40402 23390
rect 40350 23314 40402 23326
rect 45166 23378 45218 23390
rect 45166 23314 45218 23326
rect 6638 23266 6690 23278
rect 6638 23202 6690 23214
rect 6750 23266 6802 23278
rect 6750 23202 6802 23214
rect 7310 23266 7362 23278
rect 7310 23202 7362 23214
rect 8766 23266 8818 23278
rect 8766 23202 8818 23214
rect 19630 23266 19682 23278
rect 22194 23214 22206 23266
rect 22258 23214 22270 23266
rect 22978 23214 22990 23266
rect 23042 23214 23054 23266
rect 27794 23214 27806 23266
rect 27858 23214 27870 23266
rect 31266 23214 31278 23266
rect 31330 23214 31342 23266
rect 43026 23214 43038 23266
rect 43090 23214 43102 23266
rect 19630 23202 19682 23214
rect 5406 23154 5458 23166
rect 1810 23102 1822 23154
rect 1874 23102 1886 23154
rect 5406 23090 5458 23102
rect 5966 23154 6018 23166
rect 5966 23090 6018 23102
rect 7422 23154 7474 23166
rect 7422 23090 7474 23102
rect 7534 23154 7586 23166
rect 7534 23090 7586 23102
rect 7982 23154 8034 23166
rect 7982 23090 8034 23102
rect 8878 23154 8930 23166
rect 10446 23154 10498 23166
rect 10894 23154 10946 23166
rect 17950 23154 18002 23166
rect 25118 23154 25170 23166
rect 10322 23102 10334 23154
rect 10386 23102 10398 23154
rect 10658 23102 10670 23154
rect 10722 23102 10734 23154
rect 11218 23102 11230 23154
rect 11282 23102 11294 23154
rect 12114 23102 12126 23154
rect 12178 23102 12190 23154
rect 12562 23102 12574 23154
rect 12626 23102 12638 23154
rect 22754 23102 22766 23154
rect 22818 23102 22830 23154
rect 24658 23102 24670 23154
rect 24722 23102 24734 23154
rect 8878 23090 8930 23102
rect 10446 23090 10498 23102
rect 10894 23090 10946 23102
rect 17950 23090 18002 23102
rect 25118 23090 25170 23102
rect 25454 23154 25506 23166
rect 30382 23154 30434 23166
rect 27010 23102 27022 23154
rect 27074 23102 27086 23154
rect 25454 23090 25506 23102
rect 30382 23090 30434 23102
rect 30606 23154 30658 23166
rect 30606 23090 30658 23102
rect 34302 23154 34354 23166
rect 34738 23102 34750 23154
rect 34802 23102 34814 23154
rect 43698 23102 43710 23154
rect 43762 23102 43774 23154
rect 44930 23102 44942 23154
rect 44994 23102 45006 23154
rect 34302 23090 34354 23102
rect 4958 23042 5010 23054
rect 2482 22990 2494 23042
rect 2546 22990 2558 23042
rect 4610 22990 4622 23042
rect 4674 22990 4686 23042
rect 4958 22978 5010 22990
rect 8318 23042 8370 23054
rect 8318 22978 8370 22990
rect 9774 23042 9826 23054
rect 14478 23042 14530 23054
rect 13122 22990 13134 23042
rect 13186 22990 13198 23042
rect 9774 22978 9826 22990
rect 14478 22978 14530 22990
rect 17726 23042 17778 23054
rect 17726 22978 17778 22990
rect 19182 23042 19234 23054
rect 19182 22978 19234 22990
rect 20974 23042 21026 23054
rect 20974 22978 21026 22990
rect 25902 23042 25954 23054
rect 25902 22978 25954 22990
rect 26686 23042 26738 23054
rect 29922 22990 29934 23042
rect 29986 22990 29998 23042
rect 32162 22990 32174 23042
rect 32226 22990 32238 23042
rect 35410 22990 35422 23042
rect 35474 22990 35486 23042
rect 37538 22990 37550 23042
rect 37602 22990 37614 23042
rect 40898 22990 40910 23042
rect 40962 22990 40974 23042
rect 26686 22978 26738 22990
rect 5518 22930 5570 22942
rect 5518 22866 5570 22878
rect 14702 22930 14754 22942
rect 14702 22866 14754 22878
rect 18622 22930 18674 22942
rect 18622 22866 18674 22878
rect 18958 22930 19010 22942
rect 18958 22866 19010 22878
rect 24558 22930 24610 22942
rect 30930 22878 30942 22930
rect 30994 22878 31006 22930
rect 24558 22866 24610 22878
rect 1344 22762 48608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48608 22762
rect 1344 22676 48608 22710
rect 4510 22594 4562 22606
rect 16930 22542 16942 22594
rect 16994 22542 17006 22594
rect 22194 22542 22206 22594
rect 22258 22542 22270 22594
rect 4510 22530 4562 22542
rect 5742 22482 5794 22494
rect 5742 22418 5794 22430
rect 9774 22482 9826 22494
rect 9774 22418 9826 22430
rect 10222 22482 10274 22494
rect 21422 22482 21474 22494
rect 26798 22482 26850 22494
rect 17490 22430 17502 22482
rect 17554 22430 17566 22482
rect 21970 22430 21982 22482
rect 22034 22430 22046 22482
rect 25330 22430 25342 22482
rect 25394 22430 25406 22482
rect 10222 22418 10274 22430
rect 21422 22418 21474 22430
rect 26798 22418 26850 22430
rect 28254 22482 28306 22494
rect 40350 22482 40402 22494
rect 32498 22430 32510 22482
rect 32562 22430 32574 22482
rect 34626 22430 34638 22482
rect 34690 22430 34702 22482
rect 37762 22430 37774 22482
rect 37826 22430 37838 22482
rect 39890 22430 39902 22482
rect 39954 22430 39966 22482
rect 28254 22418 28306 22430
rect 40350 22418 40402 22430
rect 7870 22370 7922 22382
rect 2146 22318 2158 22370
rect 2210 22318 2222 22370
rect 7870 22306 7922 22318
rect 8206 22370 8258 22382
rect 28030 22370 28082 22382
rect 10882 22318 10894 22370
rect 10946 22318 10958 22370
rect 11666 22318 11678 22370
rect 11730 22318 11742 22370
rect 11890 22318 11902 22370
rect 11954 22318 11966 22370
rect 17602 22318 17614 22370
rect 17666 22318 17678 22370
rect 18946 22318 18958 22370
rect 19010 22318 19022 22370
rect 19954 22318 19966 22370
rect 20018 22318 20030 22370
rect 20514 22318 20526 22370
rect 20578 22318 20590 22370
rect 23090 22318 23102 22370
rect 23154 22318 23166 22370
rect 23874 22318 23886 22370
rect 23938 22318 23950 22370
rect 26114 22318 26126 22370
rect 26178 22318 26190 22370
rect 8206 22306 8258 22318
rect 28030 22306 28082 22318
rect 31054 22370 31106 22382
rect 35086 22370 35138 22382
rect 31714 22318 31726 22370
rect 31778 22318 31790 22370
rect 35970 22318 35982 22370
rect 36034 22318 36046 22370
rect 37090 22318 37102 22370
rect 37154 22318 37166 22370
rect 31054 22306 31106 22318
rect 35086 22306 35138 22318
rect 27246 22258 27298 22270
rect 27246 22194 27298 22206
rect 35758 22258 35810 22270
rect 35758 22194 35810 22206
rect 7982 22146 8034 22158
rect 29262 22146 29314 22158
rect 11106 22094 11118 22146
rect 11170 22094 11182 22146
rect 27682 22094 27694 22146
rect 27746 22094 27758 22146
rect 7982 22082 8034 22094
rect 29262 22082 29314 22094
rect 31390 22146 31442 22158
rect 31390 22082 31442 22094
rect 40238 22146 40290 22158
rect 40238 22082 40290 22094
rect 1344 21978 48608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48608 21978
rect 1344 21892 48608 21926
rect 2046 21810 2098 21822
rect 2046 21746 2098 21758
rect 2270 21810 2322 21822
rect 2270 21746 2322 21758
rect 9550 21810 9602 21822
rect 9550 21746 9602 21758
rect 11230 21810 11282 21822
rect 11230 21746 11282 21758
rect 12798 21810 12850 21822
rect 12798 21746 12850 21758
rect 24222 21810 24274 21822
rect 24222 21746 24274 21758
rect 24670 21810 24722 21822
rect 24670 21746 24722 21758
rect 30382 21810 30434 21822
rect 30382 21746 30434 21758
rect 31950 21810 32002 21822
rect 39230 21810 39282 21822
rect 38098 21758 38110 21810
rect 38162 21758 38174 21810
rect 31950 21746 32002 21758
rect 39230 21746 39282 21758
rect 1710 21698 1762 21710
rect 1710 21634 1762 21646
rect 2494 21698 2546 21710
rect 2494 21634 2546 21646
rect 2606 21698 2658 21710
rect 2606 21634 2658 21646
rect 11566 21698 11618 21710
rect 11566 21634 11618 21646
rect 17390 21698 17442 21710
rect 17390 21634 17442 21646
rect 17726 21698 17778 21710
rect 42254 21698 42306 21710
rect 35074 21646 35086 21698
rect 35138 21646 35150 21698
rect 17726 21634 17778 21646
rect 42254 21634 42306 21646
rect 3054 21586 3106 21598
rect 30830 21586 30882 21598
rect 9762 21534 9774 21586
rect 9826 21534 9838 21586
rect 12114 21534 12126 21586
rect 12178 21534 12190 21586
rect 19506 21534 19518 21586
rect 19570 21534 19582 21586
rect 20850 21534 20862 21586
rect 20914 21534 20926 21586
rect 22418 21534 22430 21586
rect 22482 21534 22494 21586
rect 25218 21534 25230 21586
rect 25282 21534 25294 21586
rect 30482 21534 30494 21586
rect 30546 21534 30558 21586
rect 3054 21522 3106 21534
rect 30830 21522 30882 21534
rect 31502 21586 31554 21598
rect 36878 21586 36930 21598
rect 41918 21586 41970 21598
rect 34178 21534 34190 21586
rect 34242 21534 34254 21586
rect 36530 21534 36542 21586
rect 36594 21534 36606 21586
rect 38322 21534 38334 21586
rect 38386 21534 38398 21586
rect 31502 21522 31554 21534
rect 36878 21522 36930 21534
rect 41918 21522 41970 21534
rect 42478 21586 42530 21598
rect 42478 21522 42530 21534
rect 14254 21474 14306 21486
rect 23438 21474 23490 21486
rect 11890 21422 11902 21474
rect 11954 21422 11966 21474
rect 18610 21422 18622 21474
rect 18674 21422 18686 21474
rect 21634 21422 21646 21474
rect 21698 21422 21710 21474
rect 14254 21410 14306 21422
rect 23438 21410 23490 21422
rect 23886 21474 23938 21486
rect 38782 21474 38834 21486
rect 26002 21422 26014 21474
rect 26066 21422 26078 21474
rect 28130 21422 28142 21474
rect 28194 21422 28206 21474
rect 23886 21410 23938 21422
rect 38782 21410 38834 21422
rect 42814 21362 42866 21374
rect 18498 21310 18510 21362
rect 18562 21310 18574 21362
rect 42814 21298 42866 21310
rect 1344 21194 48608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48608 21194
rect 1344 21108 48608 21142
rect 8206 21026 8258 21038
rect 8206 20962 8258 20974
rect 8766 21026 8818 21038
rect 8766 20962 8818 20974
rect 13694 21026 13746 21038
rect 30706 20974 30718 21026
rect 30770 20974 30782 21026
rect 35858 20974 35870 21026
rect 35922 20974 35934 21026
rect 39218 20974 39230 21026
rect 39282 20974 39294 21026
rect 13694 20962 13746 20974
rect 1822 20914 1874 20926
rect 1822 20850 1874 20862
rect 3838 20914 3890 20926
rect 3838 20850 3890 20862
rect 9326 20914 9378 20926
rect 23102 20914 23154 20926
rect 16370 20862 16382 20914
rect 16434 20862 16446 20914
rect 18498 20862 18510 20914
rect 18562 20862 18574 20914
rect 9326 20850 9378 20862
rect 23102 20850 23154 20862
rect 23886 20914 23938 20926
rect 37214 20914 37266 20926
rect 24882 20862 24894 20914
rect 24946 20862 24958 20914
rect 27010 20862 27022 20914
rect 27074 20862 27086 20914
rect 30482 20862 30494 20914
rect 30546 20862 30558 20914
rect 32274 20862 32286 20914
rect 32338 20862 32350 20914
rect 34402 20862 34414 20914
rect 34466 20862 34478 20914
rect 23886 20850 23938 20862
rect 37214 20850 37266 20862
rect 38222 20914 38274 20926
rect 40226 20862 40238 20914
rect 40290 20862 40302 20914
rect 38222 20850 38274 20862
rect 13470 20802 13522 20814
rect 15262 20802 15314 20814
rect 22878 20802 22930 20814
rect 29374 20802 29426 20814
rect 36206 20802 36258 20814
rect 14018 20750 14030 20802
rect 14082 20750 14094 20802
rect 14578 20750 14590 20802
rect 14642 20750 14654 20802
rect 15586 20750 15598 20802
rect 15650 20750 15662 20802
rect 24098 20750 24110 20802
rect 24162 20750 24174 20802
rect 27906 20750 27918 20802
rect 27970 20750 27982 20802
rect 31602 20750 31614 20802
rect 31666 20750 31678 20802
rect 13470 20738 13522 20750
rect 15262 20738 15314 20750
rect 22878 20738 22930 20750
rect 29374 20738 29426 20750
rect 36206 20738 36258 20750
rect 36430 20802 36482 20814
rect 36430 20738 36482 20750
rect 38894 20802 38946 20814
rect 42814 20802 42866 20814
rect 39442 20750 39454 20802
rect 39506 20750 39518 20802
rect 40114 20750 40126 20802
rect 40178 20750 40190 20802
rect 38894 20738 38946 20750
rect 42814 20738 42866 20750
rect 8094 20690 8146 20702
rect 8094 20626 8146 20638
rect 8878 20690 8930 20702
rect 29486 20690 29538 20702
rect 22194 20638 22206 20690
rect 22258 20638 22270 20690
rect 22530 20638 22542 20690
rect 22594 20638 22606 20690
rect 30818 20638 30830 20690
rect 30882 20638 30894 20690
rect 8878 20626 8930 20638
rect 29486 20626 29538 20638
rect 4286 20578 4338 20590
rect 4286 20514 4338 20526
rect 8206 20578 8258 20590
rect 8206 20514 8258 20526
rect 14366 20578 14418 20590
rect 14366 20514 14418 20526
rect 27694 20578 27746 20590
rect 27694 20514 27746 20526
rect 37550 20578 37602 20590
rect 37550 20514 37602 20526
rect 42478 20578 42530 20590
rect 42478 20514 42530 20526
rect 1344 20410 48608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48608 20410
rect 1344 20324 48608 20358
rect 2158 20242 2210 20254
rect 2158 20178 2210 20190
rect 22878 20242 22930 20254
rect 22878 20178 22930 20190
rect 30270 20242 30322 20254
rect 30270 20178 30322 20190
rect 31166 20242 31218 20254
rect 31166 20178 31218 20190
rect 32174 20242 32226 20254
rect 32174 20178 32226 20190
rect 39454 20242 39506 20254
rect 39454 20178 39506 20190
rect 2382 20130 2434 20142
rect 2382 20066 2434 20078
rect 3054 20130 3106 20142
rect 23550 20130 23602 20142
rect 35534 20130 35586 20142
rect 3266 20078 3278 20130
rect 3330 20078 3342 20130
rect 5730 20078 5742 20130
rect 5794 20078 5806 20130
rect 13682 20078 13694 20130
rect 13746 20078 13758 20130
rect 27682 20078 27694 20130
rect 27746 20078 27758 20130
rect 42466 20078 42478 20130
rect 42530 20078 42542 20130
rect 3054 20066 3106 20078
rect 23550 20066 23602 20078
rect 35534 20066 35586 20078
rect 3390 20018 3442 20030
rect 16382 20018 16434 20030
rect 2818 19966 2830 20018
rect 2882 19966 2894 20018
rect 8978 19966 8990 20018
rect 9042 19966 9054 20018
rect 12562 19966 12574 20018
rect 12626 19966 12638 20018
rect 13010 19966 13022 20018
rect 13074 19966 13086 20018
rect 3390 19954 3442 19966
rect 16382 19954 16434 19966
rect 19070 20018 19122 20030
rect 23214 20018 23266 20030
rect 19282 19966 19294 20018
rect 19346 19966 19358 20018
rect 19070 19954 19122 19966
rect 23214 19954 23266 19966
rect 23998 20018 24050 20030
rect 34862 20018 34914 20030
rect 26898 19966 26910 20018
rect 26962 19966 26974 20018
rect 23998 19954 24050 19966
rect 34862 19954 34914 19966
rect 35086 20018 35138 20030
rect 35086 19954 35138 19966
rect 38894 20018 38946 20030
rect 38894 19954 38946 19966
rect 39230 20018 39282 20030
rect 41794 19966 41806 20018
rect 41858 19966 41870 20018
rect 39230 19954 39282 19966
rect 26574 19906 26626 19918
rect 30158 19906 30210 19918
rect 9650 19854 9662 19906
rect 9714 19854 9726 19906
rect 11778 19854 11790 19906
rect 11842 19854 11854 19906
rect 15810 19854 15822 19906
rect 15874 19854 15886 19906
rect 20066 19854 20078 19906
rect 20130 19854 20142 19906
rect 22194 19854 22206 19906
rect 22258 19854 22270 19906
rect 29810 19854 29822 19906
rect 29874 19854 29886 19906
rect 26574 19842 26626 19854
rect 30158 19842 30210 19854
rect 31614 19906 31666 19918
rect 31614 19842 31666 19854
rect 38446 19906 38498 19918
rect 41358 19906 41410 19918
rect 39442 19854 39454 19906
rect 39506 19854 39518 19906
rect 44594 19854 44606 19906
rect 44658 19854 44670 19906
rect 38446 19842 38498 19854
rect 41358 19842 41410 19854
rect 34514 19742 34526 19794
rect 34578 19742 34590 19794
rect 1344 19626 48608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48608 19626
rect 1344 19540 48608 19574
rect 6078 19458 6130 19470
rect 22878 19458 22930 19470
rect 7970 19406 7982 19458
rect 8034 19406 8046 19458
rect 6078 19394 6130 19406
rect 22878 19394 22930 19406
rect 27022 19458 27074 19470
rect 27022 19394 27074 19406
rect 45054 19458 45106 19470
rect 45054 19394 45106 19406
rect 4846 19346 4898 19358
rect 4846 19282 4898 19294
rect 8878 19346 8930 19358
rect 8878 19282 8930 19294
rect 12798 19346 12850 19358
rect 12798 19282 12850 19294
rect 24334 19346 24386 19358
rect 24334 19282 24386 19294
rect 25454 19346 25506 19358
rect 43822 19346 43874 19358
rect 39442 19294 39454 19346
rect 39506 19294 39518 19346
rect 41570 19294 41582 19346
rect 41634 19294 41646 19346
rect 25454 19282 25506 19294
rect 43822 19282 43874 19294
rect 44382 19346 44434 19358
rect 44382 19282 44434 19294
rect 44830 19346 44882 19358
rect 44830 19282 44882 19294
rect 3950 19234 4002 19246
rect 3950 19170 4002 19182
rect 7422 19234 7474 19246
rect 7422 19170 7474 19182
rect 7646 19234 7698 19246
rect 23214 19234 23266 19246
rect 8418 19182 8430 19234
rect 8482 19182 8494 19234
rect 11330 19182 11342 19234
rect 11394 19182 11406 19234
rect 7646 19170 7698 19182
rect 23214 19170 23266 19182
rect 23886 19234 23938 19246
rect 24770 19182 24782 19234
rect 24834 19182 24846 19234
rect 34962 19182 34974 19234
rect 35026 19182 35038 19234
rect 38658 19182 38670 19234
rect 38722 19182 38734 19234
rect 23886 19170 23938 19182
rect 2270 19122 2322 19134
rect 2270 19058 2322 19070
rect 2382 19122 2434 19134
rect 2382 19058 2434 19070
rect 2830 19122 2882 19134
rect 2830 19058 2882 19070
rect 3166 19122 3218 19134
rect 3166 19058 3218 19070
rect 3390 19122 3442 19134
rect 3390 19058 3442 19070
rect 3502 19122 3554 19134
rect 3502 19058 3554 19070
rect 4062 19122 4114 19134
rect 4062 19058 4114 19070
rect 5966 19122 6018 19134
rect 5966 19058 6018 19070
rect 6526 19122 6578 19134
rect 6526 19058 6578 19070
rect 11566 19122 11618 19134
rect 11566 19058 11618 19070
rect 19966 19122 20018 19134
rect 19966 19058 20018 19070
rect 20302 19122 20354 19134
rect 20302 19058 20354 19070
rect 23438 19122 23490 19134
rect 23438 19058 23490 19070
rect 27134 19122 27186 19134
rect 27134 19058 27186 19070
rect 2046 19010 2098 19022
rect 2046 18946 2098 18958
rect 2606 19010 2658 19022
rect 2606 18946 2658 18958
rect 2942 19010 2994 19022
rect 2942 18946 2994 18958
rect 3726 19010 3778 19022
rect 3726 18946 3778 18958
rect 6078 19010 6130 19022
rect 6078 18946 6130 18958
rect 6638 19010 6690 19022
rect 6638 18946 6690 18958
rect 6862 19010 6914 19022
rect 6862 18946 6914 18958
rect 8766 19010 8818 19022
rect 8766 18946 8818 18958
rect 8990 19010 9042 19022
rect 8990 18946 9042 18958
rect 25006 19010 25058 19022
rect 25006 18946 25058 18958
rect 34750 19010 34802 19022
rect 34750 18946 34802 18958
rect 38334 19010 38386 19022
rect 45378 18958 45390 19010
rect 45442 18958 45454 19010
rect 38334 18946 38386 18958
rect 1344 18842 48608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48608 18842
rect 1344 18756 48608 18790
rect 6414 18674 6466 18686
rect 6414 18610 6466 18622
rect 7422 18674 7474 18686
rect 7422 18610 7474 18622
rect 8654 18674 8706 18686
rect 23214 18674 23266 18686
rect 11330 18622 11342 18674
rect 11394 18622 11406 18674
rect 17714 18622 17726 18674
rect 17778 18622 17790 18674
rect 23874 18622 23886 18674
rect 23938 18622 23950 18674
rect 8654 18610 8706 18622
rect 23214 18610 23266 18622
rect 5406 18562 5458 18574
rect 2482 18510 2494 18562
rect 2546 18510 2558 18562
rect 5406 18498 5458 18510
rect 7758 18562 7810 18574
rect 7758 18498 7810 18510
rect 8542 18562 8594 18574
rect 8542 18498 8594 18510
rect 9662 18562 9714 18574
rect 9662 18498 9714 18510
rect 15934 18562 15986 18574
rect 41022 18562 41074 18574
rect 24434 18510 24446 18562
rect 24498 18510 24510 18562
rect 15934 18498 15986 18510
rect 41022 18498 41074 18510
rect 44158 18562 44210 18574
rect 44158 18498 44210 18510
rect 5630 18450 5682 18462
rect 1810 18398 1822 18450
rect 1874 18398 1886 18450
rect 5630 18386 5682 18398
rect 5742 18450 5794 18462
rect 5742 18386 5794 18398
rect 5854 18450 5906 18462
rect 5854 18386 5906 18398
rect 6302 18450 6354 18462
rect 6302 18386 6354 18398
rect 6526 18450 6578 18462
rect 6526 18386 6578 18398
rect 6974 18450 7026 18462
rect 8206 18450 8258 18462
rect 7186 18398 7198 18450
rect 7250 18398 7262 18450
rect 7522 18398 7534 18450
rect 7586 18398 7598 18450
rect 6974 18386 7026 18398
rect 8206 18386 8258 18398
rect 9438 18450 9490 18462
rect 9438 18386 9490 18398
rect 9774 18450 9826 18462
rect 9774 18386 9826 18398
rect 11006 18450 11058 18462
rect 11006 18386 11058 18398
rect 11790 18450 11842 18462
rect 18062 18450 18114 18462
rect 16146 18398 16158 18450
rect 16210 18398 16222 18450
rect 11790 18386 11842 18398
rect 18062 18386 18114 18398
rect 18734 18450 18786 18462
rect 18734 18386 18786 18398
rect 19966 18450 20018 18462
rect 40350 18450 40402 18462
rect 23538 18398 23550 18450
rect 23602 18398 23614 18450
rect 24098 18398 24110 18450
rect 24162 18398 24174 18450
rect 25218 18398 25230 18450
rect 25282 18398 25294 18450
rect 26002 18398 26014 18450
rect 26066 18398 26078 18450
rect 32386 18398 32398 18450
rect 32450 18398 32462 18450
rect 39778 18398 39790 18450
rect 39842 18398 39854 18450
rect 19966 18386 20018 18398
rect 40350 18386 40402 18398
rect 44494 18450 44546 18462
rect 44494 18386 44546 18398
rect 10782 18338 10834 18350
rect 4610 18286 4622 18338
rect 4674 18286 4686 18338
rect 10782 18274 10834 18286
rect 18286 18338 18338 18350
rect 18286 18274 18338 18286
rect 20414 18338 20466 18350
rect 33182 18338 33234 18350
rect 28130 18286 28142 18338
rect 28194 18286 28206 18338
rect 29586 18286 29598 18338
rect 29650 18286 29662 18338
rect 31714 18286 31726 18338
rect 31778 18286 31790 18338
rect 20414 18274 20466 18286
rect 33182 18274 33234 18286
rect 36654 18338 36706 18350
rect 36978 18286 36990 18338
rect 37042 18286 37054 18338
rect 39106 18286 39118 18338
rect 39170 18286 39182 18338
rect 36654 18274 36706 18286
rect 8094 18226 8146 18238
rect 8094 18162 8146 18174
rect 8654 18226 8706 18238
rect 8654 18162 8706 18174
rect 40910 18226 40962 18238
rect 40910 18162 40962 18174
rect 1344 18058 48608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48608 18058
rect 1344 17972 48608 18006
rect 7422 17890 7474 17902
rect 9326 17890 9378 17902
rect 24782 17890 24834 17902
rect 8866 17838 8878 17890
rect 8930 17838 8942 17890
rect 20066 17838 20078 17890
rect 20130 17838 20142 17890
rect 7422 17826 7474 17838
rect 9326 17826 9378 17838
rect 24782 17826 24834 17838
rect 25118 17890 25170 17902
rect 25118 17826 25170 17838
rect 26238 17890 26290 17902
rect 26238 17826 26290 17838
rect 37886 17890 37938 17902
rect 37886 17826 37938 17838
rect 45278 17890 45330 17902
rect 45278 17826 45330 17838
rect 4622 17778 4674 17790
rect 4622 17714 4674 17726
rect 5742 17778 5794 17790
rect 26462 17778 26514 17790
rect 15810 17726 15822 17778
rect 15874 17726 15886 17778
rect 17938 17726 17950 17778
rect 18002 17726 18014 17778
rect 24210 17726 24222 17778
rect 24274 17726 24286 17778
rect 5742 17714 5794 17726
rect 26462 17714 26514 17726
rect 33182 17778 33234 17790
rect 37326 17778 37378 17790
rect 34290 17726 34302 17778
rect 34354 17726 34366 17778
rect 36418 17726 36430 17778
rect 36482 17726 36494 17778
rect 33182 17714 33234 17726
rect 37326 17714 37378 17726
rect 1710 17666 1762 17678
rect 1710 17602 1762 17614
rect 2270 17666 2322 17678
rect 5182 17666 5234 17678
rect 3938 17614 3950 17666
rect 4002 17614 4014 17666
rect 2270 17602 2322 17614
rect 5182 17602 5234 17614
rect 6078 17666 6130 17678
rect 6078 17602 6130 17614
rect 7534 17666 7586 17678
rect 7534 17602 7586 17614
rect 7870 17666 7922 17678
rect 7870 17602 7922 17614
rect 8318 17666 8370 17678
rect 8318 17602 8370 17614
rect 8542 17666 8594 17678
rect 20414 17666 20466 17678
rect 15138 17614 15150 17666
rect 15202 17614 15214 17666
rect 18834 17614 18846 17666
rect 18898 17614 18910 17666
rect 19170 17614 19182 17666
rect 19234 17614 19246 17666
rect 8542 17602 8594 17614
rect 20414 17602 20466 17614
rect 20638 17666 20690 17678
rect 37662 17666 37714 17678
rect 21298 17614 21310 17666
rect 21362 17614 21374 17666
rect 33506 17614 33518 17666
rect 33570 17614 33582 17666
rect 20638 17602 20690 17614
rect 37662 17602 37714 17614
rect 39342 17666 39394 17678
rect 41022 17666 41074 17678
rect 39890 17614 39902 17666
rect 39954 17614 39966 17666
rect 40562 17614 40574 17666
rect 40626 17614 40638 17666
rect 39342 17602 39394 17614
rect 41022 17602 41074 17614
rect 2046 17554 2098 17566
rect 2046 17490 2098 17502
rect 2606 17554 2658 17566
rect 2606 17490 2658 17502
rect 2830 17554 2882 17566
rect 4846 17554 4898 17566
rect 7310 17554 7362 17566
rect 3490 17502 3502 17554
rect 3554 17502 3566 17554
rect 3714 17502 3726 17554
rect 3778 17502 3790 17554
rect 6290 17502 6302 17554
rect 6354 17502 6366 17554
rect 6626 17502 6638 17554
rect 6690 17502 6702 17554
rect 2830 17490 2882 17502
rect 4846 17490 4898 17502
rect 7310 17490 7362 17502
rect 9214 17554 9266 17566
rect 24558 17554 24610 17566
rect 31054 17554 31106 17566
rect 18722 17502 18734 17554
rect 18786 17502 18798 17554
rect 22082 17502 22094 17554
rect 22146 17502 22158 17554
rect 29138 17502 29150 17554
rect 29202 17502 29214 17554
rect 29922 17502 29934 17554
rect 29986 17502 29998 17554
rect 9214 17490 9266 17502
rect 24558 17490 24610 17502
rect 31054 17490 31106 17502
rect 31390 17554 31442 17566
rect 38558 17554 38610 17566
rect 38210 17502 38222 17554
rect 38274 17502 38286 17554
rect 31390 17490 31442 17502
rect 38558 17490 38610 17502
rect 38894 17554 38946 17566
rect 45390 17554 45442 17566
rect 39666 17502 39678 17554
rect 39730 17502 39742 17554
rect 38894 17490 38946 17502
rect 45390 17490 45442 17502
rect 2494 17442 2546 17454
rect 2494 17378 2546 17390
rect 4958 17442 5010 17454
rect 4958 17378 5010 17390
rect 7758 17442 7810 17454
rect 7758 17378 7810 17390
rect 9326 17442 9378 17454
rect 9326 17378 9378 17390
rect 14702 17442 14754 17454
rect 19518 17442 19570 17454
rect 19394 17390 19406 17442
rect 19458 17390 19470 17442
rect 14702 17378 14754 17390
rect 19518 17378 19570 17390
rect 25566 17442 25618 17454
rect 26910 17442 26962 17454
rect 25890 17390 25902 17442
rect 25954 17390 25966 17442
rect 25566 17378 25618 17390
rect 26910 17378 26962 17390
rect 27358 17442 27410 17454
rect 27358 17378 27410 17390
rect 28590 17442 28642 17454
rect 28590 17378 28642 17390
rect 41470 17442 41522 17454
rect 41470 17378 41522 17390
rect 1344 17274 48608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48608 17274
rect 1344 17188 48608 17222
rect 1822 17106 1874 17118
rect 1822 17042 1874 17054
rect 5406 17106 5458 17118
rect 7758 17106 7810 17118
rect 7186 17054 7198 17106
rect 7250 17054 7262 17106
rect 5406 17042 5458 17054
rect 7758 17042 7810 17054
rect 7982 17106 8034 17118
rect 7982 17042 8034 17054
rect 15262 17106 15314 17118
rect 19294 17106 19346 17118
rect 15922 17054 15934 17106
rect 15986 17054 15998 17106
rect 19170 17054 19182 17106
rect 19234 17054 19246 17106
rect 15262 17042 15314 17054
rect 19294 17042 19346 17054
rect 20190 17106 20242 17118
rect 20190 17042 20242 17054
rect 21646 17106 21698 17118
rect 21646 17042 21698 17054
rect 30270 17106 30322 17118
rect 30270 17042 30322 17054
rect 30494 17106 30546 17118
rect 32062 17106 32114 17118
rect 31042 17054 31054 17106
rect 31106 17054 31118 17106
rect 30494 17042 30546 17054
rect 32062 17042 32114 17054
rect 33294 17106 33346 17118
rect 33294 17042 33346 17054
rect 34078 17106 34130 17118
rect 34078 17042 34130 17054
rect 35198 17106 35250 17118
rect 35198 17042 35250 17054
rect 35646 17106 35698 17118
rect 35646 17042 35698 17054
rect 38782 17106 38834 17118
rect 38782 17042 38834 17054
rect 41918 17106 41970 17118
rect 41918 17042 41970 17054
rect 5294 16994 5346 17006
rect 5294 16930 5346 16942
rect 5854 16994 5906 17006
rect 5854 16930 5906 16942
rect 6078 16994 6130 17006
rect 6078 16930 6130 16942
rect 14478 16994 14530 17006
rect 14478 16930 14530 16942
rect 14814 16994 14866 17006
rect 20974 16994 21026 17006
rect 18386 16942 18398 16994
rect 18450 16942 18462 16994
rect 14814 16930 14866 16942
rect 20974 16930 21026 16942
rect 28814 16994 28866 17006
rect 28814 16930 28866 16942
rect 29710 16994 29762 17006
rect 29710 16930 29762 16942
rect 33518 16994 33570 17006
rect 33518 16930 33570 16942
rect 33630 16994 33682 17006
rect 36194 16942 36206 16994
rect 36258 16942 36270 16994
rect 44146 16942 44158 16994
rect 44210 16942 44222 16994
rect 33630 16930 33682 16942
rect 5742 16882 5794 16894
rect 5742 16818 5794 16830
rect 6302 16882 6354 16894
rect 6302 16818 6354 16830
rect 6638 16882 6690 16894
rect 6638 16818 6690 16830
rect 6862 16882 6914 16894
rect 17838 16882 17890 16894
rect 24670 16882 24722 16894
rect 30606 16882 30658 16894
rect 38894 16882 38946 16894
rect 41806 16882 41858 16894
rect 7522 16830 7534 16882
rect 7586 16830 7598 16882
rect 11890 16830 11902 16882
rect 11954 16830 11966 16882
rect 14130 16830 14142 16882
rect 14194 16830 14206 16882
rect 18610 16830 18622 16882
rect 18674 16830 18686 16882
rect 18946 16830 18958 16882
rect 19010 16830 19022 16882
rect 21410 16830 21422 16882
rect 21474 16830 21486 16882
rect 28018 16830 28030 16882
rect 28082 16830 28094 16882
rect 36530 16830 36542 16882
rect 36594 16830 36606 16882
rect 38546 16830 38558 16882
rect 38610 16830 38622 16882
rect 39778 16830 39790 16882
rect 39842 16830 39854 16882
rect 6862 16818 6914 16830
rect 17838 16818 17890 16830
rect 24670 16818 24722 16830
rect 30606 16818 30658 16830
rect 38894 16818 38946 16830
rect 41806 16818 41858 16830
rect 42142 16882 42194 16894
rect 43474 16830 43486 16882
rect 43538 16830 43550 16882
rect 42142 16818 42194 16830
rect 8094 16770 8146 16782
rect 16270 16770 16322 16782
rect 11442 16718 11454 16770
rect 11506 16718 11518 16770
rect 8094 16706 8146 16718
rect 16270 16706 16322 16718
rect 16494 16770 16546 16782
rect 16494 16706 16546 16718
rect 22094 16770 22146 16782
rect 31614 16770 31666 16782
rect 25218 16718 25230 16770
rect 25282 16718 25294 16770
rect 27346 16718 27358 16770
rect 27410 16718 27422 16770
rect 22094 16706 22146 16718
rect 31614 16706 31666 16718
rect 41022 16770 41074 16782
rect 41022 16706 41074 16718
rect 41470 16770 41522 16782
rect 41470 16706 41522 16718
rect 43038 16770 43090 16782
rect 46274 16718 46286 16770
rect 46338 16718 46350 16770
rect 43038 16706 43090 16718
rect 29150 16658 29202 16670
rect 11554 16606 11566 16658
rect 11618 16606 11630 16658
rect 29150 16594 29202 16606
rect 29486 16658 29538 16670
rect 29486 16594 29538 16606
rect 31390 16658 31442 16670
rect 41010 16606 41022 16658
rect 41074 16655 41086 16658
rect 41458 16655 41470 16658
rect 41074 16609 41470 16655
rect 41074 16606 41086 16609
rect 41458 16606 41470 16609
rect 41522 16606 41534 16658
rect 31390 16594 31442 16606
rect 1344 16490 48608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48608 16490
rect 1344 16404 48608 16438
rect 21870 16322 21922 16334
rect 21522 16270 21534 16322
rect 21586 16270 21598 16322
rect 21870 16258 21922 16270
rect 30830 16322 30882 16334
rect 43710 16322 43762 16334
rect 31154 16270 31166 16322
rect 31218 16319 31230 16322
rect 31378 16319 31390 16322
rect 31218 16273 31390 16319
rect 31218 16270 31230 16273
rect 31378 16270 31390 16273
rect 31442 16270 31454 16322
rect 30830 16258 30882 16270
rect 43710 16258 43762 16270
rect 5742 16210 5794 16222
rect 16830 16210 16882 16222
rect 10994 16158 11006 16210
rect 11058 16158 11070 16210
rect 14242 16158 14254 16210
rect 14306 16158 14318 16210
rect 16370 16158 16382 16210
rect 16434 16158 16446 16210
rect 5742 16146 5794 16158
rect 16830 16146 16882 16158
rect 19294 16210 19346 16222
rect 19294 16146 19346 16158
rect 22542 16210 22594 16222
rect 22542 16146 22594 16158
rect 22990 16210 23042 16222
rect 22990 16146 23042 16158
rect 29710 16210 29762 16222
rect 29710 16146 29762 16158
rect 30270 16210 30322 16222
rect 30270 16146 30322 16158
rect 31390 16210 31442 16222
rect 31390 16146 31442 16158
rect 33518 16210 33570 16222
rect 36194 16158 36206 16210
rect 36258 16158 36270 16210
rect 33518 16146 33570 16158
rect 5630 16098 5682 16110
rect 22094 16098 22146 16110
rect 11106 16046 11118 16098
rect 11170 16046 11182 16098
rect 13570 16046 13582 16098
rect 13634 16046 13646 16098
rect 17826 16046 17838 16098
rect 17890 16046 17902 16098
rect 18162 16046 18174 16098
rect 18226 16046 18238 16098
rect 19730 16046 19742 16098
rect 19794 16046 19806 16098
rect 5630 16034 5682 16046
rect 22094 16034 22146 16046
rect 29486 16098 29538 16110
rect 29486 16034 29538 16046
rect 30942 16098 30994 16110
rect 30942 16034 30994 16046
rect 33742 16098 33794 16110
rect 33742 16034 33794 16046
rect 34078 16098 34130 16110
rect 35198 16098 35250 16110
rect 39678 16098 39730 16110
rect 41470 16098 41522 16110
rect 34962 16046 34974 16098
rect 35026 16046 35038 16098
rect 35858 16046 35870 16098
rect 35922 16046 35934 16098
rect 37090 16046 37102 16098
rect 37154 16046 37166 16098
rect 39330 16046 39342 16098
rect 39394 16046 39406 16098
rect 40450 16046 40462 16098
rect 40514 16046 40526 16098
rect 34078 16034 34130 16046
rect 35198 16034 35250 16046
rect 39678 16034 39730 16046
rect 41470 16034 41522 16046
rect 5966 15986 6018 15998
rect 5966 15922 6018 15934
rect 6190 15986 6242 15998
rect 6190 15922 6242 15934
rect 11790 15986 11842 15998
rect 33966 15986 34018 15998
rect 41582 15986 41634 15998
rect 17266 15934 17278 15986
rect 17330 15934 17342 15986
rect 19954 15934 19966 15986
rect 20018 15934 20030 15986
rect 20402 15934 20414 15986
rect 20466 15934 20478 15986
rect 35970 15934 35982 15986
rect 36034 15934 36046 15986
rect 36978 15934 36990 15986
rect 37042 15934 37054 15986
rect 39218 15934 39230 15986
rect 39282 15934 39294 15986
rect 11790 15922 11842 15934
rect 33966 15922 34018 15934
rect 41582 15922 41634 15934
rect 43822 15986 43874 15998
rect 43822 15922 43874 15934
rect 30830 15874 30882 15886
rect 18386 15822 18398 15874
rect 18450 15822 18462 15874
rect 18610 15822 18622 15874
rect 18674 15822 18686 15874
rect 20626 15822 20638 15874
rect 20690 15822 20702 15874
rect 29138 15822 29150 15874
rect 29202 15822 29214 15874
rect 30830 15810 30882 15822
rect 42030 15874 42082 15886
rect 42030 15810 42082 15822
rect 1344 15706 48608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48608 15706
rect 1344 15620 48608 15654
rect 12798 15538 12850 15550
rect 12798 15474 12850 15486
rect 16606 15538 16658 15550
rect 16606 15474 16658 15486
rect 18622 15538 18674 15550
rect 18622 15474 18674 15486
rect 19070 15538 19122 15550
rect 19070 15474 19122 15486
rect 23998 15538 24050 15550
rect 23998 15474 24050 15486
rect 29934 15538 29986 15550
rect 29934 15474 29986 15486
rect 34078 15538 34130 15550
rect 34078 15474 34130 15486
rect 34526 15538 34578 15550
rect 34526 15474 34578 15486
rect 37550 15538 37602 15550
rect 37550 15474 37602 15486
rect 39790 15538 39842 15550
rect 39790 15474 39842 15486
rect 41134 15538 41186 15550
rect 41134 15474 41186 15486
rect 3166 15426 3218 15438
rect 28254 15426 28306 15438
rect 10658 15374 10670 15426
rect 10722 15374 10734 15426
rect 20738 15374 20750 15426
rect 20802 15374 20814 15426
rect 21858 15374 21870 15426
rect 21922 15374 21934 15426
rect 3166 15362 3218 15374
rect 28254 15362 28306 15374
rect 33406 15426 33458 15438
rect 40014 15426 40066 15438
rect 35634 15374 35646 15426
rect 35698 15374 35710 15426
rect 33406 15362 33458 15374
rect 40014 15362 40066 15374
rect 40126 15426 40178 15438
rect 40126 15362 40178 15374
rect 41022 15426 41074 15438
rect 42354 15374 42366 15426
rect 42418 15374 42430 15426
rect 41022 15362 41074 15374
rect 3278 15314 3330 15326
rect 28590 15314 28642 15326
rect 37662 15314 37714 15326
rect 41358 15314 41410 15326
rect 9762 15262 9774 15314
rect 9826 15262 9838 15314
rect 10546 15262 10558 15314
rect 10610 15262 10622 15314
rect 11106 15262 11118 15314
rect 11170 15262 11182 15314
rect 11330 15262 11342 15314
rect 11394 15262 11406 15314
rect 12002 15262 12014 15314
rect 12066 15262 12078 15314
rect 20850 15262 20862 15314
rect 20914 15262 20926 15314
rect 22530 15262 22542 15314
rect 22594 15262 22606 15314
rect 33170 15262 33182 15314
rect 33234 15262 33246 15314
rect 35298 15262 35310 15314
rect 35362 15262 35374 15314
rect 36642 15262 36654 15314
rect 36706 15262 36718 15314
rect 38434 15262 38446 15314
rect 38498 15262 38510 15314
rect 41570 15262 41582 15314
rect 41634 15262 41646 15314
rect 3278 15250 3330 15262
rect 28590 15250 28642 15262
rect 37662 15250 37714 15262
rect 41358 15250 41410 15262
rect 3614 15202 3666 15214
rect 31166 15202 31218 15214
rect 9986 15150 9998 15202
rect 10050 15150 10062 15202
rect 22418 15150 22430 15202
rect 22482 15150 22494 15202
rect 44482 15150 44494 15202
rect 44546 15150 44558 15202
rect 3614 15138 3666 15150
rect 31166 15138 31218 15150
rect 3502 15090 3554 15102
rect 3502 15026 3554 15038
rect 11902 15090 11954 15102
rect 11902 15026 11954 15038
rect 40126 15090 40178 15102
rect 40126 15026 40178 15038
rect 1344 14922 48608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48608 14922
rect 1344 14836 48608 14870
rect 12574 14754 12626 14766
rect 20402 14702 20414 14754
rect 20466 14751 20478 14754
rect 20626 14751 20638 14754
rect 20466 14705 20638 14751
rect 20466 14702 20478 14705
rect 20626 14702 20638 14705
rect 20690 14702 20702 14754
rect 12574 14690 12626 14702
rect 2046 14642 2098 14654
rect 2046 14578 2098 14590
rect 2830 14642 2882 14654
rect 14030 14642 14082 14654
rect 19742 14642 19794 14654
rect 9986 14590 9998 14642
rect 10050 14590 10062 14642
rect 11442 14590 11454 14642
rect 11506 14590 11518 14642
rect 15922 14590 15934 14642
rect 15986 14590 15998 14642
rect 2830 14578 2882 14590
rect 14030 14578 14082 14590
rect 19742 14578 19794 14590
rect 20190 14642 20242 14654
rect 20190 14578 20242 14590
rect 20638 14642 20690 14654
rect 20638 14578 20690 14590
rect 24894 14642 24946 14654
rect 24894 14578 24946 14590
rect 28702 14642 28754 14654
rect 34974 14642 35026 14654
rect 31490 14590 31502 14642
rect 31554 14590 31566 14642
rect 33618 14590 33630 14642
rect 33682 14590 33694 14642
rect 28702 14578 28754 14590
rect 34974 14578 35026 14590
rect 35422 14642 35474 14654
rect 35422 14578 35474 14590
rect 36542 14642 36594 14654
rect 36542 14578 36594 14590
rect 37214 14642 37266 14654
rect 37214 14578 37266 14590
rect 38446 14642 38498 14654
rect 40114 14590 40126 14642
rect 40178 14590 40190 14642
rect 42242 14590 42254 14642
rect 42306 14590 42318 14642
rect 38446 14578 38498 14590
rect 2270 14530 2322 14542
rect 19070 14530 19122 14542
rect 29262 14530 29314 14542
rect 3154 14478 3166 14530
rect 3218 14478 3230 14530
rect 9874 14478 9886 14530
rect 9938 14478 9950 14530
rect 11890 14478 11902 14530
rect 11954 14478 11966 14530
rect 14914 14478 14926 14530
rect 14978 14478 14990 14530
rect 22418 14478 22430 14530
rect 22482 14478 22494 14530
rect 23314 14478 23326 14530
rect 23378 14478 23390 14530
rect 24322 14478 24334 14530
rect 24386 14478 24398 14530
rect 2270 14466 2322 14478
rect 19070 14466 19122 14478
rect 29262 14466 29314 14478
rect 30158 14530 30210 14542
rect 30158 14466 30210 14478
rect 30382 14530 30434 14542
rect 39006 14530 39058 14542
rect 34402 14478 34414 14530
rect 34466 14478 34478 14530
rect 39442 14478 39454 14530
rect 39506 14478 39518 14530
rect 30382 14466 30434 14478
rect 39006 14466 39058 14478
rect 3838 14418 3890 14430
rect 3838 14354 3890 14366
rect 12798 14418 12850 14430
rect 19182 14418 19234 14430
rect 18050 14366 18062 14418
rect 18114 14366 18126 14418
rect 18834 14366 18846 14418
rect 18898 14366 18910 14418
rect 12798 14354 12850 14366
rect 19182 14354 19234 14366
rect 22542 14418 22594 14430
rect 29374 14418 29426 14430
rect 23538 14366 23550 14418
rect 23602 14366 23614 14418
rect 22542 14354 22594 14366
rect 29374 14354 29426 14366
rect 30830 14418 30882 14430
rect 30830 14354 30882 14366
rect 42926 14418 42978 14430
rect 42926 14354 42978 14366
rect 3278 14306 3330 14318
rect 1698 14254 1710 14306
rect 1762 14254 1774 14306
rect 3278 14242 3330 14254
rect 3726 14306 3778 14318
rect 3726 14242 3778 14254
rect 4846 14306 4898 14318
rect 4846 14242 4898 14254
rect 12686 14306 12738 14318
rect 12686 14242 12738 14254
rect 13582 14306 13634 14318
rect 13582 14242 13634 14254
rect 17390 14306 17442 14318
rect 24110 14306 24162 14318
rect 22642 14254 22654 14306
rect 22706 14254 22718 14306
rect 17390 14242 17442 14254
rect 24110 14242 24162 14254
rect 29598 14306 29650 14318
rect 37998 14306 38050 14318
rect 29810 14254 29822 14306
rect 29874 14254 29886 14306
rect 29598 14242 29650 14254
rect 37998 14242 38050 14254
rect 42814 14306 42866 14318
rect 42814 14242 42866 14254
rect 1344 14138 48608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48608 14138
rect 1344 14052 48608 14086
rect 5070 13970 5122 13982
rect 5070 13906 5122 13918
rect 5518 13970 5570 13982
rect 5518 13906 5570 13918
rect 5630 13970 5682 13982
rect 5630 13906 5682 13918
rect 5742 13970 5794 13982
rect 5742 13906 5794 13918
rect 10446 13970 10498 13982
rect 10446 13906 10498 13918
rect 13022 13970 13074 13982
rect 13022 13906 13074 13918
rect 22542 13970 22594 13982
rect 24222 13970 24274 13982
rect 22642 13918 22654 13970
rect 22706 13918 22718 13970
rect 22542 13906 22594 13918
rect 24222 13906 24274 13918
rect 24670 13970 24722 13982
rect 37886 13970 37938 13982
rect 30594 13918 30606 13970
rect 30658 13918 30670 13970
rect 33618 13918 33630 13970
rect 33682 13918 33694 13970
rect 24670 13906 24722 13918
rect 37886 13906 37938 13918
rect 10222 13858 10274 13870
rect 5182 13802 5234 13814
rect 6066 13806 6078 13858
rect 6130 13806 6142 13858
rect 1810 13694 1822 13746
rect 1874 13694 1886 13746
rect 5182 13738 5234 13750
rect 6862 13802 6914 13814
rect 10222 13794 10274 13806
rect 11230 13858 11282 13870
rect 13470 13858 13522 13870
rect 12226 13806 12238 13858
rect 12290 13806 12302 13858
rect 20178 13806 20190 13858
rect 20242 13806 20254 13858
rect 21074 13806 21086 13858
rect 21138 13806 21150 13858
rect 23314 13806 23326 13858
rect 23378 13806 23390 13858
rect 27794 13806 27806 13858
rect 27858 13806 27870 13858
rect 30482 13806 30494 13858
rect 30546 13806 30558 13858
rect 31602 13806 31614 13858
rect 31666 13806 31678 13858
rect 38994 13806 39006 13858
rect 39058 13806 39070 13858
rect 41682 13806 41694 13858
rect 41746 13806 41758 13858
rect 11230 13794 11282 13806
rect 13470 13794 13522 13806
rect 5954 13694 5966 13746
rect 6018 13694 6030 13746
rect 6862 13738 6914 13750
rect 12910 13746 12962 13758
rect 17726 13746 17778 13758
rect 12562 13694 12574 13746
rect 12626 13694 12638 13746
rect 13906 13694 13918 13746
rect 13970 13694 13982 13746
rect 12910 13682 12962 13694
rect 17726 13682 17778 13694
rect 17950 13746 18002 13758
rect 17950 13682 18002 13694
rect 18846 13746 18898 13758
rect 33294 13746 33346 13758
rect 21746 13694 21758 13746
rect 21810 13694 21822 13746
rect 22306 13694 22318 13746
rect 22370 13694 22382 13746
rect 23426 13694 23438 13746
rect 23490 13694 23502 13746
rect 27122 13694 27134 13746
rect 27186 13694 27198 13746
rect 30258 13694 30270 13746
rect 30322 13694 30334 13746
rect 31266 13694 31278 13746
rect 31330 13694 31342 13746
rect 18846 13682 18898 13694
rect 33294 13682 33346 13694
rect 34078 13746 34130 13758
rect 34078 13682 34130 13694
rect 36878 13746 36930 13758
rect 36878 13682 36930 13694
rect 37102 13746 37154 13758
rect 37102 13682 37154 13694
rect 38670 13746 38722 13758
rect 39106 13694 39118 13746
rect 39170 13694 39182 13746
rect 39890 13694 39902 13746
rect 39954 13694 39966 13746
rect 40898 13694 40910 13746
rect 40962 13694 40974 13746
rect 38670 13682 38722 13694
rect 9662 13634 9714 13646
rect 2482 13582 2494 13634
rect 2546 13582 2558 13634
rect 4610 13582 4622 13634
rect 4674 13582 4686 13634
rect 9662 13570 9714 13582
rect 10334 13634 10386 13646
rect 18398 13634 18450 13646
rect 26686 13634 26738 13646
rect 33070 13634 33122 13646
rect 11554 13582 11566 13634
rect 11618 13582 11630 13634
rect 11890 13582 11902 13634
rect 11954 13582 11966 13634
rect 14690 13582 14702 13634
rect 14754 13582 14766 13634
rect 16818 13582 16830 13634
rect 16882 13582 16894 13634
rect 20514 13582 20526 13634
rect 20578 13582 20590 13634
rect 29922 13582 29934 13634
rect 29986 13582 29998 13634
rect 31378 13582 31390 13634
rect 31442 13582 31454 13634
rect 40226 13582 40238 13634
rect 40290 13582 40302 13634
rect 43810 13582 43822 13634
rect 43874 13582 43886 13634
rect 10334 13570 10386 13582
rect 18398 13570 18450 13582
rect 26686 13570 26738 13582
rect 33070 13570 33122 13582
rect 6974 13522 7026 13534
rect 6974 13458 7026 13470
rect 9550 13522 9602 13534
rect 9550 13458 9602 13470
rect 13022 13522 13074 13534
rect 13022 13458 13074 13470
rect 13582 13522 13634 13534
rect 17378 13470 17390 13522
rect 17442 13470 17454 13522
rect 37426 13470 37438 13522
rect 37490 13470 37502 13522
rect 13582 13458 13634 13470
rect 1344 13354 48608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48608 13354
rect 1344 13268 48608 13302
rect 5070 13186 5122 13198
rect 5070 13122 5122 13134
rect 5966 13186 6018 13198
rect 5966 13122 6018 13134
rect 12462 13186 12514 13198
rect 12462 13122 12514 13134
rect 30942 13186 30994 13198
rect 30942 13122 30994 13134
rect 31614 13186 31666 13198
rect 31614 13122 31666 13134
rect 35982 13186 36034 13198
rect 35982 13122 36034 13134
rect 3390 13074 3442 13086
rect 3390 13010 3442 13022
rect 6862 13074 6914 13086
rect 6862 13010 6914 13022
rect 11678 13074 11730 13086
rect 11678 13010 11730 13022
rect 14702 13074 14754 13086
rect 14702 13010 14754 13022
rect 16830 13074 16882 13086
rect 16830 13010 16882 13022
rect 17054 13074 17106 13086
rect 25118 13074 25170 13086
rect 19506 13022 19518 13074
rect 19570 13022 19582 13074
rect 22530 13022 22542 13074
rect 22594 13022 22606 13074
rect 24658 13022 24670 13074
rect 24722 13022 24734 13074
rect 17054 13010 17106 13022
rect 25118 13010 25170 13022
rect 33406 13074 33458 13086
rect 33406 13010 33458 13022
rect 34078 13074 34130 13086
rect 34078 13010 34130 13022
rect 34302 13074 34354 13086
rect 34302 13010 34354 13022
rect 35646 13074 35698 13086
rect 40574 13074 40626 13086
rect 39890 13022 39902 13074
rect 39954 13022 39966 13074
rect 35646 13010 35698 13022
rect 40574 13010 40626 13022
rect 3278 12962 3330 12974
rect 3278 12898 3330 12910
rect 3502 12962 3554 12974
rect 3502 12898 3554 12910
rect 4286 12962 4338 12974
rect 4286 12898 4338 12910
rect 4958 12962 5010 12974
rect 4958 12898 5010 12910
rect 6078 12962 6130 12974
rect 6078 12898 6130 12910
rect 6302 12962 6354 12974
rect 6302 12898 6354 12910
rect 8654 12962 8706 12974
rect 10110 12962 10162 12974
rect 12238 12962 12290 12974
rect 15374 12962 15426 12974
rect 9314 12910 9326 12962
rect 9378 12910 9390 12962
rect 10434 12910 10446 12962
rect 10498 12910 10510 12962
rect 11330 12910 11342 12962
rect 11394 12910 11406 12962
rect 14242 12910 14254 12962
rect 14306 12910 14318 12962
rect 8654 12898 8706 12910
rect 10110 12898 10162 12910
rect 12238 12898 12290 12910
rect 15374 12898 15426 12910
rect 17614 12962 17666 12974
rect 31726 12962 31778 12974
rect 20066 12910 20078 12962
rect 20130 12910 20142 12962
rect 21858 12910 21870 12962
rect 21922 12910 21934 12962
rect 25778 12910 25790 12962
rect 25842 12910 25854 12962
rect 29362 12910 29374 12962
rect 29426 12910 29438 12962
rect 17614 12898 17666 12910
rect 31726 12898 31778 12910
rect 32174 12962 32226 12974
rect 32174 12898 32226 12910
rect 36094 12962 36146 12974
rect 36978 12910 36990 12962
rect 37042 12910 37054 12962
rect 36094 12898 36146 12910
rect 3726 12850 3778 12862
rect 1698 12798 1710 12850
rect 1762 12798 1774 12850
rect 2482 12798 2494 12850
rect 2546 12798 2558 12850
rect 3726 12786 3778 12798
rect 7310 12850 7362 12862
rect 11902 12850 11954 12862
rect 9426 12798 9438 12850
rect 9490 12798 9502 12850
rect 7310 12786 7362 12798
rect 11902 12786 11954 12798
rect 15038 12850 15090 12862
rect 15038 12786 15090 12798
rect 16046 12850 16098 12862
rect 31614 12850 31666 12862
rect 16482 12798 16494 12850
rect 16546 12798 16558 12850
rect 18946 12798 18958 12850
rect 19010 12798 19022 12850
rect 19842 12798 19854 12850
rect 19906 12798 19918 12850
rect 29922 12798 29934 12850
rect 29986 12798 29998 12850
rect 37762 12798 37774 12850
rect 37826 12798 37838 12850
rect 16046 12786 16098 12798
rect 31614 12786 31666 12798
rect 4846 12738 4898 12750
rect 4846 12674 4898 12686
rect 5966 12738 6018 12750
rect 5966 12674 6018 12686
rect 7870 12738 7922 12750
rect 7870 12674 7922 12686
rect 8318 12738 8370 12750
rect 8318 12674 8370 12686
rect 9886 12738 9938 12750
rect 9886 12674 9938 12686
rect 9998 12738 10050 12750
rect 13806 12738 13858 12750
rect 12786 12686 12798 12738
rect 12850 12686 12862 12738
rect 9998 12674 10050 12686
rect 13806 12674 13858 12686
rect 15710 12738 15762 12750
rect 15710 12674 15762 12686
rect 21422 12738 21474 12750
rect 21422 12674 21474 12686
rect 26014 12738 26066 12750
rect 26014 12674 26066 12686
rect 28590 12738 28642 12750
rect 28590 12674 28642 12686
rect 29598 12738 29650 12750
rect 33730 12686 33742 12738
rect 33794 12686 33806 12738
rect 29598 12674 29650 12686
rect 1344 12570 48608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48608 12570
rect 1344 12484 48608 12518
rect 1822 12402 1874 12414
rect 1822 12338 1874 12350
rect 4510 12402 4562 12414
rect 4510 12338 4562 12350
rect 5966 12402 6018 12414
rect 5966 12338 6018 12350
rect 10670 12402 10722 12414
rect 10670 12338 10722 12350
rect 15598 12402 15650 12414
rect 15598 12338 15650 12350
rect 16830 12402 16882 12414
rect 37550 12402 37602 12414
rect 23986 12350 23998 12402
rect 24050 12350 24062 12402
rect 16830 12338 16882 12350
rect 37550 12338 37602 12350
rect 4286 12290 4338 12302
rect 18846 12290 18898 12302
rect 9538 12238 9550 12290
rect 9602 12238 9614 12290
rect 12562 12238 12574 12290
rect 12626 12238 12638 12290
rect 17714 12238 17726 12290
rect 17778 12238 17790 12290
rect 18498 12238 18510 12290
rect 18562 12238 18574 12290
rect 4286 12226 4338 12238
rect 18846 12226 18898 12238
rect 23326 12290 23378 12302
rect 28478 12290 28530 12302
rect 24434 12238 24446 12290
rect 24498 12238 24510 12290
rect 27346 12238 27358 12290
rect 27410 12238 27422 12290
rect 23326 12226 23378 12238
rect 28478 12226 28530 12238
rect 28814 12290 28866 12302
rect 30370 12238 30382 12290
rect 30434 12238 30446 12290
rect 28814 12226 28866 12238
rect 4734 12178 4786 12190
rect 4734 12114 4786 12126
rect 5182 12178 5234 12190
rect 5182 12114 5234 12126
rect 5854 12178 5906 12190
rect 18622 12178 18674 12190
rect 33182 12178 33234 12190
rect 6850 12126 6862 12178
rect 6914 12126 6926 12178
rect 8082 12126 8094 12178
rect 8146 12126 8158 12178
rect 8978 12126 8990 12178
rect 9042 12126 9054 12178
rect 9986 12126 9998 12178
rect 10050 12126 10062 12178
rect 11554 12126 11566 12178
rect 11618 12126 11630 12178
rect 12898 12126 12910 12178
rect 12962 12126 12974 12178
rect 14130 12126 14142 12178
rect 14194 12126 14206 12178
rect 15250 12126 15262 12178
rect 15314 12126 15326 12178
rect 19058 12126 19070 12178
rect 19122 12126 19134 12178
rect 23090 12126 23102 12178
rect 23154 12126 23166 12178
rect 24546 12126 24558 12178
rect 24610 12126 24622 12178
rect 28018 12126 28030 12178
rect 28082 12126 28094 12178
rect 29698 12126 29710 12178
rect 29762 12126 29774 12178
rect 33730 12126 33742 12178
rect 33794 12126 33806 12178
rect 37314 12126 37326 12178
rect 37378 12126 37390 12178
rect 5854 12114 5906 12126
rect 18622 12114 18674 12126
rect 33182 12114 33234 12126
rect 4622 12066 4674 12078
rect 4622 12002 4674 12014
rect 5070 12066 5122 12078
rect 12014 12066 12066 12078
rect 7186 12014 7198 12066
rect 7250 12014 7262 12066
rect 10210 12014 10222 12066
rect 10274 12014 10286 12066
rect 11666 12014 11678 12066
rect 11730 12014 11742 12066
rect 13682 12014 13694 12066
rect 13746 12014 13758 12066
rect 19842 12014 19854 12066
rect 19906 12014 19918 12066
rect 21970 12014 21982 12066
rect 22034 12014 22046 12066
rect 25218 12014 25230 12066
rect 25282 12014 25294 12066
rect 32498 12014 32510 12066
rect 32562 12014 32574 12066
rect 34514 12014 34526 12066
rect 34578 12014 34590 12066
rect 36642 12014 36654 12066
rect 36706 12014 36718 12066
rect 5070 12002 5122 12014
rect 12014 12002 12066 12014
rect 5630 11954 5682 11966
rect 5630 11890 5682 11902
rect 1344 11786 48608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48608 11786
rect 1344 11700 48608 11734
rect 6526 11618 6578 11630
rect 6526 11554 6578 11566
rect 8094 11618 8146 11630
rect 18498 11566 18510 11618
rect 18562 11615 18574 11618
rect 19730 11615 19742 11618
rect 18562 11569 19742 11615
rect 18562 11566 18574 11569
rect 19730 11566 19742 11569
rect 19794 11566 19806 11618
rect 23650 11566 23662 11618
rect 23714 11566 23726 11618
rect 8094 11554 8146 11566
rect 5070 11506 5122 11518
rect 4834 11454 4846 11506
rect 4898 11454 4910 11506
rect 5070 11442 5122 11454
rect 5742 11506 5794 11518
rect 5742 11442 5794 11454
rect 6862 11506 6914 11518
rect 6862 11442 6914 11454
rect 7758 11506 7810 11518
rect 7758 11442 7810 11454
rect 8654 11506 8706 11518
rect 8654 11442 8706 11454
rect 9326 11506 9378 11518
rect 14142 11506 14194 11518
rect 17838 11506 17890 11518
rect 11330 11454 11342 11506
rect 11394 11454 11406 11506
rect 15250 11454 15262 11506
rect 15314 11454 15326 11506
rect 17378 11454 17390 11506
rect 17442 11454 17454 11506
rect 9326 11442 9378 11454
rect 14142 11442 14194 11454
rect 17838 11442 17890 11454
rect 18734 11506 18786 11518
rect 18734 11442 18786 11454
rect 19182 11506 19234 11518
rect 19182 11442 19234 11454
rect 19742 11506 19794 11518
rect 19742 11442 19794 11454
rect 21870 11506 21922 11518
rect 21870 11442 21922 11454
rect 24670 11506 24722 11518
rect 24670 11442 24722 11454
rect 25118 11506 25170 11518
rect 33406 11506 33458 11518
rect 25442 11454 25454 11506
rect 25506 11454 25518 11506
rect 27570 11454 27582 11506
rect 27634 11454 27646 11506
rect 25118 11442 25170 11454
rect 33406 11442 33458 11454
rect 35086 11506 35138 11518
rect 35086 11442 35138 11454
rect 5518 11394 5570 11406
rect 5518 11330 5570 11342
rect 5854 11394 5906 11406
rect 5854 11330 5906 11342
rect 6190 11394 6242 11406
rect 6190 11330 6242 11342
rect 6638 11394 6690 11406
rect 6638 11330 6690 11342
rect 6974 11394 7026 11406
rect 6974 11330 7026 11342
rect 8318 11394 8370 11406
rect 8318 11330 8370 11342
rect 8542 11394 8594 11406
rect 21646 11394 21698 11406
rect 11442 11342 11454 11394
rect 11506 11342 11518 11394
rect 12226 11342 12238 11394
rect 12290 11342 12302 11394
rect 14466 11342 14478 11394
rect 14530 11342 14542 11394
rect 8542 11330 8594 11342
rect 21646 11330 21698 11342
rect 23102 11394 23154 11406
rect 23102 11330 23154 11342
rect 23326 11394 23378 11406
rect 23326 11330 23378 11342
rect 24110 11394 24162 11406
rect 33966 11394 34018 11406
rect 39454 11394 39506 11406
rect 28242 11342 28254 11394
rect 28306 11342 28318 11394
rect 35298 11342 35310 11394
rect 35362 11342 35374 11394
rect 24110 11330 24162 11342
rect 33966 11330 34018 11342
rect 39454 11330 39506 11342
rect 4846 11282 4898 11294
rect 4846 11218 4898 11230
rect 8766 11282 8818 11294
rect 13470 11282 13522 11294
rect 11218 11230 11230 11282
rect 11282 11230 11294 11282
rect 8766 11218 8818 11230
rect 13470 11218 13522 11230
rect 20190 11282 20242 11294
rect 20190 11218 20242 11230
rect 20526 11282 20578 11294
rect 34974 11282 35026 11294
rect 21298 11230 21310 11282
rect 21362 11230 21374 11282
rect 20526 11218 20578 11230
rect 34974 11218 35026 11230
rect 39566 11282 39618 11294
rect 39566 11218 39618 11230
rect 10782 11170 10834 11182
rect 10782 11106 10834 11118
rect 12910 11170 12962 11182
rect 12910 11106 12962 11118
rect 13582 11170 13634 11182
rect 13582 11106 13634 11118
rect 13806 11170 13858 11182
rect 13806 11106 13858 11118
rect 22766 11170 22818 11182
rect 22766 11106 22818 11118
rect 34302 11170 34354 11182
rect 34302 11106 34354 11118
rect 40014 11170 40066 11182
rect 40014 11106 40066 11118
rect 1344 11002 48608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48608 11002
rect 1344 10916 48608 10950
rect 3390 10834 3442 10846
rect 3390 10770 3442 10782
rect 3950 10834 4002 10846
rect 3950 10770 4002 10782
rect 5966 10834 6018 10846
rect 5966 10770 6018 10782
rect 10334 10834 10386 10846
rect 10334 10770 10386 10782
rect 17614 10834 17666 10846
rect 17614 10770 17666 10782
rect 30158 10834 30210 10846
rect 30158 10770 30210 10782
rect 31166 10834 31218 10846
rect 31166 10770 31218 10782
rect 31950 10834 32002 10846
rect 31950 10770 32002 10782
rect 38558 10834 38610 10846
rect 38558 10770 38610 10782
rect 39118 10834 39170 10846
rect 39118 10770 39170 10782
rect 40910 10834 40962 10846
rect 40910 10770 40962 10782
rect 34638 10722 34690 10734
rect 34638 10658 34690 10670
rect 38894 10722 38946 10734
rect 38894 10658 38946 10670
rect 39790 10722 39842 10734
rect 39790 10658 39842 10670
rect 3502 10610 3554 10622
rect 2706 10558 2718 10610
rect 2770 10558 2782 10610
rect 3502 10546 3554 10558
rect 6078 10610 6130 10622
rect 10770 10558 10782 10610
rect 10834 10558 10846 10610
rect 12114 10558 12126 10610
rect 12178 10558 12190 10610
rect 12562 10558 12574 10610
rect 12626 10558 12638 10610
rect 13570 10558 13582 10610
rect 13634 10558 13646 10610
rect 14242 10558 14254 10610
rect 14306 10558 14318 10610
rect 40114 10558 40126 10610
rect 40178 10558 40190 10610
rect 6078 10546 6130 10558
rect 2046 10498 2098 10510
rect 20974 10498 21026 10510
rect 2930 10446 2942 10498
rect 2994 10446 3006 10498
rect 13346 10446 13358 10498
rect 13410 10446 13422 10498
rect 16594 10446 16606 10498
rect 16658 10446 16670 10498
rect 2046 10434 2098 10446
rect 20974 10434 21026 10446
rect 39006 10498 39058 10510
rect 39006 10434 39058 10446
rect 41022 10498 41074 10510
rect 41022 10434 41074 10446
rect 40126 10386 40178 10398
rect 11218 10334 11230 10386
rect 11282 10334 11294 10386
rect 40126 10322 40178 10334
rect 1344 10218 48608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48608 10218
rect 1344 10132 48608 10166
rect 29934 10050 29986 10062
rect 29934 9986 29986 9998
rect 31054 10050 31106 10062
rect 31054 9986 31106 9998
rect 31166 10050 31218 10062
rect 31166 9986 31218 9998
rect 33294 10050 33346 10062
rect 33294 9986 33346 9998
rect 3054 9938 3106 9950
rect 3054 9874 3106 9886
rect 6750 9938 6802 9950
rect 6750 9874 6802 9886
rect 9550 9938 9602 9950
rect 9550 9874 9602 9886
rect 15262 9938 15314 9950
rect 15262 9874 15314 9886
rect 16830 9938 16882 9950
rect 16830 9874 16882 9886
rect 17278 9938 17330 9950
rect 17278 9874 17330 9886
rect 21870 9938 21922 9950
rect 21870 9874 21922 9886
rect 23550 9938 23602 9950
rect 23550 9874 23602 9886
rect 24222 9938 24274 9950
rect 24222 9874 24274 9886
rect 24446 9938 24498 9950
rect 24446 9874 24498 9886
rect 33854 9938 33906 9950
rect 38434 9886 38446 9938
rect 38498 9886 38510 9938
rect 40562 9886 40574 9938
rect 40626 9886 40638 9938
rect 40898 9886 40910 9938
rect 40962 9886 40974 9938
rect 43026 9886 43038 9938
rect 43090 9886 43102 9938
rect 33854 9874 33906 9886
rect 2382 9826 2434 9838
rect 2382 9762 2434 9774
rect 10110 9826 10162 9838
rect 10110 9762 10162 9774
rect 10558 9826 10610 9838
rect 13582 9826 13634 9838
rect 11554 9774 11566 9826
rect 11618 9774 11630 9826
rect 11890 9774 11902 9826
rect 11954 9774 11966 9826
rect 12450 9774 12462 9826
rect 12514 9774 12526 9826
rect 10558 9762 10610 9774
rect 13582 9762 13634 9774
rect 21646 9826 21698 9838
rect 29362 9774 29374 9826
rect 29426 9774 29438 9826
rect 30482 9774 30494 9826
rect 30546 9774 30558 9826
rect 31714 9774 31726 9826
rect 31778 9774 31790 9826
rect 32498 9774 32510 9826
rect 32562 9774 32574 9826
rect 37650 9774 37662 9826
rect 37714 9774 37726 9826
rect 43698 9774 43710 9826
rect 43762 9774 43774 9826
rect 21646 9762 21698 9774
rect 2494 9714 2546 9726
rect 14030 9714 14082 9726
rect 12562 9662 12574 9714
rect 12626 9662 12638 9714
rect 2494 9650 2546 9662
rect 14030 9650 14082 9662
rect 18286 9714 18338 9726
rect 18286 9650 18338 9662
rect 29822 9714 29874 9726
rect 29822 9650 29874 9662
rect 33406 9714 33458 9726
rect 33406 9650 33458 9662
rect 2718 9602 2770 9614
rect 2718 9538 2770 9550
rect 10446 9602 10498 9614
rect 10446 9538 10498 9550
rect 14926 9602 14978 9614
rect 14926 9538 14978 9550
rect 17950 9602 18002 9614
rect 17950 9538 18002 9550
rect 20750 9602 20802 9614
rect 28590 9602 28642 9614
rect 21298 9550 21310 9602
rect 21362 9550 21374 9602
rect 23874 9550 23886 9602
rect 23938 9550 23950 9602
rect 20750 9538 20802 9550
rect 28590 9538 28642 9550
rect 29598 9602 29650 9614
rect 29598 9538 29650 9550
rect 30718 9602 30770 9614
rect 30718 9538 30770 9550
rect 30942 9602 30994 9614
rect 30942 9538 30994 9550
rect 31278 9602 31330 9614
rect 31278 9538 31330 9550
rect 31502 9602 31554 9614
rect 31502 9538 31554 9550
rect 32286 9602 32338 9614
rect 32286 9538 32338 9550
rect 37326 9602 37378 9614
rect 37326 9538 37378 9550
rect 1344 9434 48608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48608 9434
rect 1344 9348 48608 9382
rect 2718 9266 2770 9278
rect 2718 9202 2770 9214
rect 3390 9266 3442 9278
rect 3390 9202 3442 9214
rect 4622 9266 4674 9278
rect 4622 9202 4674 9214
rect 22654 9266 22706 9278
rect 22654 9202 22706 9214
rect 26574 9266 26626 9278
rect 26574 9202 26626 9214
rect 27358 9266 27410 9278
rect 27358 9202 27410 9214
rect 28590 9266 28642 9278
rect 28590 9202 28642 9214
rect 28926 9266 28978 9278
rect 28926 9202 28978 9214
rect 30158 9266 30210 9278
rect 30158 9202 30210 9214
rect 30606 9266 30658 9278
rect 30606 9202 30658 9214
rect 30942 9266 30994 9278
rect 30942 9202 30994 9214
rect 31502 9266 31554 9278
rect 32386 9214 32398 9266
rect 32450 9214 32462 9266
rect 31502 9202 31554 9214
rect 5630 9154 5682 9166
rect 5630 9090 5682 9102
rect 5854 9154 5906 9166
rect 20862 9154 20914 9166
rect 18162 9102 18174 9154
rect 18226 9102 18238 9154
rect 5854 9090 5906 9102
rect 20862 9090 20914 9102
rect 21198 9154 21250 9166
rect 21198 9090 21250 9102
rect 23998 9154 24050 9166
rect 23998 9090 24050 9102
rect 24334 9154 24386 9166
rect 24334 9090 24386 9102
rect 29374 9154 29426 9166
rect 41022 9154 41074 9166
rect 34178 9102 34190 9154
rect 34242 9102 34254 9154
rect 29374 9090 29426 9102
rect 41022 9090 41074 9102
rect 2606 9042 2658 9054
rect 2606 8978 2658 8990
rect 2942 9042 2994 9054
rect 2942 8978 2994 8990
rect 3166 9042 3218 9054
rect 3166 8978 3218 8990
rect 3838 9042 3890 9054
rect 3838 8978 3890 8990
rect 5966 9042 6018 9054
rect 16606 9042 16658 9054
rect 6514 8990 6526 9042
rect 6578 8990 6590 9042
rect 7858 8990 7870 9042
rect 7922 8990 7934 9042
rect 8194 8990 8206 9042
rect 8258 8990 8270 9042
rect 10434 8990 10446 9042
rect 10498 8990 10510 9042
rect 10994 8990 11006 9042
rect 11058 8990 11070 9042
rect 12002 8990 12014 9042
rect 12066 8990 12078 9042
rect 12338 8990 12350 9042
rect 12402 8990 12414 9042
rect 12674 8990 12686 9042
rect 12738 8990 12750 9042
rect 14354 8990 14366 9042
rect 14418 8990 14430 9042
rect 15362 8990 15374 9042
rect 15426 8990 15438 9042
rect 5966 8978 6018 8990
rect 16606 8978 16658 8990
rect 16830 9042 16882 9054
rect 27806 9042 27858 9054
rect 32062 9042 32114 9054
rect 17490 8990 17502 9042
rect 17554 8990 17566 9042
rect 26898 8990 26910 9042
rect 26962 8990 26974 9042
rect 27122 8990 27134 9042
rect 27186 8990 27198 9042
rect 29138 8990 29150 9042
rect 29202 8990 29214 9042
rect 33394 8990 33406 9042
rect 33458 8990 33470 9042
rect 16830 8978 16882 8990
rect 27806 8978 27858 8990
rect 32062 8978 32114 8990
rect 3278 8930 3330 8942
rect 3278 8866 3330 8878
rect 4174 8930 4226 8942
rect 27022 8930 27074 8942
rect 31838 8930 31890 8942
rect 11442 8878 11454 8930
rect 11506 8878 11518 8930
rect 15138 8878 15150 8930
rect 15202 8878 15214 8930
rect 20290 8878 20302 8930
rect 20354 8878 20366 8930
rect 29026 8878 29038 8930
rect 29090 8878 29102 8930
rect 36306 8878 36318 8930
rect 36370 8878 36382 8930
rect 4174 8866 4226 8878
rect 27022 8866 27074 8878
rect 31838 8866 31890 8878
rect 6850 8766 6862 8818
rect 6914 8766 6926 8818
rect 15362 8766 15374 8818
rect 15426 8766 15438 8818
rect 16258 8766 16270 8818
rect 16322 8766 16334 8818
rect 1344 8650 48608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48608 8650
rect 1344 8564 48608 8598
rect 17950 8482 18002 8494
rect 10658 8430 10670 8482
rect 10722 8430 10734 8482
rect 18274 8430 18286 8482
rect 18338 8430 18350 8482
rect 17950 8418 18002 8430
rect 12910 8370 12962 8382
rect 4498 8318 4510 8370
rect 4562 8318 4574 8370
rect 8418 8318 8430 8370
rect 8482 8318 8494 8370
rect 11666 8318 11678 8370
rect 11730 8318 11742 8370
rect 12910 8306 12962 8318
rect 13918 8370 13970 8382
rect 17726 8370 17778 8382
rect 17154 8318 17166 8370
rect 17218 8318 17230 8370
rect 13918 8306 13970 8318
rect 17726 8306 17778 8318
rect 18846 8370 18898 8382
rect 18846 8306 18898 8318
rect 21870 8370 21922 8382
rect 21870 8306 21922 8318
rect 22430 8370 22482 8382
rect 22430 8306 22482 8318
rect 22654 8370 22706 8382
rect 37550 8370 37602 8382
rect 22978 8318 22990 8370
rect 23042 8318 23054 8370
rect 25106 8318 25118 8370
rect 25170 8318 25182 8370
rect 32274 8318 32286 8370
rect 32338 8318 32350 8370
rect 34402 8318 34414 8370
rect 34466 8318 34478 8370
rect 22654 8306 22706 8318
rect 37550 8306 37602 8318
rect 7422 8258 7474 8270
rect 35758 8258 35810 8270
rect 37326 8258 37378 8270
rect 2146 8206 2158 8258
rect 2210 8206 2222 8258
rect 5842 8206 5854 8258
rect 5906 8206 5918 8258
rect 6402 8206 6414 8258
rect 6466 8206 6478 8258
rect 7970 8206 7982 8258
rect 8034 8206 8046 8258
rect 9762 8206 9774 8258
rect 9826 8206 9838 8258
rect 10882 8206 10894 8258
rect 10946 8206 10958 8258
rect 14354 8206 14366 8258
rect 14418 8206 14430 8258
rect 25890 8206 25902 8258
rect 25954 8206 25966 8258
rect 31602 8206 31614 8258
rect 31666 8206 31678 8258
rect 36194 8206 36206 8258
rect 36258 8206 36270 8258
rect 7422 8194 7474 8206
rect 35758 8194 35810 8206
rect 37326 8194 37378 8206
rect 7086 8146 7138 8158
rect 7086 8082 7138 8094
rect 7198 8146 7250 8158
rect 27470 8146 27522 8158
rect 15026 8094 15038 8146
rect 15090 8094 15102 8146
rect 7198 8082 7250 8094
rect 27470 8082 27522 8094
rect 31166 8146 31218 8158
rect 36978 8094 36990 8146
rect 37042 8094 37054 8146
rect 31166 8082 31218 8094
rect 1822 8034 1874 8046
rect 27134 8034 27186 8046
rect 22082 7982 22094 8034
rect 22146 7982 22158 8034
rect 1822 7970 1874 7982
rect 27134 7970 27186 7982
rect 36430 8034 36482 8046
rect 36430 7970 36482 7982
rect 1344 7866 48608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48608 7866
rect 1344 7780 48608 7814
rect 2046 7698 2098 7710
rect 2046 7634 2098 7646
rect 2606 7698 2658 7710
rect 9550 7698 9602 7710
rect 7186 7646 7198 7698
rect 7250 7646 7262 7698
rect 2606 7634 2658 7646
rect 9550 7634 9602 7646
rect 15262 7698 15314 7710
rect 15262 7634 15314 7646
rect 33182 7698 33234 7710
rect 33182 7634 33234 7646
rect 35646 7698 35698 7710
rect 35646 7634 35698 7646
rect 2718 7586 2770 7598
rect 6526 7586 6578 7598
rect 9774 7586 9826 7598
rect 3266 7534 3278 7586
rect 3330 7534 3342 7586
rect 7746 7534 7758 7586
rect 7810 7534 7822 7586
rect 2718 7522 2770 7534
rect 6526 7522 6578 7534
rect 9774 7522 9826 7534
rect 9886 7586 9938 7598
rect 15598 7586 15650 7598
rect 11666 7534 11678 7586
rect 11730 7534 11742 7586
rect 20514 7534 20526 7586
rect 20578 7534 20590 7586
rect 27122 7534 27134 7586
rect 27186 7534 27198 7586
rect 36754 7534 36766 7586
rect 36818 7534 36830 7586
rect 9886 7522 9938 7534
rect 15598 7522 15650 7534
rect 2382 7474 2434 7486
rect 1810 7422 1822 7474
rect 1874 7422 1886 7474
rect 2382 7410 2434 7422
rect 3054 7474 3106 7486
rect 6638 7474 6690 7486
rect 3602 7422 3614 7474
rect 3666 7422 3678 7474
rect 4498 7422 4510 7474
rect 4562 7422 4574 7474
rect 4834 7422 4846 7474
rect 4898 7422 4910 7474
rect 3054 7410 3106 7422
rect 6638 7410 6690 7422
rect 6750 7474 6802 7486
rect 10670 7474 10722 7486
rect 7522 7422 7534 7474
rect 7586 7422 7598 7474
rect 8418 7422 8430 7474
rect 8482 7422 8494 7474
rect 10322 7422 10334 7474
rect 10386 7422 10398 7474
rect 6750 7410 6802 7422
rect 10670 7410 10722 7422
rect 10894 7474 10946 7486
rect 16046 7474 16098 7486
rect 11778 7422 11790 7474
rect 11842 7422 11854 7474
rect 14354 7422 14366 7474
rect 14418 7422 14430 7474
rect 14914 7422 14926 7474
rect 14978 7422 14990 7474
rect 19730 7422 19742 7474
rect 19794 7422 19806 7474
rect 26338 7422 26350 7474
rect 26402 7422 26414 7474
rect 29586 7422 29598 7474
rect 29650 7422 29662 7474
rect 35970 7422 35982 7474
rect 36034 7422 36046 7474
rect 10894 7410 10946 7422
rect 16046 7410 16098 7422
rect 10782 7362 10834 7374
rect 17502 7362 17554 7374
rect 7970 7310 7982 7362
rect 8034 7310 8046 7362
rect 12450 7310 12462 7362
rect 12514 7310 12526 7362
rect 10782 7298 10834 7310
rect 17502 7298 17554 7310
rect 17950 7362 18002 7374
rect 17950 7298 18002 7310
rect 19406 7362 19458 7374
rect 26014 7362 26066 7374
rect 22642 7310 22654 7362
rect 22706 7310 22718 7362
rect 29250 7310 29262 7362
rect 29314 7310 29326 7362
rect 30370 7310 30382 7362
rect 30434 7310 30446 7362
rect 32498 7310 32510 7362
rect 32562 7310 32574 7362
rect 38882 7310 38894 7362
rect 38946 7310 38958 7362
rect 19406 7298 19458 7310
rect 26014 7298 26066 7310
rect 4622 7250 4674 7262
rect 4622 7186 4674 7198
rect 5406 7250 5458 7262
rect 5406 7186 5458 7198
rect 1344 7082 48608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48608 7082
rect 1344 6996 48608 7030
rect 26898 6862 26910 6914
rect 26962 6862 26974 6914
rect 12686 6802 12738 6814
rect 3154 6750 3166 6802
rect 3218 6750 3230 6802
rect 10210 6750 10222 6802
rect 10274 6750 10286 6802
rect 12686 6738 12738 6750
rect 27470 6802 27522 6814
rect 27470 6738 27522 6750
rect 27918 6802 27970 6814
rect 27918 6738 27970 6750
rect 1710 6690 1762 6702
rect 1710 6626 1762 6638
rect 2270 6690 2322 6702
rect 3838 6690 3890 6702
rect 2930 6638 2942 6690
rect 2994 6638 3006 6690
rect 2270 6626 2322 6638
rect 3838 6626 3890 6638
rect 4398 6690 4450 6702
rect 4398 6626 4450 6638
rect 4958 6690 5010 6702
rect 7982 6690 8034 6702
rect 13358 6690 13410 6702
rect 6514 6638 6526 6690
rect 6578 6638 6590 6690
rect 8306 6638 8318 6690
rect 8370 6638 8382 6690
rect 10882 6638 10894 6690
rect 10946 6638 10958 6690
rect 11330 6638 11342 6690
rect 11394 6638 11406 6690
rect 12226 6638 12238 6690
rect 12290 6638 12302 6690
rect 4958 6626 5010 6638
rect 7982 6626 8034 6638
rect 13358 6626 13410 6638
rect 13470 6690 13522 6702
rect 13470 6626 13522 6638
rect 15150 6690 15202 6702
rect 15150 6626 15202 6638
rect 20302 6690 20354 6702
rect 27246 6690 27298 6702
rect 22194 6638 22206 6690
rect 22258 6638 22270 6690
rect 20302 6626 20354 6638
rect 27246 6626 27298 6638
rect 4510 6578 4562 6590
rect 4510 6514 4562 6526
rect 5070 6578 5122 6590
rect 8542 6578 8594 6590
rect 5954 6526 5966 6578
rect 6018 6526 6030 6578
rect 5070 6514 5122 6526
rect 8542 6514 8594 6526
rect 9326 6578 9378 6590
rect 9326 6514 9378 6526
rect 9550 6578 9602 6590
rect 30494 6578 30546 6590
rect 13682 6526 13694 6578
rect 13746 6526 13758 6578
rect 14242 6526 14254 6578
rect 14306 6526 14318 6578
rect 9550 6514 9602 6526
rect 30494 6514 30546 6526
rect 30830 6578 30882 6590
rect 30830 6514 30882 6526
rect 1822 6466 1874 6478
rect 1822 6402 1874 6414
rect 2046 6466 2098 6478
rect 2046 6402 2098 6414
rect 3950 6466 4002 6478
rect 3950 6402 4002 6414
rect 4174 6466 4226 6478
rect 9438 6466 9490 6478
rect 7298 6414 7310 6466
rect 7362 6414 7374 6466
rect 4174 6402 4226 6414
rect 9438 6402 9490 6414
rect 18622 6466 18674 6478
rect 18622 6402 18674 6414
rect 19070 6466 19122 6478
rect 19070 6402 19122 6414
rect 19518 6466 19570 6478
rect 19518 6402 19570 6414
rect 21982 6466 22034 6478
rect 21982 6402 22034 6414
rect 1344 6298 48608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48608 6298
rect 1344 6212 48608 6246
rect 2270 6130 2322 6142
rect 2270 6066 2322 6078
rect 3054 6130 3106 6142
rect 3054 6066 3106 6078
rect 4398 6130 4450 6142
rect 4398 6066 4450 6078
rect 5406 6130 5458 6142
rect 5406 6066 5458 6078
rect 7534 6130 7586 6142
rect 15486 6130 15538 6142
rect 27694 6130 27746 6142
rect 8306 6078 8318 6130
rect 8370 6078 8382 6130
rect 18386 6078 18398 6130
rect 18450 6078 18462 6130
rect 19058 6078 19070 6130
rect 19122 6127 19134 6130
rect 19282 6127 19294 6130
rect 19122 6081 19294 6127
rect 19122 6078 19134 6081
rect 19282 6078 19294 6081
rect 19346 6078 19358 6130
rect 27010 6078 27022 6130
rect 27074 6078 27086 6130
rect 7534 6066 7586 6078
rect 15486 6066 15538 6078
rect 27694 6066 27746 6078
rect 30382 6130 30434 6142
rect 31266 6078 31278 6130
rect 31330 6078 31342 6130
rect 30382 6066 30434 6078
rect 8878 6018 8930 6030
rect 14478 6018 14530 6030
rect 11218 5966 11230 6018
rect 11282 5966 11294 6018
rect 13122 5966 13134 6018
rect 13186 5966 13198 6018
rect 13794 5966 13806 6018
rect 13858 5966 13870 6018
rect 8878 5954 8930 5966
rect 14478 5954 14530 5966
rect 15038 6018 15090 6030
rect 20190 6018 20242 6030
rect 25790 6018 25842 6030
rect 30718 6018 30770 6030
rect 17714 5966 17726 6018
rect 17778 5966 17790 6018
rect 18274 5966 18286 6018
rect 18338 5966 18350 6018
rect 19282 5966 19294 6018
rect 19346 5966 19358 6018
rect 19618 5966 19630 6018
rect 19682 5966 19694 6018
rect 21522 5966 21534 6018
rect 21586 5966 21598 6018
rect 26338 5966 26350 6018
rect 26402 5966 26414 6018
rect 26674 5966 26686 6018
rect 26738 5966 26750 6018
rect 15038 5954 15090 5966
rect 20190 5954 20242 5966
rect 25790 5954 25842 5966
rect 30718 5954 30770 5966
rect 9886 5906 9938 5918
rect 7746 5854 7758 5906
rect 7810 5854 7822 5906
rect 7970 5854 7982 5906
rect 8034 5854 8046 5906
rect 9886 5842 9938 5854
rect 10110 5906 10162 5918
rect 14702 5906 14754 5918
rect 10770 5854 10782 5906
rect 10834 5854 10846 5906
rect 12226 5854 12238 5906
rect 12290 5854 12302 5906
rect 14018 5854 14030 5906
rect 14082 5854 14094 5906
rect 10110 5842 10162 5854
rect 14702 5842 14754 5854
rect 18622 5906 18674 5918
rect 18622 5842 18674 5854
rect 19966 5906 20018 5918
rect 27246 5906 27298 5918
rect 20738 5854 20750 5906
rect 20802 5854 20814 5906
rect 19966 5842 20018 5854
rect 27246 5842 27298 5854
rect 30942 5906 30994 5918
rect 30942 5842 30994 5854
rect 14926 5794 14978 5806
rect 34974 5794 35026 5806
rect 13794 5742 13806 5794
rect 13858 5742 13870 5794
rect 23650 5742 23662 5794
rect 23714 5742 23726 5794
rect 14926 5730 14978 5742
rect 34974 5730 35026 5742
rect 7422 5682 7474 5694
rect 7422 5618 7474 5630
rect 8654 5682 8706 5694
rect 8654 5618 8706 5630
rect 10446 5682 10498 5694
rect 10446 5618 10498 5630
rect 1344 5514 48608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48608 5514
rect 1344 5428 48608 5462
rect 15710 5346 15762 5358
rect 15710 5282 15762 5294
rect 34078 5346 34130 5358
rect 34078 5282 34130 5294
rect 35646 5346 35698 5358
rect 35646 5282 35698 5294
rect 37438 5346 37490 5358
rect 37438 5282 37490 5294
rect 15486 5234 15538 5246
rect 4610 5182 4622 5234
rect 4674 5182 4686 5234
rect 13458 5182 13470 5234
rect 13522 5182 13534 5234
rect 15486 5170 15538 5182
rect 20414 5234 20466 5246
rect 20414 5170 20466 5182
rect 21534 5234 21586 5246
rect 21534 5170 21586 5182
rect 23886 5234 23938 5246
rect 23886 5170 23938 5182
rect 28142 5234 28194 5246
rect 28142 5170 28194 5182
rect 32734 5234 32786 5246
rect 32734 5170 32786 5182
rect 33518 5234 33570 5246
rect 33518 5170 33570 5182
rect 34302 5234 34354 5246
rect 34302 5170 34354 5182
rect 34750 5234 34802 5246
rect 34750 5170 34802 5182
rect 35870 5234 35922 5246
rect 35870 5170 35922 5182
rect 36430 5234 36482 5246
rect 36430 5170 36482 5182
rect 37214 5234 37266 5246
rect 37214 5170 37266 5182
rect 6414 5122 6466 5134
rect 8542 5122 8594 5134
rect 12350 5122 12402 5134
rect 1698 5070 1710 5122
rect 1762 5070 1774 5122
rect 6626 5070 6638 5122
rect 6690 5070 6702 5122
rect 7522 5070 7534 5122
rect 7586 5070 7598 5122
rect 9090 5070 9102 5122
rect 9154 5070 9166 5122
rect 11218 5070 11230 5122
rect 11282 5070 11294 5122
rect 6414 5058 6466 5070
rect 8542 5058 8594 5070
rect 12350 5058 12402 5070
rect 12574 5122 12626 5134
rect 12574 5058 12626 5070
rect 12798 5122 12850 5134
rect 19854 5122 19906 5134
rect 14130 5070 14142 5122
rect 14194 5070 14206 5122
rect 14690 5070 14702 5122
rect 14754 5070 14766 5122
rect 12798 5058 12850 5070
rect 19854 5058 19906 5070
rect 21870 5122 21922 5134
rect 21870 5058 21922 5070
rect 23326 5122 23378 5134
rect 23326 5058 23378 5070
rect 24894 5122 24946 5134
rect 25790 5122 25842 5134
rect 25442 5070 25454 5122
rect 25506 5070 25518 5122
rect 24894 5058 24946 5070
rect 25790 5058 25842 5070
rect 26014 5122 26066 5134
rect 26014 5058 26066 5070
rect 26462 5122 26514 5134
rect 38110 5122 38162 5134
rect 37762 5070 37774 5122
rect 37826 5070 37838 5122
rect 26462 5058 26514 5070
rect 38110 5058 38162 5070
rect 17726 5010 17778 5022
rect 2482 4958 2494 5010
rect 2546 4958 2558 5010
rect 8978 4958 8990 5010
rect 9042 4958 9054 5010
rect 10322 4958 10334 5010
rect 10386 4958 10398 5010
rect 13794 4958 13806 5010
rect 13858 4958 13870 5010
rect 17726 4946 17778 4958
rect 18398 5010 18450 5022
rect 23438 5010 23490 5022
rect 19058 4958 19070 5010
rect 19122 4958 19134 5010
rect 19618 4958 19630 5010
rect 19682 4958 19694 5010
rect 22418 4958 22430 5010
rect 22482 4958 22494 5010
rect 23090 4958 23102 5010
rect 23154 4958 23166 5010
rect 18398 4946 18450 4958
rect 23438 4946 23490 4958
rect 5070 4898 5122 4910
rect 5070 4834 5122 4846
rect 6078 4898 6130 4910
rect 14478 4898 14530 4910
rect 16494 4898 16546 4910
rect 12002 4846 12014 4898
rect 12066 4846 12078 4898
rect 16034 4846 16046 4898
rect 16098 4846 16110 4898
rect 6078 4834 6130 4846
rect 14478 4834 14530 4846
rect 16494 4834 16546 4846
rect 17054 4898 17106 4910
rect 17054 4834 17106 4846
rect 18062 4898 18114 4910
rect 38446 4898 38498 4910
rect 19282 4846 19294 4898
rect 19346 4846 19358 4898
rect 33730 4846 33742 4898
rect 33794 4846 33806 4898
rect 35298 4846 35310 4898
rect 35362 4846 35374 4898
rect 18062 4834 18114 4846
rect 38446 4834 38498 4846
rect 1344 4730 48608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48608 4730
rect 1344 4644 48608 4678
rect 8878 4562 8930 4574
rect 8878 4498 8930 4510
rect 9662 4562 9714 4574
rect 9662 4498 9714 4510
rect 10334 4562 10386 4574
rect 10334 4498 10386 4510
rect 11006 4562 11058 4574
rect 12574 4562 12626 4574
rect 11106 4510 11118 4562
rect 11170 4510 11182 4562
rect 11006 4498 11058 4510
rect 12574 4498 12626 4510
rect 30942 4562 30994 4574
rect 30942 4498 30994 4510
rect 8430 4450 8482 4462
rect 8430 4386 8482 4398
rect 10446 4450 10498 4462
rect 12686 4450 12738 4462
rect 16382 4450 16434 4462
rect 23550 4450 23602 4462
rect 11778 4398 11790 4450
rect 11842 4398 11854 4450
rect 13906 4398 13918 4450
rect 13970 4398 13982 4450
rect 18162 4398 18174 4450
rect 18226 4398 18238 4450
rect 10446 4386 10498 4398
rect 12686 4386 12738 4398
rect 16382 4386 16434 4398
rect 23550 4386 23602 4398
rect 24670 4450 24722 4462
rect 29038 4450 29090 4462
rect 26002 4398 26014 4450
rect 26066 4398 26078 4450
rect 24670 4386 24722 4398
rect 29038 4386 29090 4398
rect 32510 4450 32562 4462
rect 33842 4398 33854 4450
rect 33906 4398 33918 4450
rect 32510 4386 32562 4398
rect 7198 4338 7250 4350
rect 23886 4338 23938 4350
rect 28814 4338 28866 4350
rect 7410 4286 7422 4338
rect 7474 4286 7486 4338
rect 10770 4286 10782 4338
rect 10834 4286 10846 4338
rect 12114 4286 12126 4338
rect 12178 4286 12190 4338
rect 13234 4286 13246 4338
rect 13298 4286 13310 4338
rect 16594 4286 16606 4338
rect 16658 4286 16670 4338
rect 17490 4286 17502 4338
rect 17554 4286 17566 4338
rect 24434 4286 24446 4338
rect 24498 4286 24510 4338
rect 25330 4286 25342 4338
rect 25394 4286 25406 4338
rect 7198 4274 7250 4286
rect 23886 4274 23938 4286
rect 28814 4274 28866 4286
rect 29934 4338 29986 4350
rect 29934 4274 29986 4286
rect 30158 4338 30210 4350
rect 32274 4286 32286 4338
rect 32338 4286 32350 4338
rect 33058 4286 33070 4338
rect 33122 4286 33134 4338
rect 39106 4286 39118 4338
rect 39170 4286 39182 4338
rect 30158 4274 30210 4286
rect 16034 4174 16046 4226
rect 16098 4174 16110 4226
rect 20290 4174 20302 4226
rect 20354 4174 20366 4226
rect 28130 4174 28142 4226
rect 28194 4174 28206 4226
rect 35970 4174 35982 4226
rect 36034 4174 36046 4226
rect 36306 4174 36318 4226
rect 36370 4174 36382 4226
rect 38434 4174 38446 4226
rect 38498 4174 38510 4226
rect 10334 4114 10386 4126
rect 10334 4050 10386 4062
rect 28478 4114 28530 4126
rect 30482 4062 30494 4114
rect 30546 4062 30558 4114
rect 28478 4050 28530 4062
rect 1344 3946 48608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48608 3946
rect 1344 3860 48608 3894
rect 14142 3778 14194 3790
rect 7410 3726 7422 3778
rect 7474 3726 7486 3778
rect 11330 3726 11342 3778
rect 11394 3726 11406 3778
rect 14142 3714 14194 3726
rect 33742 3778 33794 3790
rect 33742 3714 33794 3726
rect 5070 3666 5122 3678
rect 13022 3666 13074 3678
rect 2482 3614 2494 3666
rect 2546 3614 2558 3666
rect 4610 3614 4622 3666
rect 4674 3614 4686 3666
rect 8754 3614 8766 3666
rect 8818 3614 8830 3666
rect 10882 3614 10894 3666
rect 10946 3614 10958 3666
rect 12226 3614 12238 3666
rect 12290 3614 12302 3666
rect 5070 3602 5122 3614
rect 13022 3602 13074 3614
rect 14702 3666 14754 3678
rect 18734 3666 18786 3678
rect 15922 3614 15934 3666
rect 15986 3614 15998 3666
rect 18050 3614 18062 3666
rect 18114 3614 18126 3666
rect 14702 3602 14754 3614
rect 18734 3602 18786 3614
rect 18958 3666 19010 3678
rect 18958 3602 19010 3614
rect 19518 3666 19570 3678
rect 19518 3602 19570 3614
rect 22654 3666 22706 3678
rect 33070 3666 33122 3678
rect 23762 3614 23774 3666
rect 23826 3614 23838 3666
rect 25890 3614 25902 3666
rect 25954 3614 25966 3666
rect 29698 3614 29710 3666
rect 29762 3614 29774 3666
rect 22654 3602 22706 3614
rect 33070 3602 33122 3614
rect 33966 3666 34018 3678
rect 33966 3602 34018 3614
rect 34414 3666 34466 3678
rect 34414 3602 34466 3614
rect 36206 3666 36258 3678
rect 36978 3614 36990 3666
rect 37042 3614 37054 3666
rect 39106 3614 39118 3666
rect 39170 3614 39182 3666
rect 36206 3602 36258 3614
rect 6862 3554 6914 3566
rect 12014 3554 12066 3566
rect 1698 3502 1710 3554
rect 1762 3502 1774 3554
rect 6626 3502 6638 3554
rect 6690 3502 6702 3554
rect 8194 3502 8206 3554
rect 8258 3502 8270 3554
rect 10434 3502 10446 3554
rect 10498 3502 10510 3554
rect 11890 3502 11902 3554
rect 11954 3502 11966 3554
rect 6862 3490 6914 3502
rect 12014 3490 12066 3502
rect 13918 3554 13970 3566
rect 13918 3490 13970 3502
rect 14478 3554 14530 3566
rect 19182 3554 19234 3566
rect 15138 3502 15150 3554
rect 15202 3502 15214 3554
rect 14478 3490 14530 3502
rect 19182 3490 19234 3502
rect 19854 3554 19906 3566
rect 28478 3554 28530 3566
rect 22978 3502 22990 3554
rect 23042 3502 23054 3554
rect 32610 3502 32622 3554
rect 32674 3502 32686 3554
rect 35522 3502 35534 3554
rect 35586 3502 35598 3554
rect 39778 3502 39790 3554
rect 39842 3502 39854 3554
rect 19854 3490 19906 3502
rect 28478 3490 28530 3502
rect 6974 3442 7026 3454
rect 35758 3442 35810 3454
rect 31826 3390 31838 3442
rect 31890 3390 31902 3442
rect 33394 3390 33406 3442
rect 33458 3390 33470 3442
rect 6974 3378 7026 3390
rect 35758 3378 35810 3390
rect 20190 3330 20242 3342
rect 20190 3266 20242 3278
rect 28142 3330 28194 3342
rect 28142 3266 28194 3278
rect 1344 3162 48608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48608 3162
rect 1344 3076 48608 3110
rect 6862 2994 6914 3006
rect 6402 2942 6414 2994
rect 6466 2942 6478 2994
rect 6862 2930 6914 2942
rect 18286 2994 18338 3006
rect 18286 2930 18338 2942
rect 19182 2994 19234 3006
rect 30718 2994 30770 3006
rect 23762 2942 23774 2994
rect 23826 2942 23838 2994
rect 19182 2930 19234 2942
rect 30718 2930 30770 2942
rect 36766 2994 36818 3006
rect 36766 2930 36818 2942
rect 4162 2830 4174 2882
rect 4226 2830 4238 2882
rect 20290 2830 20302 2882
rect 20354 2830 20366 2882
rect 27906 2830 27918 2882
rect 27970 2830 27982 2882
rect 7534 2770 7586 2782
rect 3378 2718 3390 2770
rect 3442 2718 3454 2770
rect 7534 2706 7586 2718
rect 7758 2770 7810 2782
rect 23214 2770 23266 2782
rect 10098 2718 10110 2770
rect 10162 2718 10174 2770
rect 10546 2718 10558 2770
rect 10610 2718 10622 2770
rect 19618 2718 19630 2770
rect 19682 2718 19694 2770
rect 7758 2706 7810 2718
rect 23214 2706 23266 2718
rect 23438 2770 23490 2782
rect 23438 2706 23490 2718
rect 24222 2770 24274 2782
rect 24222 2706 24274 2718
rect 26798 2770 26850 2782
rect 27122 2718 27134 2770
rect 27186 2718 27198 2770
rect 30482 2718 30494 2770
rect 30546 2718 30558 2770
rect 26798 2706 26850 2718
rect 10322 2606 10334 2658
rect 10386 2606 10398 2658
rect 22418 2606 22430 2658
rect 22482 2606 22494 2658
rect 30034 2606 30046 2658
rect 30098 2606 30110 2658
rect 7310 2546 7362 2558
rect 10098 2494 10110 2546
rect 10162 2494 10174 2546
rect 7310 2482 7362 2494
rect 1344 2378 48608 2412
rect 1344 2326 4478 2378
rect 4530 2326 4582 2378
rect 4634 2326 4686 2378
rect 4738 2326 35198 2378
rect 35250 2326 35302 2378
rect 35354 2326 35406 2378
rect 35458 2326 48608 2378
rect 1344 2292 48608 2326
rect 6862 2098 6914 2110
rect 6862 2034 6914 2046
rect 1344 1594 48608 1628
rect 1344 1542 19838 1594
rect 19890 1542 19942 1594
rect 19994 1542 20046 1594
rect 20098 1542 48608 1594
rect 1344 1508 48608 1542
<< via1 >>
rect 19838 78374 19890 78426
rect 19942 78374 19994 78426
rect 20046 78374 20098 78426
rect 1822 77982 1874 78034
rect 3166 77982 3218 78034
rect 2942 77870 2994 77922
rect 4478 77590 4530 77642
rect 4582 77590 4634 77642
rect 4686 77590 4738 77642
rect 35198 77590 35250 77642
rect 35302 77590 35354 77642
rect 35406 77590 35458 77642
rect 2942 77310 2994 77362
rect 33294 77310 33346 77362
rect 1822 77198 1874 77250
rect 3166 77198 3218 77250
rect 8878 77198 8930 77250
rect 9886 77198 9938 77250
rect 30494 77198 30546 77250
rect 27806 77086 27858 77138
rect 31166 77086 31218 77138
rect 6190 76974 6242 77026
rect 6638 76974 6690 77026
rect 7310 76974 7362 77026
rect 7534 76974 7586 77026
rect 21534 76974 21586 77026
rect 28142 76974 28194 77026
rect 33742 76974 33794 77026
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 3054 76638 3106 76690
rect 3614 76638 3666 76690
rect 10110 76638 10162 76690
rect 30942 76638 30994 76690
rect 27918 76526 27970 76578
rect 33518 76526 33570 76578
rect 1822 76414 1874 76466
rect 3278 76414 3330 76466
rect 4958 76414 5010 76466
rect 5966 76414 6018 76466
rect 6302 76414 6354 76466
rect 7086 76414 7138 76466
rect 10446 76414 10498 76466
rect 11230 76414 11282 76466
rect 13022 76414 13074 76466
rect 13806 76414 13858 76466
rect 18510 76414 18562 76466
rect 21758 76414 21810 76466
rect 27134 76414 27186 76466
rect 30606 76414 30658 76466
rect 33966 76414 34018 76466
rect 8206 76302 8258 76354
rect 18174 76302 18226 76354
rect 19294 76302 19346 76354
rect 21422 76302 21474 76354
rect 22542 76302 22594 76354
rect 24670 76302 24722 76354
rect 26798 76302 26850 76354
rect 30046 76302 30098 76354
rect 33182 76302 33234 76354
rect 34750 76302 34802 76354
rect 36878 76302 36930 76354
rect 12574 76190 12626 76242
rect 15150 76190 15202 76242
rect 33630 76190 33682 76242
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 8318 75854 8370 75906
rect 12014 75854 12066 75906
rect 21310 75854 21362 75906
rect 27806 75854 27858 75906
rect 30494 75854 30546 75906
rect 4286 75742 4338 75794
rect 12686 75742 12738 75794
rect 22878 75742 22930 75794
rect 23550 75742 23602 75794
rect 24110 75742 24162 75794
rect 27470 75742 27522 75794
rect 28142 75742 28194 75794
rect 30158 75742 30210 75794
rect 30942 75742 30994 75794
rect 34190 75742 34242 75794
rect 34750 75742 34802 75794
rect 36430 75742 36482 75794
rect 3054 75630 3106 75682
rect 6190 75630 6242 75682
rect 6974 75630 7026 75682
rect 9886 75630 9938 75682
rect 10894 75630 10946 75682
rect 20750 75630 20802 75682
rect 21646 75630 21698 75682
rect 22430 75630 22482 75682
rect 22766 75630 22818 75682
rect 23102 75630 23154 75682
rect 23438 75630 23490 75682
rect 24222 75630 24274 75682
rect 24558 75630 24610 75682
rect 29262 75630 29314 75682
rect 29934 75630 29986 75682
rect 31278 75630 31330 75682
rect 32062 75630 32114 75682
rect 35310 75630 35362 75682
rect 4398 75518 4450 75570
rect 25342 75518 25394 75570
rect 28366 75518 28418 75570
rect 34526 75518 34578 75570
rect 34750 75518 34802 75570
rect 5854 75406 5906 75458
rect 9550 75406 9602 75458
rect 21422 75406 21474 75458
rect 36318 75406 36370 75458
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 4286 75070 4338 75122
rect 5742 75070 5794 75122
rect 8430 75070 8482 75122
rect 8990 75070 9042 75122
rect 25566 75070 25618 75122
rect 25342 74958 25394 75010
rect 33630 74958 33682 75010
rect 3054 74846 3106 74898
rect 4398 74846 4450 74898
rect 6078 74846 6130 74898
rect 6974 74846 7026 74898
rect 9662 74846 9714 74898
rect 10558 74846 10610 74898
rect 25230 74846 25282 74898
rect 25902 74846 25954 74898
rect 34974 74846 35026 74898
rect 24222 74734 24274 74786
rect 27582 74734 27634 74786
rect 30942 74734 30994 74786
rect 32510 74734 32562 74786
rect 33406 74734 33458 74786
rect 33742 74734 33794 74786
rect 34190 74734 34242 74786
rect 34638 74734 34690 74786
rect 35758 74734 35810 74786
rect 37886 74734 37938 74786
rect 11678 74622 11730 74674
rect 33966 74622 34018 74674
rect 34638 74622 34690 74674
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 12798 74286 12850 74338
rect 36990 74286 37042 74338
rect 10334 74174 10386 74226
rect 20750 74174 20802 74226
rect 21310 74174 21362 74226
rect 33518 74174 33570 74226
rect 35758 74174 35810 74226
rect 37102 74174 37154 74226
rect 10670 74062 10722 74114
rect 11454 74062 11506 74114
rect 17838 74062 17890 74114
rect 35646 74062 35698 74114
rect 17502 73950 17554 74002
rect 18622 73950 18674 74002
rect 21422 73950 21474 74002
rect 30270 73950 30322 74002
rect 30382 73950 30434 74002
rect 33406 73950 33458 74002
rect 35310 73950 35362 74002
rect 35982 73950 36034 74002
rect 29934 73838 29986 73890
rect 30606 73838 30658 73890
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 19406 73502 19458 73554
rect 31278 73390 31330 73442
rect 9662 73278 9714 73330
rect 10334 73278 10386 73330
rect 12238 73278 12290 73330
rect 13022 73278 13074 73330
rect 19630 73278 19682 73330
rect 25902 73278 25954 73330
rect 31950 73278 32002 73330
rect 8990 73166 9042 73218
rect 18958 73166 19010 73218
rect 25566 73166 25618 73218
rect 26686 73166 26738 73218
rect 28814 73166 28866 73218
rect 29150 73166 29202 73218
rect 33182 73166 33234 73218
rect 33854 73166 33906 73218
rect 11678 73054 11730 73106
rect 14254 73054 14306 73106
rect 19294 73054 19346 73106
rect 33070 73054 33122 73106
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 34862 72718 34914 72770
rect 35198 72718 35250 72770
rect 5070 72606 5122 72658
rect 33630 72606 33682 72658
rect 35198 72606 35250 72658
rect 1822 72494 1874 72546
rect 3166 72494 3218 72546
rect 6078 72494 6130 72546
rect 6974 72494 7026 72546
rect 9214 72494 9266 72546
rect 10110 72494 10162 72546
rect 30046 72494 30098 72546
rect 30382 72494 30434 72546
rect 30830 72494 30882 72546
rect 31502 72382 31554 72434
rect 2942 72270 2994 72322
rect 8318 72270 8370 72322
rect 8766 72270 8818 72322
rect 11454 72270 11506 72322
rect 11790 72270 11842 72322
rect 23550 72270 23602 72322
rect 29262 72270 29314 72322
rect 29822 72270 29874 72322
rect 30270 72270 30322 72322
rect 34302 72270 34354 72322
rect 34750 72270 34802 72322
rect 37102 72270 37154 72322
rect 37550 72270 37602 72322
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 5070 71934 5122 71986
rect 5518 71934 5570 71986
rect 33182 71934 33234 71986
rect 3838 71822 3890 71874
rect 23998 71822 24050 71874
rect 24110 71822 24162 71874
rect 2718 71710 2770 71762
rect 4062 71710 4114 71762
rect 6302 71710 6354 71762
rect 7086 71710 7138 71762
rect 9662 71710 9714 71762
rect 10334 71710 10386 71762
rect 20302 71710 20354 71762
rect 20750 71710 20802 71762
rect 23774 71710 23826 71762
rect 33406 71710 33458 71762
rect 34862 71710 34914 71762
rect 35086 71710 35138 71762
rect 36094 71710 36146 71762
rect 36542 71710 36594 71762
rect 37550 71710 37602 71762
rect 6078 71598 6130 71650
rect 8654 71598 8706 71650
rect 8990 71598 9042 71650
rect 21422 71598 21474 71650
rect 23550 71571 23602 71623
rect 24558 71598 24610 71650
rect 25566 71598 25618 71650
rect 26126 71598 26178 71650
rect 32510 71598 32562 71650
rect 33070 71598 33122 71650
rect 33854 71598 33906 71650
rect 34302 71598 34354 71650
rect 37998 71598 38050 71650
rect 11678 71486 11730 71538
rect 24446 71486 24498 71538
rect 25678 71486 25730 71538
rect 36206 71486 36258 71538
rect 37214 71486 37266 71538
rect 37550 71486 37602 71538
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 21646 71150 21698 71202
rect 26350 71150 26402 71202
rect 36094 71150 36146 71202
rect 3502 71038 3554 71090
rect 10334 71038 10386 71090
rect 20750 71038 20802 71090
rect 21422 71038 21474 71090
rect 23550 71038 23602 71090
rect 25678 71038 25730 71090
rect 26014 71038 26066 71090
rect 29486 71038 29538 71090
rect 32958 71038 33010 71090
rect 33854 71038 33906 71090
rect 34862 71038 34914 71090
rect 37774 71038 37826 71090
rect 39902 71038 39954 71090
rect 2382 70926 2434 70978
rect 4174 70926 4226 70978
rect 4622 70926 4674 70978
rect 6414 70926 6466 70978
rect 7198 70926 7250 70978
rect 10670 70926 10722 70978
rect 11678 70926 11730 70978
rect 22878 70926 22930 70978
rect 32846 70926 32898 70978
rect 33630 70926 33682 70978
rect 34974 70926 35026 70978
rect 35982 70926 36034 70978
rect 36430 70926 36482 70978
rect 36990 70926 37042 70978
rect 3614 70814 3666 70866
rect 5630 70814 5682 70866
rect 5966 70814 6018 70866
rect 33294 70814 33346 70866
rect 8766 70702 8818 70754
rect 13022 70702 13074 70754
rect 21422 70702 21474 70754
rect 22430 70702 22482 70754
rect 26126 70702 26178 70754
rect 26910 70702 26962 70754
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 4398 70366 4450 70418
rect 6302 70366 6354 70418
rect 16830 70366 16882 70418
rect 34078 70366 34130 70418
rect 38334 70366 38386 70418
rect 38782 70366 38834 70418
rect 4958 70254 5010 70306
rect 34414 70254 34466 70306
rect 34638 70254 34690 70306
rect 38894 70254 38946 70306
rect 5630 70142 5682 70194
rect 6750 70142 6802 70194
rect 7534 70142 7586 70194
rect 9886 70142 9938 70194
rect 10782 70142 10834 70194
rect 12350 70142 12402 70194
rect 13358 70142 13410 70194
rect 14702 70142 14754 70194
rect 17726 70142 17778 70194
rect 23102 70142 23154 70194
rect 23438 70142 23490 70194
rect 23998 70142 24050 70194
rect 25454 70142 25506 70194
rect 25790 70142 25842 70194
rect 26574 70142 26626 70194
rect 26910 70142 26962 70194
rect 28030 70142 28082 70194
rect 29038 70142 29090 70194
rect 29934 70142 29986 70194
rect 31166 70142 31218 70194
rect 35086 70142 35138 70194
rect 38446 70142 38498 70194
rect 3838 70030 3890 70082
rect 9102 70030 9154 70082
rect 18398 70030 18450 70082
rect 20526 70030 20578 70082
rect 20862 70030 20914 70082
rect 23326 70030 23378 70082
rect 24446 70030 24498 70082
rect 26014 70030 26066 70082
rect 28366 70030 28418 70082
rect 29262 70030 29314 70082
rect 29710 70030 29762 70082
rect 30718 70030 30770 70082
rect 31614 70030 31666 70082
rect 33630 70030 33682 70082
rect 34750 70030 34802 70082
rect 35870 70030 35922 70082
rect 37998 70030 38050 70082
rect 4062 69918 4114 69970
rect 11902 69918 11954 69970
rect 20974 69918 21026 69970
rect 24222 69918 24274 69970
rect 26798 69918 26850 69970
rect 28702 69918 28754 69970
rect 30270 69918 30322 69970
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 5630 69582 5682 69634
rect 35982 69582 36034 69634
rect 4622 69470 4674 69522
rect 5742 69470 5794 69522
rect 6190 69470 6242 69522
rect 6638 69470 6690 69522
rect 13022 69470 13074 69522
rect 23438 69470 23490 69522
rect 25678 69470 25730 69522
rect 27806 69470 27858 69522
rect 32510 69470 32562 69522
rect 34974 69470 35026 69522
rect 10670 69358 10722 69410
rect 11454 69358 11506 69410
rect 18734 69358 18786 69410
rect 21422 69358 21474 69410
rect 21870 69358 21922 69410
rect 22542 69358 22594 69410
rect 23102 69358 23154 69410
rect 25006 69358 25058 69410
rect 28590 69358 28642 69410
rect 29598 69358 29650 69410
rect 34862 69358 34914 69410
rect 35646 69358 35698 69410
rect 35870 69358 35922 69410
rect 37102 69358 37154 69410
rect 18510 69246 18562 69298
rect 19070 69246 19122 69298
rect 22318 69246 22370 69298
rect 30382 69246 30434 69298
rect 9438 69134 9490 69186
rect 10334 69134 10386 69186
rect 18958 69134 19010 69186
rect 24110 69134 24162 69186
rect 24558 69134 24610 69186
rect 28254 69134 28306 69186
rect 32958 69134 33010 69186
rect 34190 69134 34242 69186
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 12014 68798 12066 68850
rect 19742 68798 19794 68850
rect 23774 68798 23826 68850
rect 25342 68798 25394 68850
rect 30494 68798 30546 68850
rect 35534 68798 35586 68850
rect 2494 68686 2546 68738
rect 2942 68686 2994 68738
rect 3390 68686 3442 68738
rect 24670 68686 24722 68738
rect 28030 68686 28082 68738
rect 33070 68686 33122 68738
rect 20302 68574 20354 68626
rect 20862 68574 20914 68626
rect 21422 68574 21474 68626
rect 21982 68574 22034 68626
rect 22430 68574 22482 68626
rect 23102 68574 23154 68626
rect 27358 68574 27410 68626
rect 30718 68574 30770 68626
rect 33406 68574 33458 68626
rect 19630 68462 19682 68514
rect 24222 68462 24274 68514
rect 25790 68462 25842 68514
rect 26910 68462 26962 68514
rect 30158 68462 30210 68514
rect 35646 68462 35698 68514
rect 21870 68350 21922 68402
rect 24222 68350 24274 68402
rect 24558 68350 24610 68402
rect 24782 68350 24834 68402
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 3838 68014 3890 68066
rect 5742 68014 5794 68066
rect 10782 68014 10834 68066
rect 20302 68014 20354 68066
rect 6414 67902 6466 67954
rect 8318 67902 8370 67954
rect 16382 67902 16434 67954
rect 19630 67902 19682 67954
rect 23326 67902 23378 67954
rect 32622 67902 32674 67954
rect 34750 67902 34802 67954
rect 2942 67790 2994 67842
rect 3166 67790 3218 67842
rect 3502 67790 3554 67842
rect 6078 67790 6130 67842
rect 7646 67790 7698 67842
rect 8766 67790 8818 67842
rect 9662 67790 9714 67842
rect 16830 67790 16882 67842
rect 31838 67790 31890 67842
rect 2270 67678 2322 67730
rect 2606 67678 2658 67730
rect 17502 67678 17554 67730
rect 20414 67678 20466 67730
rect 21422 67678 21474 67730
rect 1934 67566 1986 67618
rect 3726 67566 3778 67618
rect 7198 67566 7250 67618
rect 22878 67566 22930 67618
rect 31502 67566 31554 67618
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 3726 67230 3778 67282
rect 17950 67230 18002 67282
rect 3614 67118 3666 67170
rect 6526 67118 6578 67170
rect 33630 67118 33682 67170
rect 35086 67118 35138 67170
rect 37214 67118 37266 67170
rect 39230 67118 39282 67170
rect 1822 67006 1874 67058
rect 3054 67006 3106 67058
rect 4062 67006 4114 67058
rect 5518 67006 5570 67058
rect 6862 67006 6914 67058
rect 7310 67006 7362 67058
rect 7534 67006 7586 67058
rect 10782 67006 10834 67058
rect 11678 67006 11730 67058
rect 18286 67006 18338 67058
rect 27470 67006 27522 67058
rect 35310 67006 35362 67058
rect 36990 67006 37042 67058
rect 38558 67006 38610 67058
rect 2942 66894 2994 66946
rect 4846 66894 4898 66946
rect 6078 66894 6130 66946
rect 8766 66894 8818 66946
rect 25342 66894 25394 66946
rect 27246 66894 27298 66946
rect 28030 66894 28082 66946
rect 28590 66894 28642 66946
rect 32622 66894 32674 66946
rect 33070 66894 33122 66946
rect 34190 66894 34242 66946
rect 34526 66894 34578 66946
rect 6974 66782 7026 66834
rect 9662 66782 9714 66834
rect 27806 66782 27858 66834
rect 33294 66782 33346 66834
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 2606 66446 2658 66498
rect 7198 66446 7250 66498
rect 7870 66446 7922 66498
rect 33630 66446 33682 66498
rect 34190 66446 34242 66498
rect 2942 66334 2994 66386
rect 3614 66334 3666 66386
rect 4286 66334 4338 66386
rect 4734 66334 4786 66386
rect 6750 66334 6802 66386
rect 9438 66334 9490 66386
rect 14702 66334 14754 66386
rect 25230 66334 25282 66386
rect 28478 66334 28530 66386
rect 33630 66334 33682 66386
rect 39902 66334 39954 66386
rect 2718 66222 2770 66274
rect 6638 66222 6690 66274
rect 7646 66222 7698 66274
rect 11118 66222 11170 66274
rect 12462 66222 12514 66274
rect 13470 66222 13522 66274
rect 21758 66222 21810 66274
rect 22318 66222 22370 66274
rect 25678 66222 25730 66274
rect 36206 66222 36258 66274
rect 36990 66222 37042 66274
rect 3502 66110 3554 66162
rect 8206 66110 8258 66162
rect 8542 66110 8594 66162
rect 14814 66110 14866 66162
rect 23102 66110 23154 66162
rect 26350 66110 26402 66162
rect 36430 66110 36482 66162
rect 37774 66110 37826 66162
rect 3726 65998 3778 66050
rect 4174 65998 4226 66050
rect 10222 65998 10274 66050
rect 11342 65998 11394 66050
rect 21422 65998 21474 66050
rect 21870 65998 21922 66050
rect 34078 65998 34130 66050
rect 35758 65998 35810 66050
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 7310 65662 7362 65714
rect 14366 65662 14418 65714
rect 26462 65662 26514 65714
rect 38110 65662 38162 65714
rect 25342 65550 25394 65602
rect 30494 65550 30546 65602
rect 34750 65550 34802 65602
rect 37438 65550 37490 65602
rect 2718 65438 2770 65490
rect 7758 65438 7810 65490
rect 9550 65438 9602 65490
rect 10782 65438 10834 65490
rect 12126 65438 12178 65490
rect 13134 65438 13186 65490
rect 14478 65438 14530 65490
rect 17950 65438 18002 65490
rect 21198 65438 21250 65490
rect 26686 65438 26738 65490
rect 30830 65438 30882 65490
rect 32062 65438 32114 65490
rect 33742 65438 33794 65490
rect 34190 65438 34242 65490
rect 35982 65438 36034 65490
rect 38334 65438 38386 65490
rect 39230 65438 39282 65490
rect 4062 65326 4114 65378
rect 8206 65326 8258 65378
rect 8990 65326 9042 65378
rect 12014 65326 12066 65378
rect 17614 65326 17666 65378
rect 18734 65326 18786 65378
rect 20862 65326 20914 65378
rect 21982 65326 22034 65378
rect 24110 65326 24162 65378
rect 24446 65326 24498 65378
rect 32510 65326 32562 65378
rect 39006 65326 39058 65378
rect 39678 65326 39730 65378
rect 2830 65214 2882 65266
rect 10110 65214 10162 65266
rect 24558 65214 24610 65266
rect 25454 65214 25506 65266
rect 33182 65214 33234 65266
rect 33518 65214 33570 65266
rect 38670 65214 38722 65266
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 21422 64878 21474 64930
rect 22094 64878 22146 64930
rect 36990 64878 37042 64930
rect 23550 64766 23602 64818
rect 25678 64766 25730 64818
rect 30158 64766 30210 64818
rect 32286 64766 32338 64818
rect 35758 64766 35810 64818
rect 37998 64766 38050 64818
rect 9438 64654 9490 64706
rect 10782 64654 10834 64706
rect 28590 64654 28642 64706
rect 29374 64654 29426 64706
rect 32846 64654 32898 64706
rect 37326 64654 37378 64706
rect 37550 64654 37602 64706
rect 40798 64654 40850 64706
rect 18510 64542 18562 64594
rect 21758 64542 21810 64594
rect 22430 64542 22482 64594
rect 23326 64542 23378 64594
rect 27806 64542 27858 64594
rect 33630 64542 33682 64594
rect 40126 64542 40178 64594
rect 10670 64430 10722 64482
rect 18622 64430 18674 64482
rect 20750 64430 20802 64482
rect 21534 64430 21586 64482
rect 22206 64430 22258 64482
rect 22878 64430 22930 64482
rect 23550 64430 23602 64482
rect 24110 64430 24162 64482
rect 25342 64430 25394 64482
rect 36430 64430 36482 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 5294 64094 5346 64146
rect 21982 64094 22034 64146
rect 27918 64094 27970 64146
rect 30606 64094 30658 64146
rect 30942 64094 30994 64146
rect 33854 64094 33906 64146
rect 34526 64094 34578 64146
rect 39678 64094 39730 64146
rect 22878 63982 22930 64034
rect 33518 63982 33570 64034
rect 35198 63982 35250 64034
rect 10782 63870 10834 63922
rect 12126 63870 12178 63922
rect 16830 63870 16882 63922
rect 17390 63870 17442 63922
rect 22766 63870 22818 63922
rect 28254 63870 28306 63922
rect 28702 63870 28754 63922
rect 31278 63870 31330 63922
rect 31502 63870 31554 63922
rect 32510 63870 32562 63922
rect 33182 63870 33234 63922
rect 35310 63870 35362 63922
rect 37102 63870 37154 63922
rect 37774 63870 37826 63922
rect 38558 63870 38610 63922
rect 11902 63758 11954 63810
rect 18174 63758 18226 63810
rect 20302 63758 20354 63810
rect 37662 63758 37714 63810
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 4062 63310 4114 63362
rect 4958 63310 5010 63362
rect 7758 63310 7810 63362
rect 19182 63310 19234 63362
rect 30382 63310 30434 63362
rect 4062 63198 4114 63250
rect 4510 63198 4562 63250
rect 4958 63198 5010 63250
rect 16382 63198 16434 63250
rect 18510 63198 18562 63250
rect 18958 63198 19010 63250
rect 30606 63198 30658 63250
rect 31054 63198 31106 63250
rect 31950 63198 32002 63250
rect 37550 63198 37602 63250
rect 37998 63198 38050 63250
rect 39230 63198 39282 63250
rect 5630 63086 5682 63138
rect 6414 63086 6466 63138
rect 8318 63086 8370 63138
rect 13470 63086 13522 63138
rect 14814 63086 14866 63138
rect 15598 63086 15650 63138
rect 18846 63086 18898 63138
rect 19630 63086 19682 63138
rect 32398 63086 32450 63138
rect 33966 63086 34018 63138
rect 36430 63086 36482 63138
rect 37326 63086 37378 63138
rect 38558 63086 38610 63138
rect 2718 62974 2770 63026
rect 9550 62974 9602 63026
rect 32958 62974 33010 63026
rect 35646 62974 35698 63026
rect 38782 62974 38834 63026
rect 2382 62862 2434 62914
rect 9438 62862 9490 62914
rect 14702 62862 14754 62914
rect 30046 62862 30098 62914
rect 34862 62862 34914 62914
rect 36990 62862 37042 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 3054 62526 3106 62578
rect 3726 62526 3778 62578
rect 7422 62526 7474 62578
rect 14254 62526 14306 62578
rect 35982 62526 36034 62578
rect 17726 62414 17778 62466
rect 17950 62414 18002 62466
rect 18510 62414 18562 62466
rect 18958 62414 19010 62466
rect 19630 62414 19682 62466
rect 23326 62414 23378 62466
rect 23662 62414 23714 62466
rect 23774 62414 23826 62466
rect 1934 62302 1986 62354
rect 3278 62302 3330 62354
rect 4286 62302 4338 62354
rect 4622 62302 4674 62354
rect 5182 62302 5234 62354
rect 6078 62302 6130 62354
rect 10334 62302 10386 62354
rect 11678 62302 11730 62354
rect 13022 62302 13074 62354
rect 14478 62302 14530 62354
rect 28366 62302 28418 62354
rect 31726 62302 31778 62354
rect 39118 62302 39170 62354
rect 11454 62190 11506 62242
rect 18062 62190 18114 62242
rect 29150 62190 29202 62242
rect 31278 62190 31330 62242
rect 36318 62190 36370 62242
rect 38446 62190 38498 62242
rect 4062 62078 4114 62130
rect 4734 62078 4786 62130
rect 19742 62078 19794 62130
rect 23774 62078 23826 62130
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 4286 61742 4338 61794
rect 32958 61742 33010 61794
rect 3054 61630 3106 61682
rect 5742 61630 5794 61682
rect 14702 61630 14754 61682
rect 20750 61630 20802 61682
rect 21646 61630 21698 61682
rect 23774 61630 23826 61682
rect 25902 61630 25954 61682
rect 26238 61630 26290 61682
rect 33182 61630 33234 61682
rect 33630 61630 33682 61682
rect 39566 61630 39618 61682
rect 42814 61630 42866 61682
rect 1934 61518 1986 61570
rect 3278 61518 3330 61570
rect 3950 61518 4002 61570
rect 4622 61518 4674 61570
rect 7646 61518 7698 61570
rect 9438 61518 9490 61570
rect 13470 61518 13522 61570
rect 14814 61518 14866 61570
rect 17838 61518 17890 61570
rect 22990 61518 23042 61570
rect 30046 61518 30098 61570
rect 37102 61518 37154 61570
rect 39902 61518 39954 61570
rect 5630 61406 5682 61458
rect 5854 61406 5906 61458
rect 8878 61406 8930 61458
rect 10782 61406 10834 61458
rect 18622 61406 18674 61458
rect 29710 61406 29762 61458
rect 40686 61406 40738 61458
rect 8766 61294 8818 61346
rect 10670 61294 10722 61346
rect 17502 61294 17554 61346
rect 21758 61294 21810 61346
rect 22654 61294 22706 61346
rect 26350 61294 26402 61346
rect 32622 61294 32674 61346
rect 37438 61294 37490 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 19854 60958 19906 61010
rect 20638 60958 20690 61010
rect 24558 60958 24610 61010
rect 16494 60846 16546 60898
rect 19966 60846 20018 60898
rect 32174 60846 32226 60898
rect 32510 60846 32562 60898
rect 40238 60846 40290 60898
rect 7534 60734 7586 60786
rect 8766 60734 8818 60786
rect 15374 60734 15426 60786
rect 20974 60734 21026 60786
rect 25230 60734 25282 60786
rect 33182 60734 33234 60786
rect 40910 60734 40962 60786
rect 3726 60622 3778 60674
rect 3838 60622 3890 60674
rect 5070 60622 5122 60674
rect 8654 60622 8706 60674
rect 15150 60622 15202 60674
rect 19406 60622 19458 60674
rect 21758 60622 21810 60674
rect 23886 60622 23938 60674
rect 24670 60622 24722 60674
rect 26014 60622 26066 60674
rect 28142 60622 28194 60674
rect 33854 60622 33906 60674
rect 35982 60622 36034 60674
rect 39678 60622 39730 60674
rect 40350 60622 40402 60674
rect 41694 60622 41746 60674
rect 43822 60622 43874 60674
rect 19742 60510 19794 60562
rect 24334 60510 24386 60562
rect 40014 60510 40066 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 7646 60174 7698 60226
rect 23774 60174 23826 60226
rect 26462 60174 26514 60226
rect 41246 60174 41298 60226
rect 17838 60062 17890 60114
rect 18286 60062 18338 60114
rect 23886 60062 23938 60114
rect 24894 60062 24946 60114
rect 30718 60062 30770 60114
rect 40126 60062 40178 60114
rect 42366 60062 42418 60114
rect 42814 60062 42866 60114
rect 15038 59950 15090 60002
rect 21982 59950 22034 60002
rect 24334 59950 24386 60002
rect 26798 59950 26850 60002
rect 27582 59950 27634 60002
rect 31278 59950 31330 60002
rect 41246 59950 41298 60002
rect 7086 59838 7138 59890
rect 7534 59838 7586 59890
rect 15710 59838 15762 59890
rect 21646 59838 21698 59890
rect 27022 59838 27074 59890
rect 31838 59838 31890 59890
rect 40910 59838 40962 59890
rect 6750 59726 6802 59778
rect 21758 59726 21810 59778
rect 22318 59726 22370 59778
rect 26126 59726 26178 59778
rect 27358 59726 27410 59778
rect 32734 59726 32786 59778
rect 40574 59726 40626 59778
rect 42254 59726 42306 59778
rect 42702 59726 42754 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 5854 59390 5906 59442
rect 6750 59390 6802 59442
rect 16942 59390 16994 59442
rect 18062 59390 18114 59442
rect 26014 59390 26066 59442
rect 33406 59390 33458 59442
rect 2382 59278 2434 59330
rect 12014 59278 12066 59330
rect 15598 59278 15650 59330
rect 16382 59278 16434 59330
rect 17390 59278 17442 59330
rect 27134 59278 27186 59330
rect 30606 59278 30658 59330
rect 6190 59166 6242 59218
rect 10670 59166 10722 59218
rect 12798 59166 12850 59218
rect 14254 59166 14306 59218
rect 17614 59166 17666 59218
rect 18398 59166 18450 59218
rect 21982 59166 22034 59218
rect 22430 59166 22482 59218
rect 22878 59166 22930 59218
rect 23438 59166 23490 59218
rect 26350 59166 26402 59218
rect 33070 59166 33122 59218
rect 34638 59166 34690 59218
rect 35086 59166 35138 59218
rect 4174 59054 4226 59106
rect 4622 59054 4674 59106
rect 5406 59054 5458 59106
rect 11902 59054 11954 59106
rect 14030 59054 14082 59106
rect 18846 59054 18898 59106
rect 19630 59054 19682 59106
rect 22094 59054 22146 59106
rect 22766 59054 22818 59106
rect 24334 59054 24386 59106
rect 24782 59054 24834 59106
rect 25454 59054 25506 59106
rect 29262 59054 29314 59106
rect 31054 59054 31106 59106
rect 35758 59054 35810 59106
rect 37886 59054 37938 59106
rect 2270 58942 2322 58994
rect 2606 58942 2658 58994
rect 6414 58942 6466 58994
rect 30046 58942 30098 58994
rect 30382 58942 30434 58994
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 24670 58606 24722 58658
rect 27470 58606 27522 58658
rect 29150 58606 29202 58658
rect 5070 58494 5122 58546
rect 6638 58494 6690 58546
rect 16270 58494 16322 58546
rect 18398 58494 18450 58546
rect 23774 58494 23826 58546
rect 24782 58494 24834 58546
rect 25678 58494 25730 58546
rect 31614 58494 31666 58546
rect 33742 58494 33794 58546
rect 40686 58494 40738 58546
rect 41134 58494 41186 58546
rect 1822 58382 1874 58434
rect 2718 58382 2770 58434
rect 4062 58382 4114 58434
rect 4510 58382 4562 58434
rect 6302 58382 6354 58434
rect 6526 58382 6578 58434
rect 10670 58382 10722 58434
rect 12014 58382 12066 58434
rect 13470 58382 13522 58434
rect 14814 58382 14866 58434
rect 15598 58382 15650 58434
rect 23550 58382 23602 58434
rect 24222 58382 24274 58434
rect 24558 58382 24610 58434
rect 26126 58382 26178 58434
rect 27134 58382 27186 58434
rect 27806 58382 27858 58434
rect 29486 58382 29538 58434
rect 29710 58382 29762 58434
rect 30942 58382 30994 58434
rect 34302 58382 34354 58434
rect 35646 58382 35698 58434
rect 37550 58382 37602 58434
rect 37886 58382 37938 58434
rect 18846 58270 18898 58322
rect 19294 58270 19346 58322
rect 19854 58270 19906 58322
rect 20302 58270 20354 58322
rect 28030 58270 28082 58322
rect 35870 58270 35922 58322
rect 38558 58270 38610 58322
rect 41022 58270 41074 58322
rect 4286 58158 4338 58210
rect 7198 58158 7250 58210
rect 11902 58158 11954 58210
rect 14702 58158 14754 58210
rect 19070 58158 19122 58210
rect 19406 58158 19458 58210
rect 28478 58158 28530 58210
rect 30158 58158 30210 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 2270 57822 2322 57874
rect 5294 57822 5346 57874
rect 6414 57822 6466 57874
rect 14030 57822 14082 57874
rect 17390 57822 17442 57874
rect 32286 57822 32338 57874
rect 32398 57822 32450 57874
rect 34078 57822 34130 57874
rect 35646 57822 35698 57874
rect 36094 57822 36146 57874
rect 2606 57710 2658 57762
rect 10894 57710 10946 57762
rect 17950 57710 18002 57762
rect 18734 57710 18786 57762
rect 20862 57710 20914 57762
rect 23326 57710 23378 57762
rect 31838 57710 31890 57762
rect 38558 57710 38610 57762
rect 38782 57710 38834 57762
rect 1934 57598 1986 57650
rect 3278 57598 3330 57650
rect 4174 57598 4226 57650
rect 5406 57598 5458 57650
rect 7982 57598 8034 57650
rect 8990 57598 9042 57650
rect 12126 57598 12178 57650
rect 12798 57598 12850 57650
rect 14254 57598 14306 57650
rect 18286 57598 18338 57650
rect 18510 57598 18562 57650
rect 18958 57598 19010 57650
rect 19966 57598 20018 57650
rect 20302 57598 20354 57650
rect 22430 57598 22482 57650
rect 22766 57598 22818 57650
rect 25454 57598 25506 57650
rect 25678 57598 25730 57650
rect 26798 57598 26850 57650
rect 27918 57598 27970 57650
rect 31502 57598 31554 57650
rect 32062 57598 32114 57650
rect 35310 57598 35362 57650
rect 2158 57486 2210 57538
rect 3054 57486 3106 57538
rect 11006 57486 11058 57538
rect 18846 57486 18898 57538
rect 22542 57486 22594 57538
rect 25342 57486 25394 57538
rect 26910 57486 26962 57538
rect 28590 57486 28642 57538
rect 30718 57486 30770 57538
rect 32174 57486 32226 57538
rect 33182 57486 33234 57538
rect 33742 57486 33794 57538
rect 35086 57486 35138 57538
rect 38110 57486 38162 57538
rect 38446 57486 38498 57538
rect 6862 57374 6914 57426
rect 17726 57374 17778 57426
rect 20078 57374 20130 57426
rect 26350 57374 26402 57426
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 3166 57038 3218 57090
rect 3502 57038 3554 57090
rect 5070 57038 5122 57090
rect 9550 57038 9602 57090
rect 12126 57038 12178 57090
rect 19854 57038 19906 57090
rect 25454 57038 25506 57090
rect 32062 57038 32114 57090
rect 4958 56926 5010 56978
rect 6638 56926 6690 56978
rect 25790 56926 25842 56978
rect 26238 56926 26290 56978
rect 30718 56926 30770 56978
rect 34302 56926 34354 56978
rect 34526 56926 34578 56978
rect 34974 56926 35026 56978
rect 41358 56926 41410 56978
rect 2158 56814 2210 56866
rect 2606 56814 2658 56866
rect 2942 56814 2994 56866
rect 5854 56814 5906 56866
rect 6526 56814 6578 56866
rect 7086 56814 7138 56866
rect 7534 56814 7586 56866
rect 8318 56814 8370 56866
rect 9998 56814 10050 56866
rect 10782 56814 10834 56866
rect 19406 56814 19458 56866
rect 19742 56814 19794 56866
rect 20302 56814 20354 56866
rect 22990 56814 23042 56866
rect 23326 56814 23378 56866
rect 31054 56814 31106 56866
rect 44158 56814 44210 56866
rect 5966 56702 6018 56754
rect 21310 56702 21362 56754
rect 23886 56702 23938 56754
rect 25678 56702 25730 56754
rect 29822 56702 29874 56754
rect 30158 56702 30210 56754
rect 38446 56702 38498 56754
rect 43486 56702 43538 56754
rect 4286 56590 4338 56642
rect 4734 56590 4786 56642
rect 18174 56590 18226 56642
rect 18734 56590 18786 56642
rect 22318 56590 22370 56642
rect 33966 56590 34018 56642
rect 38558 56590 38610 56642
rect 41022 56590 41074 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 7982 56254 8034 56306
rect 9662 56254 9714 56306
rect 38670 56254 38722 56306
rect 41918 56254 41970 56306
rect 42142 56254 42194 56306
rect 26014 56142 26066 56194
rect 33406 56142 33458 56194
rect 33742 56142 33794 56194
rect 6302 56030 6354 56082
rect 21870 56030 21922 56082
rect 22318 56030 22370 56082
rect 22766 56030 22818 56082
rect 23438 56030 23490 56082
rect 25230 56030 25282 56082
rect 35422 56030 35474 56082
rect 41806 56030 41858 56082
rect 42478 56030 42530 56082
rect 3166 55918 3218 55970
rect 20974 55918 21026 55970
rect 23102 55918 23154 55970
rect 24782 55918 24834 55970
rect 28142 55918 28194 55970
rect 36094 55918 36146 55970
rect 38222 55918 38274 55970
rect 41246 55918 41298 55970
rect 20974 55806 21026 55858
rect 21422 55806 21474 55858
rect 23326 55806 23378 55858
rect 41246 55806 41298 55858
rect 41582 55806 41634 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 2718 55470 2770 55522
rect 3278 55470 3330 55522
rect 17054 55470 17106 55522
rect 18062 55358 18114 55410
rect 21310 55358 21362 55410
rect 22430 55358 22482 55410
rect 33518 55358 33570 55410
rect 35646 55358 35698 55410
rect 41246 55358 41298 55410
rect 41918 55358 41970 55410
rect 42366 55358 42418 55410
rect 42814 55358 42866 55410
rect 1934 55246 1986 55298
rect 3278 55246 3330 55298
rect 4622 55246 4674 55298
rect 6638 55246 6690 55298
rect 7982 55246 8034 55298
rect 8878 55246 8930 55298
rect 17838 55246 17890 55298
rect 19518 55246 19570 55298
rect 20190 55246 20242 55298
rect 20638 55246 20690 55298
rect 24334 55246 24386 55298
rect 24782 55246 24834 55298
rect 32846 55246 32898 55298
rect 38446 55246 38498 55298
rect 3726 55134 3778 55186
rect 6190 55134 6242 55186
rect 16942 55134 16994 55186
rect 20750 55134 20802 55186
rect 21422 55134 21474 55186
rect 21646 55134 21698 55186
rect 22766 55134 22818 55186
rect 25342 55134 25394 55186
rect 39118 55134 39170 55186
rect 41582 55134 41634 55186
rect 41806 55134 41858 55186
rect 2382 55022 2434 55074
rect 2942 55022 2994 55074
rect 4174 55022 4226 55074
rect 5182 55022 5234 55074
rect 5742 55022 5794 55074
rect 5966 55022 6018 55074
rect 6078 55022 6130 55074
rect 17502 55022 17554 55074
rect 18510 55022 18562 55074
rect 24222 55022 24274 55074
rect 32398 55022 32450 55074
rect 42254 55022 42306 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 13134 54686 13186 54738
rect 19518 54686 19570 54738
rect 19630 54686 19682 54738
rect 29710 54686 29762 54738
rect 35198 54686 35250 54738
rect 41022 54686 41074 54738
rect 17390 54574 17442 54626
rect 21310 54574 21362 54626
rect 24110 54574 24162 54626
rect 25342 54574 25394 54626
rect 28030 54574 28082 54626
rect 29262 54574 29314 54626
rect 30494 54574 30546 54626
rect 38334 54574 38386 54626
rect 38894 54574 38946 54626
rect 42142 54574 42194 54626
rect 1822 54462 1874 54514
rect 3166 54462 3218 54514
rect 3614 54462 3666 54514
rect 13806 54462 13858 54514
rect 17614 54462 17666 54514
rect 19854 54462 19906 54514
rect 20078 54462 20130 54514
rect 20526 54462 20578 54514
rect 25230 54462 25282 54514
rect 25566 54462 25618 54514
rect 25902 54462 25954 54514
rect 28926 54462 28978 54514
rect 30158 54462 30210 54514
rect 34862 54462 34914 54514
rect 41358 54462 41410 54514
rect 2494 54350 2546 54402
rect 6302 54350 6354 54402
rect 14478 54350 14530 54402
rect 16606 54350 16658 54402
rect 18174 54350 18226 54402
rect 18846 54350 18898 54402
rect 19294 54350 19346 54402
rect 23438 54350 23490 54402
rect 23998 54350 24050 54402
rect 24558 54350 24610 54402
rect 27806 54350 27858 54402
rect 28590 54350 28642 54402
rect 33294 54350 33346 54402
rect 33742 54350 33794 54402
rect 38670 54350 38722 54402
rect 39006 54350 39058 54402
rect 44270 54350 44322 54402
rect 28254 54238 28306 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 7198 53902 7250 53954
rect 29710 53902 29762 53954
rect 34190 53902 34242 53954
rect 40910 53902 40962 53954
rect 2606 53790 2658 53842
rect 2942 53790 2994 53842
rect 3726 53790 3778 53842
rect 6638 53790 6690 53842
rect 7646 53790 7698 53842
rect 9438 53790 9490 53842
rect 17054 53790 17106 53842
rect 19182 53790 19234 53842
rect 23438 53790 23490 53842
rect 30942 53790 30994 53842
rect 33070 53790 33122 53842
rect 33854 53790 33906 53842
rect 41134 53790 41186 53842
rect 42142 53790 42194 53842
rect 44046 53790 44098 53842
rect 1934 53678 1986 53730
rect 3166 53678 3218 53730
rect 3614 53678 3666 53730
rect 4286 53678 4338 53730
rect 4510 53678 4562 53730
rect 6974 53678 7026 53730
rect 12686 53678 12738 53730
rect 14478 53678 14530 53730
rect 15934 53678 15986 53730
rect 16382 53678 16434 53730
rect 23326 53678 23378 53730
rect 24110 53678 24162 53730
rect 26014 53678 26066 53730
rect 26350 53678 26402 53730
rect 28590 53678 28642 53730
rect 29374 53678 29426 53730
rect 30158 53678 30210 53730
rect 33630 53678 33682 53730
rect 41022 53678 41074 53730
rect 41694 53678 41746 53730
rect 42254 53678 42306 53730
rect 5630 53566 5682 53618
rect 6526 53566 6578 53618
rect 7982 53566 8034 53618
rect 8542 53566 8594 53618
rect 13582 53566 13634 53618
rect 15038 53566 15090 53618
rect 15374 53566 15426 53618
rect 23214 53566 23266 53618
rect 24446 53566 24498 53618
rect 26910 53566 26962 53618
rect 29150 53566 29202 53618
rect 35982 53566 36034 53618
rect 38558 53566 38610 53618
rect 2046 53454 2098 53506
rect 2494 53454 2546 53506
rect 2718 53454 2770 53506
rect 3838 53454 3890 53506
rect 4846 53454 4898 53506
rect 4958 53454 5010 53506
rect 5070 53454 5122 53506
rect 5742 53454 5794 53506
rect 5966 53454 6018 53506
rect 6750 53454 6802 53506
rect 7534 53454 7586 53506
rect 7758 53454 7810 53506
rect 8430 53454 8482 53506
rect 8990 53454 9042 53506
rect 12126 53454 12178 53506
rect 12350 53454 12402 53506
rect 12574 53454 12626 53506
rect 20302 53454 20354 53506
rect 25342 53454 25394 53506
rect 34638 53454 34690 53506
rect 36318 53454 36370 53506
rect 38670 53454 38722 53506
rect 40238 53454 40290 53506
rect 43150 53454 43202 53506
rect 43934 53454 43986 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 3278 53118 3330 53170
rect 4174 53118 4226 53170
rect 5182 53118 5234 53170
rect 8430 53118 8482 53170
rect 8878 53118 8930 53170
rect 22766 53118 22818 53170
rect 23998 53118 24050 53170
rect 24110 53118 24162 53170
rect 32398 53118 32450 53170
rect 38894 53118 38946 53170
rect 42366 53118 42418 53170
rect 42814 53118 42866 53170
rect 3726 53006 3778 53058
rect 4286 53006 4338 53058
rect 4510 53006 4562 53058
rect 6190 53006 6242 53058
rect 11902 53006 11954 53058
rect 20638 53006 20690 53058
rect 23214 53006 23266 53058
rect 26014 53006 26066 53058
rect 29262 53006 29314 53058
rect 36318 53006 36370 53058
rect 2942 52894 2994 52946
rect 3502 52894 3554 52946
rect 4062 52894 4114 52946
rect 5406 52894 5458 52946
rect 5518 52894 5570 52946
rect 6750 52894 6802 52946
rect 7534 52894 7586 52946
rect 11118 52894 11170 52946
rect 19406 52894 19458 52946
rect 19966 52894 20018 52946
rect 20302 52894 20354 52946
rect 23438 52894 23490 52946
rect 23774 52894 23826 52946
rect 25230 52894 25282 52946
rect 28590 52894 28642 52946
rect 33630 52894 33682 52946
rect 35534 52894 35586 52946
rect 43150 52894 43202 52946
rect 2270 52782 2322 52834
rect 2606 52782 2658 52834
rect 3278 52782 3330 52834
rect 5294 52782 5346 52834
rect 6414 52782 6466 52834
rect 8094 52782 8146 52834
rect 14030 52782 14082 52834
rect 14478 52782 14530 52834
rect 14926 52782 14978 52834
rect 19070 52782 19122 52834
rect 24670 52782 24722 52834
rect 28142 52782 28194 52834
rect 31390 52782 31442 52834
rect 31838 52782 31890 52834
rect 33182 52782 33234 52834
rect 38446 52782 38498 52834
rect 41022 52782 41074 52834
rect 41470 52782 41522 52834
rect 43934 52782 43986 52834
rect 46062 52782 46114 52834
rect 2158 52670 2210 52722
rect 2718 52670 2770 52722
rect 5854 52670 5906 52722
rect 19630 52670 19682 52722
rect 22654 52670 22706 52722
rect 23102 52670 23154 52722
rect 32062 52670 32114 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 4062 52334 4114 52386
rect 4734 52334 4786 52386
rect 22654 52334 22706 52386
rect 35646 52334 35698 52386
rect 35982 52334 36034 52386
rect 37326 52334 37378 52386
rect 39678 52334 39730 52386
rect 42478 52334 42530 52386
rect 43598 52334 43650 52386
rect 43934 52334 43986 52386
rect 3166 52222 3218 52274
rect 7646 52222 7698 52274
rect 23214 52222 23266 52274
rect 30718 52222 30770 52274
rect 36430 52222 36482 52274
rect 38222 52222 38274 52274
rect 42142 52222 42194 52274
rect 45054 52222 45106 52274
rect 45166 52222 45218 52274
rect 2270 52110 2322 52162
rect 3502 52110 3554 52162
rect 3726 52110 3778 52162
rect 6302 52110 6354 52162
rect 12014 52110 12066 52162
rect 33518 52110 33570 52162
rect 35086 52110 35138 52162
rect 35422 52110 35474 52162
rect 37662 52110 37714 52162
rect 38334 52110 38386 52162
rect 39230 52110 39282 52162
rect 39566 52110 39618 52162
rect 40238 52110 40290 52162
rect 41134 52110 41186 52162
rect 41694 52110 41746 52162
rect 42030 52110 42082 52162
rect 42366 52110 42418 52162
rect 43934 52110 43986 52162
rect 4398 51998 4450 52050
rect 11230 51998 11282 52050
rect 22766 51998 22818 52050
rect 32734 51998 32786 52050
rect 2718 51886 2770 51938
rect 4622 51886 4674 51938
rect 11342 51886 11394 51938
rect 11566 51886 11618 51938
rect 31166 51886 31218 51938
rect 31838 51886 31890 51938
rect 32286 51886 32338 51938
rect 34526 51886 34578 51938
rect 37438 51886 37490 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 29822 51550 29874 51602
rect 30718 51550 30770 51602
rect 39902 51550 39954 51602
rect 40350 51550 40402 51602
rect 43710 51550 43762 51602
rect 44158 51550 44210 51602
rect 6974 51438 7026 51490
rect 10334 51438 10386 51490
rect 14702 51438 14754 51490
rect 20638 51438 20690 51490
rect 26574 51438 26626 51490
rect 38670 51438 38722 51490
rect 4510 51326 4562 51378
rect 4846 51326 4898 51378
rect 6302 51326 6354 51378
rect 6750 51326 6802 51378
rect 7310 51326 7362 51378
rect 7646 51326 7698 51378
rect 9662 51326 9714 51378
rect 12798 51326 12850 51378
rect 14366 51326 14418 51378
rect 19518 51326 19570 51378
rect 19854 51326 19906 51378
rect 23438 51326 23490 51378
rect 23662 51326 23714 51378
rect 26798 51326 26850 51378
rect 33070 51326 33122 51378
rect 39454 51326 39506 51378
rect 41134 51326 41186 51378
rect 41358 51326 41410 51378
rect 42142 51326 42194 51378
rect 42254 51326 42306 51378
rect 42814 51326 42866 51378
rect 3278 51214 3330 51266
rect 3726 51214 3778 51266
rect 4174 51214 4226 51266
rect 8542 51214 8594 51266
rect 12462 51214 12514 51266
rect 13470 51214 13522 51266
rect 22766 51214 22818 51266
rect 30270 51214 30322 51266
rect 31390 51214 31442 51266
rect 31838 51214 31890 51266
rect 32286 51214 32338 51266
rect 33854 51214 33906 51266
rect 35982 51214 36034 51266
rect 36542 51214 36594 51266
rect 23102 51102 23154 51154
rect 30606 51102 30658 51154
rect 31390 51102 31442 51154
rect 42702 51102 42754 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 3726 50766 3778 50818
rect 13918 50766 13970 50818
rect 27582 50766 27634 50818
rect 33854 50766 33906 50818
rect 34190 50766 34242 50818
rect 37102 50766 37154 50818
rect 37326 50766 37378 50818
rect 10782 50654 10834 50706
rect 11454 50654 11506 50706
rect 12686 50654 12738 50706
rect 14478 50654 14530 50706
rect 15822 50654 15874 50706
rect 17950 50654 18002 50706
rect 25790 50654 25842 50706
rect 27246 50654 27298 50706
rect 27806 50654 27858 50706
rect 28254 50654 28306 50706
rect 29486 50654 29538 50706
rect 32734 50654 32786 50706
rect 33294 50654 33346 50706
rect 35758 50654 35810 50706
rect 37102 50654 37154 50706
rect 37662 50654 37714 50706
rect 42030 50654 42082 50706
rect 3950 50542 4002 50594
rect 4398 50542 4450 50594
rect 4846 50542 4898 50594
rect 7310 50542 7362 50594
rect 7870 50542 7922 50594
rect 14254 50542 14306 50594
rect 18734 50542 18786 50594
rect 22542 50542 22594 50594
rect 22990 50542 23042 50594
rect 29710 50542 29762 50594
rect 30494 50542 30546 50594
rect 32398 50542 32450 50594
rect 34750 50542 34802 50594
rect 34862 50542 34914 50594
rect 35086 50542 35138 50594
rect 35310 50542 35362 50594
rect 36206 50542 36258 50594
rect 8654 50430 8706 50482
rect 23662 50430 23714 50482
rect 26238 50430 26290 50482
rect 26910 50430 26962 50482
rect 29374 50430 29426 50482
rect 31502 50430 31554 50482
rect 33966 50430 34018 50482
rect 41358 50430 41410 50482
rect 6078 50318 6130 50370
rect 14926 50318 14978 50370
rect 15486 50318 15538 50370
rect 26574 50318 26626 50370
rect 30382 50318 30434 50370
rect 34974 50318 35026 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 23662 49982 23714 50034
rect 24110 49982 24162 50034
rect 25342 49982 25394 50034
rect 29710 49982 29762 50034
rect 31054 49982 31106 50034
rect 31166 49982 31218 50034
rect 10670 49870 10722 49922
rect 14926 49870 14978 49922
rect 19294 49870 19346 49922
rect 23326 49870 23378 49922
rect 26462 49870 26514 49922
rect 31278 49870 31330 49922
rect 33966 49870 34018 49922
rect 42030 49870 42082 49922
rect 1822 49758 1874 49810
rect 5294 49758 5346 49810
rect 6862 49758 6914 49810
rect 7310 49758 7362 49810
rect 8430 49758 8482 49810
rect 9774 49758 9826 49810
rect 15598 49758 15650 49810
rect 19630 49758 19682 49810
rect 20638 49758 20690 49810
rect 25678 49758 25730 49810
rect 29710 49758 29762 49810
rect 29822 49758 29874 49810
rect 30830 49758 30882 49810
rect 31390 49758 31442 49810
rect 33070 49758 33122 49810
rect 34750 49758 34802 49810
rect 41694 49758 41746 49810
rect 42366 49758 42418 49810
rect 2494 49646 2546 49698
rect 4622 49646 4674 49698
rect 9998 49646 10050 49698
rect 11118 49646 11170 49698
rect 12798 49646 12850 49698
rect 16158 49646 16210 49698
rect 20078 49646 20130 49698
rect 20638 49646 20690 49698
rect 7758 49534 7810 49586
rect 21086 49646 21138 49698
rect 21534 49646 21586 49698
rect 23102 49646 23154 49698
rect 28590 49646 28642 49698
rect 30158 49646 30210 49698
rect 31950 49646 32002 49698
rect 32398 49646 32450 49698
rect 34078 49646 34130 49698
rect 36206 49646 36258 49698
rect 36542 49646 36594 49698
rect 41134 49646 41186 49698
rect 41918 49646 41970 49698
rect 43150 49646 43202 49698
rect 45278 49646 45330 49698
rect 21198 49534 21250 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 5966 49198 6018 49250
rect 21198 49198 21250 49250
rect 27694 49198 27746 49250
rect 28030 49198 28082 49250
rect 29822 49198 29874 49250
rect 34414 49198 34466 49250
rect 35758 49198 35810 49250
rect 42254 49198 42306 49250
rect 43038 49198 43090 49250
rect 2606 49086 2658 49138
rect 4510 49086 4562 49138
rect 6414 49086 6466 49138
rect 7982 49086 8034 49138
rect 8990 49086 9042 49138
rect 14926 49086 14978 49138
rect 18398 49086 18450 49138
rect 18734 49086 18786 49138
rect 20190 49086 20242 49138
rect 25790 49086 25842 49138
rect 28254 49086 28306 49138
rect 29262 49086 29314 49138
rect 31054 49086 31106 49138
rect 41134 49086 41186 49138
rect 41582 49086 41634 49138
rect 42590 49086 42642 49138
rect 43038 49086 43090 49138
rect 44942 49086 44994 49138
rect 2718 48974 2770 49026
rect 3278 48974 3330 49026
rect 3950 48974 4002 49026
rect 6302 48974 6354 49026
rect 6862 48974 6914 49026
rect 8206 48974 8258 49026
rect 14702 48974 14754 49026
rect 15486 48974 15538 49026
rect 19518 48974 19570 49026
rect 20078 48974 20130 49026
rect 21310 48974 21362 49026
rect 21870 48974 21922 49026
rect 22542 48974 22594 49026
rect 24446 48974 24498 49026
rect 27358 48974 27410 49026
rect 32398 48974 32450 49026
rect 33742 48974 33794 49026
rect 38334 48974 38386 49026
rect 1934 48862 1986 48914
rect 2270 48862 2322 48914
rect 7422 48862 7474 48914
rect 7646 48862 7698 48914
rect 8542 48862 8594 48914
rect 16270 48862 16322 48914
rect 20750 48862 20802 48914
rect 22654 48862 22706 48914
rect 25006 48862 25058 48914
rect 25678 48862 25730 48914
rect 30270 48862 30322 48914
rect 30382 48862 30434 48914
rect 30494 48862 30546 48914
rect 32958 48862 33010 48914
rect 33854 48862 33906 48914
rect 35870 48862 35922 48914
rect 39006 48862 39058 48914
rect 2494 48750 2546 48802
rect 3054 48750 3106 48802
rect 3166 48750 3218 48802
rect 3502 48750 3554 48802
rect 7534 48750 7586 48802
rect 8878 48750 8930 48802
rect 9102 48750 9154 48802
rect 9326 48750 9378 48802
rect 9886 48750 9938 48802
rect 10334 48750 10386 48802
rect 14030 48750 14082 48802
rect 14366 48750 14418 48802
rect 18846 48750 18898 48802
rect 23326 48750 23378 48802
rect 23886 48750 23938 48802
rect 31502 48750 31554 48802
rect 36318 48750 36370 48802
rect 37102 48750 37154 48802
rect 41694 48750 41746 48802
rect 42142 48750 42194 48802
rect 44830 48750 44882 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 2830 48414 2882 48466
rect 15150 48414 15202 48466
rect 16158 48414 16210 48466
rect 16382 48414 16434 48466
rect 24222 48414 24274 48466
rect 37662 48414 37714 48466
rect 40126 48414 40178 48466
rect 42926 48414 42978 48466
rect 1934 48078 1986 48130
rect 2382 48078 2434 48130
rect 1934 47966 1986 48018
rect 3054 48302 3106 48354
rect 9662 48302 9714 48354
rect 14142 48302 14194 48354
rect 16606 48302 16658 48354
rect 16718 48302 16770 48354
rect 18846 48302 18898 48354
rect 26798 48302 26850 48354
rect 27582 48302 27634 48354
rect 36766 48302 36818 48354
rect 38782 48302 38834 48354
rect 41246 48302 41298 48354
rect 7870 48190 7922 48242
rect 13246 48190 13298 48242
rect 13806 48190 13858 48242
rect 14366 48190 14418 48242
rect 18622 48190 18674 48242
rect 18958 48190 19010 48242
rect 19742 48190 19794 48242
rect 20302 48190 20354 48242
rect 20638 48190 20690 48242
rect 25230 48190 25282 48242
rect 28366 48190 28418 48242
rect 32510 48190 32562 48242
rect 33070 48190 33122 48242
rect 36430 48190 36482 48242
rect 41022 48190 41074 48242
rect 41582 48190 41634 48242
rect 42254 48190 42306 48242
rect 3838 48078 3890 48130
rect 8990 48078 9042 48130
rect 10446 48078 10498 48130
rect 12574 48078 12626 48130
rect 18062 48078 18114 48130
rect 21422 48078 21474 48130
rect 23550 48078 23602 48130
rect 24670 48078 24722 48130
rect 26126 48078 26178 48130
rect 28926 48078 28978 48130
rect 29598 48078 29650 48130
rect 31390 48078 31442 48130
rect 33854 48078 33906 48130
rect 35982 48078 36034 48130
rect 37214 48078 37266 48130
rect 38222 48078 38274 48130
rect 38894 48078 38946 48130
rect 39342 48078 39394 48130
rect 43374 48078 43426 48130
rect 13582 47966 13634 48018
rect 13918 47966 13970 48018
rect 19518 47966 19570 48018
rect 36990 47966 37042 48018
rect 38222 47966 38274 48018
rect 38558 47966 38610 48018
rect 40910 47966 40962 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 2942 47630 2994 47682
rect 6750 47630 6802 47682
rect 36430 47630 36482 47682
rect 2718 47518 2770 47570
rect 4174 47518 4226 47570
rect 6190 47518 6242 47570
rect 14254 47518 14306 47570
rect 16382 47518 16434 47570
rect 23998 47518 24050 47570
rect 26686 47518 26738 47570
rect 29598 47518 29650 47570
rect 29822 47518 29874 47570
rect 33182 47518 33234 47570
rect 37774 47518 37826 47570
rect 39902 47518 39954 47570
rect 40350 47518 40402 47570
rect 41134 47518 41186 47570
rect 41470 47518 41522 47570
rect 42702 47518 42754 47570
rect 42926 47518 42978 47570
rect 2494 47406 2546 47458
rect 3166 47406 3218 47458
rect 3502 47406 3554 47458
rect 3726 47406 3778 47458
rect 4062 47406 4114 47458
rect 5854 47406 5906 47458
rect 7534 47406 7586 47458
rect 9998 47406 10050 47458
rect 10334 47406 10386 47458
rect 10558 47406 10610 47458
rect 11902 47406 11954 47458
rect 13582 47406 13634 47458
rect 24446 47406 24498 47458
rect 26126 47406 26178 47458
rect 27918 47406 27970 47458
rect 28590 47406 28642 47458
rect 31502 47406 31554 47458
rect 32174 47406 32226 47458
rect 34414 47406 34466 47458
rect 34638 47406 34690 47458
rect 35870 47406 35922 47458
rect 36094 47406 36146 47458
rect 37102 47406 37154 47458
rect 40910 47406 40962 47458
rect 41694 47406 41746 47458
rect 2270 47294 2322 47346
rect 2382 47294 2434 47346
rect 9662 47294 9714 47346
rect 11230 47294 11282 47346
rect 11566 47294 11618 47346
rect 11678 47294 11730 47346
rect 12238 47294 12290 47346
rect 22094 47294 22146 47346
rect 22430 47294 22482 47346
rect 25678 47294 25730 47346
rect 26574 47294 26626 47346
rect 31390 47294 31442 47346
rect 32062 47294 32114 47346
rect 43822 47294 43874 47346
rect 4174 47182 4226 47234
rect 4398 47182 4450 47234
rect 4958 47182 5010 47234
rect 8878 47182 8930 47234
rect 9326 47182 9378 47234
rect 9774 47182 9826 47234
rect 16830 47182 16882 47234
rect 18510 47182 18562 47234
rect 19518 47182 19570 47234
rect 19966 47182 20018 47234
rect 20414 47182 20466 47234
rect 21422 47182 21474 47234
rect 29262 47182 29314 47234
rect 30158 47182 30210 47234
rect 34078 47182 34130 47234
rect 35086 47182 35138 47234
rect 35534 47182 35586 47234
rect 43262 47182 43314 47234
rect 44158 47182 44210 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 3166 46846 3218 46898
rect 4174 46846 4226 46898
rect 4510 46846 4562 46898
rect 4622 46846 4674 46898
rect 7982 46846 8034 46898
rect 8542 46846 8594 46898
rect 17614 46846 17666 46898
rect 25902 46846 25954 46898
rect 28590 46846 28642 46898
rect 31838 46846 31890 46898
rect 33854 46846 33906 46898
rect 38894 46846 38946 46898
rect 41246 46846 41298 46898
rect 4846 46734 4898 46786
rect 5518 46734 5570 46786
rect 8766 46734 8818 46786
rect 10110 46734 10162 46786
rect 10446 46734 10498 46786
rect 21534 46734 21586 46786
rect 22318 46734 22370 46786
rect 26574 46734 26626 46786
rect 28142 46734 28194 46786
rect 32398 46734 32450 46786
rect 34638 46734 34690 46786
rect 36206 46734 36258 46786
rect 37102 46734 37154 46786
rect 39006 46734 39058 46786
rect 39902 46734 39954 46786
rect 41134 46734 41186 46786
rect 43598 46734 43650 46786
rect 45950 46734 46002 46786
rect 4398 46622 4450 46674
rect 6190 46622 6242 46674
rect 6862 46622 6914 46674
rect 7198 46622 7250 46674
rect 7422 46622 7474 46674
rect 7534 46622 7586 46674
rect 8318 46622 8370 46674
rect 9662 46622 9714 46674
rect 19406 46622 19458 46674
rect 20414 46622 20466 46674
rect 21646 46622 21698 46674
rect 23998 46622 24050 46674
rect 26238 46622 26290 46674
rect 32286 46622 32338 46674
rect 34078 46622 34130 46674
rect 35534 46622 35586 46674
rect 38558 46622 38610 46674
rect 39678 46622 39730 46674
rect 41022 46622 41074 46674
rect 44718 46622 44770 46674
rect 45166 46622 45218 46674
rect 2270 46510 2322 46562
rect 2606 46510 2658 46562
rect 3614 46510 3666 46562
rect 5966 46510 6018 46562
rect 8430 46510 8482 46562
rect 9438 46510 9490 46562
rect 11118 46510 11170 46562
rect 15374 46510 15426 46562
rect 18286 46510 18338 46562
rect 18846 46510 18898 46562
rect 19854 46510 19906 46562
rect 20078 46510 20130 46562
rect 23438 46510 23490 46562
rect 29038 46510 29090 46562
rect 29822 46510 29874 46562
rect 30382 46510 30434 46562
rect 33294 46510 33346 46562
rect 37886 46510 37938 46562
rect 40350 46510 40402 46562
rect 48078 46510 48130 46562
rect 2830 46398 2882 46450
rect 17502 46398 17554 46450
rect 17838 46398 17890 46450
rect 29822 46398 29874 46450
rect 30606 46398 30658 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 2942 46062 2994 46114
rect 20414 46062 20466 46114
rect 22654 46062 22706 46114
rect 42478 46062 42530 46114
rect 43150 46062 43202 46114
rect 2158 45950 2210 46002
rect 3054 45950 3106 46002
rect 4174 45950 4226 46002
rect 9102 45950 9154 46002
rect 16830 45950 16882 46002
rect 18958 45950 19010 46002
rect 29150 45950 29202 46002
rect 33518 45950 33570 46002
rect 37774 45950 37826 46002
rect 40126 45950 40178 46002
rect 42254 45950 42306 46002
rect 43150 45950 43202 46002
rect 1934 45838 1986 45890
rect 2606 45838 2658 45890
rect 3278 45838 3330 45890
rect 3614 45838 3666 45890
rect 3726 45838 3778 45890
rect 9886 45838 9938 45890
rect 14478 45838 14530 45890
rect 16158 45838 16210 45890
rect 19294 45838 19346 45890
rect 20190 45838 20242 45890
rect 20750 45838 20802 45890
rect 22318 45838 22370 45890
rect 22990 45838 23042 45890
rect 23662 45838 23714 45890
rect 29934 45838 29986 45890
rect 30382 45838 30434 45890
rect 31278 45838 31330 45890
rect 35198 45838 35250 45890
rect 36094 45838 36146 45890
rect 39454 45838 39506 45890
rect 2382 45726 2434 45778
rect 14926 45726 14978 45778
rect 19518 45726 19570 45778
rect 23214 45726 23266 45778
rect 29374 45726 29426 45778
rect 29598 45726 29650 45778
rect 30718 45726 30770 45778
rect 34638 45726 34690 45778
rect 4622 45614 4674 45666
rect 5070 45614 5122 45666
rect 6078 45614 6130 45666
rect 6414 45614 6466 45666
rect 6862 45614 6914 45666
rect 10334 45614 10386 45666
rect 15710 45614 15762 45666
rect 21422 45614 21474 45666
rect 21870 45614 21922 45666
rect 26462 45614 26514 45666
rect 28142 45614 28194 45666
rect 28590 45614 28642 45666
rect 30158 45614 30210 45666
rect 30606 45614 30658 45666
rect 34302 45614 34354 45666
rect 37326 45614 37378 45666
rect 38222 45614 38274 45666
rect 38670 45614 38722 45666
rect 42702 45614 42754 45666
rect 43598 45614 43650 45666
rect 44046 45614 44098 45666
rect 44942 45614 44994 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 2830 45278 2882 45330
rect 19182 45278 19234 45330
rect 26910 45278 26962 45330
rect 27134 45278 27186 45330
rect 31166 45278 31218 45330
rect 32510 45278 32562 45330
rect 34302 45278 34354 45330
rect 35086 45278 35138 45330
rect 35534 45278 35586 45330
rect 39678 45278 39730 45330
rect 8094 45166 8146 45218
rect 19070 45166 19122 45218
rect 22206 45166 22258 45218
rect 23326 45166 23378 45218
rect 28030 45166 28082 45218
rect 29038 45166 29090 45218
rect 30494 45166 30546 45218
rect 31614 45166 31666 45218
rect 33070 45166 33122 45218
rect 41918 45166 41970 45218
rect 3502 45054 3554 45106
rect 12910 45054 12962 45106
rect 20974 45054 21026 45106
rect 22094 45054 22146 45106
rect 22990 45054 23042 45106
rect 25454 45054 25506 45106
rect 25678 45054 25730 45106
rect 26686 45054 26738 45106
rect 27358 45054 27410 45106
rect 27918 45054 27970 45106
rect 28254 45054 28306 45106
rect 28926 45054 28978 45106
rect 29934 45054 29986 45106
rect 30942 45054 30994 45106
rect 31390 45054 31442 45106
rect 33294 45054 33346 45106
rect 33630 45054 33682 45106
rect 37550 45054 37602 45106
rect 38110 45054 38162 45106
rect 38782 45054 38834 45106
rect 41694 45054 41746 45106
rect 42366 45054 42418 45106
rect 42926 45054 42978 45106
rect 43486 45054 43538 45106
rect 2382 44942 2434 44994
rect 16494 44942 16546 44994
rect 19630 44942 19682 44994
rect 21758 44942 21810 44994
rect 23662 44942 23714 44994
rect 24222 44942 24274 44994
rect 24670 44942 24722 44994
rect 27246 44942 27298 44994
rect 27694 44942 27746 44994
rect 29374 44942 29426 44994
rect 31278 44942 31330 44994
rect 32062 44942 32114 44994
rect 34638 44942 34690 44994
rect 35982 44942 36034 44994
rect 36766 44942 36818 44994
rect 37102 44942 37154 44994
rect 38558 44942 38610 44994
rect 39118 44942 39170 44994
rect 39342 44942 39394 44994
rect 40126 44942 40178 44994
rect 41246 44942 41298 44994
rect 44270 44942 44322 44994
rect 46398 44942 46450 44994
rect 23998 44830 24050 44882
rect 26014 44830 26066 44882
rect 28702 44830 28754 44882
rect 35534 44830 35586 44882
rect 35870 44830 35922 44882
rect 41582 44830 41634 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 21982 44494 22034 44546
rect 22542 44494 22594 44546
rect 38782 44494 38834 44546
rect 44046 44494 44098 44546
rect 6302 44382 6354 44434
rect 6750 44382 6802 44434
rect 12910 44382 12962 44434
rect 13582 44382 13634 44434
rect 16606 44382 16658 44434
rect 18622 44382 18674 44434
rect 21422 44382 21474 44434
rect 21982 44382 22034 44434
rect 23550 44382 23602 44434
rect 25678 44382 25730 44434
rect 27358 44382 27410 44434
rect 28030 44382 28082 44434
rect 33406 44382 33458 44434
rect 39902 44382 39954 44434
rect 40350 44382 40402 44434
rect 42702 44382 42754 44434
rect 43374 44382 43426 44434
rect 43710 44382 43762 44434
rect 2494 44270 2546 44322
rect 2942 44270 2994 44322
rect 3502 44270 3554 44322
rect 4398 44270 4450 44322
rect 4734 44270 4786 44322
rect 5966 44270 6018 44322
rect 6190 44270 6242 44322
rect 6526 44270 6578 44322
rect 9662 44270 9714 44322
rect 10110 44270 10162 44322
rect 16382 44270 16434 44322
rect 19182 44270 19234 44322
rect 22766 44270 22818 44322
rect 28366 44270 28418 44322
rect 29150 44270 29202 44322
rect 30606 44270 30658 44322
rect 32174 44270 32226 44322
rect 33070 44270 33122 44322
rect 34974 44270 35026 44322
rect 35422 44270 35474 44322
rect 37662 44270 37714 44322
rect 38334 44270 38386 44322
rect 39006 44270 39058 44322
rect 41582 44270 41634 44322
rect 42590 44270 42642 44322
rect 44046 44270 44098 44322
rect 2830 44158 2882 44210
rect 4174 44158 4226 44210
rect 8878 44158 8930 44210
rect 10782 44158 10834 44210
rect 15486 44158 15538 44210
rect 16046 44158 16098 44210
rect 19070 44158 19122 44210
rect 26126 44158 26178 44210
rect 26238 44158 26290 44210
rect 28478 44158 28530 44210
rect 30382 44158 30434 44210
rect 31950 44158 32002 44210
rect 32958 44158 33010 44210
rect 35982 44158 36034 44210
rect 37774 44158 37826 44210
rect 39454 44158 39506 44210
rect 40798 44158 40850 44210
rect 42814 44158 42866 44210
rect 2606 44046 2658 44098
rect 3838 44046 3890 44098
rect 15150 44046 15202 44098
rect 17054 44046 17106 44098
rect 17502 44046 17554 44098
rect 18846 44046 18898 44098
rect 20638 44046 20690 44098
rect 22430 44046 22482 44098
rect 26462 44046 26514 44098
rect 26798 44046 26850 44098
rect 28702 44046 28754 44098
rect 29262 44046 29314 44098
rect 29486 44046 29538 44098
rect 31166 44046 31218 44098
rect 35198 44046 35250 44098
rect 35310 44046 35362 44098
rect 35534 44046 35586 44098
rect 36318 44046 36370 44098
rect 37214 44046 37266 44098
rect 41246 44046 41298 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 8654 43710 8706 43762
rect 8878 43710 8930 43762
rect 9886 43710 9938 43762
rect 10334 43710 10386 43762
rect 11342 43710 11394 43762
rect 17838 43710 17890 43762
rect 41806 43710 41858 43762
rect 8206 43598 8258 43650
rect 14702 43598 14754 43650
rect 18958 43598 19010 43650
rect 22878 43598 22930 43650
rect 23998 43598 24050 43650
rect 28814 43598 28866 43650
rect 30942 43598 30994 43650
rect 34750 43598 34802 43650
rect 35534 43598 35586 43650
rect 38222 43598 38274 43650
rect 41022 43598 41074 43650
rect 42814 43598 42866 43650
rect 44270 43598 44322 43650
rect 45950 43598 46002 43650
rect 6638 43486 6690 43538
rect 7534 43486 7586 43538
rect 7870 43486 7922 43538
rect 8542 43486 8594 43538
rect 13918 43486 13970 43538
rect 18286 43486 18338 43538
rect 21422 43486 21474 43538
rect 23550 43486 23602 43538
rect 30382 43486 30434 43538
rect 32286 43486 32338 43538
rect 34638 43486 34690 43538
rect 37102 43486 37154 43538
rect 37438 43486 37490 43538
rect 43262 43486 43314 43538
rect 43710 43486 43762 43538
rect 2718 43374 2770 43426
rect 10894 43374 10946 43426
rect 11790 43374 11842 43426
rect 16830 43374 16882 43426
rect 21086 43374 21138 43426
rect 21758 43374 21810 43426
rect 25342 43374 25394 43426
rect 29262 43374 29314 43426
rect 30046 43374 30098 43426
rect 31502 43374 31554 43426
rect 31838 43374 31890 43426
rect 33182 43374 33234 43426
rect 40350 43374 40402 43426
rect 7422 43262 7474 43314
rect 10782 43262 10834 43314
rect 11454 43262 11506 43314
rect 32958 43262 33010 43314
rect 33518 43262 33570 43314
rect 33966 43262 34018 43314
rect 45838 43262 45890 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 20862 42926 20914 42978
rect 25678 42926 25730 42978
rect 26574 42926 26626 42978
rect 27806 42926 27858 42978
rect 2606 42814 2658 42866
rect 4062 42814 4114 42866
rect 6750 42814 6802 42866
rect 7198 42814 7250 42866
rect 7758 42814 7810 42866
rect 11454 42814 11506 42866
rect 16158 42814 16210 42866
rect 17614 42814 17666 42866
rect 18958 42814 19010 42866
rect 21310 42814 21362 42866
rect 26574 42814 26626 42866
rect 29262 42814 29314 42866
rect 29822 42814 29874 42866
rect 30718 42814 30770 42866
rect 31166 42814 31218 42866
rect 32958 42814 33010 42866
rect 35198 42814 35250 42866
rect 1934 42702 1986 42754
rect 2270 42702 2322 42754
rect 2494 42702 2546 42754
rect 2718 42702 2770 42754
rect 3502 42702 3554 42754
rect 4398 42702 4450 42754
rect 6190 42702 6242 42754
rect 6526 42702 6578 42754
rect 10558 42702 10610 42754
rect 13918 42702 13970 42754
rect 19294 42702 19346 42754
rect 20078 42702 20130 42754
rect 20750 42702 20802 42754
rect 27246 42702 27298 42754
rect 33294 42702 33346 42754
rect 33518 42702 33570 42754
rect 35534 42702 35586 42754
rect 35758 42702 35810 42754
rect 37550 42702 37602 42754
rect 37662 42702 37714 42754
rect 39790 42702 39842 42754
rect 40238 42702 40290 42754
rect 2942 42590 2994 42642
rect 3278 42590 3330 42642
rect 3726 42590 3778 42642
rect 4174 42590 4226 42642
rect 9886 42590 9938 42642
rect 11006 42590 11058 42642
rect 11230 42590 11282 42642
rect 11566 42590 11618 42642
rect 19406 42590 19458 42642
rect 27134 42590 27186 42642
rect 27358 42590 27410 42642
rect 33182 42590 33234 42642
rect 33966 42590 34018 42642
rect 35422 42590 35474 42642
rect 37438 42590 37490 42642
rect 38670 42590 38722 42642
rect 40686 42590 40738 42642
rect 2046 42478 2098 42530
rect 3838 42478 3890 42530
rect 4846 42478 4898 42530
rect 4958 42478 5010 42530
rect 5070 42478 5122 42530
rect 12126 42478 12178 42530
rect 12574 42478 12626 42530
rect 12910 42478 12962 42530
rect 17166 42478 17218 42530
rect 18062 42478 18114 42530
rect 18510 42478 18562 42530
rect 21422 42478 21474 42530
rect 21870 42478 21922 42530
rect 22318 42478 22370 42530
rect 26014 42478 26066 42530
rect 28254 42478 28306 42530
rect 30270 42478 30322 42530
rect 36206 42478 36258 42530
rect 36990 42478 37042 42530
rect 38222 42478 38274 42530
rect 42478 42478 42530 42530
rect 42926 42478 42978 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 2270 42142 2322 42194
rect 8990 42142 9042 42194
rect 9438 42142 9490 42194
rect 9662 42142 9714 42194
rect 10558 42142 10610 42194
rect 14814 42142 14866 42194
rect 16606 42142 16658 42194
rect 23326 42142 23378 42194
rect 28814 42142 28866 42194
rect 34974 42142 35026 42194
rect 2718 42030 2770 42082
rect 10446 42030 10498 42082
rect 17502 42030 17554 42082
rect 18622 42030 18674 42082
rect 23438 42030 23490 42082
rect 29262 42030 29314 42082
rect 30270 42030 30322 42082
rect 32286 42030 32338 42082
rect 33070 42030 33122 42082
rect 36094 42030 36146 42082
rect 37326 42030 37378 42082
rect 40126 42030 40178 42082
rect 40238 42030 40290 42082
rect 2830 41918 2882 41970
rect 3838 41918 3890 41970
rect 9774 41918 9826 41970
rect 10110 41918 10162 41970
rect 10670 41918 10722 41970
rect 11006 41918 11058 41970
rect 14478 41918 14530 41970
rect 16158 41918 16210 41970
rect 17726 41918 17778 41970
rect 18398 41918 18450 41970
rect 18734 41918 18786 41970
rect 19070 41918 19122 41970
rect 19406 41918 19458 41970
rect 21982 41918 22034 41970
rect 23102 41918 23154 41970
rect 24670 41918 24722 41970
rect 25230 41918 25282 41970
rect 29374 41918 29426 41970
rect 30046 41918 30098 41970
rect 31502 41918 31554 41970
rect 33854 41918 33906 41970
rect 35534 41918 35586 41970
rect 38670 41918 38722 41970
rect 39118 41918 39170 41970
rect 41246 41918 41298 41970
rect 41470 41918 41522 41970
rect 42254 41918 42306 41970
rect 42814 41918 42866 41970
rect 43822 41918 43874 41970
rect 7534 41806 7586 41858
rect 11790 41806 11842 41858
rect 13918 41806 13970 41858
rect 16494 41806 16546 41858
rect 19966 41806 20018 41858
rect 23886 41806 23938 41858
rect 26014 41806 26066 41858
rect 28142 41806 28194 41858
rect 30270 41806 30322 41858
rect 31838 41806 31890 41858
rect 33966 41806 34018 41858
rect 35982 41806 36034 41858
rect 43374 41806 43426 41858
rect 44606 41806 44658 41858
rect 2942 41694 2994 41746
rect 18062 41694 18114 41746
rect 22654 41694 22706 41746
rect 23662 41694 23714 41746
rect 23886 41694 23938 41746
rect 39342 41694 39394 41746
rect 39678 41694 39730 41746
rect 40238 41694 40290 41746
rect 41918 41694 41970 41746
rect 43598 41694 43650 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 25566 41358 25618 41410
rect 27470 41358 27522 41410
rect 27806 41358 27858 41410
rect 36094 41358 36146 41410
rect 44270 41358 44322 41410
rect 45166 41358 45218 41410
rect 2494 41246 2546 41298
rect 4622 41246 4674 41298
rect 8430 41246 8482 41298
rect 11454 41246 11506 41298
rect 13694 41246 13746 41298
rect 15934 41246 15986 41298
rect 17950 41246 18002 41298
rect 19966 41246 20018 41298
rect 20750 41246 20802 41298
rect 22094 41246 22146 41298
rect 24222 41246 24274 41298
rect 25790 41246 25842 41298
rect 28254 41246 28306 41298
rect 29934 41246 29986 41298
rect 32398 41246 32450 41298
rect 36318 41246 36370 41298
rect 37102 41246 37154 41298
rect 40462 41246 40514 41298
rect 41694 41246 41746 41298
rect 43822 41246 43874 41298
rect 44158 41246 44210 41298
rect 44830 41246 44882 41298
rect 1822 41134 1874 41186
rect 6526 41134 6578 41186
rect 11566 41134 11618 41186
rect 11902 41134 11954 41186
rect 12350 41134 12402 41186
rect 12462 41134 12514 41186
rect 14030 41134 14082 41186
rect 19070 41134 19122 41186
rect 21422 41134 21474 41186
rect 24670 41134 24722 41186
rect 25230 41134 25282 41186
rect 26798 41134 26850 41186
rect 26910 41134 26962 41186
rect 29710 41134 29762 41186
rect 30046 41134 30098 41186
rect 30718 41134 30770 41186
rect 33294 41134 33346 41186
rect 34414 41134 34466 41186
rect 35646 41134 35698 41186
rect 37550 41134 37602 41186
rect 38334 41134 38386 41186
rect 40910 41134 40962 41186
rect 11342 41022 11394 41074
rect 12686 41022 12738 41074
rect 27022 41022 27074 41074
rect 27582 41022 27634 41074
rect 32174 41022 32226 41074
rect 33070 41022 33122 41074
rect 35534 41022 35586 41074
rect 5070 40910 5122 40962
rect 12238 40910 12290 40962
rect 24894 40910 24946 40962
rect 26350 40910 26402 40962
rect 29262 40910 29314 40962
rect 29822 40910 29874 40962
rect 30158 40910 30210 40962
rect 34526 40910 34578 40962
rect 34638 40910 34690 40962
rect 36318 40910 36370 40962
rect 44942 40910 44994 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 2494 40574 2546 40626
rect 3614 40574 3666 40626
rect 4398 40574 4450 40626
rect 24670 40574 24722 40626
rect 28926 40574 28978 40626
rect 32510 40574 32562 40626
rect 40238 40574 40290 40626
rect 42814 40574 42866 40626
rect 5630 40462 5682 40514
rect 6302 40462 6354 40514
rect 7982 40462 8034 40514
rect 8318 40462 8370 40514
rect 9550 40462 9602 40514
rect 12238 40462 12290 40514
rect 17502 40462 17554 40514
rect 18734 40462 18786 40514
rect 18958 40462 19010 40514
rect 20526 40462 20578 40514
rect 26462 40462 26514 40514
rect 28478 40462 28530 40514
rect 29822 40462 29874 40514
rect 31950 40462 32002 40514
rect 33630 40462 33682 40514
rect 34862 40462 34914 40514
rect 40350 40462 40402 40514
rect 40910 40462 40962 40514
rect 44382 40462 44434 40514
rect 2718 40350 2770 40402
rect 3166 40350 3218 40402
rect 4846 40350 4898 40402
rect 5518 40350 5570 40402
rect 6414 40350 6466 40402
rect 7086 40350 7138 40402
rect 7646 40350 7698 40402
rect 8430 40350 8482 40402
rect 9998 40350 10050 40402
rect 11006 40350 11058 40402
rect 15374 40350 15426 40402
rect 18174 40350 18226 40402
rect 19182 40350 19234 40402
rect 19966 40350 20018 40402
rect 21758 40350 21810 40402
rect 26910 40350 26962 40402
rect 27358 40350 27410 40402
rect 29486 40350 29538 40402
rect 30158 40350 30210 40402
rect 33518 40350 33570 40402
rect 34750 40350 34802 40402
rect 36654 40350 36706 40402
rect 37438 40350 37490 40402
rect 38334 40350 38386 40402
rect 38558 40350 38610 40402
rect 39678 40350 39730 40402
rect 41022 40350 41074 40402
rect 43598 40350 43650 40402
rect 2158 40238 2210 40290
rect 2606 40238 2658 40290
rect 3726 40238 3778 40290
rect 9886 40238 9938 40290
rect 21870 40238 21922 40290
rect 35870 40238 35922 40290
rect 39454 40238 39506 40290
rect 41358 40238 41410 40290
rect 43262 40238 43314 40290
rect 46510 40238 46562 40290
rect 3838 40126 3890 40178
rect 30718 40126 30770 40178
rect 32174 40126 32226 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 5070 39790 5122 39842
rect 30158 39790 30210 39842
rect 38334 39790 38386 39842
rect 2830 39678 2882 39730
rect 3838 39678 3890 39730
rect 4510 39678 4562 39730
rect 5854 39678 5906 39730
rect 10894 39678 10946 39730
rect 13582 39678 13634 39730
rect 16830 39678 16882 39730
rect 17950 39678 18002 39730
rect 20078 39678 20130 39730
rect 28142 39678 28194 39730
rect 28590 39678 28642 39730
rect 29374 39678 29426 39730
rect 31278 39678 31330 39730
rect 35198 39678 35250 39730
rect 36430 39678 36482 39730
rect 37102 39678 37154 39730
rect 1822 39566 1874 39618
rect 4734 39566 4786 39618
rect 5742 39566 5794 39618
rect 6974 39566 7026 39618
rect 7198 39566 7250 39618
rect 12798 39566 12850 39618
rect 13918 39566 13970 39618
rect 17278 39566 17330 39618
rect 21982 39566 22034 39618
rect 23438 39566 23490 39618
rect 25902 39566 25954 39618
rect 26126 39566 26178 39618
rect 27246 39566 27298 39618
rect 33070 39566 33122 39618
rect 33406 39566 33458 39618
rect 37774 39566 37826 39618
rect 5966 39454 6018 39506
rect 14702 39454 14754 39506
rect 23550 39454 23602 39506
rect 24222 39454 24274 39506
rect 26238 39454 26290 39506
rect 27358 39454 27410 39506
rect 27582 39454 27634 39506
rect 32510 39454 32562 39506
rect 39902 39790 39954 39842
rect 45054 39790 45106 39842
rect 39902 39678 39954 39730
rect 40350 39678 40402 39730
rect 40910 39678 40962 39730
rect 41358 39678 41410 39730
rect 42142 39678 42194 39730
rect 44270 39678 44322 39730
rect 46510 39678 46562 39730
rect 41470 39566 41522 39618
rect 42590 39566 42642 39618
rect 44830 39566 44882 39618
rect 46398 39566 46450 39618
rect 33966 39454 34018 39506
rect 39118 39454 39170 39506
rect 42926 39454 42978 39506
rect 45390 39454 45442 39506
rect 45726 39454 45778 39506
rect 2046 39342 2098 39394
rect 3278 39342 3330 39394
rect 4286 39342 4338 39394
rect 20526 39342 20578 39394
rect 21422 39342 21474 39394
rect 23662 39342 23714 39394
rect 26350 39342 26402 39394
rect 26462 39342 26514 39394
rect 29934 39342 29986 39394
rect 30046 39342 30098 39394
rect 30718 39342 30770 39394
rect 34974 39342 35026 39394
rect 39454 39342 39506 39394
rect 46062 39342 46114 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 2270 39006 2322 39058
rect 2382 39006 2434 39058
rect 2494 39006 2546 39058
rect 3166 39006 3218 39058
rect 10110 39006 10162 39058
rect 10558 39006 10610 39058
rect 11454 39006 11506 39058
rect 15374 39006 15426 39058
rect 16270 39006 16322 39058
rect 20526 39006 20578 39058
rect 21086 39006 21138 39058
rect 21310 39006 21362 39058
rect 21982 39006 22034 39058
rect 31838 39006 31890 39058
rect 33182 39006 33234 39058
rect 33630 39006 33682 39058
rect 34078 39006 34130 39058
rect 38446 39006 38498 39058
rect 38894 39006 38946 39058
rect 41022 39006 41074 39058
rect 41918 39006 41970 39058
rect 42366 39006 42418 39058
rect 43486 39006 43538 39058
rect 3054 38894 3106 38946
rect 3950 38894 4002 38946
rect 20862 38894 20914 38946
rect 26462 38894 26514 38946
rect 26798 38894 26850 38946
rect 29598 38894 29650 38946
rect 30494 38894 30546 38946
rect 31950 38894 32002 38946
rect 39342 38894 39394 38946
rect 1822 38782 1874 38834
rect 2830 38782 2882 38834
rect 3502 38782 3554 38834
rect 7534 38782 7586 38834
rect 9662 38782 9714 38834
rect 11790 38782 11842 38834
rect 15710 38782 15762 38834
rect 16606 38782 16658 38834
rect 17950 38782 18002 38834
rect 21534 38782 21586 38834
rect 21646 38782 21698 38834
rect 26910 38782 26962 38834
rect 27358 38782 27410 38834
rect 28030 38782 28082 38834
rect 30830 38782 30882 38834
rect 32286 38782 32338 38834
rect 37438 38782 37490 38834
rect 39678 38782 39730 38834
rect 40014 38782 40066 38834
rect 41470 38782 41522 38834
rect 11006 38670 11058 38722
rect 12574 38670 12626 38722
rect 14702 38670 14754 38722
rect 19182 38670 19234 38722
rect 26350 38670 26402 38722
rect 28702 38670 28754 38722
rect 34638 38670 34690 38722
rect 36766 38670 36818 38722
rect 38110 38670 38162 38722
rect 42814 38670 42866 38722
rect 9550 38558 9602 38610
rect 10670 38558 10722 38610
rect 11342 38558 11394 38610
rect 15934 38558 15986 38610
rect 16158 38558 16210 38610
rect 40014 38558 40066 38610
rect 41134 38558 41186 38610
rect 41694 38558 41746 38610
rect 42478 38558 42530 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 19966 38222 20018 38274
rect 29262 38222 29314 38274
rect 29934 38222 29986 38274
rect 43822 38222 43874 38274
rect 1710 38110 1762 38162
rect 4062 38110 4114 38162
rect 10670 38110 10722 38162
rect 12350 38110 12402 38162
rect 18398 38110 18450 38162
rect 20190 38110 20242 38162
rect 24222 38110 24274 38162
rect 27246 38110 27298 38162
rect 28254 38110 28306 38162
rect 29262 38110 29314 38162
rect 29710 38110 29762 38162
rect 30718 38110 30770 38162
rect 35870 38110 35922 38162
rect 37998 38110 38050 38162
rect 40126 38110 40178 38162
rect 41358 38110 41410 38162
rect 1822 37998 1874 38050
rect 2830 37998 2882 38050
rect 3278 37998 3330 38050
rect 4398 37998 4450 38050
rect 4958 37998 5010 38050
rect 6302 37998 6354 38050
rect 7646 37998 7698 38050
rect 9438 37998 9490 38050
rect 11454 37998 11506 38050
rect 11902 37998 11954 38050
rect 12126 37998 12178 38050
rect 15374 37998 15426 38050
rect 21310 37998 21362 38050
rect 27582 37998 27634 38050
rect 27806 37998 27858 38050
rect 33294 37998 33346 38050
rect 33742 37998 33794 38050
rect 36094 37998 36146 38050
rect 37214 37998 37266 38050
rect 40910 37998 40962 38050
rect 41918 37998 41970 38050
rect 42142 37998 42194 38050
rect 42926 37998 42978 38050
rect 2158 37886 2210 37938
rect 4286 37886 4338 37938
rect 4622 37886 4674 37938
rect 6526 37886 6578 37938
rect 9998 37886 10050 37938
rect 11118 37886 11170 37938
rect 12462 37886 12514 37938
rect 22094 37886 22146 37938
rect 27246 37886 27298 37938
rect 31278 37886 31330 37938
rect 32286 37886 32338 37938
rect 34302 37886 34354 37938
rect 36430 37886 36482 37938
rect 36990 37886 37042 37938
rect 42590 37886 42642 37938
rect 44046 37886 44098 37938
rect 2270 37774 2322 37826
rect 2494 37774 2546 37826
rect 4846 37774 4898 37826
rect 5854 37774 5906 37826
rect 11342 37774 11394 37826
rect 11566 37774 11618 37826
rect 12910 37774 12962 37826
rect 13582 37774 13634 37826
rect 19630 37774 19682 37826
rect 20750 37774 20802 37826
rect 27358 37774 27410 37826
rect 30158 37774 30210 37826
rect 34974 37774 35026 37826
rect 42366 37774 42418 37826
rect 42702 37774 42754 37826
rect 43038 37774 43090 37826
rect 43150 37774 43202 37826
rect 43374 37774 43426 37826
rect 43934 37774 43986 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 5182 37438 5234 37490
rect 5630 37438 5682 37490
rect 9886 37438 9938 37490
rect 16158 37438 16210 37490
rect 17950 37438 18002 37490
rect 21198 37438 21250 37490
rect 26126 37438 26178 37490
rect 27022 37438 27074 37490
rect 28142 37438 28194 37490
rect 29598 37438 29650 37490
rect 30606 37438 30658 37490
rect 30942 37438 30994 37490
rect 32510 37438 32562 37490
rect 36766 37438 36818 37490
rect 41134 37438 41186 37490
rect 41582 37438 41634 37490
rect 7198 37326 7250 37378
rect 7534 37326 7586 37378
rect 8990 37326 9042 37378
rect 9662 37326 9714 37378
rect 9774 37326 9826 37378
rect 19070 37326 19122 37378
rect 19406 37326 19458 37378
rect 26350 37326 26402 37378
rect 27358 37326 27410 37378
rect 29262 37326 29314 37378
rect 29486 37326 29538 37378
rect 31838 37326 31890 37378
rect 33966 37326 34018 37378
rect 34750 37326 34802 37378
rect 42590 37326 42642 37378
rect 44046 37326 44098 37378
rect 2158 37214 2210 37266
rect 6078 37214 6130 37266
rect 6750 37214 6802 37266
rect 7870 37214 7922 37266
rect 8542 37214 8594 37266
rect 8654 37214 8706 37266
rect 10334 37214 10386 37266
rect 10558 37214 10610 37266
rect 19742 37214 19794 37266
rect 24670 37214 24722 37266
rect 26462 37214 26514 37266
rect 27918 37214 27970 37266
rect 28366 37214 28418 37266
rect 28590 37214 28642 37266
rect 29822 37214 29874 37266
rect 31390 37214 31442 37266
rect 33070 37214 33122 37266
rect 36206 37214 36258 37266
rect 37662 37214 37714 37266
rect 43150 37214 43202 37266
rect 45166 37214 45218 37266
rect 45726 37214 45778 37266
rect 1934 37102 1986 37154
rect 3614 37102 3666 37154
rect 8878 37102 8930 37154
rect 14366 37102 14418 37154
rect 16718 37102 16770 37154
rect 17502 37102 17554 37154
rect 18734 37102 18786 37154
rect 21758 37102 21810 37154
rect 23886 37102 23938 37154
rect 25342 37102 25394 37154
rect 25902 37102 25954 37154
rect 28254 37102 28306 37154
rect 37214 37102 37266 37154
rect 38110 37102 38162 37154
rect 16494 36990 16546 37042
rect 29710 36990 29762 37042
rect 34414 36990 34466 37042
rect 37102 36990 37154 37042
rect 37438 36990 37490 37042
rect 38110 36990 38162 37042
rect 45614 36990 45666 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 2046 36654 2098 36706
rect 3390 36654 3442 36706
rect 24894 36654 24946 36706
rect 27582 36654 27634 36706
rect 27806 36654 27858 36706
rect 38110 36654 38162 36706
rect 2382 36542 2434 36594
rect 8094 36542 8146 36594
rect 9214 36542 9266 36594
rect 11342 36542 11394 36594
rect 15710 36542 15762 36594
rect 18622 36542 18674 36594
rect 20750 36542 20802 36594
rect 26126 36542 26178 36594
rect 30830 36542 30882 36594
rect 32286 36542 32338 36594
rect 35422 36542 35474 36594
rect 36990 36542 37042 36594
rect 37998 36542 38050 36594
rect 41358 36542 41410 36594
rect 43486 36542 43538 36594
rect 45950 36542 46002 36594
rect 48078 36542 48130 36594
rect 2942 36430 2994 36482
rect 3614 36430 3666 36482
rect 6190 36430 6242 36482
rect 6750 36430 6802 36482
rect 8542 36430 8594 36482
rect 14702 36430 14754 36482
rect 17838 36430 17890 36482
rect 25118 36430 25170 36482
rect 25566 36430 25618 36482
rect 25790 36430 25842 36482
rect 26910 36430 26962 36482
rect 29598 36430 29650 36482
rect 29822 36430 29874 36482
rect 30158 36430 30210 36482
rect 30942 36430 30994 36482
rect 32622 36430 32674 36482
rect 33630 36430 33682 36482
rect 35086 36430 35138 36482
rect 35310 36430 35362 36482
rect 37214 36430 37266 36482
rect 41134 36430 41186 36482
rect 41694 36430 41746 36482
rect 45278 36430 45330 36482
rect 2606 36318 2658 36370
rect 7198 36318 7250 36370
rect 17390 36318 17442 36370
rect 23774 36318 23826 36370
rect 24110 36318 24162 36370
rect 24558 36318 24610 36370
rect 26126 36318 26178 36370
rect 27246 36318 27298 36370
rect 27470 36318 27522 36370
rect 27918 36318 27970 36370
rect 30270 36318 30322 36370
rect 31614 36318 31666 36370
rect 35758 36318 35810 36370
rect 6302 36206 6354 36258
rect 17054 36206 17106 36258
rect 21422 36206 21474 36258
rect 26014 36206 26066 36258
rect 26686 36206 26738 36258
rect 28366 36206 28418 36258
rect 29262 36206 29314 36258
rect 32958 36206 33010 36258
rect 34638 36206 34690 36258
rect 35534 36206 35586 36258
rect 36206 36206 36258 36258
rect 37550 36206 37602 36258
rect 40462 36206 40514 36258
rect 40798 36206 40850 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 2494 35870 2546 35922
rect 2606 35870 2658 35922
rect 3502 35870 3554 35922
rect 6078 35870 6130 35922
rect 10670 35870 10722 35922
rect 12686 35870 12738 35922
rect 28142 35870 28194 35922
rect 31614 35870 31666 35922
rect 32062 35870 32114 35922
rect 41358 35870 41410 35922
rect 2830 35758 2882 35810
rect 5630 35758 5682 35810
rect 6190 35758 6242 35810
rect 18174 35758 18226 35810
rect 29598 35758 29650 35810
rect 30718 35758 30770 35810
rect 37550 35758 37602 35810
rect 37886 35758 37938 35810
rect 44046 35758 44098 35810
rect 2942 35646 2994 35698
rect 5854 35646 5906 35698
rect 11342 35646 11394 35698
rect 19966 35646 20018 35698
rect 30942 35646 30994 35698
rect 31166 35646 31218 35698
rect 35198 35646 35250 35698
rect 43262 35646 43314 35698
rect 8094 35534 8146 35586
rect 8542 35534 8594 35586
rect 15934 35534 15986 35586
rect 16382 35534 16434 35586
rect 16830 35534 16882 35586
rect 20414 35534 20466 35586
rect 25566 35534 25618 35586
rect 30046 35534 30098 35586
rect 30718 35534 30770 35586
rect 32510 35534 32562 35586
rect 34750 35534 34802 35586
rect 35982 35534 36034 35586
rect 36654 35534 36706 35586
rect 42926 35534 42978 35586
rect 46174 35534 46226 35586
rect 34750 35422 34802 35474
rect 34974 35422 35026 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 2382 35086 2434 35138
rect 4846 35086 4898 35138
rect 18510 35086 18562 35138
rect 4174 34974 4226 35026
rect 8766 34974 8818 35026
rect 12798 34974 12850 35026
rect 17950 34974 18002 35026
rect 19070 34974 19122 35026
rect 19518 34974 19570 35026
rect 25790 34974 25842 35026
rect 37886 34974 37938 35026
rect 40014 34974 40066 35026
rect 44942 34974 44994 35026
rect 3054 34862 3106 34914
rect 8654 34862 8706 34914
rect 10782 34862 10834 34914
rect 11118 34862 11170 34914
rect 11454 34862 11506 34914
rect 11902 34862 11954 34914
rect 12462 34862 12514 34914
rect 14254 34862 14306 34914
rect 18846 34862 18898 34914
rect 30382 34862 30434 34914
rect 32062 34862 32114 34914
rect 37214 34862 37266 34914
rect 40798 34862 40850 34914
rect 3950 34750 4002 34802
rect 4174 34750 4226 34802
rect 4958 34750 5010 34802
rect 6974 34750 7026 34802
rect 21422 34750 21474 34802
rect 21758 34750 21810 34802
rect 31278 34750 31330 34802
rect 34414 34750 34466 34802
rect 4846 34638 4898 34690
rect 6638 34638 6690 34690
rect 7086 34638 7138 34690
rect 7198 34638 7250 34690
rect 7758 34638 7810 34690
rect 8990 34638 9042 34690
rect 10558 34638 10610 34690
rect 11118 34638 11170 34690
rect 11790 34638 11842 34690
rect 12014 34638 12066 34690
rect 13582 34638 13634 34690
rect 27022 34638 27074 34690
rect 27470 34638 27522 34690
rect 27918 34638 27970 34690
rect 29934 34638 29986 34690
rect 31726 34638 31778 34690
rect 34750 34638 34802 34690
rect 36430 34638 36482 34690
rect 40574 34638 40626 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 2830 34302 2882 34354
rect 5854 34302 5906 34354
rect 8766 34302 8818 34354
rect 26126 34302 26178 34354
rect 33630 34302 33682 34354
rect 39118 34302 39170 34354
rect 42702 34302 42754 34354
rect 4398 34190 4450 34242
rect 4846 34190 4898 34242
rect 5630 34190 5682 34242
rect 6302 34190 6354 34242
rect 7646 34190 7698 34242
rect 7982 34190 8034 34242
rect 10782 34190 10834 34242
rect 25790 34190 25842 34242
rect 29262 34190 29314 34242
rect 30158 34190 30210 34242
rect 33070 34190 33122 34242
rect 35422 34190 35474 34242
rect 39454 34190 39506 34242
rect 39678 34190 39730 34242
rect 40238 34190 40290 34242
rect 43038 34190 43090 34242
rect 43262 34190 43314 34242
rect 1934 34078 1986 34130
rect 2158 34078 2210 34130
rect 3950 34078 4002 34130
rect 4734 34078 4786 34130
rect 5518 34078 5570 34130
rect 6862 34078 6914 34130
rect 7086 34078 7138 34130
rect 8318 34078 8370 34130
rect 14366 34078 14418 34130
rect 15934 34078 15986 34130
rect 17614 34078 17666 34130
rect 24558 34078 24610 34130
rect 26462 34078 26514 34130
rect 29374 34078 29426 34130
rect 29710 34078 29762 34130
rect 34638 34078 34690 34130
rect 40126 34078 40178 34130
rect 4286 33966 4338 34018
rect 6078 33966 6130 34018
rect 6190 33966 6242 34018
rect 16382 33966 16434 34018
rect 19070 33966 19122 34018
rect 21422 33966 21474 34018
rect 21758 33966 21810 34018
rect 23886 33966 23938 34018
rect 26686 33966 26738 34018
rect 27134 33966 27186 34018
rect 28814 33966 28866 34018
rect 32510 33966 32562 34018
rect 34302 33966 34354 34018
rect 37550 33966 37602 34018
rect 2382 33854 2434 33906
rect 18398 33854 18450 33906
rect 25230 33854 25282 33906
rect 25566 33854 25618 33906
rect 33294 33854 33346 33906
rect 39790 33854 39842 33906
rect 43374 33854 43426 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 8206 33518 8258 33570
rect 14030 33518 14082 33570
rect 14366 33518 14418 33570
rect 21310 33518 21362 33570
rect 21646 33518 21698 33570
rect 34190 33518 34242 33570
rect 44830 33518 44882 33570
rect 3614 33406 3666 33458
rect 7422 33406 7474 33458
rect 8094 33406 8146 33458
rect 11454 33406 11506 33458
rect 15822 33406 15874 33458
rect 17950 33406 18002 33458
rect 20750 33406 20802 33458
rect 22542 33406 22594 33458
rect 26574 33406 26626 33458
rect 30270 33406 30322 33458
rect 33518 33406 33570 33458
rect 33966 33406 34018 33458
rect 2606 33294 2658 33346
rect 4174 33294 4226 33346
rect 6078 33294 6130 33346
rect 6302 33294 6354 33346
rect 7086 33294 7138 33346
rect 8542 33294 8594 33346
rect 15150 33294 15202 33346
rect 21870 33294 21922 33346
rect 22766 33294 22818 33346
rect 24222 33294 24274 33346
rect 25230 33294 25282 33346
rect 28254 33294 28306 33346
rect 30606 33294 30658 33346
rect 3166 33182 3218 33234
rect 7198 33182 7250 33234
rect 9326 33182 9378 33234
rect 13806 33182 13858 33234
rect 23438 33182 23490 33234
rect 23774 33182 23826 33234
rect 27358 33182 27410 33234
rect 31390 33182 31442 33234
rect 23102 33070 23154 33122
rect 24894 33070 24946 33122
rect 25566 33070 25618 33122
rect 26126 33070 26178 33122
rect 27694 33070 27746 33122
rect 35758 33406 35810 33458
rect 40014 33406 40066 33458
rect 42142 33406 42194 33458
rect 43374 33406 43426 33458
rect 44270 33406 44322 33458
rect 45166 33406 45218 33458
rect 34974 33294 35026 33346
rect 39230 33294 39282 33346
rect 42590 33294 42642 33346
rect 43262 33294 43314 33346
rect 43822 33182 43874 33234
rect 34414 33070 34466 33122
rect 34526 33070 34578 33122
rect 38894 33070 38946 33122
rect 45054 33070 45106 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4510 32734 4562 32786
rect 7310 32734 7362 32786
rect 7534 32734 7586 32786
rect 8990 32734 9042 32786
rect 9662 32734 9714 32786
rect 10558 32734 10610 32786
rect 10894 32734 10946 32786
rect 29934 32734 29986 32786
rect 32510 32734 32562 32786
rect 34526 32734 34578 32786
rect 42030 32734 42082 32786
rect 42478 32734 42530 32786
rect 2270 32622 2322 32674
rect 3166 32622 3218 32674
rect 6638 32622 6690 32674
rect 10110 32622 10162 32674
rect 12238 32622 12290 32674
rect 26014 32622 26066 32674
rect 28590 32622 28642 32674
rect 30046 32622 30098 32674
rect 30606 32622 30658 32674
rect 35870 32622 35922 32674
rect 40126 32622 40178 32674
rect 42366 32622 42418 32674
rect 43822 32622 43874 32674
rect 1710 32510 1762 32562
rect 2606 32510 2658 32562
rect 4398 32510 4450 32562
rect 6190 32510 6242 32562
rect 6302 32510 6354 32562
rect 6526 32510 6578 32562
rect 7086 32510 7138 32562
rect 7198 32510 7250 32562
rect 7422 32510 7474 32562
rect 9550 32510 9602 32562
rect 9774 32510 9826 32562
rect 10446 32510 10498 32562
rect 10670 32510 10722 32562
rect 11454 32510 11506 32562
rect 17950 32510 18002 32562
rect 25230 32510 25282 32562
rect 28478 32510 28530 32562
rect 30158 32510 30210 32562
rect 30718 32510 30770 32562
rect 31502 32510 31554 32562
rect 31838 32510 31890 32562
rect 35534 32510 35586 32562
rect 38894 32510 38946 32562
rect 39678 32510 39730 32562
rect 43038 32510 43090 32562
rect 46398 32510 46450 32562
rect 8206 32398 8258 32450
rect 14366 32398 14418 32450
rect 14814 32398 14866 32450
rect 15486 32398 15538 32450
rect 17502 32398 17554 32450
rect 18622 32398 18674 32450
rect 20750 32398 20802 32450
rect 24670 32398 24722 32450
rect 28142 32398 28194 32450
rect 33182 32398 33234 32450
rect 33742 32398 33794 32450
rect 34078 32398 34130 32450
rect 39342 32398 39394 32450
rect 45950 32398 46002 32450
rect 30494 32286 30546 32338
rect 46286 32286 46338 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 11118 31950 11170 32002
rect 11342 31950 11394 32002
rect 28254 31950 28306 32002
rect 28590 31950 28642 32002
rect 31502 31950 31554 32002
rect 38894 31950 38946 32002
rect 42590 31950 42642 32002
rect 1822 31838 1874 31890
rect 4734 31838 4786 31890
rect 11342 31838 11394 31890
rect 11678 31838 11730 31890
rect 14590 31838 14642 31890
rect 18286 31838 18338 31890
rect 18510 31838 18562 31890
rect 19966 31838 20018 31890
rect 26238 31838 26290 31890
rect 29262 31838 29314 31890
rect 30046 31838 30098 31890
rect 32734 31838 32786 31890
rect 36318 31838 36370 31890
rect 44270 31838 44322 31890
rect 45614 31838 45666 31890
rect 47742 31838 47794 31890
rect 2494 31726 2546 31778
rect 3278 31726 3330 31778
rect 3950 31726 4002 31778
rect 4398 31726 4450 31778
rect 19406 31726 19458 31778
rect 26126 31726 26178 31778
rect 26798 31726 26850 31778
rect 27470 31726 27522 31778
rect 27918 31726 27970 31778
rect 29486 31726 29538 31778
rect 30158 31726 30210 31778
rect 31054 31726 31106 31778
rect 31614 31726 31666 31778
rect 32062 31726 32114 31778
rect 33406 31726 33458 31778
rect 38670 31726 38722 31778
rect 39342 31726 39394 31778
rect 40126 31726 40178 31778
rect 41918 31726 41970 31778
rect 42702 31726 42754 31778
rect 43150 31726 43202 31778
rect 44830 31726 44882 31778
rect 2718 31614 2770 31666
rect 2942 31614 2994 31666
rect 3726 31614 3778 31666
rect 13470 31614 13522 31666
rect 17278 31614 17330 31666
rect 19182 31614 19234 31666
rect 25678 31614 25730 31666
rect 26686 31614 26738 31666
rect 28478 31614 28530 31666
rect 30942 31614 30994 31666
rect 34190 31614 34242 31666
rect 37662 31614 37714 31666
rect 38894 31614 38946 31666
rect 41806 31614 41858 31666
rect 4062 31502 4114 31554
rect 6862 31502 6914 31554
rect 13806 31502 13858 31554
rect 16942 31502 16994 31554
rect 17950 31502 18002 31554
rect 25902 31502 25954 31554
rect 26238 31502 26290 31554
rect 29934 31502 29986 31554
rect 38110 31502 38162 31554
rect 40574 31502 40626 31554
rect 41246 31502 41298 31554
rect 43710 31502 43762 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 3166 31166 3218 31218
rect 5518 31166 5570 31218
rect 6190 31166 6242 31218
rect 19070 31166 19122 31218
rect 26574 31166 26626 31218
rect 29710 31166 29762 31218
rect 30494 31166 30546 31218
rect 31278 31166 31330 31218
rect 32286 31166 32338 31218
rect 2606 31054 2658 31106
rect 2942 31054 2994 31106
rect 14142 31054 14194 31106
rect 31838 31054 31890 31106
rect 32510 31054 32562 31106
rect 33630 31054 33682 31106
rect 34638 31054 34690 31106
rect 36430 31054 36482 31106
rect 37438 31054 37490 31106
rect 43934 31054 43986 31106
rect 46398 31054 46450 31106
rect 2270 30942 2322 30994
rect 3166 30942 3218 30994
rect 4174 30942 4226 30994
rect 4622 30942 4674 30994
rect 4846 30942 4898 30994
rect 5182 30942 5234 30994
rect 5742 30942 5794 30994
rect 10670 30942 10722 30994
rect 14814 30942 14866 30994
rect 19406 30942 19458 30994
rect 20078 30942 20130 30994
rect 29150 30942 29202 30994
rect 31502 30942 31554 30994
rect 32062 30942 32114 30994
rect 33070 30942 33122 30994
rect 34750 30942 34802 30994
rect 36654 30942 36706 30994
rect 43038 30942 43090 30994
rect 43598 30942 43650 30994
rect 44382 30942 44434 30994
rect 45502 30942 45554 30994
rect 46286 30942 46338 30994
rect 4062 30830 4114 30882
rect 4734 30830 4786 30882
rect 5630 30830 5682 30882
rect 11454 30830 11506 30882
rect 12014 30830 12066 30882
rect 15374 30830 15426 30882
rect 18734 30830 18786 30882
rect 19630 30830 19682 30882
rect 20750 30830 20802 30882
rect 22878 30830 22930 30882
rect 28814 30830 28866 30882
rect 39566 30830 39618 30882
rect 41470 30830 41522 30882
rect 43374 30830 43426 30882
rect 44718 30830 44770 30882
rect 45054 30830 45106 30882
rect 2494 30718 2546 30770
rect 10558 30718 10610 30770
rect 29374 30718 29426 30770
rect 31166 30718 31218 30770
rect 32398 30718 32450 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 6414 30382 6466 30434
rect 13470 30382 13522 30434
rect 26238 30382 26290 30434
rect 29486 30382 29538 30434
rect 33966 30382 34018 30434
rect 34190 30382 34242 30434
rect 34526 30382 34578 30434
rect 34862 30382 34914 30434
rect 43150 30382 43202 30434
rect 3726 30270 3778 30322
rect 6190 30270 6242 30322
rect 7534 30270 7586 30322
rect 14478 30270 14530 30322
rect 15150 30270 15202 30322
rect 18398 30270 18450 30322
rect 19854 30270 19906 30322
rect 25230 30270 25282 30322
rect 26574 30270 26626 30322
rect 33742 30270 33794 30322
rect 40798 30270 40850 30322
rect 41246 30270 41298 30322
rect 2942 30158 2994 30210
rect 4062 30158 4114 30210
rect 5966 30158 6018 30210
rect 6302 30158 6354 30210
rect 7982 30158 8034 30210
rect 11790 30158 11842 30210
rect 13806 30158 13858 30210
rect 15598 30158 15650 30210
rect 16270 30158 16322 30210
rect 21534 30158 21586 30210
rect 22318 30158 22370 30210
rect 25902 30158 25954 30210
rect 30046 30158 30098 30210
rect 31726 30158 31778 30210
rect 35758 30158 35810 30210
rect 36206 30158 36258 30210
rect 40350 30158 40402 30210
rect 41582 30158 41634 30210
rect 42478 30158 42530 30210
rect 42814 30158 42866 30210
rect 44942 30158 44994 30210
rect 2830 30046 2882 30098
rect 4174 30046 4226 30098
rect 4958 30046 5010 30098
rect 7422 30046 7474 30098
rect 7646 30046 7698 30098
rect 10222 30046 10274 30098
rect 10670 30046 10722 30098
rect 11118 30046 11170 30098
rect 12126 30046 12178 30098
rect 14030 30046 14082 30098
rect 21310 30046 21362 30098
rect 23102 30046 23154 30098
rect 25678 30046 25730 30098
rect 30830 30046 30882 30098
rect 33518 30046 33570 30098
rect 35310 30046 35362 30098
rect 41694 30046 41746 30098
rect 9886 29934 9938 29986
rect 11006 29934 11058 29986
rect 12238 29934 12290 29986
rect 12350 29934 12402 29986
rect 12798 29934 12850 29986
rect 26126 29934 26178 29986
rect 27134 29934 27186 29986
rect 28590 29934 28642 29986
rect 32622 29934 32674 29986
rect 33294 29934 33346 29986
rect 33406 29934 33458 29986
rect 34638 29934 34690 29986
rect 37102 29934 37154 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 5630 29598 5682 29650
rect 5742 29598 5794 29650
rect 6862 29598 6914 29650
rect 6974 29598 7026 29650
rect 8206 29598 8258 29650
rect 9886 29598 9938 29650
rect 10670 29598 10722 29650
rect 20974 29598 21026 29650
rect 26462 29598 26514 29650
rect 27134 29598 27186 29650
rect 32174 29598 32226 29650
rect 33182 29598 33234 29650
rect 33630 29598 33682 29650
rect 34078 29598 34130 29650
rect 34974 29598 35026 29650
rect 35534 29598 35586 29650
rect 36654 29598 36706 29650
rect 38110 29598 38162 29650
rect 40910 29598 40962 29650
rect 41918 29598 41970 29650
rect 42366 29598 42418 29650
rect 43038 29598 43090 29650
rect 3054 29486 3106 29538
rect 7646 29486 7698 29538
rect 10558 29486 10610 29538
rect 11230 29486 11282 29538
rect 13358 29486 13410 29538
rect 16046 29486 16098 29538
rect 17390 29486 17442 29538
rect 21422 29486 21474 29538
rect 27022 29486 27074 29538
rect 29710 29486 29762 29538
rect 32398 29486 32450 29538
rect 39230 29486 39282 29538
rect 43150 29486 43202 29538
rect 45166 29486 45218 29538
rect 2270 29374 2322 29426
rect 4174 29374 4226 29426
rect 5070 29374 5122 29426
rect 5518 29374 5570 29426
rect 6414 29374 6466 29426
rect 7086 29374 7138 29426
rect 8430 29374 8482 29426
rect 8542 29374 8594 29426
rect 8654 29374 8706 29426
rect 8990 29374 9042 29426
rect 9774 29374 9826 29426
rect 10334 29374 10386 29426
rect 11006 29374 11058 29426
rect 11790 29374 11842 29426
rect 12238 29374 12290 29426
rect 12798 29374 12850 29426
rect 13246 29374 13298 29426
rect 16830 29374 16882 29426
rect 17614 29374 17666 29426
rect 20638 29374 20690 29426
rect 26014 29374 26066 29426
rect 28814 29374 28866 29426
rect 29150 29374 29202 29426
rect 31502 29374 31554 29426
rect 31950 29374 32002 29426
rect 34638 29374 34690 29426
rect 41134 29374 41186 29426
rect 41582 29374 41634 29426
rect 42926 29374 42978 29426
rect 43598 29374 43650 29426
rect 44158 29374 44210 29426
rect 44830 29374 44882 29426
rect 45502 29374 45554 29426
rect 1934 29262 1986 29314
rect 3838 29262 3890 29314
rect 5294 29262 5346 29314
rect 11902 29262 11954 29314
rect 13918 29262 13970 29314
rect 20414 29262 20466 29314
rect 21982 29262 22034 29314
rect 32174 29262 32226 29314
rect 35870 29262 35922 29314
rect 38894 29262 38946 29314
rect 41022 29262 41074 29314
rect 9886 29150 9938 29202
rect 10782 29150 10834 29202
rect 31726 29150 31778 29202
rect 39454 29150 39506 29202
rect 39790 29150 39842 29202
rect 45502 29150 45554 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 16270 28814 16322 28866
rect 16606 28814 16658 28866
rect 30158 28814 30210 28866
rect 31390 28814 31442 28866
rect 31726 28814 31778 28866
rect 33518 28814 33570 28866
rect 33966 28814 34018 28866
rect 36206 28814 36258 28866
rect 3390 28702 3442 28754
rect 6638 28702 6690 28754
rect 12686 28702 12738 28754
rect 17054 28702 17106 28754
rect 17502 28702 17554 28754
rect 24446 28702 24498 28754
rect 25902 28702 25954 28754
rect 26686 28702 26738 28754
rect 27358 28702 27410 28754
rect 27694 28702 27746 28754
rect 28254 28702 28306 28754
rect 29934 28702 29986 28754
rect 31166 28702 31218 28754
rect 31726 28702 31778 28754
rect 32622 28702 32674 28754
rect 33294 28702 33346 28754
rect 33742 28702 33794 28754
rect 38110 28702 38162 28754
rect 38446 28702 38498 28754
rect 40574 28702 40626 28754
rect 41694 28702 41746 28754
rect 42926 28702 42978 28754
rect 43374 28702 43426 28754
rect 43822 28702 43874 28754
rect 45726 28702 45778 28754
rect 47854 28702 47906 28754
rect 2942 28590 2994 28642
rect 4174 28590 4226 28642
rect 6190 28590 6242 28642
rect 6974 28590 7026 28642
rect 13582 28590 13634 28642
rect 23550 28590 23602 28642
rect 30606 28590 30658 28642
rect 34414 28590 34466 28642
rect 34862 28590 34914 28642
rect 35422 28590 35474 28642
rect 35982 28590 36034 28642
rect 36878 28590 36930 28642
rect 36990 28590 37042 28642
rect 37550 28590 37602 28642
rect 41358 28590 41410 28642
rect 41806 28590 41858 28642
rect 42254 28590 42306 28642
rect 42366 28590 42418 28642
rect 44270 28590 44322 28642
rect 44942 28590 44994 28642
rect 1934 28478 1986 28530
rect 2158 28478 2210 28530
rect 3054 28478 3106 28530
rect 11006 28478 11058 28530
rect 16046 28478 16098 28530
rect 23326 28478 23378 28530
rect 30830 28478 30882 28530
rect 31054 28478 31106 28530
rect 35310 28478 35362 28530
rect 35534 28478 35586 28530
rect 36318 28478 36370 28530
rect 2046 28366 2098 28418
rect 27806 28366 27858 28418
rect 32174 28366 32226 28418
rect 37214 28366 37266 28418
rect 37438 28366 37490 28418
rect 42030 28366 42082 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4398 28030 4450 28082
rect 5182 28030 5234 28082
rect 6302 28030 6354 28082
rect 10782 28030 10834 28082
rect 16270 28030 16322 28082
rect 16830 28030 16882 28082
rect 25678 28030 25730 28082
rect 30158 28030 30210 28082
rect 32286 28030 32338 28082
rect 33182 28030 33234 28082
rect 33630 28030 33682 28082
rect 36878 28030 36930 28082
rect 2830 27918 2882 27970
rect 3726 27918 3778 27970
rect 4734 27918 4786 27970
rect 5966 27918 6018 27970
rect 8094 27918 8146 27970
rect 8878 27918 8930 27970
rect 14142 27918 14194 27970
rect 22766 27918 22818 27970
rect 25230 27918 25282 27970
rect 25790 27918 25842 27970
rect 26574 27918 26626 27970
rect 27022 27918 27074 27970
rect 29038 27918 29090 27970
rect 30494 27918 30546 27970
rect 40014 27918 40066 27970
rect 40350 27918 40402 27970
rect 47294 27918 47346 27970
rect 2158 27806 2210 27858
rect 2718 27806 2770 27858
rect 3838 27806 3890 27858
rect 5070 27806 5122 27858
rect 5294 27806 5346 27858
rect 6302 27806 6354 27858
rect 6862 27806 6914 27858
rect 7422 27806 7474 27858
rect 7758 27806 7810 27858
rect 8766 27806 8818 27858
rect 9102 27806 9154 27858
rect 9662 27806 9714 27858
rect 10110 27806 10162 27858
rect 11118 27806 11170 27858
rect 13358 27806 13410 27858
rect 15598 27806 15650 27858
rect 17614 27806 17666 27858
rect 23438 27806 23490 27858
rect 24334 27806 24386 27858
rect 25454 27806 25506 27858
rect 27470 27806 27522 27858
rect 27694 27806 27746 27858
rect 27918 27806 27970 27858
rect 29934 27806 29986 27858
rect 35086 27806 35138 27858
rect 37550 27806 37602 27858
rect 37774 27806 37826 27858
rect 41022 27806 41074 27858
rect 3614 27694 3666 27746
rect 12014 27694 12066 27746
rect 13470 27694 13522 27746
rect 15262 27694 15314 27746
rect 18398 27694 18450 27746
rect 20526 27694 20578 27746
rect 22206 27694 22258 27746
rect 24670 27694 24722 27746
rect 26126 27694 26178 27746
rect 34414 27694 34466 27746
rect 34750 27694 34802 27746
rect 34862 27694 34914 27746
rect 35534 27694 35586 27746
rect 36430 27694 36482 27746
rect 39678 27694 39730 27746
rect 41694 27694 41746 27746
rect 43822 27694 43874 27746
rect 5294 27582 5346 27634
rect 7758 27582 7810 27634
rect 9662 27582 9714 27634
rect 37214 27582 37266 27634
rect 47182 27582 47234 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 5966 27246 6018 27298
rect 6078 27246 6130 27298
rect 6414 27246 6466 27298
rect 10222 27246 10274 27298
rect 10334 27246 10386 27298
rect 10558 27246 10610 27298
rect 10670 27246 10722 27298
rect 23550 27246 23602 27298
rect 23886 27246 23938 27298
rect 26574 27246 26626 27298
rect 27246 27246 27298 27298
rect 30270 27246 30322 27298
rect 30606 27246 30658 27298
rect 3054 27134 3106 27186
rect 4846 27134 4898 27186
rect 7422 27134 7474 27186
rect 11342 27134 11394 27186
rect 14814 27134 14866 27186
rect 23214 27134 23266 27186
rect 24110 27134 24162 27186
rect 25342 27134 25394 27186
rect 25678 27134 25730 27186
rect 26126 27134 26178 27186
rect 28254 27134 28306 27186
rect 29374 27134 29426 27186
rect 31838 27134 31890 27186
rect 32174 27134 32226 27186
rect 32622 27134 32674 27186
rect 34302 27134 34354 27186
rect 36430 27134 36482 27186
rect 36990 27134 37042 27186
rect 40574 27134 40626 27186
rect 43038 27134 43090 27186
rect 43374 27134 43426 27186
rect 2942 27022 2994 27074
rect 3950 27022 4002 27074
rect 6302 27022 6354 27074
rect 7646 27022 7698 27074
rect 21310 27022 21362 27074
rect 22206 27022 22258 27074
rect 24558 27022 24610 27074
rect 8206 26966 8258 27018
rect 25902 27022 25954 27074
rect 27806 27022 27858 27074
rect 28478 27022 28530 27074
rect 29262 27022 29314 27074
rect 29486 27022 29538 27074
rect 30830 27022 30882 27074
rect 33518 27022 33570 27074
rect 39902 27022 39954 27074
rect 43598 27022 43650 27074
rect 3278 26910 3330 26962
rect 3838 26910 3890 26962
rect 18062 26910 18114 26962
rect 18398 26910 18450 26962
rect 21422 26910 21474 26962
rect 22542 26910 22594 26962
rect 26910 26910 26962 26962
rect 29934 26910 29986 26962
rect 31278 26910 31330 26962
rect 39118 26910 39170 26962
rect 40238 26910 40290 26962
rect 40462 26910 40514 26962
rect 7758 26798 7810 26850
rect 7982 26798 8034 26850
rect 8318 26798 8370 26850
rect 8542 26798 8594 26850
rect 9214 26798 9266 26850
rect 9662 26798 9714 26850
rect 11790 26798 11842 26850
rect 22430 26798 22482 26850
rect 29710 26798 29762 26850
rect 33182 26798 33234 26850
rect 43934 26798 43986 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 2158 26462 2210 26514
rect 2606 26462 2658 26514
rect 4062 26462 4114 26514
rect 6750 26462 6802 26514
rect 8206 26462 8258 26514
rect 8878 26462 8930 26514
rect 17726 26462 17778 26514
rect 25454 26462 25506 26514
rect 26014 26462 26066 26514
rect 26686 26462 26738 26514
rect 27806 26462 27858 26514
rect 28478 26462 28530 26514
rect 37662 26462 37714 26514
rect 39902 26462 39954 26514
rect 7198 26350 7250 26402
rect 14590 26350 14642 26402
rect 15150 26350 15202 26402
rect 25566 26350 25618 26402
rect 27582 26350 27634 26402
rect 28814 26350 28866 26402
rect 29038 26350 29090 26402
rect 37326 26350 37378 26402
rect 43822 26350 43874 26402
rect 2270 26238 2322 26290
rect 3502 26238 3554 26290
rect 3726 26238 3778 26290
rect 7086 26238 7138 26290
rect 15374 26238 15426 26290
rect 21422 26238 21474 26290
rect 32286 26238 32338 26290
rect 33070 26238 33122 26290
rect 44046 26238 44098 26290
rect 3054 26126 3106 26178
rect 5630 26126 5682 26178
rect 6190 26126 6242 26178
rect 10894 26126 10946 26178
rect 18286 26126 18338 26178
rect 18734 26126 18786 26178
rect 20974 26126 21026 26178
rect 22094 26126 22146 26178
rect 24222 26126 24274 26178
rect 29150 26126 29202 26178
rect 29486 26126 29538 26178
rect 31614 26126 31666 26178
rect 35198 26126 35250 26178
rect 36654 26126 36706 26178
rect 7870 26014 7922 26066
rect 14030 26014 14082 26066
rect 18062 26014 18114 26066
rect 25454 26014 25506 26066
rect 27918 26014 27970 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 9214 25678 9266 25730
rect 9438 25678 9490 25730
rect 10446 25678 10498 25730
rect 30494 25678 30546 25730
rect 2382 25566 2434 25618
rect 8990 25566 9042 25618
rect 12574 25566 12626 25618
rect 15150 25566 15202 25618
rect 17278 25566 17330 25618
rect 20638 25566 20690 25618
rect 24558 25566 24610 25618
rect 26686 25566 26738 25618
rect 28254 25566 28306 25618
rect 29262 25566 29314 25618
rect 29710 25566 29762 25618
rect 31950 25566 32002 25618
rect 32398 25566 32450 25618
rect 45390 25566 45442 25618
rect 7982 25454 8034 25506
rect 8542 25454 8594 25506
rect 10334 25454 10386 25506
rect 11342 25454 11394 25506
rect 11678 25454 11730 25506
rect 14478 25454 14530 25506
rect 17726 25454 17778 25506
rect 23438 25454 23490 25506
rect 23886 25454 23938 25506
rect 30270 25454 30322 25506
rect 32622 25454 32674 25506
rect 45166 25454 45218 25506
rect 7870 25342 7922 25394
rect 10670 25342 10722 25394
rect 10894 25342 10946 25394
rect 11230 25342 11282 25394
rect 18510 25342 18562 25394
rect 21982 25342 22034 25394
rect 22318 25342 22370 25394
rect 30830 25342 30882 25394
rect 31166 25342 31218 25394
rect 31502 25342 31554 25394
rect 32958 25342 33010 25394
rect 8094 25230 8146 25282
rect 9326 25230 9378 25282
rect 9774 25230 9826 25282
rect 10110 25230 10162 25282
rect 14030 25230 14082 25282
rect 32846 25230 32898 25282
rect 33406 25230 33458 25282
rect 44270 25230 44322 25282
rect 44830 25230 44882 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 2942 24894 2994 24946
rect 4958 24894 5010 24946
rect 6638 24894 6690 24946
rect 7646 24894 7698 24946
rect 16494 24894 16546 24946
rect 17502 24894 17554 24946
rect 18510 24894 18562 24946
rect 29598 24894 29650 24946
rect 37214 24894 37266 24946
rect 42814 24894 42866 24946
rect 3838 24782 3890 24834
rect 4398 24782 4450 24834
rect 5630 24782 5682 24834
rect 5966 24782 6018 24834
rect 8878 24782 8930 24834
rect 10558 24782 10610 24834
rect 12798 24782 12850 24834
rect 36654 24782 36706 24834
rect 42254 24782 42306 24834
rect 43934 24782 43986 24834
rect 7422 24670 7474 24722
rect 7758 24670 7810 24722
rect 8990 24670 9042 24722
rect 9550 24670 9602 24722
rect 9774 24670 9826 24722
rect 10110 24670 10162 24722
rect 10782 24670 10834 24722
rect 11902 24670 11954 24722
rect 13246 24670 13298 24722
rect 18286 24670 18338 24722
rect 20974 24670 21026 24722
rect 22318 24670 22370 24722
rect 22990 24670 23042 24722
rect 36430 24670 36482 24722
rect 42030 24670 42082 24722
rect 43262 24670 43314 24722
rect 7198 24558 7250 24610
rect 8430 24558 8482 24610
rect 9662 24558 9714 24610
rect 13918 24558 13970 24610
rect 16046 24558 16098 24610
rect 19742 24558 19794 24610
rect 23102 24558 23154 24610
rect 24670 24558 24722 24610
rect 25454 24558 25506 24610
rect 30046 24558 30098 24610
rect 32398 24558 32450 24610
rect 46062 24558 46114 24610
rect 4622 24446 4674 24498
rect 6302 24446 6354 24498
rect 8878 24446 8930 24498
rect 20190 24446 20242 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 3950 24110 4002 24162
rect 4286 24110 4338 24162
rect 15150 24110 15202 24162
rect 21758 24110 21810 24162
rect 36990 24110 37042 24162
rect 42254 24110 42306 24162
rect 42590 24110 42642 24162
rect 2382 23998 2434 24050
rect 6750 23998 6802 24050
rect 10782 23998 10834 24050
rect 13470 23998 13522 24050
rect 15710 23998 15762 24050
rect 16830 23998 16882 24050
rect 18510 23998 18562 24050
rect 25342 23998 25394 24050
rect 27022 23998 27074 24050
rect 27694 23998 27746 24050
rect 30942 23998 30994 24050
rect 31950 23998 32002 24050
rect 32510 23998 32562 24050
rect 38558 23998 38610 24050
rect 40686 23998 40738 24050
rect 41918 23998 41970 24050
rect 42814 23998 42866 24050
rect 47742 23998 47794 24050
rect 2270 23886 2322 23938
rect 3390 23886 3442 23938
rect 6190 23886 6242 23938
rect 6526 23886 6578 23938
rect 7422 23886 7474 23938
rect 7646 23886 7698 23938
rect 7870 23886 7922 23938
rect 8542 23886 8594 23938
rect 8766 23886 8818 23938
rect 8990 23886 9042 23938
rect 9886 23886 9938 23938
rect 10894 23886 10946 23938
rect 13582 23886 13634 23938
rect 13806 23886 13858 23938
rect 14814 23886 14866 23938
rect 15486 23886 15538 23938
rect 22094 23886 22146 23938
rect 27582 23886 27634 23938
rect 27806 23886 27858 23938
rect 27918 23886 27970 23938
rect 32174 23886 32226 23938
rect 33070 23886 33122 23938
rect 41470 23886 41522 23938
rect 44270 23886 44322 23938
rect 44830 23886 44882 23938
rect 2718 23774 2770 23826
rect 3166 23774 3218 23826
rect 5070 23774 5122 23826
rect 5854 23774 5906 23826
rect 6638 23774 6690 23826
rect 8094 23774 8146 23826
rect 9214 23774 9266 23826
rect 11678 23774 11730 23826
rect 16046 23774 16098 23826
rect 16382 23774 16434 23826
rect 22318 23774 22370 23826
rect 24334 23774 24386 23826
rect 27358 23774 27410 23826
rect 37102 23774 37154 23826
rect 45614 23774 45666 23826
rect 5518 23662 5570 23714
rect 5742 23662 5794 23714
rect 6862 23662 6914 23714
rect 7310 23662 7362 23714
rect 8430 23662 8482 23714
rect 12910 23662 12962 23714
rect 22766 23662 22818 23714
rect 24894 23662 24946 23714
rect 31614 23662 31666 23714
rect 32846 23662 32898 23714
rect 38222 23662 38274 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 5070 23326 5122 23378
rect 5518 23326 5570 23378
rect 6078 23326 6130 23378
rect 6302 23326 6354 23378
rect 6414 23326 6466 23378
rect 8542 23326 8594 23378
rect 10110 23326 10162 23378
rect 15038 23326 15090 23378
rect 15486 23326 15538 23378
rect 18286 23326 18338 23378
rect 25342 23326 25394 23378
rect 25790 23326 25842 23378
rect 33182 23326 33234 23378
rect 40350 23326 40402 23378
rect 45166 23326 45218 23378
rect 6638 23214 6690 23266
rect 6750 23214 6802 23266
rect 7310 23214 7362 23266
rect 8766 23214 8818 23266
rect 19630 23214 19682 23266
rect 22206 23214 22258 23266
rect 22990 23214 23042 23266
rect 27806 23214 27858 23266
rect 31278 23214 31330 23266
rect 43038 23214 43090 23266
rect 1822 23102 1874 23154
rect 5406 23102 5458 23154
rect 5966 23102 6018 23154
rect 7422 23102 7474 23154
rect 7534 23102 7586 23154
rect 7982 23102 8034 23154
rect 8878 23102 8930 23154
rect 10334 23102 10386 23154
rect 10446 23102 10498 23154
rect 10670 23102 10722 23154
rect 10894 23102 10946 23154
rect 11230 23102 11282 23154
rect 12126 23102 12178 23154
rect 12574 23102 12626 23154
rect 17950 23102 18002 23154
rect 22766 23102 22818 23154
rect 24670 23102 24722 23154
rect 25118 23102 25170 23154
rect 25454 23102 25506 23154
rect 27022 23102 27074 23154
rect 30382 23102 30434 23154
rect 30606 23102 30658 23154
rect 34302 23102 34354 23154
rect 34750 23102 34802 23154
rect 43710 23102 43762 23154
rect 44942 23102 44994 23154
rect 2494 22990 2546 23042
rect 4622 22990 4674 23042
rect 4958 22990 5010 23042
rect 8318 22990 8370 23042
rect 9774 22990 9826 23042
rect 13134 22990 13186 23042
rect 14478 22990 14530 23042
rect 17726 22990 17778 23042
rect 19182 22990 19234 23042
rect 20974 22990 21026 23042
rect 25902 22990 25954 23042
rect 26686 22990 26738 23042
rect 29934 22990 29986 23042
rect 32174 22990 32226 23042
rect 35422 22990 35474 23042
rect 37550 22990 37602 23042
rect 40910 22990 40962 23042
rect 5518 22878 5570 22930
rect 14702 22878 14754 22930
rect 18622 22878 18674 22930
rect 18958 22878 19010 22930
rect 24558 22878 24610 22930
rect 30942 22878 30994 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 4510 22542 4562 22594
rect 16942 22542 16994 22594
rect 22206 22542 22258 22594
rect 5742 22430 5794 22482
rect 9774 22430 9826 22482
rect 10222 22430 10274 22482
rect 17502 22430 17554 22482
rect 21422 22430 21474 22482
rect 21982 22430 22034 22482
rect 25342 22430 25394 22482
rect 26798 22430 26850 22482
rect 28254 22430 28306 22482
rect 32510 22430 32562 22482
rect 34638 22430 34690 22482
rect 37774 22430 37826 22482
rect 39902 22430 39954 22482
rect 40350 22430 40402 22482
rect 2158 22318 2210 22370
rect 7870 22318 7922 22370
rect 8206 22318 8258 22370
rect 10894 22318 10946 22370
rect 11678 22318 11730 22370
rect 11902 22318 11954 22370
rect 17614 22318 17666 22370
rect 18958 22318 19010 22370
rect 19966 22318 20018 22370
rect 20526 22318 20578 22370
rect 23102 22318 23154 22370
rect 23886 22318 23938 22370
rect 26126 22318 26178 22370
rect 28030 22318 28082 22370
rect 31054 22318 31106 22370
rect 31726 22318 31778 22370
rect 35086 22318 35138 22370
rect 35982 22318 36034 22370
rect 37102 22318 37154 22370
rect 27246 22206 27298 22258
rect 35758 22206 35810 22258
rect 7982 22094 8034 22146
rect 11118 22094 11170 22146
rect 27694 22094 27746 22146
rect 29262 22094 29314 22146
rect 31390 22094 31442 22146
rect 40238 22094 40290 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 2046 21758 2098 21810
rect 2270 21758 2322 21810
rect 9550 21758 9602 21810
rect 11230 21758 11282 21810
rect 12798 21758 12850 21810
rect 24222 21758 24274 21810
rect 24670 21758 24722 21810
rect 30382 21758 30434 21810
rect 31950 21758 32002 21810
rect 38110 21758 38162 21810
rect 39230 21758 39282 21810
rect 1710 21646 1762 21698
rect 2494 21646 2546 21698
rect 2606 21646 2658 21698
rect 11566 21646 11618 21698
rect 17390 21646 17442 21698
rect 17726 21646 17778 21698
rect 35086 21646 35138 21698
rect 42254 21646 42306 21698
rect 3054 21534 3106 21586
rect 9774 21534 9826 21586
rect 12126 21534 12178 21586
rect 19518 21534 19570 21586
rect 20862 21534 20914 21586
rect 22430 21534 22482 21586
rect 25230 21534 25282 21586
rect 30494 21534 30546 21586
rect 30830 21534 30882 21586
rect 31502 21534 31554 21586
rect 34190 21534 34242 21586
rect 36542 21534 36594 21586
rect 36878 21534 36930 21586
rect 38334 21534 38386 21586
rect 41918 21534 41970 21586
rect 42478 21534 42530 21586
rect 11902 21422 11954 21474
rect 14254 21422 14306 21474
rect 18622 21422 18674 21474
rect 21646 21422 21698 21474
rect 23438 21422 23490 21474
rect 23886 21422 23938 21474
rect 26014 21422 26066 21474
rect 28142 21422 28194 21474
rect 38782 21422 38834 21474
rect 18510 21310 18562 21362
rect 42814 21310 42866 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 8206 20974 8258 21026
rect 8766 20974 8818 21026
rect 13694 20974 13746 21026
rect 30718 20974 30770 21026
rect 35870 20974 35922 21026
rect 39230 20974 39282 21026
rect 1822 20862 1874 20914
rect 3838 20862 3890 20914
rect 9326 20862 9378 20914
rect 16382 20862 16434 20914
rect 18510 20862 18562 20914
rect 23102 20862 23154 20914
rect 23886 20862 23938 20914
rect 24894 20862 24946 20914
rect 27022 20862 27074 20914
rect 30494 20862 30546 20914
rect 32286 20862 32338 20914
rect 34414 20862 34466 20914
rect 37214 20862 37266 20914
rect 38222 20862 38274 20914
rect 40238 20862 40290 20914
rect 13470 20750 13522 20802
rect 14030 20750 14082 20802
rect 14590 20750 14642 20802
rect 15262 20750 15314 20802
rect 15598 20750 15650 20802
rect 22878 20750 22930 20802
rect 24110 20750 24162 20802
rect 27918 20750 27970 20802
rect 29374 20750 29426 20802
rect 31614 20750 31666 20802
rect 36206 20750 36258 20802
rect 36430 20750 36482 20802
rect 38894 20750 38946 20802
rect 39454 20750 39506 20802
rect 40126 20750 40178 20802
rect 42814 20750 42866 20802
rect 8094 20638 8146 20690
rect 8878 20638 8930 20690
rect 22206 20638 22258 20690
rect 22542 20638 22594 20690
rect 29486 20638 29538 20690
rect 30830 20638 30882 20690
rect 4286 20526 4338 20578
rect 8206 20526 8258 20578
rect 14366 20526 14418 20578
rect 27694 20526 27746 20578
rect 37550 20526 37602 20578
rect 42478 20526 42530 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 2158 20190 2210 20242
rect 22878 20190 22930 20242
rect 30270 20190 30322 20242
rect 31166 20190 31218 20242
rect 32174 20190 32226 20242
rect 39454 20190 39506 20242
rect 2382 20078 2434 20130
rect 3054 20078 3106 20130
rect 3278 20078 3330 20130
rect 5742 20078 5794 20130
rect 13694 20078 13746 20130
rect 23550 20078 23602 20130
rect 27694 20078 27746 20130
rect 35534 20078 35586 20130
rect 42478 20078 42530 20130
rect 2830 19966 2882 20018
rect 3390 19966 3442 20018
rect 8990 19966 9042 20018
rect 12574 19966 12626 20018
rect 13022 19966 13074 20018
rect 16382 19966 16434 20018
rect 19070 19966 19122 20018
rect 19294 19966 19346 20018
rect 23214 19966 23266 20018
rect 23998 19966 24050 20018
rect 26910 19966 26962 20018
rect 34862 19966 34914 20018
rect 35086 19966 35138 20018
rect 38894 19966 38946 20018
rect 39230 19966 39282 20018
rect 41806 19966 41858 20018
rect 9662 19854 9714 19906
rect 11790 19854 11842 19906
rect 15822 19854 15874 19906
rect 20078 19854 20130 19906
rect 22206 19854 22258 19906
rect 26574 19854 26626 19906
rect 29822 19854 29874 19906
rect 30158 19854 30210 19906
rect 31614 19854 31666 19906
rect 38446 19854 38498 19906
rect 39454 19854 39506 19906
rect 41358 19854 41410 19906
rect 44606 19854 44658 19906
rect 34526 19742 34578 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 6078 19406 6130 19458
rect 7982 19406 8034 19458
rect 22878 19406 22930 19458
rect 27022 19406 27074 19458
rect 45054 19406 45106 19458
rect 4846 19294 4898 19346
rect 8878 19294 8930 19346
rect 12798 19294 12850 19346
rect 24334 19294 24386 19346
rect 25454 19294 25506 19346
rect 39454 19294 39506 19346
rect 41582 19294 41634 19346
rect 43822 19294 43874 19346
rect 44382 19294 44434 19346
rect 44830 19294 44882 19346
rect 3950 19182 4002 19234
rect 7422 19182 7474 19234
rect 7646 19182 7698 19234
rect 8430 19182 8482 19234
rect 11342 19182 11394 19234
rect 23214 19182 23266 19234
rect 23886 19182 23938 19234
rect 24782 19182 24834 19234
rect 34974 19182 35026 19234
rect 38670 19182 38722 19234
rect 2270 19070 2322 19122
rect 2382 19070 2434 19122
rect 2830 19070 2882 19122
rect 3166 19070 3218 19122
rect 3390 19070 3442 19122
rect 3502 19070 3554 19122
rect 4062 19070 4114 19122
rect 5966 19070 6018 19122
rect 6526 19070 6578 19122
rect 11566 19070 11618 19122
rect 19966 19070 20018 19122
rect 20302 19070 20354 19122
rect 23438 19070 23490 19122
rect 27134 19070 27186 19122
rect 2046 18958 2098 19010
rect 2606 18958 2658 19010
rect 2942 18958 2994 19010
rect 3726 18958 3778 19010
rect 6078 18958 6130 19010
rect 6638 18958 6690 19010
rect 6862 18958 6914 19010
rect 8766 18958 8818 19010
rect 8990 18958 9042 19010
rect 25006 18958 25058 19010
rect 34750 18958 34802 19010
rect 38334 18958 38386 19010
rect 45390 18958 45442 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 6414 18622 6466 18674
rect 7422 18622 7474 18674
rect 8654 18622 8706 18674
rect 11342 18622 11394 18674
rect 17726 18622 17778 18674
rect 23214 18622 23266 18674
rect 23886 18622 23938 18674
rect 2494 18510 2546 18562
rect 5406 18510 5458 18562
rect 7758 18510 7810 18562
rect 8542 18510 8594 18562
rect 9662 18510 9714 18562
rect 15934 18510 15986 18562
rect 24446 18510 24498 18562
rect 41022 18510 41074 18562
rect 44158 18510 44210 18562
rect 1822 18398 1874 18450
rect 5630 18398 5682 18450
rect 5742 18398 5794 18450
rect 5854 18398 5906 18450
rect 6302 18398 6354 18450
rect 6526 18398 6578 18450
rect 6974 18398 7026 18450
rect 7198 18398 7250 18450
rect 7534 18398 7586 18450
rect 8206 18398 8258 18450
rect 9438 18398 9490 18450
rect 9774 18398 9826 18450
rect 11006 18398 11058 18450
rect 11790 18398 11842 18450
rect 16158 18398 16210 18450
rect 18062 18398 18114 18450
rect 18734 18398 18786 18450
rect 19966 18398 20018 18450
rect 23550 18398 23602 18450
rect 24110 18398 24162 18450
rect 25230 18398 25282 18450
rect 26014 18398 26066 18450
rect 32398 18398 32450 18450
rect 39790 18398 39842 18450
rect 40350 18398 40402 18450
rect 44494 18398 44546 18450
rect 4622 18286 4674 18338
rect 10782 18286 10834 18338
rect 18286 18286 18338 18338
rect 20414 18286 20466 18338
rect 28142 18286 28194 18338
rect 29598 18286 29650 18338
rect 31726 18286 31778 18338
rect 33182 18286 33234 18338
rect 36654 18286 36706 18338
rect 36990 18286 37042 18338
rect 39118 18286 39170 18338
rect 8094 18174 8146 18226
rect 8654 18174 8706 18226
rect 40910 18174 40962 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 7422 17838 7474 17890
rect 8878 17838 8930 17890
rect 9326 17838 9378 17890
rect 20078 17838 20130 17890
rect 24782 17838 24834 17890
rect 25118 17838 25170 17890
rect 26238 17838 26290 17890
rect 37886 17838 37938 17890
rect 45278 17838 45330 17890
rect 4622 17726 4674 17778
rect 5742 17726 5794 17778
rect 15822 17726 15874 17778
rect 17950 17726 18002 17778
rect 24222 17726 24274 17778
rect 26462 17726 26514 17778
rect 33182 17726 33234 17778
rect 34302 17726 34354 17778
rect 36430 17726 36482 17778
rect 37326 17726 37378 17778
rect 1710 17614 1762 17666
rect 2270 17614 2322 17666
rect 3950 17614 4002 17666
rect 5182 17614 5234 17666
rect 6078 17614 6130 17666
rect 7534 17614 7586 17666
rect 7870 17614 7922 17666
rect 8318 17614 8370 17666
rect 8542 17614 8594 17666
rect 15150 17614 15202 17666
rect 18846 17614 18898 17666
rect 19182 17614 19234 17666
rect 20414 17614 20466 17666
rect 20638 17614 20690 17666
rect 21310 17614 21362 17666
rect 33518 17614 33570 17666
rect 37662 17614 37714 17666
rect 39342 17614 39394 17666
rect 39902 17614 39954 17666
rect 40574 17614 40626 17666
rect 41022 17614 41074 17666
rect 2046 17502 2098 17554
rect 2606 17502 2658 17554
rect 2830 17502 2882 17554
rect 3502 17502 3554 17554
rect 3726 17502 3778 17554
rect 4846 17502 4898 17554
rect 6302 17502 6354 17554
rect 6638 17502 6690 17554
rect 7310 17502 7362 17554
rect 9214 17502 9266 17554
rect 18734 17502 18786 17554
rect 22094 17502 22146 17554
rect 24558 17502 24610 17554
rect 29150 17502 29202 17554
rect 29934 17502 29986 17554
rect 31054 17502 31106 17554
rect 31390 17502 31442 17554
rect 38222 17502 38274 17554
rect 38558 17502 38610 17554
rect 38894 17502 38946 17554
rect 39678 17502 39730 17554
rect 45390 17502 45442 17554
rect 2494 17390 2546 17442
rect 4958 17390 5010 17442
rect 7758 17390 7810 17442
rect 9326 17390 9378 17442
rect 14702 17390 14754 17442
rect 19406 17390 19458 17442
rect 19518 17390 19570 17442
rect 25566 17390 25618 17442
rect 25902 17390 25954 17442
rect 26910 17390 26962 17442
rect 27358 17390 27410 17442
rect 28590 17390 28642 17442
rect 41470 17390 41522 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 1822 17054 1874 17106
rect 5406 17054 5458 17106
rect 7198 17054 7250 17106
rect 7758 17054 7810 17106
rect 7982 17054 8034 17106
rect 15262 17054 15314 17106
rect 15934 17054 15986 17106
rect 19182 17054 19234 17106
rect 19294 17054 19346 17106
rect 20190 17054 20242 17106
rect 21646 17054 21698 17106
rect 30270 17054 30322 17106
rect 30494 17054 30546 17106
rect 31054 17054 31106 17106
rect 32062 17054 32114 17106
rect 33294 17054 33346 17106
rect 34078 17054 34130 17106
rect 35198 17054 35250 17106
rect 35646 17054 35698 17106
rect 38782 17054 38834 17106
rect 41918 17054 41970 17106
rect 5294 16942 5346 16994
rect 5854 16942 5906 16994
rect 6078 16942 6130 16994
rect 14478 16942 14530 16994
rect 14814 16942 14866 16994
rect 18398 16942 18450 16994
rect 20974 16942 21026 16994
rect 28814 16942 28866 16994
rect 29710 16942 29762 16994
rect 33518 16942 33570 16994
rect 33630 16942 33682 16994
rect 36206 16942 36258 16994
rect 44158 16942 44210 16994
rect 5742 16830 5794 16882
rect 6302 16830 6354 16882
rect 6638 16830 6690 16882
rect 6862 16830 6914 16882
rect 7534 16830 7586 16882
rect 11902 16830 11954 16882
rect 14142 16830 14194 16882
rect 17838 16830 17890 16882
rect 18622 16830 18674 16882
rect 18958 16830 19010 16882
rect 21422 16830 21474 16882
rect 24670 16830 24722 16882
rect 28030 16830 28082 16882
rect 30606 16830 30658 16882
rect 36542 16830 36594 16882
rect 38558 16830 38610 16882
rect 38894 16830 38946 16882
rect 39790 16830 39842 16882
rect 41806 16830 41858 16882
rect 42142 16830 42194 16882
rect 43486 16830 43538 16882
rect 8094 16718 8146 16770
rect 11454 16718 11506 16770
rect 16270 16718 16322 16770
rect 16494 16718 16546 16770
rect 22094 16718 22146 16770
rect 25230 16718 25282 16770
rect 27358 16718 27410 16770
rect 31614 16718 31666 16770
rect 41022 16718 41074 16770
rect 41470 16718 41522 16770
rect 43038 16718 43090 16770
rect 46286 16718 46338 16770
rect 11566 16606 11618 16658
rect 29150 16606 29202 16658
rect 29486 16606 29538 16658
rect 31390 16606 31442 16658
rect 41022 16606 41074 16658
rect 41470 16606 41522 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 21534 16270 21586 16322
rect 21870 16270 21922 16322
rect 30830 16270 30882 16322
rect 31166 16270 31218 16322
rect 31390 16270 31442 16322
rect 43710 16270 43762 16322
rect 5742 16158 5794 16210
rect 11006 16158 11058 16210
rect 14254 16158 14306 16210
rect 16382 16158 16434 16210
rect 16830 16158 16882 16210
rect 19294 16158 19346 16210
rect 22542 16158 22594 16210
rect 22990 16158 23042 16210
rect 29710 16158 29762 16210
rect 30270 16158 30322 16210
rect 31390 16158 31442 16210
rect 33518 16158 33570 16210
rect 36206 16158 36258 16210
rect 5630 16046 5682 16098
rect 11118 16046 11170 16098
rect 13582 16046 13634 16098
rect 17838 16046 17890 16098
rect 18174 16046 18226 16098
rect 19742 16046 19794 16098
rect 22094 16046 22146 16098
rect 29486 16046 29538 16098
rect 30942 16046 30994 16098
rect 33742 16046 33794 16098
rect 34078 16046 34130 16098
rect 34974 16046 35026 16098
rect 35198 16046 35250 16098
rect 35870 16046 35922 16098
rect 37102 16046 37154 16098
rect 39342 16046 39394 16098
rect 39678 16046 39730 16098
rect 40462 16046 40514 16098
rect 41470 16046 41522 16098
rect 5966 15934 6018 15986
rect 6190 15934 6242 15986
rect 11790 15934 11842 15986
rect 17278 15934 17330 15986
rect 19966 15934 20018 15986
rect 20414 15934 20466 15986
rect 33966 15934 34018 15986
rect 35982 15934 36034 15986
rect 36990 15934 37042 15986
rect 39230 15934 39282 15986
rect 41582 15934 41634 15986
rect 43822 15934 43874 15986
rect 18398 15822 18450 15874
rect 18622 15822 18674 15874
rect 20638 15822 20690 15874
rect 29150 15822 29202 15874
rect 30830 15822 30882 15874
rect 42030 15822 42082 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 12798 15486 12850 15538
rect 16606 15486 16658 15538
rect 18622 15486 18674 15538
rect 19070 15486 19122 15538
rect 23998 15486 24050 15538
rect 29934 15486 29986 15538
rect 34078 15486 34130 15538
rect 34526 15486 34578 15538
rect 37550 15486 37602 15538
rect 39790 15486 39842 15538
rect 41134 15486 41186 15538
rect 3166 15374 3218 15426
rect 10670 15374 10722 15426
rect 20750 15374 20802 15426
rect 21870 15374 21922 15426
rect 28254 15374 28306 15426
rect 33406 15374 33458 15426
rect 35646 15374 35698 15426
rect 40014 15374 40066 15426
rect 40126 15374 40178 15426
rect 41022 15374 41074 15426
rect 42366 15374 42418 15426
rect 3278 15262 3330 15314
rect 9774 15262 9826 15314
rect 10558 15262 10610 15314
rect 11118 15262 11170 15314
rect 11342 15262 11394 15314
rect 12014 15262 12066 15314
rect 20862 15262 20914 15314
rect 22542 15262 22594 15314
rect 28590 15262 28642 15314
rect 33182 15262 33234 15314
rect 35310 15262 35362 15314
rect 36654 15262 36706 15314
rect 37662 15262 37714 15314
rect 38446 15262 38498 15314
rect 41358 15262 41410 15314
rect 41582 15262 41634 15314
rect 3614 15150 3666 15202
rect 9998 15150 10050 15202
rect 22430 15150 22482 15202
rect 31166 15150 31218 15202
rect 44494 15150 44546 15202
rect 3502 15038 3554 15090
rect 11902 15038 11954 15090
rect 40126 15038 40178 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 12574 14702 12626 14754
rect 20414 14702 20466 14754
rect 20638 14702 20690 14754
rect 2046 14590 2098 14642
rect 2830 14590 2882 14642
rect 9998 14590 10050 14642
rect 11454 14590 11506 14642
rect 14030 14590 14082 14642
rect 15934 14590 15986 14642
rect 19742 14590 19794 14642
rect 20190 14590 20242 14642
rect 20638 14590 20690 14642
rect 24894 14590 24946 14642
rect 28702 14590 28754 14642
rect 31502 14590 31554 14642
rect 33630 14590 33682 14642
rect 34974 14590 35026 14642
rect 35422 14590 35474 14642
rect 36542 14590 36594 14642
rect 37214 14590 37266 14642
rect 38446 14590 38498 14642
rect 40126 14590 40178 14642
rect 42254 14590 42306 14642
rect 2270 14478 2322 14530
rect 3166 14478 3218 14530
rect 9886 14478 9938 14530
rect 11902 14478 11954 14530
rect 14926 14478 14978 14530
rect 19070 14478 19122 14530
rect 22430 14478 22482 14530
rect 23326 14478 23378 14530
rect 24334 14478 24386 14530
rect 29262 14478 29314 14530
rect 30158 14478 30210 14530
rect 30382 14478 30434 14530
rect 34414 14478 34466 14530
rect 39006 14478 39058 14530
rect 39454 14478 39506 14530
rect 3838 14366 3890 14418
rect 12798 14366 12850 14418
rect 18062 14366 18114 14418
rect 18846 14366 18898 14418
rect 19182 14366 19234 14418
rect 22542 14366 22594 14418
rect 23550 14366 23602 14418
rect 29374 14366 29426 14418
rect 30830 14366 30882 14418
rect 42926 14366 42978 14418
rect 1710 14254 1762 14306
rect 3278 14254 3330 14306
rect 3726 14254 3778 14306
rect 4846 14254 4898 14306
rect 12686 14254 12738 14306
rect 13582 14254 13634 14306
rect 17390 14254 17442 14306
rect 22654 14254 22706 14306
rect 24110 14254 24162 14306
rect 29598 14254 29650 14306
rect 29822 14254 29874 14306
rect 37998 14254 38050 14306
rect 42814 14254 42866 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 5070 13918 5122 13970
rect 5518 13918 5570 13970
rect 5630 13918 5682 13970
rect 5742 13918 5794 13970
rect 10446 13918 10498 13970
rect 13022 13918 13074 13970
rect 22542 13918 22594 13970
rect 22654 13918 22706 13970
rect 24222 13918 24274 13970
rect 24670 13918 24722 13970
rect 30606 13918 30658 13970
rect 33630 13918 33682 13970
rect 37886 13918 37938 13970
rect 6078 13806 6130 13858
rect 5182 13750 5234 13802
rect 1822 13694 1874 13746
rect 6862 13750 6914 13802
rect 10222 13806 10274 13858
rect 11230 13806 11282 13858
rect 12238 13806 12290 13858
rect 13470 13806 13522 13858
rect 20190 13806 20242 13858
rect 21086 13806 21138 13858
rect 23326 13806 23378 13858
rect 27806 13806 27858 13858
rect 30494 13806 30546 13858
rect 31614 13806 31666 13858
rect 39006 13806 39058 13858
rect 41694 13806 41746 13858
rect 5966 13694 6018 13746
rect 12574 13694 12626 13746
rect 12910 13694 12962 13746
rect 13918 13694 13970 13746
rect 17726 13694 17778 13746
rect 17950 13694 18002 13746
rect 18846 13694 18898 13746
rect 21758 13694 21810 13746
rect 22318 13694 22370 13746
rect 23438 13694 23490 13746
rect 27134 13694 27186 13746
rect 30270 13694 30322 13746
rect 31278 13694 31330 13746
rect 33294 13694 33346 13746
rect 34078 13694 34130 13746
rect 36878 13694 36930 13746
rect 37102 13694 37154 13746
rect 38670 13694 38722 13746
rect 39118 13694 39170 13746
rect 39902 13694 39954 13746
rect 40910 13694 40962 13746
rect 2494 13582 2546 13634
rect 4622 13582 4674 13634
rect 9662 13582 9714 13634
rect 10334 13582 10386 13634
rect 11566 13582 11618 13634
rect 11902 13582 11954 13634
rect 14702 13582 14754 13634
rect 16830 13582 16882 13634
rect 18398 13582 18450 13634
rect 20526 13582 20578 13634
rect 26686 13582 26738 13634
rect 29934 13582 29986 13634
rect 31390 13582 31442 13634
rect 33070 13582 33122 13634
rect 40238 13582 40290 13634
rect 43822 13582 43874 13634
rect 6974 13470 7026 13522
rect 9550 13470 9602 13522
rect 13022 13470 13074 13522
rect 13582 13470 13634 13522
rect 17390 13470 17442 13522
rect 37438 13470 37490 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 5070 13134 5122 13186
rect 5966 13134 6018 13186
rect 12462 13134 12514 13186
rect 30942 13134 30994 13186
rect 31614 13134 31666 13186
rect 35982 13134 36034 13186
rect 3390 13022 3442 13074
rect 6862 13022 6914 13074
rect 11678 13022 11730 13074
rect 14702 13022 14754 13074
rect 16830 13022 16882 13074
rect 17054 13022 17106 13074
rect 19518 13022 19570 13074
rect 22542 13022 22594 13074
rect 24670 13022 24722 13074
rect 25118 13022 25170 13074
rect 33406 13022 33458 13074
rect 34078 13022 34130 13074
rect 34302 13022 34354 13074
rect 35646 13022 35698 13074
rect 39902 13022 39954 13074
rect 40574 13022 40626 13074
rect 3278 12910 3330 12962
rect 3502 12910 3554 12962
rect 4286 12910 4338 12962
rect 4958 12910 5010 12962
rect 6078 12910 6130 12962
rect 6302 12910 6354 12962
rect 8654 12910 8706 12962
rect 9326 12910 9378 12962
rect 10110 12910 10162 12962
rect 10446 12910 10498 12962
rect 11342 12910 11394 12962
rect 12238 12910 12290 12962
rect 14254 12910 14306 12962
rect 15374 12910 15426 12962
rect 17614 12910 17666 12962
rect 20078 12910 20130 12962
rect 21870 12910 21922 12962
rect 25790 12910 25842 12962
rect 29374 12910 29426 12962
rect 31726 12910 31778 12962
rect 32174 12910 32226 12962
rect 36094 12910 36146 12962
rect 36990 12910 37042 12962
rect 1710 12798 1762 12850
rect 2494 12798 2546 12850
rect 3726 12798 3778 12850
rect 7310 12798 7362 12850
rect 9438 12798 9490 12850
rect 11902 12798 11954 12850
rect 15038 12798 15090 12850
rect 16046 12798 16098 12850
rect 16494 12798 16546 12850
rect 18958 12798 19010 12850
rect 19854 12798 19906 12850
rect 29934 12798 29986 12850
rect 31614 12798 31666 12850
rect 37774 12798 37826 12850
rect 4846 12686 4898 12738
rect 5966 12686 6018 12738
rect 7870 12686 7922 12738
rect 8318 12686 8370 12738
rect 9886 12686 9938 12738
rect 9998 12686 10050 12738
rect 12798 12686 12850 12738
rect 13806 12686 13858 12738
rect 15710 12686 15762 12738
rect 21422 12686 21474 12738
rect 26014 12686 26066 12738
rect 28590 12686 28642 12738
rect 29598 12686 29650 12738
rect 33742 12686 33794 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 1822 12350 1874 12402
rect 4510 12350 4562 12402
rect 5966 12350 6018 12402
rect 10670 12350 10722 12402
rect 15598 12350 15650 12402
rect 16830 12350 16882 12402
rect 23998 12350 24050 12402
rect 37550 12350 37602 12402
rect 4286 12238 4338 12290
rect 9550 12238 9602 12290
rect 12574 12238 12626 12290
rect 17726 12238 17778 12290
rect 18510 12238 18562 12290
rect 18846 12238 18898 12290
rect 23326 12238 23378 12290
rect 24446 12238 24498 12290
rect 27358 12238 27410 12290
rect 28478 12238 28530 12290
rect 28814 12238 28866 12290
rect 30382 12238 30434 12290
rect 4734 12126 4786 12178
rect 5182 12126 5234 12178
rect 5854 12126 5906 12178
rect 6862 12126 6914 12178
rect 8094 12126 8146 12178
rect 8990 12126 9042 12178
rect 9998 12126 10050 12178
rect 11566 12126 11618 12178
rect 12910 12126 12962 12178
rect 14142 12126 14194 12178
rect 15262 12126 15314 12178
rect 18622 12126 18674 12178
rect 19070 12126 19122 12178
rect 23102 12126 23154 12178
rect 24558 12126 24610 12178
rect 28030 12126 28082 12178
rect 29710 12126 29762 12178
rect 33182 12126 33234 12178
rect 33742 12126 33794 12178
rect 37326 12126 37378 12178
rect 4622 12014 4674 12066
rect 5070 12014 5122 12066
rect 7198 12014 7250 12066
rect 10222 12014 10274 12066
rect 11678 12014 11730 12066
rect 12014 12014 12066 12066
rect 13694 12014 13746 12066
rect 19854 12014 19906 12066
rect 21982 12014 22034 12066
rect 25230 12014 25282 12066
rect 32510 12014 32562 12066
rect 34526 12014 34578 12066
rect 36654 12014 36706 12066
rect 5630 11902 5682 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 6526 11566 6578 11618
rect 8094 11566 8146 11618
rect 18510 11566 18562 11618
rect 19742 11566 19794 11618
rect 23662 11566 23714 11618
rect 4846 11454 4898 11506
rect 5070 11454 5122 11506
rect 5742 11454 5794 11506
rect 6862 11454 6914 11506
rect 7758 11454 7810 11506
rect 8654 11454 8706 11506
rect 9326 11454 9378 11506
rect 11342 11454 11394 11506
rect 14142 11454 14194 11506
rect 15262 11454 15314 11506
rect 17390 11454 17442 11506
rect 17838 11454 17890 11506
rect 18734 11454 18786 11506
rect 19182 11454 19234 11506
rect 19742 11454 19794 11506
rect 21870 11454 21922 11506
rect 24670 11454 24722 11506
rect 25118 11454 25170 11506
rect 25454 11454 25506 11506
rect 27582 11454 27634 11506
rect 33406 11454 33458 11506
rect 35086 11454 35138 11506
rect 5518 11342 5570 11394
rect 5854 11342 5906 11394
rect 6190 11342 6242 11394
rect 6638 11342 6690 11394
rect 6974 11342 7026 11394
rect 8318 11342 8370 11394
rect 8542 11342 8594 11394
rect 11454 11342 11506 11394
rect 12238 11342 12290 11394
rect 14478 11342 14530 11394
rect 21646 11342 21698 11394
rect 23102 11342 23154 11394
rect 23326 11342 23378 11394
rect 24110 11342 24162 11394
rect 28254 11342 28306 11394
rect 33966 11342 34018 11394
rect 35310 11342 35362 11394
rect 39454 11342 39506 11394
rect 4846 11230 4898 11282
rect 8766 11230 8818 11282
rect 11230 11230 11282 11282
rect 13470 11230 13522 11282
rect 20190 11230 20242 11282
rect 20526 11230 20578 11282
rect 21310 11230 21362 11282
rect 34974 11230 35026 11282
rect 39566 11230 39618 11282
rect 10782 11118 10834 11170
rect 12910 11118 12962 11170
rect 13582 11118 13634 11170
rect 13806 11118 13858 11170
rect 22766 11118 22818 11170
rect 34302 11118 34354 11170
rect 40014 11118 40066 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 3390 10782 3442 10834
rect 3950 10782 4002 10834
rect 5966 10782 6018 10834
rect 10334 10782 10386 10834
rect 17614 10782 17666 10834
rect 30158 10782 30210 10834
rect 31166 10782 31218 10834
rect 31950 10782 32002 10834
rect 38558 10782 38610 10834
rect 39118 10782 39170 10834
rect 40910 10782 40962 10834
rect 34638 10670 34690 10722
rect 38894 10670 38946 10722
rect 39790 10670 39842 10722
rect 2718 10558 2770 10610
rect 3502 10558 3554 10610
rect 6078 10558 6130 10610
rect 10782 10558 10834 10610
rect 12126 10558 12178 10610
rect 12574 10558 12626 10610
rect 13582 10558 13634 10610
rect 14254 10558 14306 10610
rect 40126 10558 40178 10610
rect 2046 10446 2098 10498
rect 2942 10446 2994 10498
rect 13358 10446 13410 10498
rect 16606 10446 16658 10498
rect 20974 10446 21026 10498
rect 39006 10446 39058 10498
rect 41022 10446 41074 10498
rect 11230 10334 11282 10386
rect 40126 10334 40178 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 29934 9998 29986 10050
rect 31054 9998 31106 10050
rect 31166 9998 31218 10050
rect 33294 9998 33346 10050
rect 3054 9886 3106 9938
rect 6750 9886 6802 9938
rect 9550 9886 9602 9938
rect 15262 9886 15314 9938
rect 16830 9886 16882 9938
rect 17278 9886 17330 9938
rect 21870 9886 21922 9938
rect 23550 9886 23602 9938
rect 24222 9886 24274 9938
rect 24446 9886 24498 9938
rect 33854 9886 33906 9938
rect 38446 9886 38498 9938
rect 40574 9886 40626 9938
rect 40910 9886 40962 9938
rect 43038 9886 43090 9938
rect 2382 9774 2434 9826
rect 10110 9774 10162 9826
rect 10558 9774 10610 9826
rect 11566 9774 11618 9826
rect 11902 9774 11954 9826
rect 12462 9774 12514 9826
rect 13582 9774 13634 9826
rect 21646 9774 21698 9826
rect 29374 9774 29426 9826
rect 30494 9774 30546 9826
rect 31726 9774 31778 9826
rect 32510 9774 32562 9826
rect 37662 9774 37714 9826
rect 43710 9774 43762 9826
rect 2494 9662 2546 9714
rect 12574 9662 12626 9714
rect 14030 9662 14082 9714
rect 18286 9662 18338 9714
rect 29822 9662 29874 9714
rect 33406 9662 33458 9714
rect 2718 9550 2770 9602
rect 10446 9550 10498 9602
rect 14926 9550 14978 9602
rect 17950 9550 18002 9602
rect 20750 9550 20802 9602
rect 21310 9550 21362 9602
rect 23886 9550 23938 9602
rect 28590 9550 28642 9602
rect 29598 9550 29650 9602
rect 30718 9550 30770 9602
rect 30942 9550 30994 9602
rect 31278 9550 31330 9602
rect 31502 9550 31554 9602
rect 32286 9550 32338 9602
rect 37326 9550 37378 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 2718 9214 2770 9266
rect 3390 9214 3442 9266
rect 4622 9214 4674 9266
rect 22654 9214 22706 9266
rect 26574 9214 26626 9266
rect 27358 9214 27410 9266
rect 28590 9214 28642 9266
rect 28926 9214 28978 9266
rect 30158 9214 30210 9266
rect 30606 9214 30658 9266
rect 30942 9214 30994 9266
rect 31502 9214 31554 9266
rect 32398 9214 32450 9266
rect 5630 9102 5682 9154
rect 5854 9102 5906 9154
rect 18174 9102 18226 9154
rect 20862 9102 20914 9154
rect 21198 9102 21250 9154
rect 23998 9102 24050 9154
rect 24334 9102 24386 9154
rect 29374 9102 29426 9154
rect 34190 9102 34242 9154
rect 41022 9102 41074 9154
rect 2606 8990 2658 9042
rect 2942 8990 2994 9042
rect 3166 8990 3218 9042
rect 3838 8990 3890 9042
rect 5966 8990 6018 9042
rect 6526 8990 6578 9042
rect 7870 8990 7922 9042
rect 8206 8990 8258 9042
rect 10446 8990 10498 9042
rect 11006 8990 11058 9042
rect 12014 8990 12066 9042
rect 12350 8990 12402 9042
rect 12686 8990 12738 9042
rect 14366 8990 14418 9042
rect 15374 8990 15426 9042
rect 16606 8990 16658 9042
rect 16830 8990 16882 9042
rect 17502 8990 17554 9042
rect 26910 8990 26962 9042
rect 27134 8990 27186 9042
rect 27806 8990 27858 9042
rect 29150 8990 29202 9042
rect 32062 8990 32114 9042
rect 33406 8990 33458 9042
rect 3278 8878 3330 8930
rect 4174 8878 4226 8930
rect 11454 8878 11506 8930
rect 15150 8878 15202 8930
rect 20302 8878 20354 8930
rect 27022 8878 27074 8930
rect 29038 8878 29090 8930
rect 31838 8878 31890 8930
rect 36318 8878 36370 8930
rect 6862 8766 6914 8818
rect 15374 8766 15426 8818
rect 16270 8766 16322 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 10670 8430 10722 8482
rect 17950 8430 18002 8482
rect 18286 8430 18338 8482
rect 4510 8318 4562 8370
rect 8430 8318 8482 8370
rect 11678 8318 11730 8370
rect 12910 8318 12962 8370
rect 13918 8318 13970 8370
rect 17166 8318 17218 8370
rect 17726 8318 17778 8370
rect 18846 8318 18898 8370
rect 21870 8318 21922 8370
rect 22430 8318 22482 8370
rect 22654 8318 22706 8370
rect 22990 8318 23042 8370
rect 25118 8318 25170 8370
rect 32286 8318 32338 8370
rect 34414 8318 34466 8370
rect 37550 8318 37602 8370
rect 2158 8206 2210 8258
rect 5854 8206 5906 8258
rect 6414 8206 6466 8258
rect 7422 8206 7474 8258
rect 7982 8206 8034 8258
rect 9774 8206 9826 8258
rect 10894 8206 10946 8258
rect 14366 8206 14418 8258
rect 25902 8206 25954 8258
rect 31614 8206 31666 8258
rect 35758 8206 35810 8258
rect 36206 8206 36258 8258
rect 37326 8206 37378 8258
rect 7086 8094 7138 8146
rect 7198 8094 7250 8146
rect 15038 8094 15090 8146
rect 27470 8094 27522 8146
rect 31166 8094 31218 8146
rect 36990 8094 37042 8146
rect 1822 7982 1874 8034
rect 22094 7982 22146 8034
rect 27134 7982 27186 8034
rect 36430 7982 36482 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 2046 7646 2098 7698
rect 2606 7646 2658 7698
rect 7198 7646 7250 7698
rect 9550 7646 9602 7698
rect 15262 7646 15314 7698
rect 33182 7646 33234 7698
rect 35646 7646 35698 7698
rect 2718 7534 2770 7586
rect 3278 7534 3330 7586
rect 6526 7534 6578 7586
rect 7758 7534 7810 7586
rect 9774 7534 9826 7586
rect 9886 7534 9938 7586
rect 11678 7534 11730 7586
rect 15598 7534 15650 7586
rect 20526 7534 20578 7586
rect 27134 7534 27186 7586
rect 36766 7534 36818 7586
rect 1822 7422 1874 7474
rect 2382 7422 2434 7474
rect 3054 7422 3106 7474
rect 3614 7422 3666 7474
rect 4510 7422 4562 7474
rect 4846 7422 4898 7474
rect 6638 7422 6690 7474
rect 6750 7422 6802 7474
rect 7534 7422 7586 7474
rect 8430 7422 8482 7474
rect 10334 7422 10386 7474
rect 10670 7422 10722 7474
rect 10894 7422 10946 7474
rect 11790 7422 11842 7474
rect 14366 7422 14418 7474
rect 14926 7422 14978 7474
rect 16046 7422 16098 7474
rect 19742 7422 19794 7474
rect 26350 7422 26402 7474
rect 29598 7422 29650 7474
rect 35982 7422 36034 7474
rect 7982 7310 8034 7362
rect 10782 7310 10834 7362
rect 12462 7310 12514 7362
rect 17502 7310 17554 7362
rect 17950 7310 18002 7362
rect 19406 7310 19458 7362
rect 22654 7310 22706 7362
rect 26014 7310 26066 7362
rect 29262 7310 29314 7362
rect 30382 7310 30434 7362
rect 32510 7310 32562 7362
rect 38894 7310 38946 7362
rect 4622 7198 4674 7250
rect 5406 7198 5458 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 26910 6862 26962 6914
rect 3166 6750 3218 6802
rect 10222 6750 10274 6802
rect 12686 6750 12738 6802
rect 27470 6750 27522 6802
rect 27918 6750 27970 6802
rect 1710 6638 1762 6690
rect 2270 6638 2322 6690
rect 2942 6638 2994 6690
rect 3838 6638 3890 6690
rect 4398 6638 4450 6690
rect 4958 6638 5010 6690
rect 6526 6638 6578 6690
rect 7982 6638 8034 6690
rect 8318 6638 8370 6690
rect 10894 6638 10946 6690
rect 11342 6638 11394 6690
rect 12238 6638 12290 6690
rect 13358 6638 13410 6690
rect 13470 6638 13522 6690
rect 15150 6638 15202 6690
rect 20302 6638 20354 6690
rect 22206 6638 22258 6690
rect 27246 6638 27298 6690
rect 4510 6526 4562 6578
rect 5070 6526 5122 6578
rect 5966 6526 6018 6578
rect 8542 6526 8594 6578
rect 9326 6526 9378 6578
rect 9550 6526 9602 6578
rect 13694 6526 13746 6578
rect 14254 6526 14306 6578
rect 30494 6526 30546 6578
rect 30830 6526 30882 6578
rect 1822 6414 1874 6466
rect 2046 6414 2098 6466
rect 3950 6414 4002 6466
rect 4174 6414 4226 6466
rect 7310 6414 7362 6466
rect 9438 6414 9490 6466
rect 18622 6414 18674 6466
rect 19070 6414 19122 6466
rect 19518 6414 19570 6466
rect 21982 6414 22034 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 2270 6078 2322 6130
rect 3054 6078 3106 6130
rect 4398 6078 4450 6130
rect 5406 6078 5458 6130
rect 7534 6078 7586 6130
rect 8318 6078 8370 6130
rect 15486 6078 15538 6130
rect 18398 6078 18450 6130
rect 19070 6078 19122 6130
rect 19294 6078 19346 6130
rect 27022 6078 27074 6130
rect 27694 6078 27746 6130
rect 30382 6078 30434 6130
rect 31278 6078 31330 6130
rect 8878 5966 8930 6018
rect 11230 5966 11282 6018
rect 13134 5966 13186 6018
rect 13806 5966 13858 6018
rect 14478 5966 14530 6018
rect 15038 5966 15090 6018
rect 17726 5966 17778 6018
rect 18286 5966 18338 6018
rect 19294 5966 19346 6018
rect 19630 5966 19682 6018
rect 20190 5966 20242 6018
rect 21534 5966 21586 6018
rect 25790 5966 25842 6018
rect 26350 5966 26402 6018
rect 26686 5966 26738 6018
rect 30718 5966 30770 6018
rect 7758 5854 7810 5906
rect 7982 5854 8034 5906
rect 9886 5854 9938 5906
rect 10110 5854 10162 5906
rect 10782 5854 10834 5906
rect 12238 5854 12290 5906
rect 14030 5854 14082 5906
rect 14702 5854 14754 5906
rect 18622 5854 18674 5906
rect 19966 5854 20018 5906
rect 20750 5854 20802 5906
rect 27246 5854 27298 5906
rect 30942 5854 30994 5906
rect 13806 5742 13858 5794
rect 14926 5742 14978 5794
rect 23662 5742 23714 5794
rect 34974 5742 35026 5794
rect 7422 5630 7474 5682
rect 8654 5630 8706 5682
rect 10446 5630 10498 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 15710 5294 15762 5346
rect 34078 5294 34130 5346
rect 35646 5294 35698 5346
rect 37438 5294 37490 5346
rect 4622 5182 4674 5234
rect 13470 5182 13522 5234
rect 15486 5182 15538 5234
rect 20414 5182 20466 5234
rect 21534 5182 21586 5234
rect 23886 5182 23938 5234
rect 28142 5182 28194 5234
rect 32734 5182 32786 5234
rect 33518 5182 33570 5234
rect 34302 5182 34354 5234
rect 34750 5182 34802 5234
rect 35870 5182 35922 5234
rect 36430 5182 36482 5234
rect 37214 5182 37266 5234
rect 1710 5070 1762 5122
rect 6414 5070 6466 5122
rect 6638 5070 6690 5122
rect 7534 5070 7586 5122
rect 8542 5070 8594 5122
rect 9102 5070 9154 5122
rect 11230 5070 11282 5122
rect 12350 5070 12402 5122
rect 12574 5070 12626 5122
rect 12798 5070 12850 5122
rect 14142 5070 14194 5122
rect 14702 5070 14754 5122
rect 19854 5070 19906 5122
rect 21870 5070 21922 5122
rect 23326 5070 23378 5122
rect 24894 5070 24946 5122
rect 25454 5070 25506 5122
rect 25790 5070 25842 5122
rect 26014 5070 26066 5122
rect 26462 5070 26514 5122
rect 37774 5070 37826 5122
rect 38110 5070 38162 5122
rect 2494 4958 2546 5010
rect 8990 4958 9042 5010
rect 10334 4958 10386 5010
rect 13806 4958 13858 5010
rect 17726 4958 17778 5010
rect 18398 4958 18450 5010
rect 19070 4958 19122 5010
rect 19630 4958 19682 5010
rect 22430 4958 22482 5010
rect 23102 4958 23154 5010
rect 23438 4958 23490 5010
rect 5070 4846 5122 4898
rect 6078 4846 6130 4898
rect 12014 4846 12066 4898
rect 14478 4846 14530 4898
rect 16046 4846 16098 4898
rect 16494 4846 16546 4898
rect 17054 4846 17106 4898
rect 18062 4846 18114 4898
rect 19294 4846 19346 4898
rect 33742 4846 33794 4898
rect 35310 4846 35362 4898
rect 38446 4846 38498 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 8878 4510 8930 4562
rect 9662 4510 9714 4562
rect 10334 4510 10386 4562
rect 11006 4510 11058 4562
rect 11118 4510 11170 4562
rect 12574 4510 12626 4562
rect 30942 4510 30994 4562
rect 8430 4398 8482 4450
rect 10446 4398 10498 4450
rect 11790 4398 11842 4450
rect 12686 4398 12738 4450
rect 13918 4398 13970 4450
rect 16382 4398 16434 4450
rect 18174 4398 18226 4450
rect 23550 4398 23602 4450
rect 24670 4398 24722 4450
rect 26014 4398 26066 4450
rect 29038 4398 29090 4450
rect 32510 4398 32562 4450
rect 33854 4398 33906 4450
rect 7198 4286 7250 4338
rect 7422 4286 7474 4338
rect 10782 4286 10834 4338
rect 12126 4286 12178 4338
rect 13246 4286 13298 4338
rect 16606 4286 16658 4338
rect 17502 4286 17554 4338
rect 23886 4286 23938 4338
rect 24446 4286 24498 4338
rect 25342 4286 25394 4338
rect 28814 4286 28866 4338
rect 29934 4286 29986 4338
rect 30158 4286 30210 4338
rect 32286 4286 32338 4338
rect 33070 4286 33122 4338
rect 39118 4286 39170 4338
rect 16046 4174 16098 4226
rect 20302 4174 20354 4226
rect 28142 4174 28194 4226
rect 35982 4174 36034 4226
rect 36318 4174 36370 4226
rect 38446 4174 38498 4226
rect 10334 4062 10386 4114
rect 28478 4062 28530 4114
rect 30494 4062 30546 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 7422 3726 7474 3778
rect 11342 3726 11394 3778
rect 14142 3726 14194 3778
rect 33742 3726 33794 3778
rect 2494 3614 2546 3666
rect 4622 3614 4674 3666
rect 5070 3614 5122 3666
rect 8766 3614 8818 3666
rect 10894 3614 10946 3666
rect 12238 3614 12290 3666
rect 13022 3614 13074 3666
rect 14702 3614 14754 3666
rect 15934 3614 15986 3666
rect 18062 3614 18114 3666
rect 18734 3614 18786 3666
rect 18958 3614 19010 3666
rect 19518 3614 19570 3666
rect 22654 3614 22706 3666
rect 23774 3614 23826 3666
rect 25902 3614 25954 3666
rect 29710 3614 29762 3666
rect 33070 3614 33122 3666
rect 33966 3614 34018 3666
rect 34414 3614 34466 3666
rect 36206 3614 36258 3666
rect 36990 3614 37042 3666
rect 39118 3614 39170 3666
rect 1710 3502 1762 3554
rect 6638 3502 6690 3554
rect 6862 3502 6914 3554
rect 8206 3502 8258 3554
rect 10446 3502 10498 3554
rect 11902 3502 11954 3554
rect 12014 3502 12066 3554
rect 13918 3502 13970 3554
rect 14478 3502 14530 3554
rect 15150 3502 15202 3554
rect 19182 3502 19234 3554
rect 19854 3502 19906 3554
rect 22990 3502 23042 3554
rect 28478 3502 28530 3554
rect 32622 3502 32674 3554
rect 35534 3502 35586 3554
rect 39790 3502 39842 3554
rect 6974 3390 7026 3442
rect 31838 3390 31890 3442
rect 33406 3390 33458 3442
rect 35758 3390 35810 3442
rect 20190 3278 20242 3330
rect 28142 3278 28194 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 6414 2942 6466 2994
rect 6862 2942 6914 2994
rect 18286 2942 18338 2994
rect 19182 2942 19234 2994
rect 23774 2942 23826 2994
rect 30718 2942 30770 2994
rect 36766 2942 36818 2994
rect 4174 2830 4226 2882
rect 20302 2830 20354 2882
rect 27918 2830 27970 2882
rect 3390 2718 3442 2770
rect 7534 2718 7586 2770
rect 7758 2718 7810 2770
rect 10110 2718 10162 2770
rect 10558 2718 10610 2770
rect 19630 2718 19682 2770
rect 23214 2718 23266 2770
rect 23438 2718 23490 2770
rect 24222 2718 24274 2770
rect 26798 2718 26850 2770
rect 27134 2718 27186 2770
rect 30494 2718 30546 2770
rect 10334 2606 10386 2658
rect 22430 2606 22482 2658
rect 30046 2606 30098 2658
rect 7310 2494 7362 2546
rect 10110 2494 10162 2546
rect 4478 2326 4530 2378
rect 4582 2326 4634 2378
rect 4686 2326 4738 2378
rect 35198 2326 35250 2378
rect 35302 2326 35354 2378
rect 35406 2326 35458 2378
rect 6862 2046 6914 2098
rect 19838 1542 19890 1594
rect 19942 1542 19994 1594
rect 20046 1542 20098 1594
<< metal2 >>
rect 19836 78428 20100 78438
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 19836 78362 20100 78372
rect 1820 78034 1876 78046
rect 1820 77982 1822 78034
rect 1874 77982 1876 78034
rect 1820 77250 1876 77982
rect 3164 78034 3220 78046
rect 3164 77982 3166 78034
rect 3218 77982 3220 78034
rect 2940 77922 2996 77934
rect 2940 77870 2942 77922
rect 2994 77870 2996 77922
rect 2940 77364 2996 77870
rect 2940 77362 3108 77364
rect 2940 77310 2942 77362
rect 2994 77310 3108 77362
rect 2940 77308 3108 77310
rect 2940 77298 2996 77308
rect 1820 77198 1822 77250
rect 1874 77198 1876 77250
rect 1820 76466 1876 77198
rect 3052 76692 3108 77308
rect 3164 77252 3220 77982
rect 4476 77644 4740 77654
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4476 77578 4740 77588
rect 35196 77644 35460 77654
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35196 77578 35460 77588
rect 33292 77364 33348 77374
rect 33292 77362 33572 77364
rect 33292 77310 33294 77362
rect 33346 77310 33572 77362
rect 33292 77308 33572 77310
rect 33292 77298 33348 77308
rect 3164 77250 3332 77252
rect 3164 77198 3166 77250
rect 3218 77198 3332 77250
rect 3164 77196 3332 77198
rect 3164 77186 3220 77196
rect 3052 76598 3108 76636
rect 1820 76414 1822 76466
rect 1874 76414 1876 76466
rect 1820 72546 1876 76414
rect 3276 76466 3332 77196
rect 8876 77250 8932 77262
rect 8876 77198 8878 77250
rect 8930 77198 8932 77250
rect 6188 77028 6244 77038
rect 6636 77028 6692 77038
rect 7308 77028 7364 77038
rect 7532 77028 7588 77038
rect 6188 77026 7532 77028
rect 6188 76974 6190 77026
rect 6242 76974 6638 77026
rect 6690 76974 7310 77026
rect 7362 76974 7532 77026
rect 6188 76972 7532 76974
rect 3276 76414 3278 76466
rect 3330 76414 3332 76466
rect 3052 75682 3108 75694
rect 3052 75630 3054 75682
rect 3106 75630 3108 75682
rect 3052 74898 3108 75630
rect 3276 75684 3332 76414
rect 3276 75618 3332 75628
rect 3388 76916 3444 76926
rect 3052 74846 3054 74898
rect 3106 74846 3108 74898
rect 3052 74228 3108 74846
rect 1820 72494 1822 72546
rect 1874 72494 1876 72546
rect 1820 70980 1876 72494
rect 2828 74172 3108 74228
rect 2716 71764 2772 71774
rect 2828 71764 2884 74172
rect 3164 72546 3220 72558
rect 3164 72494 3166 72546
rect 3218 72494 3220 72546
rect 3164 72436 3220 72494
rect 3164 72370 3220 72380
rect 2940 72322 2996 72334
rect 2940 72270 2942 72322
rect 2994 72270 2996 72322
rect 2940 72212 2996 72270
rect 2940 72146 2996 72156
rect 2716 71762 2884 71764
rect 2716 71710 2718 71762
rect 2770 71710 2884 71762
rect 2716 71708 2884 71710
rect 1820 70914 1876 70924
rect 2380 70980 2436 70990
rect 2380 70886 2436 70924
rect 2716 70980 2772 71708
rect 2716 70914 2772 70924
rect 3388 68964 3444 76860
rect 3612 76692 3668 76702
rect 3612 76598 3668 76636
rect 4284 76692 4340 76702
rect 4284 75794 4340 76636
rect 4956 76692 5012 76702
rect 6188 76692 6244 76972
rect 6636 76962 6692 76972
rect 4956 76466 5012 76636
rect 4956 76414 4958 76466
rect 5010 76414 5012 76466
rect 4956 76402 5012 76414
rect 5852 76636 6244 76692
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 4284 75742 4286 75794
rect 4338 75742 4340 75794
rect 4284 75124 4340 75742
rect 4284 75058 4340 75068
rect 4396 75684 4452 75694
rect 4396 75570 4452 75628
rect 4396 75518 4398 75570
rect 4450 75518 4452 75570
rect 4396 74900 4452 75518
rect 5852 75458 5908 76636
rect 5964 76468 6020 76478
rect 6300 76468 6356 76478
rect 5964 76466 6356 76468
rect 5964 76414 5966 76466
rect 6018 76414 6302 76466
rect 6354 76414 6356 76466
rect 5964 76412 6356 76414
rect 5964 76402 6020 76412
rect 5852 75406 5854 75458
rect 5906 75406 5908 75458
rect 4956 75124 5012 75134
rect 5740 75124 5796 75134
rect 5852 75124 5908 75406
rect 5012 75068 5124 75124
rect 4956 75058 5012 75068
rect 4172 74898 4452 74900
rect 4172 74846 4398 74898
rect 4450 74846 4452 74898
rect 4172 74844 4452 74846
rect 4172 73948 4228 74844
rect 4396 74834 4452 74844
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 4060 73892 4228 73948
rect 4060 72436 4116 73892
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 3500 72212 3556 72222
rect 3500 71090 3556 72156
rect 3500 71038 3502 71090
rect 3554 71038 3556 71090
rect 3500 71026 3556 71038
rect 3724 71988 3780 71998
rect 3948 71988 4004 71998
rect 3612 70868 3668 70878
rect 3612 70774 3668 70812
rect 3724 69300 3780 71932
rect 3836 71932 3948 71988
rect 3836 71874 3892 71932
rect 3948 71922 4004 71932
rect 3836 71822 3838 71874
rect 3890 71822 3892 71874
rect 3836 71810 3892 71822
rect 4060 71762 4116 72380
rect 5068 72658 5124 75068
rect 5796 75068 5908 75124
rect 6188 75682 6244 76412
rect 6300 76402 6356 76412
rect 6972 76468 7028 76972
rect 7308 76962 7364 76972
rect 7532 76934 7588 76972
rect 8204 77028 8260 77038
rect 7084 76468 7140 76478
rect 6972 76466 7140 76468
rect 6972 76414 7086 76466
rect 7138 76414 7140 76466
rect 6972 76412 7140 76414
rect 6188 75630 6190 75682
rect 6242 75630 6244 75682
rect 5740 75030 5796 75068
rect 5068 72606 5070 72658
rect 5122 72606 5124 72658
rect 5068 71988 5124 72606
rect 6076 74900 6132 74910
rect 6188 74900 6244 75630
rect 6076 74898 6244 74900
rect 6076 74846 6078 74898
rect 6130 74846 6244 74898
rect 6076 74844 6244 74846
rect 6972 75682 7028 76412
rect 7084 76402 7140 76412
rect 8204 76354 8260 76972
rect 8876 77028 8932 77198
rect 8876 76962 8932 76972
rect 9884 77250 9940 77262
rect 9884 77198 9886 77250
rect 9938 77198 9940 77250
rect 8204 76302 8206 76354
rect 8258 76302 8260 76354
rect 8204 75908 8260 76302
rect 8316 75908 8372 75918
rect 8204 75906 8484 75908
rect 8204 75854 8318 75906
rect 8370 75854 8484 75906
rect 8204 75852 8484 75854
rect 8316 75814 8372 75852
rect 6972 75630 6974 75682
rect 7026 75630 7028 75682
rect 6972 74898 7028 75630
rect 8428 75124 8484 75852
rect 9884 75684 9940 77198
rect 30492 77252 30548 77262
rect 30492 77158 30548 77196
rect 31276 77252 31332 77262
rect 27804 77138 27860 77150
rect 31164 77140 31220 77150
rect 27804 77086 27806 77138
rect 27858 77086 27860 77138
rect 10108 77028 10164 77038
rect 10108 76690 10164 76972
rect 10108 76638 10110 76690
rect 10162 76638 10164 76690
rect 10108 76626 10164 76638
rect 11228 77028 11284 77038
rect 10444 76468 10500 76478
rect 11228 76468 11284 76972
rect 21532 77026 21588 77038
rect 21532 76974 21534 77026
rect 21586 76974 21588 77026
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 13020 76468 13076 76478
rect 10444 75684 10500 76412
rect 10892 76466 11508 76468
rect 10892 76414 11230 76466
rect 11282 76414 11508 76466
rect 10892 76412 11508 76414
rect 10892 75684 10948 76412
rect 11228 76402 11284 76412
rect 9884 75682 10500 75684
rect 9884 75630 9886 75682
rect 9938 75630 10500 75682
rect 9884 75628 10500 75630
rect 10556 75682 10948 75684
rect 10556 75630 10894 75682
rect 10946 75630 10948 75682
rect 10556 75628 10948 75630
rect 9548 75458 9604 75470
rect 9548 75406 9550 75458
rect 9602 75406 9604 75458
rect 8988 75124 9044 75134
rect 9548 75124 9604 75406
rect 8428 75122 9604 75124
rect 8428 75070 8430 75122
rect 8482 75070 8990 75122
rect 9042 75070 9604 75122
rect 8428 75068 9604 75070
rect 8428 75058 8484 75068
rect 6972 74846 6974 74898
rect 7026 74846 7028 74898
rect 6076 72548 6132 74844
rect 6972 72548 7028 74846
rect 8988 73218 9044 75068
rect 8988 73166 8990 73218
rect 9042 73166 9044 73218
rect 6076 72546 6356 72548
rect 6076 72494 6078 72546
rect 6130 72494 6356 72546
rect 6076 72492 6356 72494
rect 6076 72482 6132 72492
rect 5516 71988 5572 71998
rect 5124 71986 5572 71988
rect 5124 71934 5518 71986
rect 5570 71934 5572 71986
rect 5124 71932 5572 71934
rect 5068 71894 5124 71932
rect 5516 71922 5572 71932
rect 4060 71710 4062 71762
rect 4114 71710 4116 71762
rect 4060 70868 4116 71710
rect 6300 71764 6356 72492
rect 6972 72546 7140 72548
rect 6972 72494 6974 72546
rect 7026 72494 7140 72546
rect 6972 72492 7140 72494
rect 6972 72482 7028 72492
rect 7084 71764 7140 72492
rect 8316 72324 8372 72334
rect 8764 72324 8820 72334
rect 8316 72322 8820 72324
rect 8316 72270 8318 72322
rect 8370 72270 8766 72322
rect 8818 72270 8820 72322
rect 8316 72268 8820 72270
rect 8316 72258 8372 72268
rect 6300 71762 6468 71764
rect 6300 71710 6302 71762
rect 6354 71710 6468 71762
rect 6300 71708 6468 71710
rect 6300 71698 6356 71708
rect 6076 71652 6132 71662
rect 5964 71650 6132 71652
rect 5964 71598 6078 71650
rect 6130 71598 6132 71650
rect 5964 71596 6132 71598
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 4172 70980 4228 70990
rect 4620 70980 4676 70990
rect 4172 70886 4228 70924
rect 4396 70978 4676 70980
rect 4396 70926 4622 70978
rect 4674 70926 4676 70978
rect 4396 70924 4676 70926
rect 4060 70802 4116 70812
rect 4396 70418 4452 70924
rect 4620 70914 4676 70924
rect 5628 70868 5684 70878
rect 5628 70774 5684 70812
rect 5964 70866 6020 71596
rect 6076 71586 6132 71596
rect 5964 70814 5966 70866
rect 6018 70814 6020 70866
rect 4396 70366 4398 70418
rect 4450 70366 4452 70418
rect 4396 70354 4452 70366
rect 4956 70306 5012 70318
rect 4956 70254 4958 70306
rect 5010 70254 5012 70306
rect 3836 70082 3892 70094
rect 3836 70030 3838 70082
rect 3890 70030 3892 70082
rect 3836 69524 3892 70030
rect 4060 69972 4116 69982
rect 4956 69972 5012 70254
rect 4060 69970 5012 69972
rect 4060 69918 4062 69970
rect 4114 69918 5012 69970
rect 4060 69916 5012 69918
rect 4060 69906 4116 69916
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 3836 69458 3892 69468
rect 4284 69524 4340 69534
rect 3724 69244 4228 69300
rect 3388 68908 3556 68964
rect 2492 68740 2548 68750
rect 2940 68740 2996 68750
rect 3388 68740 3444 68750
rect 2492 68738 2772 68740
rect 2492 68686 2494 68738
rect 2546 68686 2772 68738
rect 2492 68684 2772 68686
rect 2492 68674 2548 68684
rect 2268 67732 2324 67742
rect 2604 67732 2660 67742
rect 2268 67730 2660 67732
rect 2268 67678 2270 67730
rect 2322 67678 2606 67730
rect 2658 67678 2660 67730
rect 2268 67676 2660 67678
rect 2268 67666 2324 67676
rect 2604 67666 2660 67676
rect 1932 67618 1988 67630
rect 1932 67566 1934 67618
rect 1986 67566 1988 67618
rect 1932 67228 1988 67566
rect 1820 67172 1988 67228
rect 2604 67508 2660 67518
rect 1820 67058 1876 67172
rect 1820 67006 1822 67058
rect 1874 67006 1876 67058
rect 1820 66994 1876 67006
rect 2492 67060 2548 67070
rect 2492 65268 2548 67004
rect 2604 66498 2660 67452
rect 2604 66446 2606 66498
rect 2658 66446 2660 66498
rect 2604 66434 2660 66446
rect 2716 66274 2772 68684
rect 2716 66222 2718 66274
rect 2770 66222 2772 66274
rect 2716 66210 2772 66222
rect 2828 68738 2996 68740
rect 2828 68686 2942 68738
rect 2994 68686 2996 68738
rect 2828 68684 2996 68686
rect 2716 65492 2772 65502
rect 2828 65492 2884 68684
rect 2940 68674 2996 68684
rect 3276 68738 3444 68740
rect 3276 68686 3390 68738
rect 3442 68686 3444 68738
rect 3276 68684 3444 68686
rect 2940 67844 2996 67854
rect 2940 67508 2996 67788
rect 2940 67442 2996 67452
rect 3164 67842 3220 67854
rect 3164 67790 3166 67842
rect 3218 67790 3220 67842
rect 3164 67172 3220 67790
rect 3164 67106 3220 67116
rect 3052 67060 3108 67070
rect 3052 66966 3108 67004
rect 2940 66948 2996 66958
rect 2940 66854 2996 66892
rect 3276 66612 3332 68684
rect 3388 68674 3444 68684
rect 3500 68068 3556 68908
rect 2940 66556 3332 66612
rect 3388 68012 3556 68068
rect 3836 68068 3892 68078
rect 3836 68066 4116 68068
rect 3836 68014 3838 68066
rect 3890 68014 4116 68066
rect 3836 68012 4116 68014
rect 2940 66386 2996 66556
rect 2940 66334 2942 66386
rect 2994 66334 2996 66386
rect 2940 66322 2996 66334
rect 2716 65490 2884 65492
rect 2716 65438 2718 65490
rect 2770 65438 2884 65490
rect 2716 65436 2884 65438
rect 2716 65426 2772 65436
rect 2828 65268 2884 65278
rect 2492 65266 2884 65268
rect 2492 65214 2830 65266
rect 2882 65214 2884 65266
rect 2492 65212 2884 65214
rect 2828 65202 2884 65212
rect 3052 63252 3108 63262
rect 2716 63028 2772 63038
rect 2716 62934 2772 62972
rect 2380 62916 2436 62926
rect 1932 62914 2436 62916
rect 1932 62862 2382 62914
rect 2434 62862 2436 62914
rect 1932 62860 2436 62862
rect 1932 62354 1988 62860
rect 2380 62850 2436 62860
rect 1932 62302 1934 62354
rect 1986 62302 1988 62354
rect 1932 61570 1988 62302
rect 3052 62578 3108 63196
rect 3052 62526 3054 62578
rect 3106 62526 3108 62578
rect 3052 61682 3108 62526
rect 3052 61630 3054 61682
rect 3106 61630 3108 61682
rect 3052 61618 3108 61630
rect 3276 62354 3332 62366
rect 3276 62302 3278 62354
rect 3330 62302 3332 62354
rect 1932 61518 1934 61570
rect 1986 61518 1988 61570
rect 1932 61506 1988 61518
rect 3276 61570 3332 62302
rect 3276 61518 3278 61570
rect 3330 61518 3332 61570
rect 3276 60676 3332 61518
rect 3276 60610 3332 60620
rect 2380 59330 2436 59342
rect 2380 59278 2382 59330
rect 2434 59278 2436 59330
rect 2268 58996 2324 59006
rect 1820 58994 2324 58996
rect 1820 58942 2270 58994
rect 2322 58942 2324 58994
rect 1820 58940 2324 58942
rect 1820 58434 1876 58940
rect 2268 58930 2324 58940
rect 1820 58382 1822 58434
rect 1874 58382 1876 58434
rect 1820 58370 1876 58382
rect 2268 57876 2324 57886
rect 2380 57876 2436 59278
rect 2268 57874 2436 57876
rect 2268 57822 2270 57874
rect 2322 57822 2436 57874
rect 2268 57820 2436 57822
rect 2604 58994 2660 59006
rect 2604 58942 2606 58994
rect 2658 58942 2660 58994
rect 2268 57810 2324 57820
rect 2604 57764 2660 58942
rect 2716 58436 2772 58446
rect 2716 58342 2772 58380
rect 2604 57762 3220 57764
rect 2604 57710 2606 57762
rect 2658 57710 3220 57762
rect 2604 57708 3220 57710
rect 2604 57698 2660 57708
rect 1932 57652 1988 57662
rect 1932 57558 1988 57596
rect 2156 57538 2212 57550
rect 2156 57486 2158 57538
rect 2210 57486 2212 57538
rect 2156 56868 2212 57486
rect 3052 57540 3108 57550
rect 3052 57446 3108 57484
rect 3164 57090 3220 57708
rect 3276 57652 3332 57662
rect 3276 57558 3332 57596
rect 3164 57038 3166 57090
rect 3218 57038 3220 57090
rect 3164 57026 3220 57038
rect 2604 56868 2660 56878
rect 2940 56868 2996 56878
rect 2156 56866 2940 56868
rect 2156 56814 2158 56866
rect 2210 56814 2606 56866
rect 2658 56814 2940 56866
rect 2156 56812 2940 56814
rect 2156 56802 2212 56812
rect 2604 56802 2660 56812
rect 2716 55522 2772 56812
rect 2940 56774 2996 56812
rect 2716 55470 2718 55522
rect 2770 55470 2772 55522
rect 1932 55300 1988 55310
rect 1820 55244 1932 55300
rect 1820 54514 1876 55244
rect 1932 55206 1988 55244
rect 1820 54462 1822 54514
rect 1874 54462 1876 54514
rect 1820 54450 1876 54462
rect 2380 55074 2436 55086
rect 2380 55022 2382 55074
rect 2434 55022 2436 55074
rect 1932 54404 1988 54414
rect 1932 53730 1988 54348
rect 2380 53956 2436 55022
rect 2604 54740 2660 54750
rect 2492 54404 2548 54414
rect 2492 54310 2548 54348
rect 2380 53900 2548 53956
rect 1932 53678 1934 53730
rect 1986 53678 1988 53730
rect 1932 53666 1988 53678
rect 2044 53506 2100 53518
rect 2044 53454 2046 53506
rect 2098 53454 2100 53506
rect 2044 51044 2100 53454
rect 2492 53506 2548 53900
rect 2604 53842 2660 54684
rect 2604 53790 2606 53842
rect 2658 53790 2660 53842
rect 2604 53778 2660 53790
rect 2492 53454 2494 53506
rect 2546 53454 2548 53506
rect 2268 52836 2324 52874
rect 2268 52770 2324 52780
rect 2044 50978 2100 50988
rect 2156 52722 2212 52734
rect 2156 52670 2158 52722
rect 2210 52670 2212 52722
rect 2156 50820 2212 52670
rect 1708 50764 2212 50820
rect 2268 52612 2324 52622
rect 2268 52162 2324 52556
rect 2268 52110 2270 52162
rect 2322 52110 2324 52162
rect 1596 42084 1652 42094
rect 1596 40628 1652 42028
rect 1708 40740 1764 50764
rect 2268 50428 2324 52110
rect 2492 51940 2548 53454
rect 2716 53506 2772 55470
rect 3164 55970 3220 55982
rect 3164 55918 3166 55970
rect 3218 55918 3220 55970
rect 2940 55074 2996 55086
rect 2940 55022 2942 55074
rect 2994 55022 2996 55074
rect 2940 53844 2996 55022
rect 3164 54514 3220 55918
rect 3276 55522 3332 55534
rect 3276 55470 3278 55522
rect 3330 55470 3332 55522
rect 3276 55298 3332 55470
rect 3276 55246 3278 55298
rect 3330 55246 3332 55298
rect 3276 55234 3332 55246
rect 3164 54462 3166 54514
rect 3218 54462 3220 54514
rect 3164 54450 3220 54462
rect 3276 54516 3332 54526
rect 2940 53842 3108 53844
rect 2940 53790 2942 53842
rect 2994 53790 3108 53842
rect 2940 53788 3108 53790
rect 2940 53778 2996 53788
rect 2716 53454 2718 53506
rect 2770 53454 2772 53506
rect 2604 52834 2660 52846
rect 2604 52782 2606 52834
rect 2658 52782 2660 52834
rect 2604 52724 2660 52782
rect 2604 52658 2660 52668
rect 2716 52722 2772 53454
rect 2716 52670 2718 52722
rect 2770 52670 2772 52722
rect 2716 52658 2772 52670
rect 2940 52946 2996 52958
rect 2940 52894 2942 52946
rect 2994 52894 2996 52946
rect 2716 51940 2772 51950
rect 2492 51884 2716 51940
rect 2716 51846 2772 51884
rect 2044 50372 2324 50428
rect 2716 50484 2772 50494
rect 2940 50484 2996 52894
rect 2772 50428 2996 50484
rect 1820 49812 1876 49822
rect 1820 49718 1876 49756
rect 1932 48916 1988 48926
rect 1932 48822 1988 48860
rect 1932 48132 1988 48142
rect 2044 48132 2100 50372
rect 2492 49698 2548 49710
rect 2492 49646 2494 49698
rect 2546 49646 2548 49698
rect 2492 49140 2548 49646
rect 2604 49140 2660 49150
rect 2492 49138 2660 49140
rect 2492 49086 2606 49138
rect 2658 49086 2660 49138
rect 2492 49084 2660 49086
rect 2604 49074 2660 49084
rect 1932 48130 2100 48132
rect 1932 48078 1934 48130
rect 1986 48078 2100 48130
rect 1932 48076 2100 48078
rect 2156 49028 2212 49038
rect 1932 48018 1988 48076
rect 1932 47966 1934 48018
rect 1986 47966 1988 48018
rect 1932 47954 1988 47966
rect 1932 47796 1988 47806
rect 1932 46116 1988 47740
rect 2156 47124 2212 48972
rect 2716 49026 2772 50428
rect 3052 49476 3108 53788
rect 3164 53732 3220 53742
rect 3164 53638 3220 53676
rect 3276 53170 3332 54460
rect 3276 53118 3278 53170
rect 3330 53118 3332 53170
rect 3276 53106 3332 53118
rect 3276 52836 3332 52846
rect 3276 52742 3332 52780
rect 3388 52388 3444 68012
rect 3836 68002 3892 68012
rect 3500 67844 3556 67854
rect 3500 67750 3556 67788
rect 3724 67618 3780 67630
rect 3724 67566 3726 67618
rect 3778 67566 3780 67618
rect 3724 67282 3780 67566
rect 3724 67230 3726 67282
rect 3778 67230 3780 67282
rect 3724 67218 3780 67230
rect 3612 67172 3668 67182
rect 3612 66386 3668 67116
rect 4060 67058 4116 68012
rect 4060 67006 4062 67058
rect 4114 67006 4116 67058
rect 4060 66994 4116 67006
rect 4172 66836 4228 69244
rect 3612 66334 3614 66386
rect 3666 66334 3668 66386
rect 3612 66322 3668 66334
rect 4060 66780 4228 66836
rect 3500 66164 3556 66174
rect 3500 66162 3668 66164
rect 3500 66110 3502 66162
rect 3554 66110 3668 66162
rect 3500 66108 3668 66110
rect 3500 66098 3556 66108
rect 3500 65828 3556 65838
rect 3500 58884 3556 65772
rect 3612 65380 3668 66108
rect 3724 66052 3780 66062
rect 3724 65958 3780 65996
rect 4060 65940 4116 66780
rect 4284 66388 4340 69468
rect 4620 69524 4676 69534
rect 4620 69430 4676 69468
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 4956 68068 5012 69916
rect 5628 70194 5684 70206
rect 5628 70142 5630 70194
rect 5682 70142 5684 70194
rect 5628 69634 5684 70142
rect 5628 69582 5630 69634
rect 5682 69582 5684 69634
rect 5628 69570 5684 69582
rect 5740 69524 5796 69534
rect 5740 69430 5796 69468
rect 4956 68002 5012 68012
rect 5740 68068 5796 68078
rect 5740 67974 5796 68012
rect 5964 67844 6020 70814
rect 6412 70978 6468 71708
rect 7084 71762 7252 71764
rect 7084 71710 7086 71762
rect 7138 71710 7252 71762
rect 7084 71708 7252 71710
rect 7084 71698 7140 71708
rect 6412 70926 6414 70978
rect 6466 70926 6468 70978
rect 6300 70420 6356 70430
rect 6412 70420 6468 70926
rect 7196 70980 7252 71708
rect 8652 71652 8708 71662
rect 8764 71652 8820 72268
rect 8988 71652 9044 73166
rect 9660 74900 9716 74910
rect 9884 74900 9940 75628
rect 10556 74900 10612 75628
rect 10892 75618 10948 75628
rect 11452 75908 11508 76412
rect 13020 76374 13076 76412
rect 13804 76466 13860 76478
rect 13804 76414 13806 76466
rect 13858 76414 13860 76466
rect 12572 76244 12628 76254
rect 12012 75908 12068 75918
rect 12572 75908 12628 76188
rect 13804 76244 13860 76414
rect 18508 76468 18564 76478
rect 21532 76468 21588 76974
rect 21756 76468 21812 76478
rect 21532 76412 21756 76468
rect 18172 76356 18228 76366
rect 18508 76356 18564 76412
rect 21756 76374 21812 76412
rect 27132 76466 27188 76478
rect 27132 76414 27134 76466
rect 27186 76414 27188 76466
rect 18172 76354 18564 76356
rect 18172 76302 18174 76354
rect 18226 76302 18564 76354
rect 18172 76300 18564 76302
rect 19292 76354 19348 76366
rect 19292 76302 19294 76354
rect 19346 76302 19348 76354
rect 13804 76178 13860 76188
rect 15148 76244 15204 76254
rect 15148 76150 15204 76188
rect 11452 75906 12740 75908
rect 11452 75854 12014 75906
rect 12066 75854 12740 75906
rect 11452 75852 12740 75854
rect 9660 74898 9940 74900
rect 9660 74846 9662 74898
rect 9714 74846 9940 74898
rect 9660 74844 9940 74846
rect 10332 74898 10612 74900
rect 10332 74846 10558 74898
rect 10610 74846 10612 74898
rect 10332 74844 10612 74846
rect 9660 74004 9716 74844
rect 9660 73330 9716 73948
rect 10332 74226 10388 74844
rect 10556 74834 10612 74844
rect 10332 74174 10334 74226
rect 10386 74174 10388 74226
rect 10332 73332 10388 74174
rect 11452 74676 11508 75852
rect 12012 75842 12068 75852
rect 12684 75796 12740 75852
rect 12684 75794 12852 75796
rect 12684 75742 12686 75794
rect 12738 75742 12852 75794
rect 12684 75740 12852 75742
rect 12684 75730 12740 75740
rect 11676 74676 11732 74686
rect 11452 74674 11732 74676
rect 11452 74622 11678 74674
rect 11730 74622 11732 74674
rect 11452 74620 11732 74622
rect 10668 74114 10724 74126
rect 10668 74062 10670 74114
rect 10722 74062 10724 74114
rect 10668 74004 10724 74062
rect 11452 74114 11508 74620
rect 11452 74062 11454 74114
rect 11506 74062 11508 74114
rect 11452 74050 11508 74062
rect 10668 73938 10724 73948
rect 9660 73278 9662 73330
rect 9714 73278 9716 73330
rect 9212 72546 9268 72558
rect 9212 72494 9214 72546
rect 9266 72494 9268 72546
rect 9212 71764 9268 72494
rect 9660 71764 9716 73278
rect 10108 73330 10388 73332
rect 10108 73278 10334 73330
rect 10386 73278 10388 73330
rect 10108 73276 10388 73278
rect 10108 72548 10164 73276
rect 10332 73266 10388 73276
rect 11676 73106 11732 74620
rect 12796 74340 12852 75740
rect 12796 74338 12964 74340
rect 12796 74286 12798 74338
rect 12850 74286 12964 74338
rect 12796 74284 12964 74286
rect 12796 74274 12852 74284
rect 12236 73892 12292 73902
rect 12236 73330 12292 73836
rect 12236 73278 12238 73330
rect 12290 73278 12292 73330
rect 12236 73266 12292 73278
rect 12908 73332 12964 74284
rect 17836 74116 17892 74126
rect 18172 74116 18228 76300
rect 19292 75908 19348 76302
rect 21420 76356 21476 76366
rect 21420 76262 21476 76300
rect 22540 76356 22596 76366
rect 23548 76356 23604 76366
rect 24668 76356 24724 76366
rect 22540 76354 22932 76356
rect 22540 76302 22542 76354
rect 22594 76302 22932 76354
rect 22540 76300 22932 76302
rect 22540 76290 22596 76300
rect 19292 75842 19348 75852
rect 21308 75908 21364 75918
rect 21308 75814 21364 75852
rect 22876 75794 22932 76300
rect 22876 75742 22878 75794
rect 22930 75742 22932 75794
rect 22876 75730 22932 75742
rect 23548 75794 23604 76300
rect 23548 75742 23550 75794
rect 23602 75742 23604 75794
rect 23548 75730 23604 75742
rect 24108 76354 24724 76356
rect 24108 76302 24670 76354
rect 24722 76302 24724 76354
rect 24108 76300 24724 76302
rect 24108 75794 24164 76300
rect 24668 76290 24724 76300
rect 26796 76356 26852 76366
rect 27132 76356 27188 76414
rect 26796 76354 27188 76356
rect 26796 76302 26798 76354
rect 26850 76302 27188 76354
rect 26796 76300 27188 76302
rect 24108 75742 24110 75794
rect 24162 75742 24164 75794
rect 24108 75730 24164 75742
rect 24556 75796 24612 75806
rect 20748 75684 20804 75694
rect 20636 75628 20748 75684
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 17836 74114 18228 74116
rect 17836 74062 17838 74114
rect 17890 74062 18228 74114
rect 17836 74060 18228 74062
rect 17500 74004 17556 74014
rect 17836 74004 17892 74060
rect 17388 74002 17892 74004
rect 17388 73950 17502 74002
rect 17554 73950 17892 74002
rect 17388 73948 17892 73950
rect 18620 74004 18676 74014
rect 18620 74002 19460 74004
rect 18620 73950 18622 74002
rect 18674 73950 19460 74002
rect 18620 73948 19460 73950
rect 13020 73332 13076 73342
rect 12908 73330 13076 73332
rect 12908 73278 13022 73330
rect 13074 73278 13076 73330
rect 12908 73276 13076 73278
rect 11676 73054 11678 73106
rect 11730 73054 11732 73106
rect 10108 72546 10388 72548
rect 10108 72494 10110 72546
rect 10162 72494 10388 72546
rect 10108 72492 10388 72494
rect 10108 72482 10164 72492
rect 9212 71762 9716 71764
rect 9212 71710 9662 71762
rect 9714 71710 9716 71762
rect 9212 71708 9716 71710
rect 8652 71650 9044 71652
rect 8652 71598 8654 71650
rect 8706 71598 8990 71650
rect 9042 71598 9044 71650
rect 8652 71596 9044 71598
rect 8652 71586 8708 71596
rect 7196 70978 7588 70980
rect 7196 70926 7198 70978
rect 7250 70926 7588 70978
rect 7196 70924 7588 70926
rect 7196 70914 7252 70924
rect 6300 70418 6804 70420
rect 6300 70366 6302 70418
rect 6354 70366 6804 70418
rect 6300 70364 6804 70366
rect 6300 70354 6356 70364
rect 6636 70196 6692 70206
rect 6188 69524 6244 69534
rect 6244 69468 6580 69524
rect 6188 69430 6244 69468
rect 6412 67954 6468 67966
rect 6412 67902 6414 67954
rect 6466 67902 6468 67954
rect 6076 67844 6132 67854
rect 5964 67788 6076 67844
rect 5516 67058 5572 67070
rect 5516 67006 5518 67058
rect 5570 67006 5572 67058
rect 4844 66948 4900 66958
rect 5516 66948 5572 67006
rect 4844 66854 4900 66892
rect 5292 66892 5516 66948
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 4732 66388 4788 66398
rect 4284 66386 4788 66388
rect 4284 66334 4286 66386
rect 4338 66334 4734 66386
rect 4786 66334 4788 66386
rect 4284 66332 4788 66334
rect 4172 66052 4228 66062
rect 4172 65958 4228 65996
rect 3612 65314 3668 65324
rect 3836 65884 4116 65940
rect 3724 63028 3780 63038
rect 3724 62578 3780 62972
rect 3724 62526 3726 62578
rect 3778 62526 3780 62578
rect 3724 62514 3780 62526
rect 3836 61348 3892 65884
rect 3948 65380 4004 65390
rect 4060 65380 4116 65390
rect 4004 65378 4116 65380
rect 4004 65326 4062 65378
rect 4114 65326 4116 65378
rect 4004 65324 4116 65326
rect 3948 61796 4004 65324
rect 4060 65314 4116 65324
rect 4284 65156 4340 66332
rect 4732 66322 4788 66332
rect 4060 65100 4340 65156
rect 4476 65100 4740 65110
rect 4060 63362 4116 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 5292 64146 5348 66892
rect 5516 66882 5572 66892
rect 5292 64094 5294 64146
rect 5346 64094 5348 64146
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 4060 63310 4062 63362
rect 4114 63310 4116 63362
rect 4060 63250 4116 63310
rect 4956 63362 5012 63374
rect 4956 63310 4958 63362
rect 5010 63310 5012 63362
rect 4060 63198 4062 63250
rect 4114 63198 4116 63250
rect 4060 63186 4116 63198
rect 4508 63252 4564 63262
rect 4508 63158 4564 63196
rect 4956 63250 5012 63310
rect 4956 63198 4958 63250
rect 5010 63198 5012 63250
rect 4284 62356 4340 62366
rect 4620 62356 4676 62366
rect 4956 62356 5012 63198
rect 5292 63252 5348 64094
rect 5292 63186 5348 63196
rect 5628 63138 5684 63150
rect 5628 63086 5630 63138
rect 5682 63086 5684 63138
rect 4284 62354 5012 62356
rect 4284 62302 4286 62354
rect 4338 62302 4622 62354
rect 4674 62302 5012 62354
rect 4284 62300 5012 62302
rect 4284 62290 4340 62300
rect 4620 62290 4676 62300
rect 4060 62132 4116 62142
rect 4732 62132 4788 62170
rect 4060 62130 4228 62132
rect 4060 62078 4062 62130
rect 4114 62078 4228 62130
rect 4060 62076 4228 62078
rect 4060 62066 4116 62076
rect 3948 61730 4004 61740
rect 4060 61908 4116 61918
rect 3500 58818 3556 58828
rect 3612 61292 3892 61348
rect 3948 61570 4004 61582
rect 3948 61518 3950 61570
rect 4002 61518 4004 61570
rect 3500 57428 3556 57438
rect 3500 57090 3556 57372
rect 3500 57038 3502 57090
rect 3554 57038 3556 57090
rect 3500 57026 3556 57038
rect 3612 54740 3668 61292
rect 3724 60676 3780 60686
rect 3724 60582 3780 60620
rect 3836 60676 3892 60686
rect 3948 60676 4004 61518
rect 3836 60674 4004 60676
rect 3836 60622 3838 60674
rect 3890 60622 4004 60674
rect 3836 60620 4004 60622
rect 3836 59220 3892 60620
rect 3724 59164 3892 59220
rect 3724 55412 3780 59164
rect 4060 59108 4116 61852
rect 4172 61796 4228 62076
rect 4732 62066 4788 62076
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 4284 61796 4340 61806
rect 4172 61794 4340 61796
rect 4172 61742 4286 61794
rect 4338 61742 4340 61794
rect 4172 61740 4340 61742
rect 4284 61460 4340 61740
rect 4284 61394 4340 61404
rect 4620 61796 4676 61806
rect 4620 61570 4676 61740
rect 4620 61518 4622 61570
rect 4674 61518 4676 61570
rect 3724 55346 3780 55356
rect 3836 59052 4116 59108
rect 4172 60676 4228 60686
rect 4172 59106 4228 60620
rect 4620 60676 4676 61518
rect 4620 60610 4676 60620
rect 4956 60564 5012 62300
rect 5180 62354 5236 62366
rect 5180 62302 5182 62354
rect 5234 62302 5236 62354
rect 5180 61684 5236 62302
rect 5628 61684 5684 63086
rect 5852 62132 5908 62142
rect 5740 61684 5796 61694
rect 5180 61682 5796 61684
rect 5180 61630 5742 61682
rect 5794 61630 5796 61682
rect 5180 61628 5796 61630
rect 5740 61618 5796 61628
rect 5628 61460 5684 61470
rect 5628 61366 5684 61404
rect 5852 61458 5908 62076
rect 5852 61406 5854 61458
rect 5906 61406 5908 61458
rect 5852 61394 5908 61406
rect 5964 61236 6020 67788
rect 6076 67750 6132 67788
rect 6412 67284 6468 67902
rect 6412 67218 6468 67228
rect 6524 67172 6580 69468
rect 6636 69522 6692 70140
rect 6748 70194 6804 70364
rect 6748 70142 6750 70194
rect 6802 70142 6804 70194
rect 6748 70130 6804 70142
rect 7532 70196 7588 70924
rect 7532 70102 7588 70140
rect 8764 70754 8820 71596
rect 8988 71586 9044 71596
rect 8764 70702 8766 70754
rect 8818 70702 8820 70754
rect 8764 70084 8820 70702
rect 9660 70196 9716 71708
rect 10332 71762 10388 72492
rect 11452 72324 11508 72334
rect 11676 72324 11732 73054
rect 13020 73108 13076 73276
rect 11788 72324 11844 72334
rect 11452 72322 11844 72324
rect 11452 72270 11454 72322
rect 11506 72270 11790 72322
rect 11842 72270 11844 72322
rect 11452 72268 11844 72270
rect 11452 72258 11508 72268
rect 10332 71710 10334 71762
rect 10386 71710 10388 71762
rect 10332 71090 10388 71710
rect 10332 71038 10334 71090
rect 10386 71038 10388 71090
rect 10332 71026 10388 71038
rect 11676 71540 11732 71550
rect 11788 71540 11844 72268
rect 11676 71538 11844 71540
rect 11676 71486 11678 71538
rect 11730 71486 11844 71538
rect 11676 71484 11844 71486
rect 10668 70978 10724 70990
rect 10668 70926 10670 70978
rect 10722 70926 10724 70978
rect 9884 70196 9940 70206
rect 9660 70140 9884 70196
rect 9884 70102 9940 70140
rect 10668 70196 10724 70926
rect 11676 70978 11732 71484
rect 11676 70926 11678 70978
rect 11730 70926 11732 70978
rect 9100 70084 9156 70094
rect 8764 70082 9156 70084
rect 8764 70030 9102 70082
rect 9154 70030 9156 70082
rect 8764 70028 9156 70030
rect 6636 69470 6638 69522
rect 6690 69470 6692 69522
rect 6636 69458 6692 69470
rect 9100 69188 9156 70028
rect 10668 69410 10724 70140
rect 10668 69358 10670 69410
rect 10722 69358 10724 69410
rect 9436 69188 9492 69198
rect 9100 69186 9492 69188
rect 9100 69134 9438 69186
rect 9490 69134 9492 69186
rect 9100 69132 9492 69134
rect 8316 67956 8372 67966
rect 8316 67862 8372 67900
rect 9436 67956 9492 69132
rect 10332 69188 10388 69198
rect 10332 68068 10388 69132
rect 10332 68002 10388 68012
rect 7644 67844 7700 67854
rect 7644 67750 7700 67788
rect 8764 67842 8820 67854
rect 8764 67790 8766 67842
rect 8818 67790 8820 67842
rect 7196 67618 7252 67630
rect 7196 67566 7198 67618
rect 7250 67566 7252 67618
rect 7196 67284 7252 67566
rect 7196 67218 7252 67228
rect 6524 67170 6916 67172
rect 6524 67118 6526 67170
rect 6578 67118 6916 67170
rect 6524 67116 6916 67118
rect 6524 67106 6580 67116
rect 6860 67058 6916 67116
rect 7308 67060 7364 67070
rect 6860 67006 6862 67058
rect 6914 67006 6916 67058
rect 6076 66948 6132 66958
rect 6076 66854 6132 66892
rect 6748 66948 6804 66958
rect 6748 66386 6804 66892
rect 6748 66334 6750 66386
rect 6802 66334 6804 66386
rect 6636 66274 6692 66286
rect 6636 66222 6638 66274
rect 6690 66222 6692 66274
rect 6636 65380 6692 66222
rect 6748 65492 6804 66334
rect 6860 66276 6916 67006
rect 7196 67058 7364 67060
rect 7196 67006 7310 67058
rect 7362 67006 7364 67058
rect 7196 67004 7364 67006
rect 6972 66836 7028 66846
rect 6972 66742 7028 66780
rect 7196 66500 7252 67004
rect 7308 66994 7364 67004
rect 7532 67058 7588 67070
rect 7532 67006 7534 67058
rect 7586 67006 7588 67058
rect 7532 66836 7588 67006
rect 8764 67060 8820 67790
rect 9436 67844 9492 67900
rect 9660 67844 9716 67854
rect 9436 67842 9716 67844
rect 9436 67790 9662 67842
rect 9714 67790 9716 67842
rect 9436 67788 9716 67790
rect 8764 66946 8820 67004
rect 8764 66894 8766 66946
rect 8818 66894 8820 66946
rect 8764 66882 8820 66894
rect 7532 66770 7588 66780
rect 9660 66834 9716 67788
rect 10668 67060 10724 69358
rect 10780 70194 10836 70206
rect 10780 70142 10782 70194
rect 10834 70142 10836 70194
rect 10780 69188 10836 70142
rect 10780 69122 10836 69132
rect 11452 69410 11508 69422
rect 11452 69358 11454 69410
rect 11506 69358 11508 69410
rect 11452 69188 11508 69358
rect 11452 69122 11508 69132
rect 11676 68852 11732 70926
rect 13020 70754 13076 73052
rect 14252 73108 14308 73118
rect 14252 73014 14308 73052
rect 13020 70702 13022 70754
rect 13074 70702 13076 70754
rect 12348 70196 12404 70206
rect 12348 70102 12404 70140
rect 11900 69970 11956 69982
rect 11900 69918 11902 69970
rect 11954 69918 11956 69970
rect 11900 69188 11956 69918
rect 13020 69522 13076 70702
rect 16828 70644 16884 70654
rect 16828 70418 16884 70588
rect 16828 70366 16830 70418
rect 16882 70366 16884 70418
rect 13356 70196 13412 70206
rect 13356 70102 13412 70140
rect 14700 70196 14756 70206
rect 13020 69470 13022 69522
rect 13074 69470 13076 69522
rect 13020 69458 13076 69470
rect 11900 69122 11956 69132
rect 12012 68852 12068 68862
rect 11676 68850 12068 68852
rect 11676 68798 12014 68850
rect 12066 68798 12068 68850
rect 11676 68796 12068 68798
rect 12012 68786 12068 68796
rect 10668 66994 10724 67004
rect 10780 68068 10836 68078
rect 10780 67058 10836 68012
rect 10780 67006 10782 67058
rect 10834 67006 10836 67058
rect 9660 66782 9662 66834
rect 9714 66782 9716 66834
rect 7868 66500 7924 66510
rect 7196 66498 7924 66500
rect 7196 66446 7198 66498
rect 7250 66446 7870 66498
rect 7922 66446 7924 66498
rect 7196 66444 7924 66446
rect 7196 66434 7252 66444
rect 7868 66434 7924 66444
rect 9436 66386 9492 66398
rect 9436 66334 9438 66386
rect 9490 66334 9492 66386
rect 6860 66210 6916 66220
rect 7308 66276 7364 66286
rect 7308 65714 7364 66220
rect 7644 66276 7700 66286
rect 7644 66182 7700 66220
rect 8204 66164 8260 66174
rect 8540 66164 8596 66174
rect 8204 66162 8596 66164
rect 8204 66110 8206 66162
rect 8258 66110 8542 66162
rect 8594 66110 8596 66162
rect 8204 66108 8596 66110
rect 8204 66098 8260 66108
rect 8540 66098 8596 66108
rect 7308 65662 7310 65714
rect 7362 65662 7364 65714
rect 7308 65650 7364 65662
rect 6748 65426 6804 65436
rect 7756 65492 7812 65502
rect 7756 65398 7812 65436
rect 9436 65492 9492 66334
rect 9660 66052 9716 66782
rect 9660 65986 9716 65996
rect 10220 66052 10276 66062
rect 10220 65958 10276 65996
rect 10780 66052 10836 67006
rect 11676 67060 11732 67070
rect 11676 66966 11732 67004
rect 14700 66388 14756 70140
rect 16380 67956 16436 67966
rect 16828 67956 16884 70366
rect 16380 67954 16884 67956
rect 16380 67902 16382 67954
rect 16434 67902 16884 67954
rect 16380 67900 16884 67902
rect 16380 67890 16436 67900
rect 14364 66386 14756 66388
rect 14364 66334 14702 66386
rect 14754 66334 14756 66386
rect 14364 66332 14756 66334
rect 10780 65986 10836 65996
rect 11116 66274 11172 66286
rect 11116 66222 11118 66274
rect 11170 66222 11172 66274
rect 6636 65314 6692 65324
rect 8204 65380 8260 65390
rect 7756 63364 7812 63374
rect 7420 63362 7812 63364
rect 7420 63310 7758 63362
rect 7810 63310 7812 63362
rect 7420 63308 7812 63310
rect 6076 63252 6132 63262
rect 6076 62354 6132 63196
rect 6412 63252 6468 63262
rect 6412 63138 6468 63196
rect 6412 63086 6414 63138
rect 6466 63086 6468 63138
rect 6412 63074 6468 63086
rect 7420 63252 7476 63308
rect 7756 63298 7812 63308
rect 7420 62580 7476 63196
rect 7420 62486 7476 62524
rect 6076 62302 6078 62354
rect 6130 62302 6132 62354
rect 6076 62290 6132 62302
rect 8204 62188 8260 65324
rect 8988 65380 9044 65390
rect 8988 65286 9044 65324
rect 9436 64706 9492 65436
rect 9548 65490 9604 65502
rect 9548 65438 9550 65490
rect 9602 65438 9604 65490
rect 9548 65380 9604 65438
rect 10780 65492 10836 65502
rect 10836 65436 10948 65492
rect 10780 65398 10836 65436
rect 9548 65314 9604 65324
rect 9436 64654 9438 64706
rect 9490 64654 9492 64706
rect 9436 64642 9492 64654
rect 10108 65266 10164 65278
rect 10108 65214 10110 65266
rect 10162 65214 10164 65266
rect 10108 64708 10164 65214
rect 10108 64642 10164 64652
rect 10780 64708 10836 64718
rect 10780 64614 10836 64652
rect 10668 64484 10724 64494
rect 10668 64390 10724 64428
rect 10780 63924 10836 63934
rect 10892 63924 10948 65436
rect 11116 65380 11172 66222
rect 12460 66274 12516 66286
rect 13468 66276 13524 66286
rect 12460 66222 12462 66274
rect 12514 66222 12516 66274
rect 11116 64708 11172 65324
rect 11116 64642 11172 64652
rect 11340 66052 11396 66062
rect 11340 64484 11396 65996
rect 12124 65490 12180 65502
rect 12124 65438 12126 65490
rect 12178 65438 12180 65490
rect 12012 65378 12068 65390
rect 12012 65326 12014 65378
rect 12066 65326 12068 65378
rect 11452 64484 11508 64494
rect 11340 64428 11452 64484
rect 10556 63922 10948 63924
rect 10556 63870 10782 63922
rect 10834 63870 10948 63922
rect 10556 63868 10948 63870
rect 7868 62132 8260 62188
rect 8316 63138 8372 63150
rect 8316 63086 8318 63138
rect 8370 63086 8372 63138
rect 7644 61572 7700 61582
rect 5740 61180 6020 61236
rect 7532 61516 7644 61572
rect 5068 60676 5124 60686
rect 5068 60582 5124 60620
rect 4956 60452 5012 60508
rect 4476 60396 4740 60406
rect 4956 60396 5124 60452
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 4172 59054 4174 59106
rect 4226 59054 4228 59106
rect 3724 55188 3780 55198
rect 3724 55094 3780 55132
rect 3612 54674 3668 54684
rect 3612 54516 3668 54526
rect 3612 54422 3668 54460
rect 3612 53844 3668 53854
rect 3612 53730 3668 53788
rect 3724 53844 3780 53854
rect 3836 53844 3892 59052
rect 3724 53842 3892 53844
rect 3724 53790 3726 53842
rect 3778 53790 3892 53842
rect 3724 53788 3892 53790
rect 3948 58884 4004 58894
rect 3724 53778 3780 53788
rect 3612 53678 3614 53730
rect 3666 53678 3668 53730
rect 3612 53666 3668 53678
rect 3724 53508 3780 53518
rect 3724 53058 3780 53452
rect 3724 53006 3726 53058
rect 3778 53006 3780 53058
rect 3500 52946 3556 52958
rect 3500 52894 3502 52946
rect 3554 52894 3556 52946
rect 3500 52724 3556 52894
rect 3500 52658 3556 52668
rect 3724 52388 3780 53006
rect 3388 52332 3668 52388
rect 3164 52276 3220 52286
rect 3164 52274 3556 52276
rect 3164 52222 3166 52274
rect 3218 52222 3556 52274
rect 3164 52220 3556 52222
rect 3164 52210 3220 52220
rect 3500 52162 3556 52220
rect 3500 52110 3502 52162
rect 3554 52110 3556 52162
rect 3276 51940 3332 51950
rect 2716 48974 2718 49026
rect 2770 48974 2772 49026
rect 2716 48962 2772 48974
rect 2828 49420 3108 49476
rect 3164 51268 3220 51278
rect 2268 48916 2324 48926
rect 2268 48822 2324 48860
rect 2492 48804 2548 48814
rect 2492 48802 2660 48804
rect 2492 48750 2494 48802
rect 2546 48750 2660 48802
rect 2492 48748 2660 48750
rect 2492 48738 2548 48748
rect 2380 48132 2436 48142
rect 2380 48038 2436 48076
rect 2492 48020 2548 48030
rect 2268 47460 2324 47470
rect 2268 47346 2324 47404
rect 2492 47458 2548 47964
rect 2492 47406 2494 47458
rect 2546 47406 2548 47458
rect 2492 47394 2548 47406
rect 2268 47294 2270 47346
rect 2322 47294 2324 47346
rect 2268 47282 2324 47294
rect 2380 47348 2436 47358
rect 2380 47254 2436 47292
rect 2156 47068 2324 47124
rect 2268 46564 2324 47068
rect 2604 46788 2660 48748
rect 2828 48692 2884 49420
rect 2716 48636 2884 48692
rect 2940 49252 2996 49262
rect 2716 47796 2772 48636
rect 2716 47730 2772 47740
rect 2828 48468 2884 48478
rect 2716 47572 2772 47582
rect 2828 47572 2884 48412
rect 2940 47682 2996 49196
rect 3052 49028 3108 49038
rect 3164 49028 3220 51212
rect 3276 51266 3332 51884
rect 3276 51214 3278 51266
rect 3330 51214 3332 51266
rect 3276 50372 3332 51214
rect 3276 50306 3332 50316
rect 3388 51044 3444 51054
rect 3108 48972 3220 49028
rect 3276 49028 3332 49038
rect 3052 48962 3108 48972
rect 3276 48934 3332 48972
rect 2940 47630 2942 47682
rect 2994 47630 2996 47682
rect 2940 47618 2996 47630
rect 3052 48802 3108 48814
rect 3052 48750 3054 48802
rect 3106 48750 3108 48802
rect 3052 48354 3108 48750
rect 3052 48302 3054 48354
rect 3106 48302 3108 48354
rect 2716 47570 2884 47572
rect 2716 47518 2718 47570
rect 2770 47518 2884 47570
rect 2716 47516 2884 47518
rect 2716 47506 2772 47516
rect 2940 47012 2996 47022
rect 2604 46732 2772 46788
rect 2604 46564 2660 46574
rect 2268 46562 2604 46564
rect 2268 46510 2270 46562
rect 2322 46510 2604 46562
rect 2268 46508 2604 46510
rect 2268 46498 2324 46508
rect 2604 46470 2660 46508
rect 2156 46340 2212 46350
rect 2716 46340 2772 46732
rect 1932 46060 2100 46116
rect 1932 45892 1988 45902
rect 1820 45890 1988 45892
rect 1820 45838 1934 45890
rect 1986 45838 1988 45890
rect 1820 45836 1988 45838
rect 1820 41412 1876 45836
rect 1932 45826 1988 45836
rect 2044 44548 2100 46060
rect 2156 46002 2212 46284
rect 2492 46284 2772 46340
rect 2828 46450 2884 46462
rect 2828 46398 2830 46450
rect 2882 46398 2884 46450
rect 2156 45950 2158 46002
rect 2210 45950 2212 46002
rect 2156 45938 2212 45950
rect 2380 46116 2436 46126
rect 2380 45778 2436 46060
rect 2380 45726 2382 45778
rect 2434 45726 2436 45778
rect 2380 44996 2436 45726
rect 2492 45108 2548 46284
rect 2828 46116 2884 46398
rect 2940 46340 2996 46956
rect 3052 46564 3108 48302
rect 3164 48802 3220 48814
rect 3164 48750 3166 48802
rect 3218 48750 3220 48802
rect 3164 48020 3220 48750
rect 3164 47954 3220 47964
rect 3276 48132 3332 48142
rect 3164 47460 3220 47470
rect 3164 46898 3220 47404
rect 3164 46846 3166 46898
rect 3218 46846 3220 46898
rect 3164 46834 3220 46846
rect 3276 46676 3332 48076
rect 3276 46610 3332 46620
rect 3052 46498 3108 46508
rect 2940 46274 2996 46284
rect 2940 46116 2996 46126
rect 2828 46060 2940 46116
rect 2940 46022 2996 46060
rect 3052 46002 3108 46014
rect 3052 45950 3054 46002
rect 3106 45950 3108 46002
rect 2604 45892 2660 45902
rect 3052 45892 3108 45950
rect 2604 45890 3108 45892
rect 2604 45838 2606 45890
rect 2658 45838 3108 45890
rect 2604 45836 3108 45838
rect 3276 45892 3332 45902
rect 2604 45826 2660 45836
rect 3276 45798 3332 45836
rect 3052 45556 3108 45566
rect 2828 45332 2884 45342
rect 2828 45330 2996 45332
rect 2828 45278 2830 45330
rect 2882 45278 2996 45330
rect 2828 45276 2996 45278
rect 2828 45266 2884 45276
rect 2492 45052 2884 45108
rect 2380 44902 2436 44940
rect 2044 44482 2100 44492
rect 2492 44324 2548 44334
rect 2492 44230 2548 44268
rect 2828 44212 2884 45052
rect 2940 44996 2996 45276
rect 2940 44930 2996 44940
rect 2940 44324 2996 44334
rect 2940 44230 2996 44268
rect 2828 44118 2884 44156
rect 2604 44100 2660 44110
rect 1932 44098 2660 44100
rect 1932 44046 2606 44098
rect 2658 44046 2660 44098
rect 1932 44044 2660 44046
rect 1932 42756 1988 44044
rect 2604 44034 2660 44044
rect 2940 43988 2996 43998
rect 2716 43426 2772 43438
rect 2716 43374 2718 43426
rect 2770 43374 2772 43426
rect 2268 42812 2548 42868
rect 1932 42754 2212 42756
rect 1932 42702 1934 42754
rect 1986 42702 2212 42754
rect 1932 42700 2212 42702
rect 1932 42690 1988 42700
rect 2044 42530 2100 42542
rect 2044 42478 2046 42530
rect 2098 42478 2100 42530
rect 2044 41636 2100 42478
rect 2044 41570 2100 41580
rect 1820 41356 2100 41412
rect 1820 41188 1876 41198
rect 1820 41094 1876 41132
rect 2044 40964 2100 41356
rect 2156 41076 2212 42700
rect 2268 42754 2324 42812
rect 2268 42702 2270 42754
rect 2322 42702 2324 42754
rect 2268 42690 2324 42702
rect 2492 42754 2548 42812
rect 2492 42702 2494 42754
rect 2546 42702 2548 42754
rect 2492 42690 2548 42702
rect 2604 42866 2660 42878
rect 2604 42814 2606 42866
rect 2658 42814 2660 42866
rect 2380 42644 2436 42654
rect 2268 42196 2324 42206
rect 2380 42196 2436 42588
rect 2268 42194 2436 42196
rect 2268 42142 2270 42194
rect 2322 42142 2436 42194
rect 2268 42140 2436 42142
rect 2268 42130 2324 42140
rect 2604 41972 2660 42814
rect 2716 42754 2772 43374
rect 2716 42702 2718 42754
rect 2770 42702 2772 42754
rect 2716 42690 2772 42702
rect 2940 42644 2996 43932
rect 2940 42550 2996 42588
rect 3052 42196 3108 45500
rect 3388 45108 3444 50988
rect 3500 50596 3556 52110
rect 3500 50530 3556 50540
rect 3500 50372 3556 50382
rect 3500 48802 3556 50316
rect 3500 48750 3502 48802
rect 3554 48750 3556 48802
rect 3500 48132 3556 48750
rect 3500 48066 3556 48076
rect 3500 47460 3556 47470
rect 3500 47366 3556 47404
rect 3612 47012 3668 52332
rect 3724 52322 3780 52332
rect 3836 53506 3892 53518
rect 3836 53454 3838 53506
rect 3890 53454 3892 53506
rect 3724 52164 3780 52174
rect 3724 52070 3780 52108
rect 3724 51268 3780 51278
rect 3724 51174 3780 51212
rect 3724 50818 3780 50830
rect 3724 50766 3726 50818
rect 3778 50766 3780 50818
rect 3724 50484 3780 50766
rect 3724 50418 3780 50428
rect 3836 49924 3892 53454
rect 3948 51044 4004 58828
rect 4060 58436 4116 58446
rect 4060 58342 4116 58380
rect 4172 58212 4228 59054
rect 4620 59106 4676 59118
rect 4620 59054 4622 59106
rect 4674 59054 4676 59106
rect 4620 58996 4676 59054
rect 4284 58940 4676 58996
rect 4284 58436 4340 58940
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 5068 58546 5124 60396
rect 5740 59220 5796 61180
rect 7532 60788 7588 61516
rect 7644 61478 7700 61516
rect 7084 60786 7588 60788
rect 7084 60734 7534 60786
rect 7586 60734 7588 60786
rect 7084 60732 7588 60734
rect 5852 60564 5908 60574
rect 5852 59442 5908 60508
rect 5852 59390 5854 59442
rect 5906 59390 5908 59442
rect 5852 59332 5908 59390
rect 6300 59892 6356 59902
rect 5852 59276 6244 59332
rect 5740 59164 5908 59220
rect 5404 59108 5460 59118
rect 5068 58494 5070 58546
rect 5122 58494 5124 58546
rect 5068 58482 5124 58494
rect 5180 59106 5460 59108
rect 5180 59054 5406 59106
rect 5458 59054 5460 59106
rect 5180 59052 5460 59054
rect 4284 58370 4340 58380
rect 4508 58434 4564 58446
rect 4508 58382 4510 58434
rect 4562 58382 4564 58434
rect 4060 58156 4228 58212
rect 4284 58210 4340 58222
rect 4284 58158 4286 58210
rect 4338 58158 4340 58210
rect 4060 57540 4116 58156
rect 4172 57652 4228 57662
rect 4284 57652 4340 58158
rect 4172 57650 4340 57652
rect 4172 57598 4174 57650
rect 4226 57598 4340 57650
rect 4172 57596 4340 57598
rect 4172 57586 4228 57596
rect 4060 57474 4116 57484
rect 4508 57428 4564 58382
rect 4508 57362 4564 57372
rect 5180 57652 5236 59052
rect 5404 59042 5460 59052
rect 5740 58996 5796 59006
rect 5628 58940 5740 58996
rect 5292 58436 5348 58446
rect 5292 57876 5348 58380
rect 5292 57782 5348 57820
rect 5180 57316 5236 57596
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 4956 57260 5236 57316
rect 5404 57650 5460 57662
rect 5404 57598 5406 57650
rect 5458 57598 5460 57650
rect 4956 56978 5012 57260
rect 5404 57204 5460 57598
rect 5068 57148 5460 57204
rect 5068 57090 5124 57148
rect 5068 57038 5070 57090
rect 5122 57038 5124 57090
rect 5068 57026 5124 57038
rect 4956 56926 4958 56978
rect 5010 56926 5012 56978
rect 4284 56644 4340 56654
rect 4060 56642 4340 56644
rect 4060 56590 4286 56642
rect 4338 56590 4340 56642
rect 4060 56588 4340 56590
rect 4060 55188 4116 56588
rect 4284 56578 4340 56588
rect 4732 56644 4788 56654
rect 4732 56642 4900 56644
rect 4732 56590 4734 56642
rect 4786 56590 4900 56642
rect 4732 56588 4900 56590
rect 4732 56578 4788 56588
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4172 55412 4228 55422
rect 4228 55356 4340 55412
rect 4172 55346 4228 55356
rect 4060 53172 4116 55132
rect 4172 55076 4228 55086
rect 4172 53956 4228 55020
rect 4284 53956 4340 55356
rect 4620 55300 4676 55310
rect 4620 55206 4676 55244
rect 4732 55076 4788 55086
rect 4844 55076 4900 56588
rect 4788 55020 4900 55076
rect 4732 55010 4788 55020
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4508 53956 4564 53966
rect 4284 53900 4452 53956
rect 4172 53890 4228 53900
rect 4060 52946 4116 53116
rect 4172 53732 4228 53742
rect 4172 53170 4228 53676
rect 4284 53730 4340 53742
rect 4284 53678 4286 53730
rect 4338 53678 4340 53730
rect 4284 53620 4340 53678
rect 4284 53554 4340 53564
rect 4172 53118 4174 53170
rect 4226 53118 4228 53170
rect 4172 53106 4228 53118
rect 4284 53060 4340 53070
rect 4284 52966 4340 53004
rect 4060 52894 4062 52946
rect 4114 52894 4116 52946
rect 4060 52612 4116 52894
rect 4060 52546 4116 52556
rect 4172 52836 4228 52846
rect 4060 52388 4116 52398
rect 4060 52294 4116 52332
rect 4172 51268 4228 52780
rect 4396 52724 4452 53900
rect 4508 53730 4564 53900
rect 4956 53732 5012 56926
rect 5628 55468 5684 58940
rect 5740 58930 5796 58940
rect 5852 57092 5908 59164
rect 5740 57036 5908 57092
rect 5740 56532 5796 57036
rect 5964 56980 6020 59276
rect 6188 59218 6244 59276
rect 6188 59166 6190 59218
rect 6242 59166 6244 59218
rect 6188 59154 6244 59166
rect 6300 58996 6356 59836
rect 7084 59890 7140 60732
rect 7532 60722 7588 60732
rect 7644 60788 7700 60798
rect 7644 60226 7700 60732
rect 7644 60174 7646 60226
rect 7698 60174 7700 60226
rect 7644 60162 7700 60174
rect 7084 59838 7086 59890
rect 7138 59838 7140 59890
rect 7084 59826 7140 59838
rect 7532 59892 7588 59902
rect 7532 59798 7588 59836
rect 6748 59778 6804 59790
rect 6748 59726 6750 59778
rect 6802 59726 6804 59778
rect 6748 59442 6804 59726
rect 6748 59390 6750 59442
rect 6802 59390 6804 59442
rect 6748 59378 6804 59390
rect 6300 58434 6356 58940
rect 6412 58996 6468 59006
rect 6412 58994 6692 58996
rect 6412 58942 6414 58994
rect 6466 58942 6692 58994
rect 6412 58940 6692 58942
rect 6412 58930 6468 58940
rect 6636 58546 6692 58940
rect 6636 58494 6638 58546
rect 6690 58494 6692 58546
rect 6300 58382 6302 58434
rect 6354 58382 6356 58434
rect 6300 58370 6356 58382
rect 6524 58436 6580 58446
rect 6524 58342 6580 58380
rect 6412 57876 6468 57886
rect 6412 57782 6468 57820
rect 5852 56924 6020 56980
rect 6636 56978 6692 58494
rect 7196 58436 7252 58446
rect 7196 58212 7252 58380
rect 7196 58210 7364 58212
rect 7196 58158 7198 58210
rect 7250 58158 7364 58210
rect 7196 58156 7364 58158
rect 7196 58146 7252 58156
rect 6748 57876 6804 57886
rect 6748 57428 6804 57820
rect 7308 57540 7364 58156
rect 6860 57428 6916 57438
rect 6748 57426 6916 57428
rect 6748 57374 6862 57426
rect 6914 57374 6916 57426
rect 6748 57372 6916 57374
rect 6860 57362 6916 57372
rect 6636 56926 6638 56978
rect 6690 56926 6692 56978
rect 5852 56868 5908 56924
rect 6636 56914 6692 56926
rect 6748 56980 6804 56990
rect 6524 56868 6580 56878
rect 5852 56774 5908 56812
rect 5964 56866 6580 56868
rect 5964 56814 6526 56866
rect 6578 56814 6580 56866
rect 5964 56812 6580 56814
rect 5964 56754 6020 56812
rect 6524 56802 6580 56812
rect 5964 56702 5966 56754
rect 6018 56702 6020 56754
rect 5964 56690 6020 56702
rect 5740 56476 6020 56532
rect 5628 55412 5908 55468
rect 5180 55074 5236 55086
rect 5180 55022 5182 55074
rect 5234 55022 5236 55074
rect 5180 54964 5236 55022
rect 5740 55076 5796 55086
rect 5740 54982 5796 55020
rect 5180 54898 5236 54908
rect 5852 53844 5908 55412
rect 5964 55074 6020 56476
rect 6300 56082 6356 56094
rect 6300 56030 6302 56082
rect 6354 56030 6356 56082
rect 6188 55188 6244 55198
rect 6188 55094 6244 55132
rect 5964 55022 5966 55074
rect 6018 55022 6020 55074
rect 5964 54964 6020 55022
rect 6076 55076 6132 55086
rect 6076 54982 6132 55020
rect 5964 54628 6020 54908
rect 5964 54572 6244 54628
rect 5852 53788 6132 53844
rect 4508 53678 4510 53730
rect 4562 53678 4564 53730
rect 4508 53058 4564 53678
rect 4508 53006 4510 53058
rect 4562 53006 4564 53058
rect 4508 52948 4564 53006
rect 4508 52882 4564 52892
rect 4732 53676 5012 53732
rect 4172 51174 4228 51212
rect 4284 52668 4452 52724
rect 4732 52724 4788 53676
rect 5516 53620 5572 53630
rect 4844 53506 4900 53518
rect 4844 53454 4846 53506
rect 4898 53454 4900 53506
rect 4844 53396 4900 53454
rect 4844 53330 4900 53340
rect 4956 53506 5012 53518
rect 4956 53454 4958 53506
rect 5010 53454 5012 53506
rect 4956 53172 5012 53454
rect 5068 53508 5124 53518
rect 5068 53506 5348 53508
rect 5068 53454 5070 53506
rect 5122 53454 5348 53506
rect 5068 53452 5348 53454
rect 5068 53442 5124 53452
rect 5180 53172 5236 53182
rect 4956 53170 5236 53172
rect 4956 53118 5182 53170
rect 5234 53118 5236 53170
rect 4956 53116 5236 53118
rect 5180 53106 5236 53116
rect 5292 53172 5348 53452
rect 5292 53106 5348 53116
rect 5404 52946 5460 52958
rect 5404 52894 5406 52946
rect 5458 52894 5460 52946
rect 5292 52834 5348 52846
rect 5292 52782 5294 52834
rect 5346 52782 5348 52834
rect 4732 52668 5012 52724
rect 3948 50988 4228 51044
rect 3948 50596 4004 50606
rect 3948 50428 4004 50540
rect 3948 50372 4116 50428
rect 3948 49924 4004 49934
rect 3836 49868 3948 49924
rect 3948 49858 4004 49868
rect 3948 49700 4004 49710
rect 3948 49026 4004 49644
rect 3948 48974 3950 49026
rect 4002 48974 4004 49026
rect 3948 48356 4004 48974
rect 3612 46946 3668 46956
rect 3724 48300 4004 48356
rect 4060 48468 4116 50372
rect 3724 47458 3780 48300
rect 3724 47406 3726 47458
rect 3778 47406 3780 47458
rect 3612 46676 3668 46686
rect 3612 46562 3668 46620
rect 3612 46510 3614 46562
rect 3666 46510 3668 46562
rect 3500 46116 3556 46126
rect 3612 46116 3668 46510
rect 3556 46060 3668 46116
rect 3724 46116 3780 47406
rect 3500 46050 3556 46060
rect 3724 46050 3780 46060
rect 3836 48130 3892 48142
rect 3836 48078 3838 48130
rect 3890 48078 3892 48130
rect 3612 45892 3668 45902
rect 3612 45798 3668 45836
rect 3724 45892 3780 45902
rect 3836 45892 3892 48078
rect 4060 47460 4116 48412
rect 4172 47570 4228 50988
rect 4284 49252 4340 52668
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4844 52500 4900 52510
rect 4732 52388 4788 52398
rect 4844 52388 4900 52444
rect 4732 52386 4900 52388
rect 4732 52334 4734 52386
rect 4786 52334 4900 52386
rect 4732 52332 4900 52334
rect 4732 52322 4788 52332
rect 4396 52050 4452 52062
rect 4396 51998 4398 52050
rect 4450 51998 4452 52050
rect 4396 51940 4452 51998
rect 4620 51940 4676 51950
rect 4396 51874 4452 51884
rect 4508 51938 4676 51940
rect 4508 51886 4622 51938
rect 4674 51886 4676 51938
rect 4508 51884 4676 51886
rect 4508 51378 4564 51884
rect 4620 51874 4676 51884
rect 4508 51326 4510 51378
rect 4562 51326 4564 51378
rect 4508 51268 4564 51326
rect 4508 51202 4564 51212
rect 4844 51378 4900 51390
rect 4844 51326 4846 51378
rect 4898 51326 4900 51378
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4844 50820 4900 51326
rect 4732 50764 4900 50820
rect 4396 50594 4452 50606
rect 4396 50542 4398 50594
rect 4450 50542 4452 50594
rect 4396 49700 4452 50542
rect 4732 50484 4788 50764
rect 4844 50596 4900 50606
rect 4844 50502 4900 50540
rect 4732 50418 4788 50428
rect 4844 49924 4900 49934
rect 4620 49700 4676 49710
rect 4452 49698 4676 49700
rect 4452 49646 4622 49698
rect 4674 49646 4676 49698
rect 4452 49644 4676 49646
rect 4396 49634 4452 49644
rect 4620 49634 4676 49644
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4284 49028 4340 49196
rect 4508 49140 4564 49150
rect 4508 49046 4564 49084
rect 4284 48962 4340 48972
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4172 47518 4174 47570
rect 4226 47518 4228 47570
rect 4172 47506 4228 47518
rect 4620 47684 4676 47694
rect 4620 47460 4676 47628
rect 4060 47366 4116 47404
rect 4284 47404 4676 47460
rect 4172 47236 4228 47246
rect 3724 45890 3892 45892
rect 3724 45838 3726 45890
rect 3778 45838 3892 45890
rect 3724 45836 3892 45838
rect 3948 47234 4228 47236
rect 3948 47182 4174 47234
rect 4226 47182 4228 47234
rect 3948 47180 4228 47182
rect 3724 45826 3780 45836
rect 3500 45108 3556 45118
rect 3388 45106 3556 45108
rect 3388 45054 3502 45106
rect 3554 45054 3556 45106
rect 3388 45052 3556 45054
rect 3500 45042 3556 45052
rect 3836 44996 3892 45006
rect 3388 44324 3444 44334
rect 3500 44324 3556 44334
rect 3052 42130 3108 42140
rect 3276 44268 3388 44324
rect 3444 44322 3556 44324
rect 3444 44270 3502 44322
rect 3554 44270 3556 44322
rect 3444 44268 3556 44270
rect 3276 42642 3332 44268
rect 3388 44230 3444 44268
rect 3500 44258 3556 44268
rect 3500 44100 3556 44110
rect 3500 42754 3556 44044
rect 3836 44100 3892 44940
rect 3836 44006 3892 44044
rect 3948 43092 4004 47180
rect 4172 47170 4228 47180
rect 4060 47012 4116 47022
rect 4060 43204 4116 46956
rect 4172 46900 4228 46910
rect 4284 46900 4340 47404
rect 4396 47236 4452 47246
rect 4396 47234 4564 47236
rect 4396 47182 4398 47234
rect 4450 47182 4564 47234
rect 4396 47180 4564 47182
rect 4396 47170 4452 47180
rect 4172 46898 4340 46900
rect 4172 46846 4174 46898
rect 4226 46846 4340 46898
rect 4172 46844 4340 46846
rect 4508 46898 4564 47180
rect 4508 46846 4510 46898
rect 4562 46846 4564 46898
rect 4172 46834 4228 46844
rect 4508 46834 4564 46846
rect 4620 46898 4676 47404
rect 4844 47012 4900 49868
rect 4956 47460 5012 52668
rect 5292 52276 5348 52782
rect 5292 52210 5348 52220
rect 5292 49812 5348 49822
rect 5292 49718 5348 49756
rect 4956 47404 5236 47460
rect 4956 47236 5012 47246
rect 4956 47124 5012 47180
rect 4956 47068 5124 47124
rect 4844 46956 5012 47012
rect 4620 46846 4622 46898
rect 4674 46846 4676 46898
rect 4620 46834 4676 46846
rect 4844 46786 4900 46798
rect 4844 46734 4846 46786
rect 4898 46734 4900 46786
rect 4396 46676 4452 46686
rect 4284 46674 4452 46676
rect 4284 46622 4398 46674
rect 4450 46622 4452 46674
rect 4284 46620 4452 46622
rect 4284 46564 4340 46620
rect 4396 46610 4452 46620
rect 4844 46676 4900 46734
rect 4844 46610 4900 46620
rect 4172 46004 4228 46014
rect 4284 46004 4340 46508
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4172 46002 4340 46004
rect 4172 45950 4174 46002
rect 4226 45950 4340 46002
rect 4172 45948 4340 45950
rect 4396 46116 4452 46126
rect 4172 45556 4228 45948
rect 4396 45892 4452 46060
rect 4172 45490 4228 45500
rect 4284 45836 4452 45892
rect 4060 43138 4116 43148
rect 4172 45332 4228 45342
rect 4172 44210 4228 45276
rect 4284 44324 4340 45836
rect 4620 45666 4676 45678
rect 4620 45614 4622 45666
rect 4674 45614 4676 45666
rect 4620 44996 4676 45614
rect 4620 44930 4676 44940
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4396 44324 4452 44334
rect 4284 44322 4452 44324
rect 4284 44270 4398 44322
rect 4450 44270 4452 44322
rect 4284 44268 4452 44270
rect 4172 44158 4174 44210
rect 4226 44158 4228 44210
rect 3500 42702 3502 42754
rect 3554 42702 3556 42754
rect 3500 42690 3556 42702
rect 3612 43036 4004 43092
rect 3276 42590 3278 42642
rect 3330 42590 3332 42642
rect 3276 42196 3332 42590
rect 3276 42130 3332 42140
rect 3388 42420 3444 42430
rect 2492 41916 2660 41972
rect 2716 42082 2772 42094
rect 2716 42030 2718 42082
rect 2770 42030 2772 42082
rect 2492 41298 2548 41916
rect 2492 41246 2494 41298
rect 2546 41246 2548 41298
rect 2492 41234 2548 41246
rect 2604 41636 2660 41646
rect 2716 41636 2772 42030
rect 2828 41972 2884 41982
rect 2828 41878 2884 41916
rect 2940 41748 2996 41758
rect 2940 41654 2996 41692
rect 2716 41580 2884 41636
rect 2156 41020 2548 41076
rect 2044 40908 2436 40964
rect 1708 40684 2324 40740
rect 1596 40572 1764 40628
rect 1708 38836 1764 40572
rect 2156 40292 2212 40302
rect 1820 40290 2212 40292
rect 1820 40238 2158 40290
rect 2210 40238 2212 40290
rect 1820 40236 2212 40238
rect 1820 39620 1876 40236
rect 2156 40226 2212 40236
rect 1820 39618 1988 39620
rect 1820 39566 1822 39618
rect 1874 39566 1988 39618
rect 1820 39564 1988 39566
rect 1820 39554 1876 39564
rect 1596 38780 1764 38836
rect 1820 38834 1876 38846
rect 1820 38782 1822 38834
rect 1874 38782 1876 38834
rect 1596 37940 1652 38780
rect 1820 38668 1876 38782
rect 1708 38612 1876 38668
rect 1708 38162 1764 38612
rect 1708 38110 1710 38162
rect 1762 38110 1764 38162
rect 1708 38098 1764 38110
rect 1820 38052 1876 38062
rect 1596 37884 1764 37940
rect 1708 33124 1764 37884
rect 1820 36932 1876 37996
rect 1932 37492 1988 39564
rect 1932 37426 1988 37436
rect 2044 39394 2100 39406
rect 2044 39342 2046 39394
rect 2098 39342 2100 39394
rect 2044 37268 2100 39342
rect 2268 39058 2324 40684
rect 2268 39006 2270 39058
rect 2322 39006 2324 39058
rect 2268 38052 2324 39006
rect 2380 39058 2436 40908
rect 2492 40626 2548 41020
rect 2492 40574 2494 40626
rect 2546 40574 2548 40626
rect 2492 40562 2548 40574
rect 2604 40516 2660 41580
rect 2828 40628 2884 41580
rect 2828 40562 2884 40572
rect 3164 41412 3220 41422
rect 2604 40450 2660 40460
rect 2380 39006 2382 39058
rect 2434 39006 2436 39058
rect 2380 38994 2436 39006
rect 2492 40404 2548 40414
rect 2492 39058 2548 40348
rect 2716 40402 2772 40414
rect 2716 40350 2718 40402
rect 2770 40350 2772 40402
rect 2604 40292 2660 40302
rect 2604 40198 2660 40236
rect 2716 39396 2772 40350
rect 3164 40402 3220 41356
rect 3164 40350 3166 40402
rect 3218 40350 3220 40402
rect 3164 40338 3220 40350
rect 3388 40292 3444 42364
rect 3612 41972 3668 43036
rect 4060 42868 4116 42878
rect 3724 42866 4116 42868
rect 3724 42814 4062 42866
rect 4114 42814 4116 42866
rect 3724 42812 4116 42814
rect 3724 42642 3780 42812
rect 4060 42802 4116 42812
rect 4172 42868 4228 44158
rect 4172 42802 4228 42812
rect 4284 44100 4340 44110
rect 3724 42590 3726 42642
rect 3778 42590 3780 42642
rect 3724 42578 3780 42590
rect 3948 42644 4004 42654
rect 3612 41906 3668 41916
rect 3836 42530 3892 42542
rect 3836 42478 3838 42530
rect 3890 42478 3892 42530
rect 3836 41970 3892 42478
rect 3836 41918 3838 41970
rect 3890 41918 3892 41970
rect 3836 41906 3892 41918
rect 3948 41748 4004 42588
rect 4172 42644 4228 42654
rect 4172 42550 4228 42588
rect 3388 40226 3444 40236
rect 3500 41692 4004 41748
rect 4060 42420 4116 42430
rect 4284 42420 4340 44044
rect 4396 43428 4452 44268
rect 4732 44324 4788 44334
rect 4732 44230 4788 44268
rect 4508 43428 4564 43438
rect 4396 43372 4508 43428
rect 4508 43362 4564 43372
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4396 42754 4452 42766
rect 4396 42702 4398 42754
rect 4450 42702 4452 42754
rect 4396 42420 4452 42702
rect 4956 42756 5012 46956
rect 5068 45666 5124 47068
rect 5180 46788 5236 47404
rect 5180 46722 5236 46732
rect 5068 45614 5070 45666
rect 5122 45614 5124 45666
rect 5068 45444 5124 45614
rect 5068 45378 5124 45388
rect 5404 44548 5460 52894
rect 5516 52946 5572 53564
rect 5516 52894 5518 52946
rect 5570 52894 5572 52946
rect 5516 52882 5572 52894
rect 5628 53618 5684 53630
rect 5628 53566 5630 53618
rect 5682 53566 5684 53618
rect 5628 52500 5684 53566
rect 5852 53620 5908 53630
rect 5908 53564 6020 53620
rect 5852 53554 5908 53564
rect 5740 53508 5796 53518
rect 5740 53414 5796 53452
rect 5964 53506 6020 53564
rect 5964 53454 5966 53506
rect 6018 53454 6020 53506
rect 5964 53442 6020 53454
rect 6076 53396 6132 53788
rect 6076 53330 6132 53340
rect 6188 53058 6244 54572
rect 6188 53006 6190 53058
rect 6242 53006 6244 53058
rect 6188 52994 6244 53006
rect 6300 54402 6356 56030
rect 6748 55468 6804 56924
rect 7084 56868 7140 56878
rect 7084 56774 7140 56812
rect 6748 55412 6916 55468
rect 6636 55300 6692 55310
rect 6636 55206 6692 55244
rect 6300 54350 6302 54402
rect 6354 54350 6356 54402
rect 5628 52434 5684 52444
rect 5852 52724 5908 52734
rect 5852 50484 5908 52668
rect 6300 52162 6356 54350
rect 6636 53844 6692 53854
rect 6860 53844 6916 55412
rect 7196 55076 7252 55086
rect 7196 53954 7252 55020
rect 7196 53902 7198 53954
rect 7250 53902 7252 53954
rect 7196 53890 7252 53902
rect 6636 53842 6916 53844
rect 6636 53790 6638 53842
rect 6690 53790 6916 53842
rect 6636 53788 6916 53790
rect 6636 53778 6692 53788
rect 6972 53732 7028 53742
rect 6972 53730 7140 53732
rect 6972 53678 6974 53730
rect 7026 53678 7140 53730
rect 6972 53676 7140 53678
rect 6972 53666 7028 53676
rect 6524 53620 6580 53630
rect 6524 53526 6580 53564
rect 6748 53508 6804 53518
rect 6748 53414 6804 53452
rect 6972 53396 7028 53406
rect 6748 52946 6804 52958
rect 6748 52894 6750 52946
rect 6802 52894 6804 52946
rect 6300 52110 6302 52162
rect 6354 52110 6356 52162
rect 6300 52098 6356 52110
rect 6412 52834 6468 52846
rect 6412 52782 6414 52834
rect 6466 52782 6468 52834
rect 6412 52164 6468 52782
rect 6748 52836 6804 52894
rect 6860 52836 6916 52846
rect 6748 52780 6860 52836
rect 6860 52770 6916 52780
rect 6468 52108 6804 52164
rect 6412 52098 6468 52108
rect 6300 51380 6356 51390
rect 6356 51324 6468 51380
rect 6300 51286 6356 51324
rect 6300 50596 6356 50606
rect 6076 50484 6132 50494
rect 5852 50428 6076 50484
rect 6076 50370 6132 50428
rect 6076 50318 6078 50370
rect 6130 50318 6132 50370
rect 6076 49812 6132 50318
rect 6076 49746 6132 49756
rect 6300 49364 6356 50540
rect 6412 49812 6468 51324
rect 6748 51378 6804 52108
rect 6972 51490 7028 53340
rect 6972 51438 6974 51490
rect 7026 51438 7028 51490
rect 6972 51426 7028 51438
rect 6748 51326 6750 51378
rect 6802 51326 6804 51378
rect 6748 50428 6804 51326
rect 6748 50372 7028 50428
rect 6860 49812 6916 49822
rect 6412 49810 6916 49812
rect 6412 49758 6862 49810
rect 6914 49758 6916 49810
rect 6412 49756 6916 49758
rect 6300 49308 6580 49364
rect 5964 49252 6020 49262
rect 5964 49158 6020 49196
rect 6300 49026 6356 49308
rect 6300 48974 6302 49026
rect 6354 48974 6356 49026
rect 6300 48962 6356 48974
rect 6412 49140 6468 49150
rect 6412 48804 6468 49084
rect 6188 48748 6468 48804
rect 6188 47572 6244 48748
rect 5964 47570 6244 47572
rect 5964 47518 6190 47570
rect 6242 47518 6244 47570
rect 5964 47516 6244 47518
rect 5852 47460 5908 47470
rect 5852 47366 5908 47404
rect 5516 46788 5572 46798
rect 5516 46694 5572 46732
rect 5964 46562 6020 47516
rect 6188 47506 6244 47516
rect 5964 46510 5966 46562
rect 6018 46510 6020 46562
rect 5964 46498 6020 46510
rect 6188 46674 6244 46686
rect 6188 46622 6190 46674
rect 6242 46622 6244 46674
rect 6188 46564 6244 46622
rect 6076 45668 6132 45678
rect 5404 44492 5796 44548
rect 4956 42700 5236 42756
rect 5180 42644 5236 42700
rect 5180 42588 5348 42644
rect 4844 42532 4900 42542
rect 2828 39732 2884 39742
rect 2828 39638 2884 39676
rect 3052 39732 3108 39742
rect 2716 39330 2772 39340
rect 2492 39006 2494 39058
rect 2546 39006 2548 39058
rect 2492 38052 2548 39006
rect 3052 38946 3108 39676
rect 3500 39732 3556 41692
rect 3612 41300 3668 41310
rect 3612 40626 3668 41244
rect 3612 40574 3614 40626
rect 3666 40574 3668 40626
rect 3612 40516 3668 40574
rect 3612 40450 3668 40460
rect 3724 40628 3780 40638
rect 3724 40290 3780 40572
rect 3724 40238 3726 40290
rect 3778 40238 3780 40290
rect 3724 40226 3780 40238
rect 3836 40180 3892 40190
rect 3836 40178 4004 40180
rect 3836 40126 3838 40178
rect 3890 40126 4004 40178
rect 3836 40124 4004 40126
rect 3836 40114 3892 40124
rect 3500 39666 3556 39676
rect 3836 39844 3892 39854
rect 3836 39730 3892 39788
rect 3836 39678 3838 39730
rect 3890 39678 3892 39730
rect 3836 39666 3892 39678
rect 3276 39620 3332 39630
rect 3164 39564 3276 39620
rect 3164 39058 3220 39564
rect 3276 39554 3332 39564
rect 3164 39006 3166 39058
rect 3218 39006 3220 39058
rect 3164 38994 3220 39006
rect 3276 39396 3332 39406
rect 3052 38894 3054 38946
rect 3106 38894 3108 38946
rect 3052 38882 3108 38894
rect 2828 38834 2884 38846
rect 3276 38836 3332 39340
rect 3948 38946 4004 40124
rect 3948 38894 3950 38946
rect 4002 38894 4004 38946
rect 3948 38882 4004 38894
rect 2828 38782 2830 38834
rect 2882 38782 2884 38834
rect 2268 37996 2436 38052
rect 2156 37940 2212 37950
rect 2156 37846 2212 37884
rect 2268 37826 2324 37838
rect 2268 37774 2270 37826
rect 2322 37774 2324 37826
rect 2268 37380 2324 37774
rect 2268 37314 2324 37324
rect 2156 37268 2212 37278
rect 2044 37266 2212 37268
rect 2044 37214 2158 37266
rect 2210 37214 2212 37266
rect 2044 37212 2212 37214
rect 2156 37202 2212 37212
rect 1932 37154 1988 37166
rect 1932 37102 1934 37154
rect 1986 37102 1988 37154
rect 1932 37044 1988 37102
rect 2380 37044 2436 37996
rect 2716 38612 2772 38622
rect 2716 38052 2772 38556
rect 2828 38276 2884 38782
rect 3164 38780 3332 38836
rect 3500 38834 3556 38846
rect 3500 38782 3502 38834
rect 3554 38782 3556 38834
rect 2828 38220 2996 38276
rect 2828 38052 2884 38062
rect 2716 37996 2828 38052
rect 2492 37986 2548 37996
rect 2828 37958 2884 37996
rect 1932 36988 2436 37044
rect 2492 37826 2548 37838
rect 2492 37774 2494 37826
rect 2546 37774 2548 37826
rect 2492 37044 2548 37774
rect 2940 37380 2996 38220
rect 2940 37314 2996 37324
rect 1820 36876 2100 36932
rect 2044 36706 2100 36876
rect 2044 36654 2046 36706
rect 2098 36654 2100 36706
rect 1932 36372 1988 36382
rect 1932 34130 1988 36316
rect 2044 36260 2100 36654
rect 2044 36194 2100 36204
rect 2156 36036 2212 36988
rect 2492 36978 2548 36988
rect 1932 34078 1934 34130
rect 1986 34078 1988 34130
rect 1932 33348 1988 34078
rect 1932 33282 1988 33292
rect 2044 35980 2212 36036
rect 2268 36820 2324 36830
rect 1708 33068 1988 33124
rect 1708 32564 1764 32574
rect 1708 31948 1764 32508
rect 1708 31892 1876 31948
rect 1820 31890 1876 31892
rect 1820 31838 1822 31890
rect 1874 31838 1876 31890
rect 1820 31826 1876 31838
rect 1932 31332 1988 33068
rect 1932 31266 1988 31276
rect 2044 30996 2100 35980
rect 2268 35140 2324 36764
rect 3164 36820 3220 38780
rect 3500 38668 3556 38782
rect 3500 38612 3892 38668
rect 3276 38050 3332 38062
rect 3276 37998 3278 38050
rect 3330 37998 3332 38050
rect 3276 37828 3332 37998
rect 3500 38052 3556 38062
rect 3276 37772 3444 37828
rect 3164 36754 3220 36764
rect 3276 37604 3332 37614
rect 2380 36596 2436 36606
rect 2380 36594 2996 36596
rect 2380 36542 2382 36594
rect 2434 36542 2996 36594
rect 2380 36540 2996 36542
rect 2380 36530 2436 36540
rect 2604 36372 2660 36382
rect 2604 36278 2660 36316
rect 2492 36260 2548 36270
rect 2492 35924 2548 36204
rect 2492 35830 2548 35868
rect 2604 35924 2660 35934
rect 2716 35924 2772 36540
rect 2940 36482 2996 36540
rect 2940 36430 2942 36482
rect 2994 36430 2996 36482
rect 2940 36418 2996 36430
rect 2604 35922 2772 35924
rect 2604 35870 2606 35922
rect 2658 35870 2772 35922
rect 2604 35868 2772 35870
rect 2604 35858 2660 35868
rect 2828 35812 2884 35822
rect 2716 35810 2884 35812
rect 2716 35758 2830 35810
rect 2882 35758 2884 35810
rect 2716 35756 2884 35758
rect 2380 35140 2436 35150
rect 2268 35138 2436 35140
rect 2268 35086 2382 35138
rect 2434 35086 2436 35138
rect 2268 35084 2436 35086
rect 2380 35074 2436 35084
rect 2716 34244 2772 35756
rect 2828 35746 2884 35756
rect 2940 35700 2996 35710
rect 2940 35698 3220 35700
rect 2940 35646 2942 35698
rect 2994 35646 3220 35698
rect 2940 35644 3220 35646
rect 2940 35634 2996 35644
rect 3052 34916 3108 34926
rect 2828 34914 3108 34916
rect 2828 34862 3054 34914
rect 3106 34862 3108 34914
rect 2828 34860 3108 34862
rect 2828 34354 2884 34860
rect 3052 34850 3108 34860
rect 2828 34302 2830 34354
rect 2882 34302 2884 34354
rect 2828 34290 2884 34302
rect 2156 34188 2772 34244
rect 2156 34130 2212 34188
rect 2156 34078 2158 34130
rect 2210 34078 2212 34130
rect 2156 34066 2212 34078
rect 1820 30940 2100 30996
rect 2268 32674 2324 34188
rect 2380 33908 2436 33918
rect 3164 33908 3220 35644
rect 2380 33906 3220 33908
rect 2380 33854 2382 33906
rect 2434 33854 3220 33906
rect 2380 33852 3220 33854
rect 2380 33842 2436 33852
rect 2268 32622 2270 32674
rect 2322 32622 2324 32674
rect 2268 30994 2324 32622
rect 2492 33348 2548 33358
rect 2492 31780 2548 33292
rect 2604 33346 2660 33358
rect 2604 33294 2606 33346
rect 2658 33294 2660 33346
rect 2604 32562 2660 33294
rect 3164 33234 3220 33852
rect 3164 33182 3166 33234
rect 3218 33182 3220 33234
rect 3164 32676 3220 33182
rect 2604 32510 2606 32562
rect 2658 32510 2660 32562
rect 2604 31948 2660 32510
rect 2940 32674 3220 32676
rect 2940 32622 3166 32674
rect 3218 32622 3220 32674
rect 2940 32620 3220 32622
rect 2604 31892 2772 31948
rect 2492 31778 2660 31780
rect 2492 31726 2494 31778
rect 2546 31726 2660 31778
rect 2492 31724 2660 31726
rect 2492 31714 2548 31724
rect 2604 31106 2660 31724
rect 2604 31054 2606 31106
rect 2658 31054 2660 31106
rect 2604 31042 2660 31054
rect 2716 31666 2772 31892
rect 2940 31668 2996 32620
rect 3164 32610 3220 32620
rect 3276 31948 3332 37548
rect 3388 37044 3444 37772
rect 3388 36978 3444 36988
rect 3388 36708 3444 36718
rect 3500 36708 3556 37996
rect 3724 37380 3780 37390
rect 3388 36706 3556 36708
rect 3388 36654 3390 36706
rect 3442 36654 3556 36706
rect 3388 36652 3556 36654
rect 3612 37154 3668 37166
rect 3612 37102 3614 37154
rect 3666 37102 3668 37154
rect 3388 36642 3444 36652
rect 3612 36484 3668 37102
rect 3612 36390 3668 36428
rect 3500 35924 3556 35934
rect 3500 35830 3556 35868
rect 3612 34244 3668 34254
rect 3612 33458 3668 34188
rect 3724 34132 3780 37324
rect 3836 36484 3892 38612
rect 4060 38162 4116 42364
rect 4172 42364 4452 42420
rect 4620 42530 4900 42532
rect 4620 42478 4846 42530
rect 4898 42478 4900 42530
rect 4620 42476 4900 42478
rect 4172 39396 4228 42364
rect 4620 42084 4676 42476
rect 4844 42466 4900 42476
rect 4956 42530 5012 42542
rect 4956 42478 4958 42530
rect 5010 42478 5012 42530
rect 4956 42308 5012 42478
rect 5068 42532 5124 42542
rect 5068 42530 5236 42532
rect 5068 42478 5070 42530
rect 5122 42478 5236 42530
rect 5068 42476 5236 42478
rect 5068 42466 5124 42476
rect 4956 42252 5124 42308
rect 4956 42084 5012 42094
rect 4620 42028 4900 42084
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4620 41300 4676 41310
rect 4620 41206 4676 41244
rect 4396 40628 4452 40638
rect 4844 40628 4900 42028
rect 4396 40626 4900 40628
rect 4396 40574 4398 40626
rect 4450 40574 4900 40626
rect 4396 40572 4900 40574
rect 4396 40562 4452 40572
rect 4844 40402 4900 40414
rect 4844 40350 4846 40402
rect 4898 40350 4900 40402
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4508 39844 4564 39854
rect 4508 39730 4564 39788
rect 4508 39678 4510 39730
rect 4562 39678 4564 39730
rect 4508 39666 4564 39678
rect 4732 39618 4788 39630
rect 4732 39566 4734 39618
rect 4786 39566 4788 39618
rect 4172 39330 4228 39340
rect 4284 39394 4340 39406
rect 4284 39342 4286 39394
rect 4338 39342 4340 39394
rect 4284 39172 4340 39342
rect 4284 39106 4340 39116
rect 4732 38612 4788 39566
rect 4844 39620 4900 40350
rect 4844 39554 4900 39564
rect 4956 38668 5012 42028
rect 5068 41412 5124 42252
rect 5068 41346 5124 41356
rect 5068 40964 5124 40974
rect 5068 40870 5124 40908
rect 5068 39844 5124 39854
rect 5180 39844 5236 42476
rect 5068 39842 5236 39844
rect 5068 39790 5070 39842
rect 5122 39790 5236 39842
rect 5068 39788 5236 39790
rect 5068 39778 5124 39788
rect 5292 39732 5348 42588
rect 5628 40740 5684 40750
rect 5628 40514 5684 40684
rect 5628 40462 5630 40514
rect 5682 40462 5684 40514
rect 5628 40450 5684 40462
rect 5292 39666 5348 39676
rect 5516 40402 5572 40414
rect 5516 40350 5518 40402
rect 5570 40350 5572 40402
rect 4732 38546 4788 38556
rect 4844 38612 5012 38668
rect 5180 38612 5236 38622
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4060 38110 4062 38162
rect 4114 38110 4116 38162
rect 4060 38098 4116 38110
rect 4396 38052 4452 38062
rect 4284 37938 4340 37950
rect 4284 37886 4286 37938
rect 4338 37886 4340 37938
rect 4284 37492 4340 37886
rect 4284 37426 4340 37436
rect 4396 37380 4452 37996
rect 4620 37940 4676 37950
rect 4620 37846 4676 37884
rect 4844 37828 4900 38612
rect 5068 38556 5180 38612
rect 4956 38052 5012 38062
rect 5068 38052 5124 38556
rect 5180 38546 5236 38556
rect 5012 37996 5124 38052
rect 4956 37958 5012 37996
rect 4844 37826 5012 37828
rect 4844 37774 4846 37826
rect 4898 37774 5012 37826
rect 4844 37772 5012 37774
rect 4844 37762 4900 37772
rect 4396 37314 4452 37324
rect 4476 36876 4740 36886
rect 4284 36820 4340 36830
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 3836 36418 3892 36428
rect 4060 36708 4116 36718
rect 3948 34802 4004 34814
rect 3948 34750 3950 34802
rect 4002 34750 4004 34802
rect 3948 34356 4004 34750
rect 3948 34290 4004 34300
rect 3948 34132 4004 34142
rect 3724 34130 4004 34132
rect 3724 34078 3950 34130
rect 4002 34078 4004 34130
rect 3724 34076 4004 34078
rect 3948 33572 4004 34076
rect 3948 33506 4004 33516
rect 3612 33406 3614 33458
rect 3666 33406 3668 33458
rect 3612 33394 3668 33406
rect 2716 31614 2718 31666
rect 2770 31614 2772 31666
rect 2268 30942 2270 30994
rect 2322 30942 2324 30994
rect 1820 26068 1876 30940
rect 2268 29426 2324 30942
rect 2492 30770 2548 30782
rect 2492 30718 2494 30770
rect 2546 30718 2548 30770
rect 2492 30100 2548 30718
rect 2716 30100 2772 31614
rect 2828 31666 2996 31668
rect 2828 31614 2942 31666
rect 2994 31614 2996 31666
rect 2828 31612 2996 31614
rect 2828 30324 2884 31612
rect 2940 31602 2996 31612
rect 3164 31892 3332 31948
rect 3948 32340 4004 32350
rect 3052 31332 3108 31342
rect 2828 30258 2884 30268
rect 2940 31106 2996 31118
rect 2940 31054 2942 31106
rect 2994 31054 2996 31106
rect 2940 30210 2996 31054
rect 3052 30996 3108 31276
rect 3164 31220 3220 31892
rect 3276 31780 3332 31790
rect 3276 31686 3332 31724
rect 3948 31778 4004 32284
rect 3948 31726 3950 31778
rect 4002 31726 4004 31778
rect 3948 31714 4004 31726
rect 3724 31668 3780 31678
rect 3164 31154 3220 31164
rect 3612 31666 3780 31668
rect 3612 31614 3726 31666
rect 3778 31614 3780 31666
rect 3612 31612 3780 31614
rect 3164 30996 3220 31006
rect 3052 30994 3220 30996
rect 3052 30942 3166 30994
rect 3218 30942 3220 30994
rect 3052 30940 3220 30942
rect 2940 30158 2942 30210
rect 2994 30158 2996 30210
rect 2828 30100 2884 30110
rect 2492 30098 2884 30100
rect 2492 30046 2830 30098
rect 2882 30046 2884 30098
rect 2492 30044 2884 30046
rect 2268 29374 2270 29426
rect 2322 29374 2324 29426
rect 2268 29362 2324 29374
rect 1932 29314 1988 29326
rect 1932 29262 1934 29314
rect 1986 29262 1988 29314
rect 1932 28756 1988 29262
rect 1932 28530 1988 28700
rect 2828 28644 2884 30044
rect 2940 29428 2996 30158
rect 2940 29362 2996 29372
rect 3052 29538 3108 29550
rect 3052 29486 3054 29538
rect 3106 29486 3108 29538
rect 2940 28644 2996 28654
rect 2828 28642 2996 28644
rect 2828 28590 2942 28642
rect 2994 28590 2996 28642
rect 2828 28588 2996 28590
rect 1932 28478 1934 28530
rect 1986 28478 1988 28530
rect 1932 28466 1988 28478
rect 2156 28530 2212 28542
rect 2156 28478 2158 28530
rect 2210 28478 2212 28530
rect 2044 28418 2100 28430
rect 2044 28366 2046 28418
rect 2098 28366 2100 28418
rect 2044 28196 2100 28366
rect 2156 28420 2212 28478
rect 2156 28354 2212 28364
rect 2044 28140 2884 28196
rect 2716 27972 2772 27982
rect 2156 27860 2212 27870
rect 2156 27766 2212 27804
rect 2716 27858 2772 27916
rect 2828 27970 2884 28140
rect 2828 27918 2830 27970
rect 2882 27918 2884 27970
rect 2828 27906 2884 27918
rect 2716 27806 2718 27858
rect 2770 27806 2772 27858
rect 2716 27794 2772 27806
rect 2604 27636 2660 27646
rect 2156 27524 2212 27534
rect 2156 26514 2212 27468
rect 2604 26516 2660 27580
rect 2940 27074 2996 28588
rect 2940 27022 2942 27074
rect 2994 27022 2996 27074
rect 2940 27010 2996 27022
rect 3052 28530 3108 29486
rect 3052 28478 3054 28530
rect 3106 28478 3108 28530
rect 3052 27186 3108 28478
rect 3164 28308 3220 30940
rect 3388 30996 3444 31006
rect 3388 29764 3444 30940
rect 3388 28754 3444 29708
rect 3388 28702 3390 28754
rect 3442 28702 3444 28754
rect 3164 28252 3332 28308
rect 3164 28084 3220 28094
rect 3164 27860 3220 28028
rect 3164 27794 3220 27804
rect 3276 27636 3332 28252
rect 3052 27134 3054 27186
rect 3106 27134 3108 27186
rect 2156 26462 2158 26514
rect 2210 26462 2212 26514
rect 2156 26450 2212 26462
rect 2492 26514 2660 26516
rect 2492 26462 2606 26514
rect 2658 26462 2660 26514
rect 2492 26460 2660 26462
rect 2268 26292 2324 26302
rect 2268 26198 2324 26236
rect 1820 26012 1988 26068
rect 1820 23154 1876 23166
rect 1820 23102 1822 23154
rect 1874 23102 1876 23154
rect 1708 22708 1764 22718
rect 1708 21700 1764 22652
rect 1820 22484 1876 23102
rect 1820 22418 1876 22428
rect 1708 21698 1876 21700
rect 1708 21646 1710 21698
rect 1762 21646 1876 21698
rect 1708 21644 1876 21646
rect 1708 21634 1764 21644
rect 1820 20914 1876 21644
rect 1820 20862 1822 20914
rect 1874 20862 1876 20914
rect 1820 20850 1876 20862
rect 1932 20188 1988 26012
rect 2380 25620 2436 25630
rect 2492 25620 2548 26460
rect 2604 26450 2660 26460
rect 3052 26292 3108 27134
rect 3052 26178 3108 26236
rect 3052 26126 3054 26178
rect 3106 26126 3108 26178
rect 3052 26114 3108 26126
rect 3164 27580 3332 27636
rect 3164 25956 3220 27580
rect 3276 26964 3332 26974
rect 3276 26870 3332 26908
rect 2380 25618 2548 25620
rect 2380 25566 2382 25618
rect 2434 25566 2548 25618
rect 2380 25564 2548 25566
rect 2828 25900 3220 25956
rect 2380 25554 2436 25564
rect 2380 24948 2436 24958
rect 2380 24050 2436 24892
rect 2380 23998 2382 24050
rect 2434 23998 2436 24050
rect 2380 23986 2436 23998
rect 2268 23940 2324 23950
rect 2268 23846 2324 23884
rect 2716 23828 2772 23838
rect 2604 23826 2772 23828
rect 2604 23774 2718 23826
rect 2770 23774 2772 23826
rect 2604 23772 2772 23774
rect 2492 23044 2548 23054
rect 2268 23042 2548 23044
rect 2268 22990 2494 23042
rect 2546 22990 2548 23042
rect 2268 22988 2548 22990
rect 2156 22372 2212 22382
rect 2044 22370 2212 22372
rect 2044 22318 2158 22370
rect 2210 22318 2212 22370
rect 2044 22316 2212 22318
rect 2044 21810 2100 22316
rect 2156 22306 2212 22316
rect 2044 21758 2046 21810
rect 2098 21758 2100 21810
rect 2044 21746 2100 21758
rect 2268 21810 2324 22988
rect 2492 22978 2548 22988
rect 2268 21758 2270 21810
rect 2322 21758 2324 21810
rect 2268 21746 2324 21758
rect 2492 21698 2548 21710
rect 2492 21646 2494 21698
rect 2546 21646 2548 21698
rect 2492 21588 2548 21646
rect 2604 21698 2660 23772
rect 2716 23762 2772 23772
rect 2604 21646 2606 21698
rect 2658 21646 2660 21698
rect 2604 21634 2660 21646
rect 2268 21532 2492 21588
rect 2156 20244 2212 20254
rect 2268 20244 2324 21532
rect 2492 21522 2548 21532
rect 2828 21476 2884 25900
rect 2156 20242 2324 20244
rect 2156 20190 2158 20242
rect 2210 20190 2324 20242
rect 2156 20188 2324 20190
rect 2604 21420 2884 21476
rect 2940 24948 2996 24958
rect 2604 20188 2660 21420
rect 2940 20188 2996 24892
rect 3388 24836 3444 28702
rect 3612 27746 3668 31612
rect 3724 31602 3780 31612
rect 4060 31554 4116 36652
rect 4284 35140 4340 36764
rect 4844 36596 4900 36606
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4284 35084 4452 35140
rect 4172 35028 4228 35038
rect 4172 35026 4340 35028
rect 4172 34974 4174 35026
rect 4226 34974 4340 35026
rect 4172 34972 4340 34974
rect 4172 34962 4228 34972
rect 4172 34804 4228 34814
rect 4172 34710 4228 34748
rect 4284 34018 4340 34972
rect 4396 34242 4452 35084
rect 4844 35138 4900 36540
rect 4844 35086 4846 35138
rect 4898 35086 4900 35138
rect 4844 35074 4900 35086
rect 4956 35028 5012 37772
rect 5180 37492 5236 37502
rect 5180 37398 5236 37436
rect 5516 36596 5572 40350
rect 5740 40292 5796 44492
rect 5964 44322 6020 44334
rect 5964 44270 5966 44322
rect 6018 44270 6020 44322
rect 5964 43988 6020 44270
rect 6076 43988 6132 45612
rect 6188 44436 6244 46508
rect 6188 44322 6244 44380
rect 6300 46676 6356 46686
rect 6300 44434 6356 46620
rect 6412 45668 6468 45678
rect 6524 45668 6580 49308
rect 6860 49026 6916 49756
rect 6972 49140 7028 50372
rect 6972 49074 7028 49084
rect 6860 48974 6862 49026
rect 6914 48974 6916 49026
rect 6748 48020 6804 48030
rect 6748 47684 6804 47964
rect 6748 47590 6804 47628
rect 6860 46900 6916 48974
rect 7084 47796 7140 53676
rect 7308 51604 7364 57484
rect 7532 56868 7588 56878
rect 7532 56774 7588 56812
rect 7868 55468 7924 62132
rect 8316 61572 8372 63086
rect 9548 63026 9604 63038
rect 9548 62974 9550 63026
rect 9602 62974 9604 63026
rect 9436 62914 9492 62926
rect 9436 62862 9438 62914
rect 9490 62862 9492 62914
rect 8316 61506 8372 61516
rect 8652 62580 8708 62590
rect 8652 61348 8708 62524
rect 9436 62580 9492 62862
rect 9436 62514 9492 62524
rect 9436 61572 9492 61582
rect 9436 61478 9492 61516
rect 8876 61460 8932 61470
rect 8764 61348 8820 61358
rect 8652 61346 8820 61348
rect 8652 61294 8766 61346
rect 8818 61294 8820 61346
rect 8652 61292 8820 61294
rect 8652 60676 8708 61292
rect 8764 61282 8820 61292
rect 8764 60788 8820 60798
rect 8876 60788 8932 61404
rect 9548 61460 9604 62974
rect 10332 62356 10388 62366
rect 10556 62356 10612 63868
rect 10780 63858 10836 63868
rect 10332 62354 10612 62356
rect 10332 62302 10334 62354
rect 10386 62302 10612 62354
rect 10332 62300 10612 62302
rect 10332 62290 10388 62300
rect 9548 61394 9604 61404
rect 8820 60732 8932 60788
rect 8764 60694 8820 60732
rect 8652 60582 8708 60620
rect 10556 59220 10612 62300
rect 11452 63700 11508 64428
rect 12012 64484 12068 65326
rect 12012 64418 12068 64428
rect 12124 65380 12180 65438
rect 12460 65492 12516 66222
rect 13356 66274 13524 66276
rect 13356 66222 13470 66274
rect 13522 66222 13524 66274
rect 13356 66220 13524 66222
rect 12460 65426 12516 65436
rect 13020 65492 13076 65502
rect 13132 65492 13188 65502
rect 13356 65492 13412 66220
rect 13468 66210 13524 66220
rect 13076 65490 13412 65492
rect 13076 65438 13134 65490
rect 13186 65438 13412 65490
rect 13076 65436 13412 65438
rect 14364 65714 14420 66332
rect 14700 66322 14756 66332
rect 14364 65662 14366 65714
rect 14418 65662 14420 65714
rect 12124 64036 12180 65324
rect 11452 62242 11508 63644
rect 11452 62190 11454 62242
rect 11506 62190 11508 62242
rect 10780 61460 10836 61470
rect 10780 61366 10836 61404
rect 10668 61346 10724 61358
rect 10668 61294 10670 61346
rect 10722 61294 10724 61346
rect 10668 60676 10724 61294
rect 11452 60676 11508 62190
rect 11676 63980 12180 64036
rect 11676 62354 11732 63980
rect 12124 63924 12180 63980
rect 12124 63830 12180 63868
rect 11900 63810 11956 63822
rect 11900 63758 11902 63810
rect 11954 63758 11956 63810
rect 11788 63700 11844 63710
rect 11900 63700 11956 63758
rect 11844 63644 11956 63700
rect 11788 63634 11844 63644
rect 11676 62302 11678 62354
rect 11730 62302 11732 62354
rect 11676 61572 11732 62302
rect 13020 62354 13076 65436
rect 13132 65426 13188 65436
rect 13020 62302 13022 62354
rect 13074 62302 13076 62354
rect 13020 62188 13076 62302
rect 13468 63138 13524 63150
rect 13468 63086 13470 63138
rect 13522 63086 13524 63138
rect 13468 62188 13524 63086
rect 14252 62580 14308 62590
rect 14364 62580 14420 65662
rect 14812 66162 14868 66174
rect 14812 66110 14814 66162
rect 14866 66110 14868 66162
rect 14252 62578 14420 62580
rect 14252 62526 14254 62578
rect 14306 62526 14420 62578
rect 14252 62524 14420 62526
rect 14476 65492 14532 65502
rect 14812 65492 14868 66110
rect 14476 65490 14868 65492
rect 14476 65438 14478 65490
rect 14530 65438 14868 65490
rect 14476 65436 14868 65438
rect 14476 63924 14532 65436
rect 14476 63140 14532 63868
rect 16380 63252 16436 63262
rect 16380 63158 16436 63196
rect 14812 63140 14868 63150
rect 14476 63138 14868 63140
rect 14476 63086 14814 63138
rect 14866 63086 14868 63138
rect 14476 63084 14868 63086
rect 14252 62188 14308 62524
rect 14476 62354 14532 63084
rect 14476 62302 14478 62354
rect 14530 62302 14532 62354
rect 14476 62290 14532 62302
rect 14700 62914 14756 62926
rect 14700 62862 14702 62914
rect 14754 62862 14756 62914
rect 13020 62132 13524 62188
rect 11676 61516 11956 61572
rect 11676 60676 11732 60686
rect 11452 60620 11676 60676
rect 10668 60610 10724 60620
rect 11676 60564 11732 60620
rect 11676 60508 11844 60564
rect 10668 59220 10724 59230
rect 10556 59164 10668 59220
rect 10668 58434 10724 59164
rect 11788 59108 11844 60508
rect 11900 59332 11956 61516
rect 13468 61570 13524 62132
rect 13468 61518 13470 61570
rect 13522 61518 13524 61570
rect 13468 61506 13524 61518
rect 14140 62132 14308 62188
rect 14140 61684 14196 62132
rect 14700 61684 14756 62862
rect 14140 61682 14756 61684
rect 14140 61630 14702 61682
rect 14754 61630 14756 61682
rect 14140 61628 14756 61630
rect 12012 59332 12068 59342
rect 11900 59276 12012 59332
rect 11900 59108 11956 59118
rect 11788 59106 11956 59108
rect 11788 59054 11902 59106
rect 11954 59054 11956 59106
rect 11788 59052 11956 59054
rect 10668 58382 10670 58434
rect 10722 58382 10724 58434
rect 10668 58370 10724 58382
rect 10892 58436 10948 58446
rect 7756 55412 7924 55468
rect 7980 57876 8036 57886
rect 7980 57650 8036 57820
rect 10892 57762 10948 58380
rect 10892 57710 10894 57762
rect 10946 57710 10948 57762
rect 10892 57698 10948 57710
rect 11900 58210 11956 59052
rect 12012 58436 12068 59276
rect 12012 58342 12068 58380
rect 12124 59220 12180 59230
rect 11900 58158 11902 58210
rect 11954 58158 11956 58210
rect 11900 57876 11956 58158
rect 7980 57598 7982 57650
rect 8034 57598 8036 57650
rect 7980 57092 8036 57598
rect 8988 57650 9044 57662
rect 8988 57598 8990 57650
rect 9042 57598 9044 57650
rect 7980 56306 8036 57036
rect 8316 57092 8372 57102
rect 8316 56866 8372 57036
rect 8316 56814 8318 56866
rect 8370 56814 8372 56866
rect 8316 56802 8372 56814
rect 8988 56868 9044 57598
rect 11004 57538 11060 57550
rect 11004 57486 11006 57538
rect 11058 57486 11060 57538
rect 9548 57092 9604 57102
rect 10780 57092 10836 57102
rect 11004 57092 11060 57486
rect 9604 57036 9716 57092
rect 9548 56998 9604 57036
rect 7980 56254 7982 56306
rect 8034 56254 8036 56306
rect 7980 55524 8036 56254
rect 8988 55468 9044 56812
rect 9660 56306 9716 57036
rect 10836 57036 11060 57092
rect 11900 57092 11956 57820
rect 12124 57650 12180 59164
rect 12124 57598 12126 57650
rect 12178 57598 12180 57650
rect 12124 57586 12180 57598
rect 12796 59220 12852 59230
rect 12796 57650 12852 59164
rect 13244 59220 13300 59230
rect 13300 59164 13412 59220
rect 13244 59154 13300 59164
rect 13356 58436 13412 59164
rect 14028 59108 14084 59118
rect 14140 59108 14196 61628
rect 14700 61618 14756 61628
rect 14812 61570 14868 63084
rect 14812 61518 14814 61570
rect 14866 61518 14868 61570
rect 14812 61506 14868 61518
rect 15596 63140 15652 63150
rect 15372 60788 15428 60798
rect 15260 60786 15428 60788
rect 15260 60734 15374 60786
rect 15426 60734 15428 60786
rect 15260 60732 15428 60734
rect 15148 60676 15204 60686
rect 15260 60676 15316 60732
rect 15372 60722 15428 60732
rect 15148 60674 15316 60676
rect 15148 60622 15150 60674
rect 15202 60622 15316 60674
rect 15148 60620 15316 60622
rect 15148 60610 15204 60620
rect 15036 60002 15092 60014
rect 15036 59950 15038 60002
rect 15090 59950 15092 60002
rect 14028 59106 14196 59108
rect 14028 59054 14030 59106
rect 14082 59054 14196 59106
rect 14028 59052 14196 59054
rect 14252 59332 14308 59342
rect 14252 59218 14308 59276
rect 14252 59166 14254 59218
rect 14306 59166 14308 59218
rect 13468 58436 13524 58446
rect 13356 58434 13524 58436
rect 13356 58382 13470 58434
rect 13522 58382 13524 58434
rect 13356 58380 13524 58382
rect 13468 58370 13524 58380
rect 14028 57876 14084 59052
rect 14028 57782 14084 57820
rect 12796 57598 12798 57650
rect 12850 57598 12852 57650
rect 12796 57586 12852 57598
rect 14252 57650 14308 59166
rect 14812 59332 14868 59342
rect 14812 58434 14868 59276
rect 15036 59108 15092 59950
rect 15036 59042 15092 59052
rect 14812 58382 14814 58434
rect 14866 58382 14868 58434
rect 14812 58370 14868 58382
rect 14700 58210 14756 58222
rect 14700 58158 14702 58210
rect 14754 58158 14756 58210
rect 14700 57876 14756 58158
rect 14700 57810 14756 57820
rect 14252 57598 14254 57650
rect 14306 57598 14308 57650
rect 14252 57586 14308 57598
rect 12124 57092 12180 57102
rect 11900 57036 12124 57092
rect 9996 56868 10052 56878
rect 9996 56774 10052 56812
rect 10780 56866 10836 57036
rect 12124 56998 12180 57036
rect 10780 56814 10782 56866
rect 10834 56814 10836 56866
rect 10780 56802 10836 56814
rect 9660 56254 9662 56306
rect 9714 56254 9716 56306
rect 9660 56242 9716 56254
rect 7644 53844 7700 53854
rect 7644 53750 7700 53788
rect 7532 53506 7588 53518
rect 7532 53454 7534 53506
rect 7586 53454 7588 53506
rect 7532 53172 7588 53454
rect 7532 53106 7588 53116
rect 7756 53506 7812 55412
rect 7980 55298 8036 55468
rect 7980 55246 7982 55298
rect 8034 55246 8036 55298
rect 7980 55234 8036 55246
rect 8876 55412 9044 55468
rect 8876 55298 8932 55412
rect 8876 55246 8878 55298
rect 8930 55246 8932 55298
rect 8876 55234 8932 55246
rect 13132 55076 13188 55086
rect 13132 54740 13188 55020
rect 12684 54738 13188 54740
rect 12684 54686 13134 54738
rect 13186 54686 13188 54738
rect 12684 54684 13188 54686
rect 7980 53956 8036 53966
rect 7980 53618 8036 53900
rect 9436 53956 9492 53966
rect 9436 53842 9492 53900
rect 9436 53790 9438 53842
rect 9490 53790 9492 53842
rect 9436 53778 9492 53790
rect 12684 53732 12740 54684
rect 13132 54674 13188 54684
rect 13804 54514 13860 54526
rect 13804 54462 13806 54514
rect 13858 54462 13860 54514
rect 13804 54404 13860 54462
rect 13804 54338 13860 54348
rect 14476 54404 14532 54414
rect 14476 54402 15092 54404
rect 14476 54350 14478 54402
rect 14530 54350 15092 54402
rect 14476 54348 15092 54350
rect 14476 54338 14532 54348
rect 14476 53732 14532 53742
rect 12684 53730 12964 53732
rect 12684 53678 12686 53730
rect 12738 53678 12964 53730
rect 12684 53676 12964 53678
rect 12684 53666 12740 53676
rect 7980 53566 7982 53618
rect 8034 53566 8036 53618
rect 7980 53554 8036 53566
rect 8540 53618 8596 53630
rect 8540 53566 8542 53618
rect 8594 53566 8596 53618
rect 7756 53454 7758 53506
rect 7810 53454 7812 53506
rect 7756 53172 7812 53454
rect 8428 53508 8484 53518
rect 8540 53508 8596 53566
rect 8988 53508 9044 53518
rect 8540 53506 9044 53508
rect 8540 53454 8990 53506
rect 9042 53454 9044 53506
rect 8540 53452 9044 53454
rect 8428 53414 8484 53452
rect 8876 53284 8932 53294
rect 7644 53060 7700 53070
rect 7196 51548 7364 51604
rect 7532 52946 7588 52958
rect 7532 52894 7534 52946
rect 7586 52894 7588 52946
rect 7196 48020 7252 51548
rect 7308 51378 7364 51390
rect 7308 51326 7310 51378
rect 7362 51326 7364 51378
rect 7308 51268 7364 51326
rect 7532 51380 7588 52894
rect 7644 52274 7700 53004
rect 7644 52222 7646 52274
rect 7698 52222 7700 52274
rect 7644 52210 7700 52222
rect 7644 51380 7700 51390
rect 7588 51378 7700 51380
rect 7588 51326 7646 51378
rect 7698 51326 7700 51378
rect 7588 51324 7700 51326
rect 7532 51314 7588 51324
rect 7644 51314 7700 51324
rect 7308 51202 7364 51212
rect 7308 50596 7364 50606
rect 7644 50596 7700 50606
rect 7308 50502 7364 50540
rect 7420 50540 7644 50596
rect 7308 49810 7364 49822
rect 7308 49758 7310 49810
rect 7362 49758 7364 49810
rect 7308 49140 7364 49758
rect 7308 49074 7364 49084
rect 7420 49140 7476 50540
rect 7644 50530 7700 50540
rect 7756 49586 7812 53116
rect 8428 53172 8484 53182
rect 8428 53078 8484 53116
rect 8876 53170 8932 53228
rect 8876 53118 8878 53170
rect 8930 53118 8932 53170
rect 8876 53106 8932 53118
rect 8092 52836 8148 52846
rect 7868 50594 7924 50606
rect 7868 50542 7870 50594
rect 7922 50542 7924 50594
rect 7868 50484 7924 50542
rect 7868 50418 7924 50428
rect 8092 49700 8148 52780
rect 8988 52052 9044 53452
rect 12124 53508 12180 53518
rect 12348 53508 12404 53518
rect 12124 53284 12180 53452
rect 11676 53228 12180 53284
rect 12236 53506 12404 53508
rect 12236 53454 12350 53506
rect 12402 53454 12404 53506
rect 12236 53452 12404 53454
rect 11116 52946 11172 52958
rect 11116 52894 11118 52946
rect 11170 52894 11172 52946
rect 8988 51986 9044 51996
rect 9660 52052 9716 52062
rect 9660 51378 9716 51996
rect 11116 52052 11172 52894
rect 11116 51986 11172 51996
rect 11228 52050 11284 52062
rect 11228 51998 11230 52050
rect 11282 51998 11284 52050
rect 10444 51940 10500 51950
rect 10332 51884 10444 51940
rect 10332 51490 10388 51884
rect 10444 51874 10500 51884
rect 10332 51438 10334 51490
rect 10386 51438 10388 51490
rect 10332 51426 10388 51438
rect 9660 51326 9662 51378
rect 9714 51326 9716 51378
rect 8540 51268 8596 51278
rect 8540 51174 8596 51212
rect 8652 50484 8708 50494
rect 9660 50484 9716 51326
rect 10780 50708 10836 50718
rect 8652 50482 9044 50484
rect 8652 50430 8654 50482
rect 8706 50430 9044 50482
rect 8652 50428 9044 50430
rect 8652 50418 8708 50428
rect 8428 49812 8484 49822
rect 8092 49634 8148 49644
rect 8316 49810 8484 49812
rect 8316 49758 8430 49810
rect 8482 49758 8484 49810
rect 8316 49756 8484 49758
rect 7756 49534 7758 49586
rect 7810 49534 7812 49586
rect 7756 49522 7812 49534
rect 7980 49140 8036 49150
rect 7420 49138 8036 49140
rect 7420 49086 7982 49138
rect 8034 49086 8036 49138
rect 7420 49084 8036 49086
rect 7420 48914 7476 49084
rect 7980 49074 8036 49084
rect 8204 49026 8260 49038
rect 8204 48974 8206 49026
rect 8258 48974 8260 49026
rect 7420 48862 7422 48914
rect 7474 48862 7476 48914
rect 7420 48850 7476 48862
rect 7644 48916 7700 48926
rect 8204 48916 8260 48974
rect 7644 48914 8260 48916
rect 7644 48862 7646 48914
rect 7698 48862 8260 48914
rect 7644 48860 8260 48862
rect 7644 48850 7700 48860
rect 7532 48804 7588 48814
rect 7532 48710 7588 48748
rect 7196 47954 7252 47964
rect 7868 48242 7924 48254
rect 7868 48190 7870 48242
rect 7922 48190 7924 48242
rect 7084 47740 7812 47796
rect 7532 47458 7588 47470
rect 7532 47406 7534 47458
rect 7586 47406 7588 47458
rect 7532 46900 7588 47406
rect 6860 46844 7588 46900
rect 6860 46674 6916 46844
rect 6860 46622 6862 46674
rect 6914 46622 6916 46674
rect 6860 46610 6916 46622
rect 7196 46674 7252 46686
rect 7196 46622 7198 46674
rect 7250 46622 7252 46674
rect 7196 46564 7252 46622
rect 7196 46498 7252 46508
rect 7420 46674 7476 46686
rect 7420 46622 7422 46674
rect 7474 46622 7476 46674
rect 6468 45612 6580 45668
rect 6860 45668 6916 45678
rect 6412 45574 6468 45612
rect 6860 45574 6916 45612
rect 7420 45668 7476 46622
rect 7420 45602 7476 45612
rect 7532 46674 7588 46686
rect 7532 46622 7534 46674
rect 7586 46622 7588 46674
rect 6300 44382 6302 44434
rect 6354 44382 6356 44434
rect 6300 44370 6356 44382
rect 6748 44436 6804 44446
rect 6748 44342 6804 44380
rect 7420 44436 7476 44446
rect 6188 44270 6190 44322
rect 6242 44270 6244 44322
rect 6188 44258 6244 44270
rect 6524 44324 6580 44334
rect 5964 43932 6076 43988
rect 6076 43922 6132 43932
rect 6412 43092 6468 43102
rect 5628 40236 5796 40292
rect 6188 42756 6244 42766
rect 5628 37490 5684 40236
rect 5852 39732 5908 39742
rect 5852 39638 5908 39676
rect 5740 39618 5796 39630
rect 5740 39566 5742 39618
rect 5794 39566 5796 39618
rect 5740 38612 5796 39566
rect 5964 39506 6020 39518
rect 5964 39454 5966 39506
rect 6018 39454 6020 39506
rect 5964 39172 6020 39454
rect 6076 39172 6132 39182
rect 5964 39116 6076 39172
rect 6076 39106 6132 39116
rect 5740 38546 5796 38556
rect 5852 38276 5908 38286
rect 5852 37826 5908 38220
rect 5852 37774 5854 37826
rect 5906 37774 5908 37826
rect 5852 37762 5908 37774
rect 6188 37492 6244 42700
rect 6300 40514 6356 40526
rect 6300 40462 6302 40514
rect 6354 40462 6356 40514
rect 6300 38612 6356 40462
rect 6412 40404 6468 43036
rect 6524 42754 6580 44268
rect 6860 43988 6916 43998
rect 6524 42702 6526 42754
rect 6578 42702 6580 42754
rect 6524 42690 6580 42702
rect 6636 43538 6692 43550
rect 6636 43486 6638 43538
rect 6690 43486 6692 43538
rect 6524 42420 6580 42430
rect 6524 41186 6580 42364
rect 6636 41860 6692 43486
rect 6748 42868 6804 42878
rect 6748 42774 6804 42812
rect 6748 41860 6804 41870
rect 6636 41804 6748 41860
rect 6748 41794 6804 41804
rect 6524 41134 6526 41186
rect 6578 41134 6580 41186
rect 6524 41122 6580 41134
rect 6412 40402 6692 40404
rect 6412 40350 6414 40402
rect 6466 40350 6692 40402
rect 6412 40348 6692 40350
rect 6412 40338 6468 40348
rect 6300 38276 6356 38556
rect 6300 38210 6356 38220
rect 5628 37438 5630 37490
rect 5682 37438 5684 37490
rect 5628 37426 5684 37438
rect 5852 37436 6244 37492
rect 6300 38050 6356 38062
rect 6300 37998 6302 38050
rect 6354 37998 6356 38050
rect 5740 36596 5796 36606
rect 5516 36530 5572 36540
rect 5628 36540 5740 36596
rect 5628 35810 5684 36540
rect 5740 36530 5796 36540
rect 5628 35758 5630 35810
rect 5682 35758 5684 35810
rect 5628 35746 5684 35758
rect 5852 35700 5908 37436
rect 6076 37266 6132 37278
rect 6076 37214 6078 37266
rect 6130 37214 6132 37266
rect 4956 34962 5012 34972
rect 5740 35698 5908 35700
rect 5740 35646 5854 35698
rect 5906 35646 5908 35698
rect 5740 35644 5908 35646
rect 4956 34802 5012 34814
rect 4956 34750 4958 34802
rect 5010 34750 5012 34802
rect 4396 34190 4398 34242
rect 4450 34190 4452 34242
rect 4396 34178 4452 34190
rect 4844 34690 4900 34702
rect 4844 34638 4846 34690
rect 4898 34638 4900 34690
rect 4844 34244 4900 34638
rect 4844 34150 4900 34188
rect 4284 33966 4286 34018
rect 4338 33966 4340 34018
rect 4284 33954 4340 33966
rect 4732 34130 4788 34142
rect 4732 34078 4734 34130
rect 4786 34078 4788 34130
rect 4732 33908 4788 34078
rect 4732 33852 4900 33908
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4508 33572 4564 33582
rect 4172 33348 4228 33358
rect 4228 33292 4452 33348
rect 4172 33254 4228 33292
rect 4396 32562 4452 33292
rect 4508 32786 4564 33516
rect 4508 32734 4510 32786
rect 4562 32734 4564 32786
rect 4508 32722 4564 32734
rect 4844 32564 4900 33852
rect 4396 32510 4398 32562
rect 4450 32510 4452 32562
rect 4396 32498 4452 32510
rect 4508 32508 4900 32564
rect 4508 32340 4564 32508
rect 4060 31502 4062 31554
rect 4114 31502 4116 31554
rect 4060 31490 4116 31502
rect 4284 32284 4564 32340
rect 4172 30996 4228 31006
rect 4172 30902 4228 30940
rect 4060 30882 4116 30894
rect 4060 30830 4062 30882
rect 4114 30830 4116 30882
rect 3612 27694 3614 27746
rect 3666 27694 3668 27746
rect 3612 27682 3668 27694
rect 3724 30322 3780 30334
rect 3724 30270 3726 30322
rect 3778 30270 3780 30322
rect 3724 30212 3780 30270
rect 3724 27970 3780 30156
rect 4060 30210 4116 30830
rect 4060 30158 4062 30210
rect 4114 30158 4116 30210
rect 3836 29314 3892 29326
rect 3836 29262 3838 29314
rect 3890 29262 3892 29314
rect 3836 28196 3892 29262
rect 3836 28130 3892 28140
rect 4060 28084 4116 30158
rect 4172 30098 4228 30110
rect 4172 30046 4174 30098
rect 4226 30046 4228 30098
rect 4172 29988 4228 30046
rect 4172 29922 4228 29932
rect 4060 28018 4116 28028
rect 4172 29428 4228 29438
rect 4172 28642 4228 29372
rect 4172 28590 4174 28642
rect 4226 28590 4228 28642
rect 3724 27918 3726 27970
rect 3778 27918 3780 27970
rect 3724 27524 3780 27918
rect 3724 27458 3780 27468
rect 3836 27860 3892 27870
rect 4172 27860 4228 28590
rect 3836 27858 4228 27860
rect 3836 27806 3838 27858
rect 3890 27806 4228 27858
rect 3836 27804 4228 27806
rect 3836 27412 3892 27804
rect 3836 27356 4004 27412
rect 3836 27300 3892 27356
rect 3500 27244 3892 27300
rect 3500 26290 3556 27244
rect 3948 27074 4004 27356
rect 3948 27022 3950 27074
rect 4002 27022 4004 27074
rect 3948 27010 4004 27022
rect 4172 27300 4228 27310
rect 3500 26238 3502 26290
rect 3554 26238 3556 26290
rect 3500 26226 3556 26238
rect 3724 26964 3780 26974
rect 3836 26962 3892 26974
rect 3836 26910 3838 26962
rect 3890 26910 3892 26962
rect 3836 26908 3892 26910
rect 3724 26852 3892 26908
rect 3724 26290 3780 26852
rect 4060 26516 4116 26526
rect 4060 26422 4116 26460
rect 3724 26238 3726 26290
rect 3778 26238 3780 26290
rect 3724 26226 3780 26238
rect 4172 25060 4228 27244
rect 3388 23938 3444 24780
rect 3388 23886 3390 23938
rect 3442 23886 3444 23938
rect 3388 23874 3444 23886
rect 3724 25004 4228 25060
rect 3164 23828 3220 23838
rect 3164 23826 3332 23828
rect 3164 23774 3166 23826
rect 3218 23774 3332 23826
rect 3164 23772 3332 23774
rect 3164 23762 3220 23772
rect 3052 21588 3108 21598
rect 3052 21494 3108 21532
rect 1932 20132 2100 20188
rect 2156 20178 2212 20188
rect 2044 19236 2100 20132
rect 2268 19348 2324 20188
rect 2380 20132 2660 20188
rect 2716 20132 2996 20188
rect 3052 20132 3108 20142
rect 2380 20130 2436 20132
rect 2380 20078 2382 20130
rect 2434 20078 2436 20130
rect 2380 20066 2436 20078
rect 2268 19292 2436 19348
rect 2044 19180 2212 19236
rect 1932 19012 1988 19022
rect 1820 18452 1876 18462
rect 1932 18452 1988 18956
rect 2044 19010 2100 19022
rect 2044 18958 2046 19010
rect 2098 18958 2100 19010
rect 2044 18676 2100 18958
rect 2044 18610 2100 18620
rect 1820 18450 1988 18452
rect 1820 18398 1822 18450
rect 1874 18398 1988 18450
rect 1820 18396 1988 18398
rect 1820 18386 1876 18396
rect 1708 17780 1764 17790
rect 1708 17666 1764 17724
rect 1708 17614 1710 17666
rect 1762 17614 1764 17666
rect 1708 17108 1764 17614
rect 1820 17108 1876 17118
rect 1708 17106 1876 17108
rect 1708 17054 1822 17106
rect 1874 17054 1876 17106
rect 1708 17052 1876 17054
rect 1820 17042 1876 17052
rect 1708 14306 1764 14318
rect 1708 14254 1710 14306
rect 1762 14254 1764 14306
rect 1708 13524 1764 14254
rect 1708 13458 1764 13468
rect 1820 14308 1876 14318
rect 1932 14308 1988 18396
rect 2044 17892 2100 17902
rect 2044 17554 2100 17836
rect 2044 17502 2046 17554
rect 2098 17502 2100 17554
rect 2044 17490 2100 17502
rect 2044 14644 2100 14654
rect 2044 14550 2100 14588
rect 1876 14252 1988 14308
rect 1820 13746 1876 14252
rect 1820 13694 1822 13746
rect 1874 13694 1876 13746
rect 1708 12852 1764 12862
rect 1708 12758 1764 12796
rect 1820 12628 1876 13694
rect 1708 12572 1876 12628
rect 1932 12852 1988 12862
rect 1708 6916 1764 12572
rect 1820 12404 1876 12414
rect 1932 12404 1988 12796
rect 1820 12402 1988 12404
rect 1820 12350 1822 12402
rect 1874 12350 1988 12402
rect 1820 12348 1988 12350
rect 1820 12338 1876 12348
rect 2156 12292 2212 19180
rect 2268 19122 2324 19134
rect 2268 19070 2270 19122
rect 2322 19070 2324 19122
rect 2268 17666 2324 19070
rect 2268 17614 2270 17666
rect 2322 17614 2324 17666
rect 2268 17602 2324 17614
rect 2380 19122 2436 19292
rect 2380 19070 2382 19122
rect 2434 19070 2436 19122
rect 2268 14530 2324 14542
rect 2268 14478 2270 14530
rect 2322 14478 2324 14530
rect 2268 14196 2324 14478
rect 2268 14130 2324 14140
rect 2380 12964 2436 19070
rect 2716 19124 2772 20132
rect 3052 20038 3108 20076
rect 3276 20130 3332 23772
rect 3724 20916 3780 25004
rect 3836 24834 3892 24846
rect 3836 24782 3838 24834
rect 3890 24782 3892 24834
rect 3836 21140 3892 24782
rect 3948 24612 4004 24622
rect 3948 24162 4004 24556
rect 3948 24110 3950 24162
rect 4002 24110 4004 24162
rect 3948 24098 4004 24110
rect 4284 24162 4340 32284
rect 4844 32228 4900 32238
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4620 32004 4676 32014
rect 4396 31892 4452 31902
rect 4396 31778 4452 31836
rect 4396 31726 4398 31778
rect 4450 31726 4452 31778
rect 4396 31714 4452 31726
rect 4620 30994 4676 31948
rect 4732 31892 4788 31902
rect 4844 31892 4900 32172
rect 4732 31890 4900 31892
rect 4732 31838 4734 31890
rect 4786 31838 4900 31890
rect 4732 31836 4900 31838
rect 4732 31826 4788 31836
rect 4620 30942 4622 30994
rect 4674 30942 4676 30994
rect 4620 30930 4676 30942
rect 4844 30996 4900 31006
rect 4844 30902 4900 30940
rect 4732 30882 4788 30894
rect 4732 30830 4734 30882
rect 4786 30830 4788 30882
rect 4732 30772 4788 30830
rect 4732 30716 4900 30772
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4732 29428 4788 29438
rect 4844 29428 4900 30716
rect 4956 30324 5012 34750
rect 5628 34804 5684 34814
rect 5628 34244 5684 34748
rect 5628 34150 5684 34188
rect 5516 34132 5572 34142
rect 5404 34130 5572 34132
rect 5404 34078 5518 34130
rect 5570 34078 5572 34130
rect 5404 34076 5572 34078
rect 5292 31220 5348 31230
rect 5068 31108 5124 31118
rect 5124 31052 5236 31108
rect 5068 31042 5124 31052
rect 5180 30994 5236 31052
rect 5180 30942 5182 30994
rect 5234 30942 5236 30994
rect 5180 30930 5236 30942
rect 4956 30258 5012 30268
rect 4956 30100 5012 30110
rect 5292 30100 5348 31164
rect 4956 30098 5348 30100
rect 4956 30046 4958 30098
rect 5010 30046 5348 30098
rect 4956 30044 5348 30046
rect 4956 30034 5012 30044
rect 5068 29428 5124 29438
rect 4844 29426 5124 29428
rect 4844 29374 5070 29426
rect 5122 29374 5124 29426
rect 4844 29372 5124 29374
rect 4732 29204 4788 29372
rect 5068 29362 5124 29372
rect 5292 29314 5348 29326
rect 5292 29262 5294 29314
rect 5346 29262 5348 29314
rect 4732 29148 4900 29204
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4732 28196 4788 28206
rect 4396 28084 4452 28094
rect 4396 27636 4452 28028
rect 4732 27970 4788 28140
rect 4732 27918 4734 27970
rect 4786 27918 4788 27970
rect 4732 27906 4788 27918
rect 4396 27570 4452 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4844 27186 4900 29148
rect 5180 28084 5236 28094
rect 5292 28084 5348 29262
rect 5180 28082 5348 28084
rect 5180 28030 5182 28082
rect 5234 28030 5348 28082
rect 5180 28028 5348 28030
rect 5180 28018 5236 28028
rect 5068 27858 5124 27870
rect 5292 27860 5348 27898
rect 5068 27806 5070 27858
rect 5122 27806 5124 27858
rect 5068 27412 5124 27806
rect 5068 27346 5124 27356
rect 5180 27804 5292 27860
rect 5180 27188 5236 27804
rect 5292 27794 5348 27804
rect 5292 27636 5348 27646
rect 5292 27542 5348 27580
rect 4844 27134 4846 27186
rect 4898 27134 4900 27186
rect 4844 26628 4900 27134
rect 4844 26562 4900 26572
rect 4956 27132 5236 27188
rect 4956 26516 5012 27132
rect 5404 27076 5460 34076
rect 5516 34066 5572 34076
rect 5740 32004 5796 35644
rect 5852 35634 5908 35644
rect 5964 36708 6020 36718
rect 5852 34356 5908 34366
rect 5964 34356 6020 36652
rect 6076 35922 6132 37214
rect 6188 37156 6244 37166
rect 6188 36596 6244 37100
rect 6188 36482 6244 36540
rect 6188 36430 6190 36482
rect 6242 36430 6244 36482
rect 6188 36418 6244 36430
rect 6076 35870 6078 35922
rect 6130 35870 6132 35922
rect 6076 35858 6132 35870
rect 6188 36260 6244 36270
rect 6188 35810 6244 36204
rect 6300 36258 6356 37998
rect 6524 37940 6580 37950
rect 6300 36206 6302 36258
rect 6354 36206 6356 36258
rect 6300 36194 6356 36206
rect 6412 37938 6580 37940
rect 6412 37886 6526 37938
rect 6578 37886 6580 37938
rect 6412 37884 6580 37886
rect 6188 35758 6190 35810
rect 6242 35758 6244 35810
rect 6188 35746 6244 35758
rect 5852 34354 6020 34356
rect 5852 34302 5854 34354
rect 5906 34302 6020 34354
rect 5852 34300 6020 34302
rect 5852 34290 5908 34300
rect 6300 34244 6356 34254
rect 6076 34020 6132 34030
rect 6076 33926 6132 33964
rect 6188 34018 6244 34030
rect 6188 33966 6190 34018
rect 6242 33966 6244 34018
rect 6076 33348 6132 33358
rect 6188 33348 6244 33966
rect 6300 33684 6356 34188
rect 6300 33618 6356 33628
rect 6076 33346 6244 33348
rect 6076 33294 6078 33346
rect 6130 33294 6244 33346
rect 6076 33292 6244 33294
rect 6300 33460 6356 33470
rect 6300 33346 6356 33404
rect 6300 33294 6302 33346
rect 6354 33294 6356 33346
rect 6076 33282 6132 33292
rect 6300 33236 6356 33294
rect 6188 33180 6356 33236
rect 6188 32562 6244 33180
rect 6188 32510 6190 32562
rect 6242 32510 6244 32562
rect 6188 32498 6244 32510
rect 6300 32562 6356 32574
rect 6300 32510 6302 32562
rect 6354 32510 6356 32562
rect 5740 31938 5796 31948
rect 6300 31556 6356 32510
rect 6300 31490 6356 31500
rect 6188 31332 6244 31342
rect 5516 31220 5572 31230
rect 5516 31126 5572 31164
rect 6188 31218 6244 31276
rect 6188 31166 6190 31218
rect 6242 31166 6244 31218
rect 6188 31154 6244 31166
rect 5740 30996 5796 31006
rect 5740 30902 5796 30940
rect 5628 30882 5684 30894
rect 5628 30830 5630 30882
rect 5682 30830 5684 30882
rect 5628 30548 5684 30830
rect 5628 30492 6132 30548
rect 6076 30324 6132 30492
rect 6412 30434 6468 37884
rect 6524 37874 6580 37884
rect 6524 36484 6580 36494
rect 6524 33572 6580 36428
rect 6636 34916 6692 40348
rect 6748 37266 6804 37278
rect 6748 37214 6750 37266
rect 6802 37214 6804 37266
rect 6748 36708 6804 37214
rect 6860 37044 6916 43932
rect 7420 43540 7476 44380
rect 7532 44324 7588 46622
rect 7756 46004 7812 47740
rect 7868 46116 7924 48190
rect 7980 46900 8036 48860
rect 8316 48132 8372 49756
rect 8428 49746 8484 49756
rect 8988 49138 9044 50428
rect 9660 50418 9716 50428
rect 10556 50706 10836 50708
rect 10556 50654 10782 50706
rect 10834 50654 10836 50706
rect 10556 50652 10836 50654
rect 10556 50596 10612 50652
rect 10780 50642 10836 50652
rect 8988 49086 8990 49138
rect 9042 49086 9044 49138
rect 8988 49074 9044 49086
rect 9772 49810 9828 49822
rect 9772 49758 9774 49810
rect 9826 49758 9828 49810
rect 9772 49700 9828 49758
rect 8540 48916 8596 48926
rect 8540 48822 8596 48860
rect 9100 48916 9156 48926
rect 8876 48804 8932 48814
rect 8876 48710 8932 48748
rect 9100 48802 9156 48860
rect 9100 48750 9102 48802
rect 9154 48750 9156 48802
rect 8316 48066 8372 48076
rect 8876 48468 8932 48478
rect 8876 47234 8932 48412
rect 9100 48244 9156 48750
rect 9324 48802 9380 48814
rect 9324 48750 9326 48802
rect 9378 48750 9380 48802
rect 9324 48468 9380 48750
rect 9324 48402 9380 48412
rect 9660 48356 9716 48366
rect 9660 48262 9716 48300
rect 9100 48188 9492 48244
rect 8988 48130 9044 48142
rect 8988 48078 8990 48130
rect 9042 48078 9044 48130
rect 8988 47460 9044 48078
rect 9044 47404 9268 47460
rect 8988 47394 9044 47404
rect 8876 47182 8878 47234
rect 8930 47182 8932 47234
rect 8540 46900 8596 46910
rect 7980 46898 8596 46900
rect 7980 46846 7982 46898
rect 8034 46846 8542 46898
rect 8594 46846 8596 46898
rect 7980 46844 8596 46846
rect 7980 46834 8036 46844
rect 8540 46834 8596 46844
rect 8764 46788 8820 46798
rect 8876 46788 8932 47182
rect 8764 46786 8932 46788
rect 8764 46734 8766 46786
rect 8818 46734 8932 46786
rect 8764 46732 8932 46734
rect 8316 46676 8372 46686
rect 8316 46582 8372 46620
rect 8428 46562 8484 46574
rect 8428 46510 8430 46562
rect 8482 46510 8484 46562
rect 7868 46060 8148 46116
rect 7756 45948 8036 46004
rect 7532 44258 7588 44268
rect 7532 43540 7588 43550
rect 7420 43538 7588 43540
rect 7420 43486 7534 43538
rect 7586 43486 7588 43538
rect 7420 43484 7588 43486
rect 7420 43314 7476 43326
rect 7420 43262 7422 43314
rect 7474 43262 7476 43314
rect 7196 43092 7252 43102
rect 7196 42866 7252 43036
rect 7196 42814 7198 42866
rect 7250 42814 7252 42866
rect 7196 42802 7252 42814
rect 7420 42756 7476 43262
rect 7420 42690 7476 42700
rect 7084 42532 7140 42542
rect 7084 40964 7140 42476
rect 7532 42308 7588 43484
rect 7868 43538 7924 43550
rect 7868 43486 7870 43538
rect 7922 43486 7924 43538
rect 7756 42980 7812 42990
rect 7756 42866 7812 42924
rect 7756 42814 7758 42866
rect 7810 42814 7812 42866
rect 7532 42252 7700 42308
rect 7532 41860 7588 41870
rect 7308 41748 7364 41758
rect 7364 41692 7476 41748
rect 7308 41682 7364 41692
rect 6972 40908 7140 40964
rect 6972 40180 7028 40908
rect 7084 40740 7140 40750
rect 7084 40404 7140 40684
rect 7084 40402 7252 40404
rect 7084 40350 7086 40402
rect 7138 40350 7252 40402
rect 7084 40348 7252 40350
rect 7084 40338 7140 40348
rect 6972 40124 7140 40180
rect 6860 36978 6916 36988
rect 6972 39618 7028 39630
rect 6972 39566 6974 39618
rect 7026 39566 7028 39618
rect 6748 36642 6804 36652
rect 6748 36484 6804 36494
rect 6748 36390 6804 36428
rect 6972 35924 7028 39566
rect 6972 35858 7028 35868
rect 7084 35308 7140 40124
rect 7196 39618 7252 40348
rect 7196 39566 7198 39618
rect 7250 39566 7252 39618
rect 7196 38052 7252 39566
rect 7196 37378 7252 37996
rect 7196 37326 7198 37378
rect 7250 37326 7252 37378
rect 7196 37314 7252 37326
rect 7308 37604 7364 37614
rect 7308 37156 7364 37548
rect 7196 37100 7364 37156
rect 7196 36372 7252 37100
rect 7420 37044 7476 41692
rect 7532 38834 7588 41804
rect 7644 41188 7700 42252
rect 7644 41122 7700 41132
rect 7756 40516 7812 42814
rect 7868 40628 7924 43486
rect 7868 40562 7924 40572
rect 7756 40450 7812 40460
rect 7980 40514 8036 45948
rect 8092 45218 8148 46060
rect 8428 46004 8484 46510
rect 8428 45938 8484 45948
rect 8092 45166 8094 45218
rect 8146 45166 8148 45218
rect 8092 42420 8148 45166
rect 8652 43876 8708 43886
rect 8764 43876 8820 46732
rect 9100 46004 9156 46014
rect 9100 45910 9156 45948
rect 8708 43820 8820 43876
rect 8652 43762 8708 43820
rect 8652 43710 8654 43762
rect 8706 43710 8708 43762
rect 8652 43698 8708 43710
rect 8092 42354 8148 42364
rect 8204 43650 8260 43662
rect 8204 43598 8206 43650
rect 8258 43598 8260 43650
rect 7980 40462 7982 40514
rect 8034 40462 8036 40514
rect 7980 40450 8036 40462
rect 7532 38782 7534 38834
rect 7586 38782 7588 38834
rect 7532 38770 7588 38782
rect 7644 40402 7700 40414
rect 7644 40350 7646 40402
rect 7698 40350 7700 40402
rect 7644 38668 7700 40350
rect 8092 38724 8148 38734
rect 7644 38612 7812 38668
rect 7532 38276 7588 38286
rect 7532 37940 7588 38220
rect 7644 38052 7700 38062
rect 7644 37958 7700 37996
rect 7532 37378 7588 37884
rect 7532 37326 7534 37378
rect 7586 37326 7588 37378
rect 7532 37156 7588 37326
rect 7532 37090 7588 37100
rect 7196 36278 7252 36316
rect 7308 36988 7476 37044
rect 6636 34850 6692 34860
rect 6748 35252 7140 35308
rect 6636 34692 6692 34702
rect 6748 34692 6804 35252
rect 6972 34804 7028 34814
rect 6972 34710 7028 34748
rect 6636 34690 6804 34692
rect 6636 34638 6638 34690
rect 6690 34638 6804 34690
rect 6636 34636 6804 34638
rect 7084 34690 7140 34702
rect 7084 34638 7086 34690
rect 7138 34638 7140 34690
rect 6636 34244 6692 34636
rect 7084 34356 7140 34638
rect 7196 34692 7252 34702
rect 7196 34598 7252 34636
rect 6636 34178 6692 34188
rect 6860 34300 7140 34356
rect 6860 34130 6916 34300
rect 6860 34078 6862 34130
rect 6914 34078 6916 34130
rect 6860 34066 6916 34078
rect 7084 34130 7140 34142
rect 7084 34078 7086 34130
rect 7138 34078 7140 34130
rect 7084 33572 7140 34078
rect 6524 33516 6692 33572
rect 6636 32674 6692 33516
rect 7084 33506 7140 33516
rect 7196 34020 7252 34030
rect 6972 33460 7028 33470
rect 6636 32622 6638 32674
rect 6690 32622 6692 32674
rect 6524 32564 6580 32574
rect 6524 32470 6580 32508
rect 6636 32116 6692 32622
rect 6636 32050 6692 32060
rect 6748 32788 6804 32798
rect 6748 31948 6804 32732
rect 6412 30382 6414 30434
rect 6466 30382 6468 30434
rect 6412 30370 6468 30382
rect 6524 31892 6804 31948
rect 6972 32228 7028 33404
rect 7084 33346 7140 33358
rect 7084 33294 7086 33346
rect 7138 33294 7140 33346
rect 7084 32788 7140 33294
rect 7196 33234 7252 33964
rect 7196 33182 7198 33234
rect 7250 33182 7252 33234
rect 7196 33170 7252 33182
rect 7084 32722 7140 32732
rect 7308 32786 7364 36988
rect 7756 36932 7812 38612
rect 7868 38612 8148 38668
rect 7868 37268 7924 38612
rect 8204 37268 8260 43598
rect 8540 43538 8596 43550
rect 8540 43486 8542 43538
rect 8594 43486 8596 43538
rect 8540 42868 8596 43486
rect 8764 43540 8820 43820
rect 8876 44210 8932 44222
rect 8876 44158 8878 44210
rect 8930 44158 8932 44210
rect 8876 43762 8932 44158
rect 8876 43710 8878 43762
rect 8930 43710 8932 43762
rect 8876 43698 8932 43710
rect 8764 43484 9044 43540
rect 8540 42802 8596 42812
rect 8428 42644 8484 42654
rect 8428 41298 8484 42588
rect 8988 42196 9044 43484
rect 9212 42980 9268 47404
rect 9436 47348 9492 48188
rect 9660 47348 9716 47358
rect 9436 47346 9716 47348
rect 9436 47294 9662 47346
rect 9714 47294 9716 47346
rect 9436 47292 9716 47294
rect 9324 47234 9380 47246
rect 9324 47182 9326 47234
rect 9378 47182 9380 47234
rect 9324 47012 9380 47182
rect 9324 46946 9380 46956
rect 9660 46674 9716 47292
rect 9772 47234 9828 49644
rect 9996 49698 10052 49710
rect 9996 49646 9998 49698
rect 10050 49646 10052 49698
rect 9996 48916 10052 49646
rect 9996 48850 10052 48860
rect 9884 48802 9940 48814
rect 9884 48750 9886 48802
rect 9938 48750 9940 48802
rect 9884 48468 9940 48750
rect 9884 48402 9940 48412
rect 10332 48802 10388 48814
rect 10332 48750 10334 48802
rect 10386 48750 10388 48802
rect 10332 48580 10388 48750
rect 10556 48580 10612 50540
rect 11228 50428 11284 51998
rect 11452 52052 11508 52062
rect 11340 51938 11396 51950
rect 11340 51886 11342 51938
rect 11394 51886 11396 51938
rect 11340 51828 11396 51886
rect 11340 50596 11396 51772
rect 11452 50708 11508 51996
rect 11564 51940 11620 51950
rect 11564 51846 11620 51884
rect 11452 50614 11508 50652
rect 11340 50530 11396 50540
rect 10668 50372 11284 50428
rect 10668 49922 10724 50372
rect 10668 49870 10670 49922
rect 10722 49870 10724 49922
rect 10668 49858 10724 49870
rect 11116 49700 11172 49710
rect 11116 49606 11172 49644
rect 11676 48692 11732 53228
rect 12236 53172 12292 53452
rect 12348 53442 12404 53452
rect 12572 53508 12628 53518
rect 12572 53414 12628 53452
rect 11900 53116 12292 53172
rect 11900 53058 11956 53116
rect 11900 53006 11902 53058
rect 11954 53006 11956 53058
rect 11900 52994 11956 53006
rect 12012 52162 12068 52174
rect 12012 52110 12014 52162
rect 12066 52110 12068 52162
rect 12012 51828 12068 52110
rect 12012 51762 12068 51772
rect 12796 51380 12852 51390
rect 12460 51378 12852 51380
rect 12460 51326 12798 51378
rect 12850 51326 12852 51378
rect 12460 51324 12852 51326
rect 12460 51266 12516 51324
rect 12796 51314 12852 51324
rect 12460 51214 12462 51266
rect 12514 51214 12516 51266
rect 12460 51202 12516 51214
rect 12684 50708 12740 50718
rect 12684 50614 12740 50652
rect 12796 49700 12852 49710
rect 12796 49606 12852 49644
rect 11004 48636 11732 48692
rect 10332 48524 10724 48580
rect 10332 48356 10388 48524
rect 10332 48290 10388 48300
rect 10444 48132 10500 48142
rect 10500 48076 10612 48132
rect 10444 48038 10500 48076
rect 9996 47460 10052 47470
rect 10332 47460 10388 47470
rect 9996 47458 10388 47460
rect 9996 47406 9998 47458
rect 10050 47406 10334 47458
rect 10386 47406 10388 47458
rect 9996 47404 10388 47406
rect 9996 47394 10052 47404
rect 10332 47394 10388 47404
rect 10556 47458 10612 48076
rect 10556 47406 10558 47458
rect 10610 47406 10612 47458
rect 9772 47182 9774 47234
rect 9826 47182 9828 47234
rect 9772 47012 9828 47182
rect 9772 46788 9828 46956
rect 10108 46788 10164 46798
rect 9772 46732 10108 46788
rect 10108 46694 10164 46732
rect 10444 46788 10500 46798
rect 10556 46788 10612 47406
rect 10444 46786 10612 46788
rect 10444 46734 10446 46786
rect 10498 46734 10612 46786
rect 10444 46732 10612 46734
rect 9660 46622 9662 46674
rect 9714 46622 9716 46674
rect 9660 46610 9716 46622
rect 9436 46564 9492 46574
rect 9212 42914 9268 42924
rect 9324 46562 9492 46564
rect 9324 46510 9438 46562
rect 9490 46510 9492 46562
rect 9324 46508 9492 46510
rect 8988 42102 9044 42140
rect 8428 41246 8430 41298
rect 8482 41246 8484 41298
rect 8428 41234 8484 41246
rect 8540 40964 8596 40974
rect 8316 40514 8372 40526
rect 8316 40462 8318 40514
rect 8370 40462 8372 40514
rect 8316 40404 8372 40462
rect 8316 40338 8372 40348
rect 8428 40402 8484 40414
rect 8428 40350 8430 40402
rect 8482 40350 8484 40402
rect 8428 38052 8484 40350
rect 8428 37986 8484 37996
rect 8540 37604 8596 40908
rect 9324 40516 9380 46508
rect 9436 46498 9492 46508
rect 9884 45890 9940 45902
rect 9884 45838 9886 45890
rect 9938 45838 9940 45890
rect 9884 45668 9940 45838
rect 10332 45668 10388 45678
rect 9884 45666 10388 45668
rect 9884 45614 10334 45666
rect 10386 45614 10388 45666
rect 9884 45612 10388 45614
rect 9660 44322 9716 44334
rect 9660 44270 9662 44322
rect 9714 44270 9716 44322
rect 9660 43764 9716 44270
rect 10108 44324 10164 44334
rect 10332 44324 10388 45612
rect 10108 44322 10388 44324
rect 10108 44270 10110 44322
rect 10162 44270 10388 44322
rect 10108 44268 10388 44270
rect 9884 43764 9940 43774
rect 10108 43764 10164 44268
rect 10444 44212 10500 46732
rect 9660 43762 10108 43764
rect 9660 43710 9886 43762
rect 9938 43710 10108 43762
rect 9660 43708 10108 43710
rect 9884 43698 9940 43708
rect 10108 43698 10164 43708
rect 10220 44156 10500 44212
rect 9884 42644 9940 42654
rect 9436 42642 9940 42644
rect 9436 42590 9886 42642
rect 9938 42590 9940 42642
rect 9436 42588 9940 42590
rect 9436 42194 9492 42588
rect 9884 42578 9940 42588
rect 9436 42142 9438 42194
rect 9490 42142 9492 42194
rect 9436 42130 9492 42142
rect 9660 42196 9716 42206
rect 9660 42102 9716 42140
rect 9772 41970 9828 41982
rect 9772 41918 9774 41970
rect 9826 41918 9828 41970
rect 9548 40516 9604 40526
rect 9772 40516 9828 41918
rect 10108 41972 10164 41982
rect 10108 41878 10164 41916
rect 7868 37266 8148 37268
rect 7868 37214 7870 37266
rect 7922 37214 8148 37266
rect 7868 37212 8148 37214
rect 7868 37202 7924 37212
rect 7644 36876 7812 36932
rect 7532 36372 7588 36382
rect 7420 35924 7476 35934
rect 7420 33458 7476 35868
rect 7532 33796 7588 36316
rect 7644 34242 7700 36876
rect 8092 36594 8148 37212
rect 8204 37202 8260 37212
rect 8428 37548 8596 37604
rect 8764 40460 9492 40516
rect 8092 36542 8094 36594
rect 8146 36542 8148 36594
rect 8092 36530 8148 36542
rect 8204 37044 8260 37054
rect 8092 35588 8148 35598
rect 8204 35588 8260 36988
rect 8428 36484 8484 37548
rect 8540 37380 8596 37390
rect 8540 37266 8596 37324
rect 8540 37214 8542 37266
rect 8594 37214 8596 37266
rect 8540 37202 8596 37214
rect 8652 37266 8708 37278
rect 8652 37214 8654 37266
rect 8706 37214 8708 37266
rect 8652 37044 8708 37214
rect 8652 36978 8708 36988
rect 8540 36484 8596 36494
rect 8428 36482 8596 36484
rect 8428 36430 8542 36482
rect 8594 36430 8596 36482
rect 8428 36428 8596 36430
rect 8092 35586 8260 35588
rect 8092 35534 8094 35586
rect 8146 35534 8260 35586
rect 8092 35532 8260 35534
rect 8540 35586 8596 36428
rect 8540 35534 8542 35586
rect 8594 35534 8596 35586
rect 7644 34190 7646 34242
rect 7698 34190 7700 34242
rect 7644 34178 7700 34190
rect 7756 34692 7812 34702
rect 8092 34692 8148 35532
rect 7812 34636 8148 34692
rect 8204 34916 8260 34926
rect 7532 33730 7588 33740
rect 7420 33406 7422 33458
rect 7474 33406 7476 33458
rect 7420 33394 7476 33406
rect 7532 33572 7588 33582
rect 7308 32734 7310 32786
rect 7362 32734 7364 32786
rect 7308 32722 7364 32734
rect 7532 32786 7588 33516
rect 7532 32734 7534 32786
rect 7586 32734 7588 32786
rect 7532 32722 7588 32734
rect 7084 32564 7140 32574
rect 7084 32470 7140 32508
rect 7196 32564 7252 32574
rect 7196 32562 7364 32564
rect 7196 32510 7198 32562
rect 7250 32510 7364 32562
rect 7196 32508 7364 32510
rect 7196 32498 7252 32508
rect 6188 30324 6244 30334
rect 6076 30322 6244 30324
rect 6076 30270 6190 30322
rect 6242 30270 6244 30322
rect 6076 30268 6244 30270
rect 6188 30258 6244 30268
rect 5964 30212 6020 30222
rect 5964 30118 6020 30156
rect 6300 30210 6356 30222
rect 6300 30158 6302 30210
rect 6354 30158 6356 30210
rect 5628 30100 5684 30110
rect 5628 29650 5684 30044
rect 5628 29598 5630 29650
rect 5682 29598 5684 29650
rect 5628 29586 5684 29598
rect 5740 29764 5796 29774
rect 5740 29650 5796 29708
rect 5740 29598 5742 29650
rect 5794 29598 5796 29650
rect 5740 29586 5796 29598
rect 4956 26450 5012 26460
rect 5068 27020 5460 27076
rect 5516 29426 5572 29438
rect 5516 29374 5518 29426
rect 5570 29374 5572 29426
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4956 24948 5012 24958
rect 5068 24948 5124 27020
rect 5516 26908 5572 29374
rect 6188 28644 6244 28654
rect 6076 28084 6132 28094
rect 5964 27972 6020 27982
rect 4956 24946 5124 24948
rect 4956 24894 4958 24946
rect 5010 24894 5124 24946
rect 4956 24892 5124 24894
rect 5404 26852 5572 26908
rect 5628 27970 6020 27972
rect 5628 27918 5966 27970
rect 6018 27918 6020 27970
rect 5628 27916 6020 27918
rect 4956 24882 5012 24892
rect 4396 24836 4452 24846
rect 4396 24742 4452 24780
rect 4620 24500 4676 24510
rect 4620 24498 4900 24500
rect 4620 24446 4622 24498
rect 4674 24446 4900 24498
rect 4620 24444 4900 24446
rect 4620 24434 4676 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 24110 4286 24162
rect 4338 24110 4340 24162
rect 4284 24098 4340 24110
rect 3836 21074 3892 21084
rect 4284 23380 4340 23390
rect 3836 20916 3892 20926
rect 3276 20078 3278 20130
rect 3330 20078 3332 20130
rect 2828 20020 2884 20030
rect 2828 20018 2996 20020
rect 2828 19966 2830 20018
rect 2882 19966 2996 20018
rect 2828 19964 2996 19966
rect 2828 19954 2884 19964
rect 2940 19236 2996 19964
rect 3276 19572 3332 20078
rect 3388 20914 3892 20916
rect 3388 20862 3838 20914
rect 3890 20862 3892 20914
rect 3388 20860 3892 20862
rect 3388 20020 3444 20860
rect 3836 20850 3892 20860
rect 3388 19926 3444 19964
rect 4284 20578 4340 23324
rect 4844 23268 4900 24444
rect 5404 24164 5460 26852
rect 5628 26404 5684 27916
rect 5964 27906 6020 27916
rect 5740 27636 5796 27646
rect 5796 27580 6020 27636
rect 5740 27570 5796 27580
rect 5964 27298 6020 27580
rect 5964 27246 5966 27298
rect 6018 27246 6020 27298
rect 5964 27234 6020 27246
rect 6076 27300 6132 28028
rect 6076 27206 6132 27244
rect 6188 26908 6244 28588
rect 6300 28082 6356 30158
rect 6412 29764 6468 29774
rect 6412 29426 6468 29708
rect 6412 29374 6414 29426
rect 6466 29374 6468 29426
rect 6412 29362 6468 29374
rect 6300 28030 6302 28082
rect 6354 28030 6356 28082
rect 6300 28018 6356 28030
rect 6412 28868 6468 28878
rect 6412 27972 6468 28812
rect 6300 27860 6356 27870
rect 6412 27860 6468 27916
rect 6300 27858 6468 27860
rect 6300 27806 6302 27858
rect 6354 27806 6468 27858
rect 6300 27804 6468 27806
rect 6300 27794 6356 27804
rect 6412 27298 6468 27804
rect 6412 27246 6414 27298
rect 6466 27246 6468 27298
rect 6412 27234 6468 27246
rect 5292 24108 5460 24164
rect 5516 26348 5684 26404
rect 6076 26852 6244 26908
rect 6300 27074 6356 27086
rect 6300 27022 6302 27074
rect 6354 27022 6356 27074
rect 5068 24052 5124 24062
rect 5068 23828 5124 23996
rect 4956 23826 5124 23828
rect 4956 23774 5070 23826
rect 5122 23774 5124 23826
rect 4956 23772 5124 23774
rect 4956 23380 5012 23772
rect 5068 23762 5124 23772
rect 5292 23716 5348 24108
rect 5516 23940 5572 26348
rect 5628 26178 5684 26190
rect 5628 26126 5630 26178
rect 5682 26126 5684 26178
rect 5628 25060 5684 26126
rect 5628 24994 5684 25004
rect 5628 24834 5684 24846
rect 5628 24782 5630 24834
rect 5682 24782 5684 24834
rect 5628 24052 5684 24782
rect 5964 24836 6020 24846
rect 5964 24742 6020 24780
rect 5628 23986 5684 23996
rect 5292 23650 5348 23660
rect 5404 23884 5572 23940
rect 4956 23314 5012 23324
rect 5068 23492 5124 23502
rect 5404 23492 5460 23884
rect 5852 23826 5908 23838
rect 5852 23774 5854 23826
rect 5906 23774 5908 23826
rect 5516 23716 5572 23726
rect 5740 23716 5796 23726
rect 5516 23714 5684 23716
rect 5516 23662 5518 23714
rect 5570 23662 5684 23714
rect 5516 23660 5684 23662
rect 5516 23650 5572 23660
rect 5068 23378 5124 23436
rect 5068 23326 5070 23378
rect 5122 23326 5124 23378
rect 5068 23314 5124 23326
rect 5180 23436 5460 23492
rect 5628 23492 5684 23660
rect 5740 23622 5796 23660
rect 4844 23202 4900 23212
rect 4620 23044 4676 23054
rect 4956 23044 5012 23054
rect 4620 23042 5012 23044
rect 4620 22990 4622 23042
rect 4674 22990 4958 23042
rect 5010 22990 5012 23042
rect 4620 22988 5012 22990
rect 4620 22978 4676 22988
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4508 22596 4564 22606
rect 4508 22502 4564 22540
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4284 20526 4286 20578
rect 4338 20526 4340 20578
rect 4284 20132 4340 20526
rect 3276 19516 3556 19572
rect 3500 19236 3556 19516
rect 2940 19180 3108 19236
rect 2828 19124 2884 19134
rect 2716 19122 2884 19124
rect 2716 19070 2830 19122
rect 2882 19070 2884 19122
rect 2716 19068 2884 19070
rect 2604 19010 2660 19022
rect 2604 18958 2606 19010
rect 2658 18958 2660 19010
rect 2492 18564 2548 18574
rect 2604 18564 2660 18958
rect 2828 18676 2884 19068
rect 2828 18610 2884 18620
rect 2940 19010 2996 19022
rect 2940 18958 2942 19010
rect 2994 18958 2996 19010
rect 2492 18562 2660 18564
rect 2492 18510 2494 18562
rect 2546 18510 2660 18562
rect 2492 18508 2660 18510
rect 2716 18564 2772 18574
rect 2492 18498 2548 18508
rect 2604 17556 2660 17566
rect 2716 17556 2772 18508
rect 2940 18452 2996 18958
rect 2604 17554 2772 17556
rect 2604 17502 2606 17554
rect 2658 17502 2772 17554
rect 2604 17500 2772 17502
rect 2828 17554 2884 17566
rect 2828 17502 2830 17554
rect 2882 17502 2884 17554
rect 2604 17490 2660 17500
rect 2492 17442 2548 17454
rect 2492 17390 2494 17442
rect 2546 17390 2548 17442
rect 2492 17332 2548 17390
rect 2828 17332 2884 17502
rect 2492 17276 2884 17332
rect 2828 14644 2884 17276
rect 2940 17332 2996 18396
rect 3052 17892 3108 19180
rect 3164 19124 3220 19134
rect 3388 19124 3444 19134
rect 3164 19122 3444 19124
rect 3164 19070 3166 19122
rect 3218 19070 3390 19122
rect 3442 19070 3444 19122
rect 3164 19068 3444 19070
rect 3164 19058 3220 19068
rect 3388 19058 3444 19068
rect 3500 19122 3556 19180
rect 3948 19236 4004 19246
rect 3948 19142 4004 19180
rect 3500 19070 3502 19122
rect 3554 19070 3556 19122
rect 3500 19058 3556 19070
rect 4060 19122 4116 19134
rect 4060 19070 4062 19122
rect 4114 19070 4116 19122
rect 3724 19010 3780 19022
rect 3724 18958 3726 19010
rect 3778 18958 3780 19010
rect 3724 18564 3780 18958
rect 3724 18498 3780 18508
rect 3948 18676 4004 18686
rect 3500 18228 3556 18238
rect 3052 17836 3220 17892
rect 2940 17266 2996 17276
rect 3164 15426 3220 17836
rect 3388 17556 3444 17566
rect 3164 15374 3166 15426
rect 3218 15374 3220 15426
rect 3164 15362 3220 15374
rect 3276 17332 3332 17342
rect 3388 17332 3444 17500
rect 3500 17554 3556 18172
rect 3948 17780 4004 18620
rect 4060 18228 4116 19070
rect 4284 18788 4340 20076
rect 4844 20132 4900 20142
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4844 19346 4900 20076
rect 4844 19294 4846 19346
rect 4898 19294 4900 19346
rect 4844 19012 4900 19294
rect 4844 18946 4900 18956
rect 4284 18732 4900 18788
rect 4620 18338 4676 18350
rect 4620 18286 4622 18338
rect 4674 18286 4676 18338
rect 4060 18162 4116 18172
rect 4508 18228 4564 18238
rect 4620 18228 4676 18286
rect 4564 18172 4676 18228
rect 4508 18162 4564 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4844 17892 4900 18732
rect 4956 18452 5012 22988
rect 5180 18676 5236 23436
rect 5628 23426 5684 23436
rect 5852 23492 5908 23774
rect 5852 23426 5908 23436
rect 5964 23716 6020 23726
rect 6076 23716 6132 26852
rect 6188 26180 6244 26190
rect 6188 24724 6244 26124
rect 6300 25060 6356 27022
rect 6300 24994 6356 25004
rect 6524 24948 6580 31892
rect 6860 31556 6916 31566
rect 6860 31462 6916 31500
rect 6972 29876 7028 32172
rect 7308 30324 7364 32508
rect 7420 32562 7476 32574
rect 7420 32510 7422 32562
rect 7474 32510 7476 32562
rect 7420 30772 7476 32510
rect 7420 30706 7476 30716
rect 7532 30324 7588 30334
rect 7308 30322 7588 30324
rect 7308 30270 7534 30322
rect 7586 30270 7588 30322
rect 7308 30268 7588 30270
rect 7532 30258 7588 30268
rect 7420 30100 7476 30110
rect 6860 29820 7028 29876
rect 7308 30098 7476 30100
rect 7308 30046 7422 30098
rect 7474 30046 7476 30098
rect 7308 30044 7476 30046
rect 6860 29652 6916 29820
rect 6860 29558 6916 29596
rect 6972 29652 7028 29662
rect 7308 29652 7364 30044
rect 7420 30034 7476 30044
rect 7644 30100 7700 30110
rect 7644 30006 7700 30044
rect 6972 29650 7364 29652
rect 6972 29598 6974 29650
rect 7026 29598 7364 29650
rect 6972 29596 7364 29598
rect 7532 29652 7588 29662
rect 7588 29596 7700 29652
rect 6972 29586 7028 29596
rect 7532 29586 7588 29596
rect 7644 29538 7700 29596
rect 7644 29486 7646 29538
rect 7698 29486 7700 29538
rect 7644 29474 7700 29486
rect 7084 29428 7140 29438
rect 7084 29334 7140 29372
rect 6636 28756 6692 28766
rect 6636 27972 6692 28700
rect 6972 28644 7028 28654
rect 6972 28550 7028 28588
rect 7532 28084 7588 28094
rect 7756 28084 7812 34636
rect 7980 34242 8036 34254
rect 7980 34190 7982 34242
rect 8034 34190 8036 34242
rect 7980 34020 8036 34190
rect 7980 33954 8036 33964
rect 8204 33570 8260 34860
rect 8316 34132 8372 34142
rect 8316 34038 8372 34076
rect 8204 33518 8206 33570
rect 8258 33518 8260 33570
rect 8204 33506 8260 33518
rect 8092 33460 8148 33470
rect 8092 33366 8148 33404
rect 8540 33348 8596 35534
rect 8764 35026 8820 40460
rect 9436 40292 9492 40460
rect 9548 40514 9828 40516
rect 9548 40462 9550 40514
rect 9602 40462 9828 40514
rect 9548 40460 9828 40462
rect 9548 40450 9604 40460
rect 9996 40404 10052 40414
rect 9884 40292 9940 40302
rect 9436 40290 9940 40292
rect 9436 40238 9886 40290
rect 9938 40238 9940 40290
rect 9436 40236 9940 40238
rect 9884 40226 9940 40236
rect 9996 40068 10052 40348
rect 9884 40012 10052 40068
rect 10108 40292 10164 40302
rect 9660 38836 9716 38846
rect 9660 38742 9716 38780
rect 9548 38610 9604 38622
rect 9548 38558 9550 38610
rect 9602 38558 9604 38610
rect 9436 38052 9492 38062
rect 9436 37958 9492 37996
rect 9548 37604 9604 38558
rect 9884 37716 9940 40012
rect 9996 39620 10052 39630
rect 9996 39060 10052 39564
rect 9996 37938 10052 39004
rect 9996 37886 9998 37938
rect 10050 37886 10052 37938
rect 9996 37874 10052 37886
rect 10108 39058 10164 40236
rect 10108 39006 10110 39058
rect 10162 39006 10164 39058
rect 9884 37660 10052 37716
rect 9548 37538 9604 37548
rect 9884 37492 9940 37502
rect 9884 37398 9940 37436
rect 8988 37380 9044 37390
rect 9660 37380 9716 37390
rect 8988 37378 9716 37380
rect 8988 37326 8990 37378
rect 9042 37326 9662 37378
rect 9714 37326 9716 37378
rect 8988 37324 9716 37326
rect 8988 37314 9044 37324
rect 8876 37154 8932 37166
rect 8876 37102 8878 37154
rect 8930 37102 8932 37154
rect 8876 36932 8932 37102
rect 8876 36876 9268 36932
rect 8764 34974 8766 35026
rect 8818 34974 8820 35026
rect 8764 34962 8820 34974
rect 8876 36708 8932 36718
rect 8652 34916 8708 34926
rect 8652 34822 8708 34860
rect 8764 34356 8820 34366
rect 8876 34356 8932 36652
rect 9212 36594 9268 36876
rect 9212 36542 9214 36594
rect 9266 36542 9268 36594
rect 9212 36530 9268 36542
rect 9324 34916 9380 37324
rect 9660 37314 9716 37324
rect 9772 37380 9828 37390
rect 9772 37286 9828 37324
rect 9996 36708 10052 37660
rect 9996 36642 10052 36652
rect 9324 34850 9380 34860
rect 10108 34804 10164 39006
rect 10220 38836 10276 44156
rect 10332 43876 10388 43886
rect 10332 43762 10388 43820
rect 10332 43710 10334 43762
rect 10386 43710 10388 43762
rect 10332 43652 10388 43710
rect 10332 43586 10388 43596
rect 10556 43764 10612 43774
rect 10444 43428 10500 43438
rect 10332 42980 10388 42990
rect 10332 39620 10388 42924
rect 10332 39554 10388 39564
rect 10444 42082 10500 43372
rect 10556 42754 10612 43708
rect 10668 42868 10724 48524
rect 10780 44210 10836 44222
rect 10780 44158 10782 44210
rect 10834 44158 10836 44210
rect 10780 43314 10836 44158
rect 10892 43428 10948 43438
rect 10892 43334 10948 43372
rect 10780 43262 10782 43314
rect 10834 43262 10836 43314
rect 10780 43250 10836 43262
rect 10780 42980 10836 42990
rect 11004 42980 11060 48636
rect 11676 48468 11732 48478
rect 11228 47348 11284 47358
rect 11564 47348 11620 47358
rect 11228 47346 11620 47348
rect 11228 47294 11230 47346
rect 11282 47294 11566 47346
rect 11618 47294 11620 47346
rect 11228 47292 11620 47294
rect 11228 47282 11284 47292
rect 11564 47282 11620 47292
rect 11676 47348 11732 48412
rect 12908 48468 12964 53676
rect 14028 53730 14532 53732
rect 14028 53678 14478 53730
rect 14530 53678 14532 53730
rect 14028 53676 14532 53678
rect 13580 53618 13636 53630
rect 13580 53566 13582 53618
rect 13634 53566 13636 53618
rect 13580 53508 13636 53566
rect 13580 53442 13636 53452
rect 14028 52834 14084 53676
rect 14476 53666 14532 53676
rect 15036 53618 15092 54348
rect 15036 53566 15038 53618
rect 15090 53566 15092 53618
rect 15036 53554 15092 53566
rect 14028 52782 14030 52834
rect 14082 52782 14084 52834
rect 14028 52770 14084 52782
rect 14476 52834 14532 52846
rect 14476 52782 14478 52834
rect 14530 52782 14532 52834
rect 14476 52052 14532 52782
rect 14476 51986 14532 51996
rect 14924 52836 14980 52846
rect 14924 51716 14980 52780
rect 14588 51660 14980 51716
rect 14364 51380 14420 51390
rect 14028 51378 14420 51380
rect 14028 51326 14366 51378
rect 14418 51326 14420 51378
rect 14028 51324 14420 51326
rect 13468 51266 13524 51278
rect 13468 51214 13470 51266
rect 13522 51214 13524 51266
rect 12908 48402 12964 48412
rect 13244 50708 13300 50718
rect 13244 48244 13300 50652
rect 13468 49812 13524 51214
rect 13916 50820 13972 50830
rect 14028 50820 14084 51324
rect 14364 51314 14420 51324
rect 13916 50818 14084 50820
rect 13916 50766 13918 50818
rect 13970 50766 14084 50818
rect 13916 50764 14084 50766
rect 13916 50754 13972 50764
rect 14476 50708 14532 50718
rect 14476 50614 14532 50652
rect 14252 50596 14308 50606
rect 14252 50502 14308 50540
rect 13468 49746 13524 49756
rect 14028 48804 14084 48814
rect 13916 48748 14028 48804
rect 13804 48244 13860 48254
rect 13244 48242 13860 48244
rect 13244 48190 13246 48242
rect 13298 48190 13806 48242
rect 13858 48190 13860 48242
rect 13244 48188 13860 48190
rect 13244 48178 13300 48188
rect 12572 48132 12628 48142
rect 11900 48130 12628 48132
rect 11900 48078 12574 48130
rect 12626 48078 12628 48130
rect 11900 48076 12628 48078
rect 11900 47458 11956 48076
rect 12572 48066 12628 48076
rect 11900 47406 11902 47458
rect 11954 47406 11956 47458
rect 11900 47394 11956 47406
rect 13580 48018 13636 48030
rect 13580 47966 13582 48018
rect 13634 47966 13636 48018
rect 13580 47458 13636 47966
rect 13580 47406 13582 47458
rect 13634 47406 13636 47458
rect 13580 47394 13636 47406
rect 11676 47254 11732 47292
rect 12236 47348 12292 47358
rect 12236 47254 12292 47292
rect 10836 42924 11060 42980
rect 11116 46788 11172 46798
rect 11116 46562 11172 46732
rect 11116 46510 11118 46562
rect 11170 46510 11172 46562
rect 10780 42914 10836 42924
rect 10668 42802 10724 42812
rect 10556 42702 10558 42754
rect 10610 42702 10612 42754
rect 10556 42420 10612 42702
rect 11004 42644 11060 42654
rect 10556 42354 10612 42364
rect 10668 42642 11060 42644
rect 10668 42590 11006 42642
rect 11058 42590 11060 42642
rect 10668 42588 11060 42590
rect 10556 42196 10612 42206
rect 10668 42196 10724 42588
rect 11004 42578 11060 42588
rect 11116 42420 11172 46510
rect 13468 45892 13524 45902
rect 12908 45106 12964 45118
rect 12908 45054 12910 45106
rect 12962 45054 12964 45106
rect 12908 44434 12964 45054
rect 12908 44382 12910 44434
rect 12962 44382 12964 44434
rect 12908 44370 12964 44382
rect 11340 43764 11396 43774
rect 11340 43670 11396 43708
rect 11788 43426 11844 43438
rect 11788 43374 11790 43426
rect 11842 43374 11844 43426
rect 11452 43314 11508 43326
rect 11452 43262 11454 43314
rect 11506 43262 11508 43314
rect 11452 42866 11508 43262
rect 11452 42814 11454 42866
rect 11506 42814 11508 42866
rect 11452 42802 11508 42814
rect 11228 42642 11284 42654
rect 11564 42644 11620 42654
rect 11228 42590 11230 42642
rect 11282 42590 11284 42642
rect 11228 42532 11284 42590
rect 11228 42466 11284 42476
rect 11340 42642 11620 42644
rect 11340 42590 11566 42642
rect 11618 42590 11620 42642
rect 11340 42588 11620 42590
rect 10556 42194 10724 42196
rect 10556 42142 10558 42194
rect 10610 42142 10724 42194
rect 10556 42140 10724 42142
rect 10780 42364 11172 42420
rect 10556 42130 10612 42140
rect 10444 42030 10446 42082
rect 10498 42030 10500 42082
rect 10332 38836 10388 38846
rect 10220 38780 10332 38836
rect 10332 38770 10388 38780
rect 10444 38724 10500 42030
rect 10668 41970 10724 41982
rect 10668 41918 10670 41970
rect 10722 41918 10724 41970
rect 10668 40964 10724 41918
rect 10668 40898 10724 40908
rect 10668 39172 10724 39182
rect 10556 39060 10612 39070
rect 10556 38966 10612 39004
rect 10444 38658 10500 38668
rect 10668 38610 10724 39116
rect 10668 38558 10670 38610
rect 10722 38558 10724 38610
rect 10668 38162 10724 38558
rect 10668 38110 10670 38162
rect 10722 38110 10724 38162
rect 10668 38098 10724 38110
rect 10332 38052 10388 38062
rect 10332 37268 10388 37996
rect 10556 37268 10612 37278
rect 10332 37266 10500 37268
rect 10332 37214 10334 37266
rect 10386 37214 10500 37266
rect 10332 37212 10500 37214
rect 10332 37202 10388 37212
rect 10444 37044 10500 37212
rect 10556 37174 10612 37212
rect 10444 36988 10724 37044
rect 10108 34738 10164 34748
rect 10220 35924 10276 35934
rect 8988 34692 9044 34702
rect 8988 34690 9268 34692
rect 8988 34638 8990 34690
rect 9042 34638 9268 34690
rect 8988 34636 9268 34638
rect 8988 34626 9044 34636
rect 8764 34354 8932 34356
rect 8764 34302 8766 34354
rect 8818 34302 8932 34354
rect 8764 34300 8932 34302
rect 8764 33460 8820 34300
rect 8820 33404 9044 33460
rect 8764 33394 8820 33404
rect 8204 33346 8596 33348
rect 8204 33294 8542 33346
rect 8594 33294 8596 33346
rect 8204 33292 8596 33294
rect 8204 32452 8260 33292
rect 8540 33282 8596 33292
rect 8988 32786 9044 33404
rect 8988 32734 8990 32786
rect 9042 32734 9044 32786
rect 8988 32676 9044 32734
rect 8988 32610 9044 32620
rect 8092 32396 8204 32452
rect 7980 30212 8036 30222
rect 7980 30118 8036 30156
rect 8092 28196 8148 32396
rect 8204 32358 8260 32396
rect 9212 30772 9268 34636
rect 10220 34580 10276 35868
rect 10668 35922 10724 36988
rect 10668 35870 10670 35922
rect 10722 35870 10724 35922
rect 10668 35858 10724 35870
rect 10780 35308 10836 42364
rect 11004 42196 11060 42206
rect 11004 41972 11060 42140
rect 10892 41970 11060 41972
rect 10892 41918 11006 41970
rect 11058 41918 11060 41970
rect 10892 41916 11060 41918
rect 10892 39732 10948 41916
rect 11004 41906 11060 41916
rect 11340 41074 11396 42588
rect 11564 42578 11620 42588
rect 11788 42532 11844 43374
rect 13468 43092 13524 45836
rect 13580 44436 13636 44446
rect 13692 44436 13748 48188
rect 13804 48178 13860 48188
rect 13580 44434 13748 44436
rect 13580 44382 13582 44434
rect 13634 44382 13748 44434
rect 13580 44380 13748 44382
rect 13916 48018 13972 48748
rect 14028 48710 14084 48748
rect 14364 48802 14420 48814
rect 14364 48750 14366 48802
rect 14418 48750 14420 48802
rect 13916 47966 13918 48018
rect 13970 47966 13972 48018
rect 13580 43764 13636 44380
rect 13636 43708 13748 43764
rect 13580 43698 13636 43708
rect 13468 43026 13524 43036
rect 11788 42466 11844 42476
rect 12124 42530 12180 42542
rect 12124 42478 12126 42530
rect 12178 42478 12180 42530
rect 12124 41972 12180 42478
rect 12124 41906 12180 41916
rect 12572 42532 12628 42542
rect 11788 41860 11844 41870
rect 11452 41858 11844 41860
rect 11452 41806 11790 41858
rect 11842 41806 11844 41858
rect 11452 41804 11844 41806
rect 11452 41298 11508 41804
rect 11788 41794 11844 41804
rect 11452 41246 11454 41298
rect 11506 41246 11508 41298
rect 11452 41234 11508 41246
rect 11564 41188 11620 41198
rect 11564 41094 11620 41132
rect 11900 41188 11956 41198
rect 12348 41188 12404 41198
rect 11900 41186 12404 41188
rect 11900 41134 11902 41186
rect 11954 41134 12350 41186
rect 12402 41134 12404 41186
rect 11900 41132 12404 41134
rect 11900 41122 11956 41132
rect 12348 41122 12404 41132
rect 12460 41188 12516 41198
rect 12572 41188 12628 42476
rect 12908 42530 12964 42542
rect 12908 42478 12910 42530
rect 12962 42478 12964 42530
rect 12460 41186 12628 41188
rect 12460 41134 12462 41186
rect 12514 41134 12628 41186
rect 12460 41132 12628 41134
rect 12684 41972 12740 41982
rect 12684 41188 12740 41916
rect 12908 41972 12964 42478
rect 12908 41906 12964 41916
rect 13692 41298 13748 43708
rect 13916 43540 13972 47966
rect 14140 48354 14196 48366
rect 14140 48302 14142 48354
rect 14194 48302 14196 48354
rect 14140 47572 14196 48302
rect 14364 48242 14420 48750
rect 14364 48190 14366 48242
rect 14418 48190 14420 48242
rect 14364 48178 14420 48190
rect 14252 47572 14308 47582
rect 14140 47570 14308 47572
rect 14140 47518 14254 47570
rect 14306 47518 14308 47570
rect 14140 47516 14308 47518
rect 14252 47506 14308 47516
rect 13916 43446 13972 43484
rect 14476 46564 14532 46574
rect 14476 45890 14532 46508
rect 14476 45838 14478 45890
rect 14530 45838 14532 45890
rect 13916 42754 13972 42766
rect 13916 42702 13918 42754
rect 13970 42702 13972 42754
rect 13916 41858 13972 42702
rect 14476 42532 14532 45838
rect 14476 42466 14532 42476
rect 13916 41806 13918 41858
rect 13970 41806 13972 41858
rect 13916 41794 13972 41806
rect 14476 41972 14532 41982
rect 13692 41246 13694 41298
rect 13746 41246 13748 41298
rect 13692 41234 13748 41246
rect 12460 41122 12516 41132
rect 11340 41022 11342 41074
rect 11394 41022 11396 41074
rect 11340 40964 11396 41022
rect 12684 41074 12740 41132
rect 12684 41022 12686 41074
rect 12738 41022 12740 41074
rect 12684 41010 12740 41022
rect 13580 41188 13636 41198
rect 11340 40898 11396 40908
rect 12236 40964 12292 40974
rect 12236 40514 12292 40908
rect 12236 40462 12238 40514
rect 12290 40462 12292 40514
rect 11004 40404 11060 40414
rect 11004 40310 11060 40348
rect 10892 39730 11508 39732
rect 10892 39678 10894 39730
rect 10946 39678 11508 39730
rect 10892 39676 11508 39678
rect 10892 39666 10948 39676
rect 11452 39060 11508 39676
rect 11452 39058 11844 39060
rect 11452 39006 11454 39058
rect 11506 39006 11844 39058
rect 11452 39004 11844 39006
rect 11452 38994 11508 39004
rect 11788 38834 11844 39004
rect 11788 38782 11790 38834
rect 11842 38782 11844 38834
rect 11788 38770 11844 38782
rect 12124 38836 12180 38846
rect 11004 38722 11060 38734
rect 11004 38670 11006 38722
rect 11058 38670 11060 38722
rect 11004 37492 11060 38670
rect 11340 38610 11396 38622
rect 11340 38558 11342 38610
rect 11394 38558 11396 38610
rect 11116 38052 11172 38062
rect 11116 37938 11172 37996
rect 11116 37886 11118 37938
rect 11170 37886 11172 37938
rect 11116 37874 11172 37886
rect 11340 37828 11396 38558
rect 11452 38052 11508 38062
rect 11900 38052 11956 38062
rect 11452 38050 11956 38052
rect 11452 37998 11454 38050
rect 11506 37998 11902 38050
rect 11954 37998 11956 38050
rect 11452 37996 11956 37998
rect 11452 37986 11508 37996
rect 11900 37986 11956 37996
rect 12124 38050 12180 38780
rect 12124 37998 12126 38050
rect 12178 37998 12180 38050
rect 12124 37986 12180 37998
rect 12236 37940 12292 40462
rect 13580 40516 13636 41132
rect 14028 41188 14084 41198
rect 14028 41094 14084 41132
rect 13580 39730 13636 40460
rect 13580 39678 13582 39730
rect 13634 39678 13636 39730
rect 12796 39618 12852 39630
rect 12796 39566 12798 39618
rect 12850 39566 12852 39618
rect 12572 38722 12628 38734
rect 12572 38670 12574 38722
rect 12626 38670 12628 38722
rect 12572 38668 12628 38670
rect 12348 38612 12628 38668
rect 12796 38668 12852 39566
rect 12796 38612 13188 38668
rect 12348 38162 12404 38612
rect 12348 38110 12350 38162
rect 12402 38110 12404 38162
rect 12348 38098 12404 38110
rect 12908 38052 12964 38062
rect 12460 37940 12516 37950
rect 12236 37938 12516 37940
rect 12236 37886 12462 37938
rect 12514 37886 12516 37938
rect 12236 37884 12516 37886
rect 11564 37828 11620 37838
rect 11340 37826 11508 37828
rect 11340 37774 11342 37826
rect 11394 37774 11508 37826
rect 11340 37772 11508 37774
rect 11340 37762 11396 37772
rect 11004 35924 11060 37436
rect 11004 35858 11060 35868
rect 11340 36594 11396 36606
rect 11340 36542 11342 36594
rect 11394 36542 11396 36594
rect 11340 35698 11396 36542
rect 11452 35812 11508 37772
rect 11564 37734 11620 37772
rect 12460 37828 12516 37884
rect 12460 37762 12516 37772
rect 12908 37826 12964 37996
rect 12908 37774 12910 37826
rect 12962 37774 12964 37826
rect 12908 37044 12964 37774
rect 12908 36978 12964 36988
rect 13132 37044 13188 38612
rect 13580 38052 13636 39678
rect 14028 40404 14084 40414
rect 13916 39620 13972 39630
rect 13916 39526 13972 39564
rect 13580 37986 13636 37996
rect 13692 38724 13748 38734
rect 13580 37826 13636 37838
rect 13580 37774 13582 37826
rect 13634 37774 13636 37826
rect 13580 37044 13636 37774
rect 13132 36988 13636 37044
rect 11452 35746 11508 35756
rect 12684 35924 12740 35934
rect 11340 35646 11342 35698
rect 11394 35646 11396 35698
rect 11340 35634 11396 35646
rect 12684 35700 12740 35868
rect 12684 35634 12740 35644
rect 12908 35812 12964 35822
rect 10556 35252 11172 35308
rect 10556 34692 10612 35252
rect 10892 35028 10948 35038
rect 10556 34598 10612 34636
rect 10780 34916 10836 34926
rect 10780 34692 10836 34860
rect 10108 34524 10276 34580
rect 9324 33236 9380 33246
rect 9324 33234 9716 33236
rect 9324 33182 9326 33234
rect 9378 33182 9716 33234
rect 9324 33180 9716 33182
rect 9324 33170 9380 33180
rect 9660 32786 9716 33180
rect 10108 32900 10164 34524
rect 9660 32734 9662 32786
rect 9714 32734 9716 32786
rect 9660 32722 9716 32734
rect 9996 32844 10164 32900
rect 10780 34242 10836 34636
rect 10780 34190 10782 34242
rect 10834 34190 10836 34242
rect 9772 32676 9828 32686
rect 9548 32564 9604 32574
rect 9548 32470 9604 32508
rect 9772 32562 9828 32620
rect 9772 32510 9774 32562
rect 9826 32510 9828 32562
rect 9772 32498 9828 32510
rect 9996 32452 10052 32844
rect 10556 32788 10612 32798
rect 10108 32786 10612 32788
rect 10108 32734 10558 32786
rect 10610 32734 10612 32786
rect 10108 32732 10612 32734
rect 10108 32674 10164 32732
rect 10556 32722 10612 32732
rect 10108 32622 10110 32674
rect 10162 32622 10164 32674
rect 10108 32610 10164 32622
rect 10444 32564 10500 32574
rect 10444 32470 10500 32508
rect 10668 32562 10724 32574
rect 10668 32510 10670 32562
rect 10722 32510 10724 32562
rect 9996 32396 10164 32452
rect 9212 30716 9380 30772
rect 8204 30100 8260 30110
rect 8204 29650 8260 30044
rect 8204 29598 8206 29650
rect 8258 29598 8260 29650
rect 8204 29586 8260 29598
rect 8540 29652 8596 29662
rect 8092 28130 8148 28140
rect 8428 29426 8484 29438
rect 8428 29374 8430 29426
rect 8482 29374 8484 29426
rect 7588 28028 7700 28084
rect 7756 28028 7924 28084
rect 7532 28018 7588 28028
rect 6636 27906 6692 27916
rect 6860 27860 6916 27870
rect 6636 27300 6692 27310
rect 6636 26516 6692 27244
rect 6860 27076 6916 27804
rect 7420 27860 7476 27870
rect 7644 27860 7700 28028
rect 7756 27860 7812 27870
rect 7644 27858 7812 27860
rect 7644 27806 7758 27858
rect 7810 27806 7812 27858
rect 7644 27804 7812 27806
rect 7420 27766 7476 27804
rect 7756 27794 7812 27804
rect 7756 27636 7812 27646
rect 6860 27010 6916 27020
rect 7308 27634 7812 27636
rect 7308 27582 7758 27634
rect 7810 27582 7812 27634
rect 7308 27580 7812 27582
rect 6748 26516 6804 26526
rect 6636 26460 6748 26516
rect 6748 26422 6804 26460
rect 7196 26402 7252 26414
rect 7196 26350 7198 26402
rect 7250 26350 7252 26402
rect 7084 26290 7140 26302
rect 7084 26238 7086 26290
rect 7138 26238 7140 26290
rect 6636 24948 6692 24958
rect 6524 24946 6692 24948
rect 6524 24894 6638 24946
rect 6690 24894 6692 24946
rect 6524 24892 6692 24894
rect 6636 24882 6692 24892
rect 7084 24836 7140 26238
rect 7196 26180 7252 26350
rect 7196 26114 7252 26124
rect 7084 24770 7140 24780
rect 7196 25060 7252 25070
rect 6300 24724 6356 24734
rect 6188 24668 6300 24724
rect 6300 24658 6356 24668
rect 7196 24610 7252 25004
rect 7196 24558 7198 24610
rect 7250 24558 7252 24610
rect 6300 24500 6356 24510
rect 6972 24500 7028 24510
rect 6300 24498 6804 24500
rect 6300 24446 6302 24498
rect 6354 24446 6804 24498
rect 6300 24444 6804 24446
rect 6300 24434 6356 24444
rect 6748 24050 6804 24444
rect 6748 23998 6750 24050
rect 6802 23998 6804 24050
rect 6748 23986 6804 23998
rect 6188 23940 6244 23950
rect 6524 23940 6580 23950
rect 6188 23938 6356 23940
rect 6188 23886 6190 23938
rect 6242 23886 6356 23938
rect 6188 23884 6356 23886
rect 6188 23874 6244 23884
rect 6076 23660 6244 23716
rect 5516 23380 5572 23390
rect 5292 23378 5572 23380
rect 5292 23326 5518 23378
rect 5570 23326 5572 23378
rect 5292 23324 5572 23326
rect 5964 23380 6020 23660
rect 6076 23380 6132 23390
rect 5964 23378 6132 23380
rect 5964 23326 6078 23378
rect 6130 23326 6132 23378
rect 5964 23324 6132 23326
rect 5292 19908 5348 23324
rect 5516 23314 5572 23324
rect 6076 23314 6132 23324
rect 5404 23154 5460 23166
rect 5964 23156 6020 23166
rect 5404 23102 5406 23154
rect 5458 23102 5460 23154
rect 5404 23044 5460 23102
rect 5404 22978 5460 22988
rect 5628 23154 6020 23156
rect 5628 23102 5966 23154
rect 6018 23102 6020 23154
rect 5628 23100 6020 23102
rect 5516 22932 5572 22942
rect 5628 22932 5684 23100
rect 5964 23090 6020 23100
rect 5516 22930 5684 22932
rect 5516 22878 5518 22930
rect 5570 22878 5684 22930
rect 5516 22876 5684 22878
rect 5516 22866 5572 22876
rect 5740 22484 5796 22494
rect 5740 20132 5796 22428
rect 5740 20038 5796 20076
rect 5292 19852 6132 19908
rect 5964 19684 6020 19694
rect 4956 18386 5012 18396
rect 5068 18620 5236 18676
rect 5740 19628 5964 19684
rect 4732 17836 4900 17892
rect 4620 17780 4676 17790
rect 3948 17778 4676 17780
rect 3948 17726 4622 17778
rect 4674 17726 4676 17778
rect 3948 17724 4676 17726
rect 3948 17666 4004 17724
rect 4620 17714 4676 17724
rect 3948 17614 3950 17666
rect 4002 17614 4004 17666
rect 3948 17602 4004 17614
rect 3500 17502 3502 17554
rect 3554 17502 3556 17554
rect 3500 17490 3556 17502
rect 3724 17556 3780 17594
rect 3724 17490 3780 17500
rect 3332 17276 3444 17332
rect 4732 17332 4788 17836
rect 4844 17556 4900 17566
rect 4844 17462 4900 17500
rect 4956 17444 5012 17454
rect 4956 17350 5012 17388
rect 4732 17276 4900 17332
rect 3276 15314 3332 17276
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 3276 15262 3278 15314
rect 3330 15262 3332 15314
rect 3276 15250 3332 15262
rect 3388 15260 3668 15316
rect 2828 14550 2884 14588
rect 3164 14530 3220 14542
rect 3164 14478 3166 14530
rect 3218 14478 3220 14530
rect 3164 14196 3220 14478
rect 3164 14130 3220 14140
rect 3276 14306 3332 14318
rect 3276 14254 3278 14306
rect 3330 14254 3332 14306
rect 2492 13634 2548 13646
rect 2492 13582 2494 13634
rect 2546 13582 2548 13634
rect 2492 13076 2548 13582
rect 3276 13636 3332 14254
rect 3388 13748 3444 15260
rect 3612 15202 3668 15260
rect 3612 15150 3614 15202
rect 3666 15150 3668 15202
rect 3612 15138 3668 15150
rect 4844 15148 4900 17276
rect 5068 17108 5124 18620
rect 5404 18564 5460 18574
rect 5404 18470 5460 18508
rect 5180 18452 5236 18462
rect 5180 17666 5236 18396
rect 5628 18450 5684 18462
rect 5628 18398 5630 18450
rect 5682 18398 5684 18450
rect 5404 17780 5460 17790
rect 5180 17614 5182 17666
rect 5234 17614 5236 17666
rect 5180 17602 5236 17614
rect 5292 17724 5404 17780
rect 5068 17042 5124 17052
rect 5292 16994 5348 17724
rect 5404 17714 5460 17724
rect 5404 17332 5460 17342
rect 5404 17106 5460 17276
rect 5404 17054 5406 17106
rect 5458 17054 5460 17106
rect 5404 17042 5460 17054
rect 5292 16942 5294 16994
rect 5346 16942 5348 16994
rect 5292 16930 5348 16942
rect 5628 16100 5684 18398
rect 5740 18450 5796 19628
rect 5964 19618 6020 19628
rect 6076 19458 6132 19852
rect 6076 19406 6078 19458
rect 6130 19406 6132 19458
rect 6076 19394 6132 19406
rect 5964 19122 6020 19134
rect 5964 19070 5966 19122
rect 6018 19070 6020 19122
rect 5740 18398 5742 18450
rect 5794 18398 5796 18450
rect 5740 18386 5796 18398
rect 5852 18676 5908 18686
rect 5852 18450 5908 18620
rect 5852 18398 5854 18450
rect 5906 18398 5908 18450
rect 5852 18004 5908 18398
rect 5964 18116 6020 19070
rect 6076 19012 6132 19022
rect 6076 18918 6132 18956
rect 6188 18228 6244 23660
rect 6300 23378 6356 23884
rect 6524 23846 6580 23884
rect 6636 23828 6692 23838
rect 6636 23734 6692 23772
rect 6860 23716 6916 23726
rect 6972 23716 7028 24444
rect 7196 24388 7252 24558
rect 7196 24322 7252 24332
rect 7308 24164 7364 27580
rect 7756 27570 7812 27580
rect 7420 27188 7476 27198
rect 7420 27094 7476 27132
rect 7756 27188 7812 27198
rect 7868 27188 7924 28028
rect 8092 27972 8148 27982
rect 8092 27878 8148 27916
rect 7812 27132 7924 27188
rect 7756 27122 7812 27132
rect 7644 27076 7700 27086
rect 8428 27076 8484 29374
rect 8540 29426 8596 29596
rect 8540 29374 8542 29426
rect 8594 29374 8596 29426
rect 8540 29362 8596 29374
rect 8652 29426 8708 29438
rect 8652 29374 8654 29426
rect 8706 29374 8708 29426
rect 7644 26982 7700 27020
rect 8204 27020 8428 27076
rect 8204 27018 8260 27020
rect 7532 26964 7588 26974
rect 8204 26966 8206 27018
rect 8258 26966 8260 27018
rect 8428 27010 8484 27020
rect 8204 26954 8260 26966
rect 7420 24724 7476 24734
rect 7420 24630 7476 24668
rect 6916 23660 7028 23716
rect 7084 24108 7364 24164
rect 7420 24276 7476 24286
rect 6860 23622 6916 23660
rect 6524 23604 6580 23614
rect 6300 23326 6302 23378
rect 6354 23326 6356 23378
rect 6300 23314 6356 23326
rect 6412 23492 6468 23502
rect 6412 23378 6468 23436
rect 6412 23326 6414 23378
rect 6466 23326 6468 23378
rect 6412 23314 6468 23326
rect 6300 22932 6356 22942
rect 6300 18788 6356 22876
rect 6524 19460 6580 23548
rect 6748 23492 6804 23502
rect 6636 23266 6692 23278
rect 6636 23214 6638 23266
rect 6690 23214 6692 23266
rect 6636 19684 6692 23214
rect 6748 23266 6804 23436
rect 6748 23214 6750 23266
rect 6802 23214 6804 23266
rect 6748 23044 6804 23214
rect 6748 22978 6804 22988
rect 6636 19618 6692 19628
rect 6524 19404 6692 19460
rect 6636 19236 6692 19404
rect 6636 19180 6804 19236
rect 6524 19124 6580 19134
rect 6300 18722 6356 18732
rect 6412 19122 6580 19124
rect 6412 19070 6526 19122
rect 6578 19070 6580 19122
rect 6412 19068 6580 19070
rect 6412 18674 6468 19068
rect 6524 19058 6580 19068
rect 6636 19010 6692 19022
rect 6636 18958 6638 19010
rect 6690 18958 6692 19010
rect 6636 18900 6692 18958
rect 6412 18622 6414 18674
rect 6466 18622 6468 18674
rect 6412 18610 6468 18622
rect 6524 18844 6692 18900
rect 6524 18676 6580 18844
rect 6748 18788 6804 19180
rect 6860 19012 6916 19022
rect 6860 18918 6916 18956
rect 6524 18610 6580 18620
rect 6636 18732 6804 18788
rect 6300 18452 6356 18462
rect 6300 18358 6356 18396
rect 6524 18452 6580 18462
rect 6524 18358 6580 18396
rect 6636 18228 6692 18732
rect 6972 18452 7028 18462
rect 6972 18358 7028 18396
rect 6188 18172 6468 18228
rect 5964 18060 6132 18116
rect 5852 17938 5908 17948
rect 6076 17892 6132 18060
rect 5964 17836 6132 17892
rect 6188 18004 6244 18014
rect 5740 17780 5796 17790
rect 5740 17686 5796 17724
rect 5740 17108 5796 17118
rect 5796 17052 5908 17108
rect 5740 17042 5796 17052
rect 5852 16994 5908 17052
rect 5852 16942 5854 16994
rect 5906 16942 5908 16994
rect 5852 16930 5908 16942
rect 5740 16882 5796 16894
rect 5740 16830 5742 16882
rect 5794 16830 5796 16882
rect 5740 16210 5796 16830
rect 5964 16436 6020 17836
rect 6076 17668 6132 17678
rect 6076 17574 6132 17612
rect 6076 16996 6132 17006
rect 6076 16902 6132 16940
rect 5740 16158 5742 16210
rect 5794 16158 5796 16210
rect 5740 16146 5796 16158
rect 5852 16380 6020 16436
rect 6076 16772 6132 16782
rect 5516 16098 5684 16100
rect 5516 16046 5630 16098
rect 5682 16046 5684 16098
rect 5516 16044 5684 16046
rect 3500 15090 3556 15102
rect 4844 15092 5012 15148
rect 3500 15038 3502 15090
rect 3554 15038 3556 15090
rect 3500 14532 3556 15038
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 3500 14476 3892 14532
rect 3836 14418 3892 14476
rect 3836 14366 3838 14418
rect 3890 14366 3892 14418
rect 3724 14306 3780 14318
rect 3724 14254 3726 14306
rect 3778 14254 3780 14306
rect 3724 14196 3780 14254
rect 3724 14130 3780 14140
rect 3388 13692 3668 13748
rect 3276 13580 3444 13636
rect 3052 13524 3108 13534
rect 3108 13468 3332 13524
rect 3052 13458 3108 13468
rect 2492 13010 2548 13020
rect 2380 12898 2436 12908
rect 2828 12964 2884 12974
rect 2492 12852 2548 12862
rect 2492 12758 2548 12796
rect 1932 12236 2212 12292
rect 1820 8034 1876 8046
rect 1820 7982 1822 8034
rect 1874 7982 1876 8034
rect 1820 7924 1876 7982
rect 1932 8036 1988 12236
rect 2716 10836 2772 10846
rect 2716 10610 2772 10780
rect 2716 10558 2718 10610
rect 2770 10558 2772 10610
rect 2716 10546 2772 10558
rect 2044 10500 2100 10510
rect 2044 10498 2436 10500
rect 2044 10446 2046 10498
rect 2098 10446 2436 10498
rect 2044 10444 2436 10446
rect 2044 10434 2100 10444
rect 2380 9826 2436 10444
rect 2828 10164 2884 12908
rect 3276 12962 3332 13468
rect 3388 13300 3444 13580
rect 3388 13244 3556 13300
rect 3388 13076 3444 13086
rect 3388 12982 3444 13020
rect 3276 12910 3278 12962
rect 3330 12910 3332 12962
rect 3276 12898 3332 12910
rect 3500 12962 3556 13244
rect 3500 12910 3502 12962
rect 3554 12910 3556 12962
rect 3500 11844 3556 12910
rect 3276 11788 3556 11844
rect 2940 10500 2996 10510
rect 3276 10500 3332 11788
rect 3388 10836 3444 10846
rect 3388 10742 3444 10780
rect 2940 10498 3332 10500
rect 2940 10446 2942 10498
rect 2994 10446 3332 10498
rect 2940 10444 3332 10446
rect 3500 10612 3556 10622
rect 3612 10612 3668 13692
rect 3836 13636 3892 14366
rect 4844 14308 4900 14318
rect 4844 14214 4900 14252
rect 4620 13636 4676 13646
rect 3836 13634 4676 13636
rect 3836 13582 4622 13634
rect 4674 13582 4676 13634
rect 3836 13580 4676 13582
rect 4620 13570 4676 13580
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4956 13188 5012 15092
rect 4732 13132 5012 13188
rect 5068 13972 5124 13982
rect 5516 13972 5572 16044
rect 5628 16034 5684 16044
rect 5852 15876 5908 16380
rect 5068 13970 5572 13972
rect 5068 13918 5070 13970
rect 5122 13918 5518 13970
rect 5570 13918 5572 13970
rect 5068 13916 5572 13918
rect 5068 13186 5124 13916
rect 5516 13906 5572 13916
rect 5628 15820 5908 15876
rect 5964 15988 6020 15998
rect 6076 15988 6132 16716
rect 5964 15986 6132 15988
rect 5964 15934 5966 15986
rect 6018 15934 6132 15986
rect 5964 15932 6132 15934
rect 6188 15986 6244 17948
rect 6300 17556 6356 17566
rect 6300 17462 6356 17500
rect 6188 15934 6190 15986
rect 6242 15934 6244 15986
rect 5628 13970 5684 15820
rect 5964 14084 6020 15932
rect 5628 13918 5630 13970
rect 5682 13918 5684 13970
rect 5628 13906 5684 13918
rect 5740 14028 6020 14084
rect 5740 13970 5796 14028
rect 5740 13918 5742 13970
rect 5794 13918 5796 13970
rect 5068 13134 5070 13186
rect 5122 13134 5124 13186
rect 3724 12964 3780 12974
rect 3724 12850 3780 12908
rect 4284 12964 4340 12974
rect 4284 12870 4340 12908
rect 3724 12798 3726 12850
rect 3778 12798 3780 12850
rect 3724 12786 3780 12798
rect 4732 12516 4788 13132
rect 5068 13122 5124 13134
rect 5180 13802 5236 13814
rect 5180 13750 5182 13802
rect 5234 13750 5236 13802
rect 4956 12964 5012 12974
rect 4956 12870 5012 12908
rect 4844 12738 4900 12750
rect 4844 12686 4846 12738
rect 4898 12686 4900 12738
rect 4844 12628 4900 12686
rect 5180 12740 5236 13750
rect 5740 13524 5796 13918
rect 5964 13860 6020 13870
rect 5964 13746 6020 13804
rect 5964 13694 5966 13746
rect 6018 13694 6020 13746
rect 5964 13682 6020 13694
rect 6076 13858 6132 13870
rect 6076 13806 6078 13858
rect 6130 13806 6132 13858
rect 5180 12674 5236 12684
rect 5404 13468 5796 13524
rect 4844 12572 5124 12628
rect 5068 12516 5124 12572
rect 4732 12460 5012 12516
rect 5068 12460 5348 12516
rect 4508 12404 4564 12414
rect 4508 12402 4900 12404
rect 4508 12350 4510 12402
rect 4562 12350 4900 12402
rect 4508 12348 4900 12350
rect 4508 12338 4564 12348
rect 4284 12292 4340 12302
rect 4284 12198 4340 12236
rect 4732 12180 4788 12190
rect 4732 12086 4788 12124
rect 4620 12068 4676 12078
rect 4620 11974 4676 12012
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 3948 11620 4004 11630
rect 3948 10836 4004 11564
rect 4844 11506 4900 12348
rect 4844 11454 4846 11506
rect 4898 11454 4900 11506
rect 4844 11442 4900 11454
rect 4844 11284 4900 11294
rect 4844 11190 4900 11228
rect 3948 10742 4004 10780
rect 3500 10610 3668 10612
rect 3500 10558 3502 10610
rect 3554 10558 3668 10610
rect 3500 10556 3668 10558
rect 2940 10434 2996 10444
rect 2380 9774 2382 9826
rect 2434 9774 2436 9826
rect 2380 9762 2436 9774
rect 2492 10108 3108 10164
rect 2492 9714 2548 10108
rect 3052 9938 3108 10108
rect 3052 9886 3054 9938
rect 3106 9886 3108 9938
rect 3052 9874 3108 9886
rect 2492 9662 2494 9714
rect 2546 9662 2548 9714
rect 2492 9604 2548 9662
rect 2716 9604 2772 9614
rect 2268 9548 2548 9604
rect 2604 9602 2772 9604
rect 2604 9550 2718 9602
rect 2770 9550 2772 9602
rect 2604 9548 2772 9550
rect 2156 8260 2212 8270
rect 1932 7970 1988 7980
rect 2044 8258 2212 8260
rect 2044 8206 2158 8258
rect 2210 8206 2212 8258
rect 2044 8204 2212 8206
rect 1820 7474 1876 7868
rect 2044 7698 2100 8204
rect 2156 8194 2212 8204
rect 2044 7646 2046 7698
rect 2098 7646 2100 7698
rect 2044 7634 2100 7646
rect 2268 7588 2324 9548
rect 2604 9268 2660 9548
rect 2716 9538 2772 9548
rect 1820 7422 1822 7474
rect 1874 7422 1876 7474
rect 1820 7410 1876 7422
rect 2156 7532 2324 7588
rect 2492 9212 2660 9268
rect 2716 9268 2772 9278
rect 3164 9268 3220 10444
rect 3500 9492 3556 10556
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4956 9940 5012 12460
rect 5180 12292 5236 12302
rect 5180 12178 5236 12236
rect 5180 12126 5182 12178
rect 5234 12126 5236 12178
rect 5180 12114 5236 12126
rect 5068 12068 5124 12078
rect 5068 11974 5124 12012
rect 5068 11508 5124 11518
rect 5068 11414 5124 11452
rect 5292 10612 5348 12460
rect 5404 11956 5460 13468
rect 6076 13412 6132 13806
rect 6188 13636 6244 15934
rect 6188 13570 6244 13580
rect 6300 16882 6356 16894
rect 6300 16830 6302 16882
rect 6354 16830 6356 16882
rect 5404 11890 5460 11900
rect 5516 13356 6132 13412
rect 5516 11508 5572 13356
rect 5964 13188 6020 13198
rect 6300 13188 6356 16830
rect 6412 13300 6468 18172
rect 6524 18172 6692 18228
rect 6524 14084 6580 18172
rect 6636 17554 6692 17566
rect 6636 17502 6638 17554
rect 6690 17502 6692 17554
rect 6636 17444 6692 17502
rect 6748 17556 6804 17566
rect 6804 17500 6916 17556
rect 6748 17490 6804 17500
rect 6636 16884 6692 17388
rect 6636 16790 6692 16828
rect 6860 16882 6916 17500
rect 6860 16830 6862 16882
rect 6914 16830 6916 16882
rect 6636 16660 6692 16670
rect 6636 14308 6692 16604
rect 6860 14420 6916 16830
rect 6860 14354 6916 14364
rect 6636 14242 6692 14252
rect 7084 14084 7140 24108
rect 7420 23938 7476 24220
rect 7420 23886 7422 23938
rect 7474 23886 7476 23938
rect 7420 23874 7476 23886
rect 7308 23716 7364 23726
rect 7308 23622 7364 23660
rect 7532 23492 7588 26908
rect 7756 26852 7812 26862
rect 7644 26628 7700 26638
rect 7644 24946 7700 26572
rect 7756 25620 7812 26796
rect 7980 26852 8036 26862
rect 8316 26852 8372 26862
rect 7980 26850 8148 26852
rect 7980 26798 7982 26850
rect 8034 26798 8148 26850
rect 7980 26796 8148 26798
rect 7980 26786 8036 26796
rect 7868 26066 7924 26078
rect 7868 26014 7870 26066
rect 7922 26014 7924 26066
rect 7868 25732 7924 26014
rect 7868 25666 7924 25676
rect 8092 25620 8148 26796
rect 8316 26758 8372 26796
rect 8540 26850 8596 26862
rect 8540 26798 8542 26850
rect 8594 26798 8596 26850
rect 8316 26628 8372 26638
rect 8204 26572 8316 26628
rect 8204 26514 8260 26572
rect 8316 26562 8372 26572
rect 8204 26462 8206 26514
rect 8258 26462 8260 26514
rect 8204 26450 8260 26462
rect 8092 25564 8260 25620
rect 7756 25554 7812 25564
rect 7980 25508 8036 25546
rect 7980 25442 8036 25452
rect 7868 25396 7924 25406
rect 7868 25302 7924 25340
rect 8092 25284 8148 25294
rect 8092 25190 8148 25228
rect 7644 24894 7646 24946
rect 7698 24894 7700 24946
rect 7644 24836 7700 24894
rect 7644 24500 7700 24780
rect 7644 24434 7700 24444
rect 7756 24722 7812 24734
rect 8204 24724 8260 25564
rect 8540 25506 8596 26798
rect 8540 25454 8542 25506
rect 8594 25454 8596 25506
rect 8540 25442 8596 25454
rect 7756 24670 7758 24722
rect 7810 24670 7812 24722
rect 7756 24164 7812 24670
rect 7980 24668 8260 24724
rect 7756 24098 7812 24108
rect 7868 24388 7924 24398
rect 7868 24052 7924 24332
rect 7196 23436 7588 23492
rect 7644 23938 7700 23950
rect 7644 23886 7646 23938
rect 7698 23886 7700 23938
rect 7644 23492 7700 23886
rect 7868 23938 7924 23996
rect 7868 23886 7870 23938
rect 7922 23886 7924 23938
rect 7868 23874 7924 23886
rect 7196 22484 7252 23436
rect 7644 23426 7700 23436
rect 7756 23716 7812 23726
rect 7308 23268 7364 23278
rect 7308 23174 7364 23212
rect 7420 23156 7476 23166
rect 7420 23062 7476 23100
rect 7532 23156 7588 23166
rect 7756 23156 7812 23660
rect 7532 23154 7812 23156
rect 7532 23102 7534 23154
rect 7586 23102 7812 23154
rect 7532 23100 7812 23102
rect 7868 23492 7924 23502
rect 7532 23090 7588 23100
rect 7196 22418 7252 22428
rect 7868 22370 7924 23436
rect 7980 23154 8036 24668
rect 8428 24610 8484 24622
rect 8428 24558 8430 24610
rect 8482 24558 8484 24610
rect 8428 24388 8484 24558
rect 8428 24322 8484 24332
rect 8316 24164 8372 24174
rect 8204 24052 8260 24062
rect 8092 23826 8148 23838
rect 8092 23774 8094 23826
rect 8146 23774 8148 23826
rect 8092 23604 8148 23774
rect 8092 23538 8148 23548
rect 7980 23102 7982 23154
rect 8034 23102 8036 23154
rect 7980 23090 8036 23102
rect 7868 22318 7870 22370
rect 7922 22318 7924 22370
rect 7868 22306 7924 22318
rect 8204 22370 8260 23996
rect 8316 23492 8372 24108
rect 8540 24164 8596 24174
rect 8540 23938 8596 24108
rect 8540 23886 8542 23938
rect 8594 23886 8596 23938
rect 8540 23874 8596 23886
rect 8428 23716 8484 23726
rect 8428 23622 8484 23660
rect 8652 23492 8708 29374
rect 8988 29426 9044 29438
rect 8988 29374 8990 29426
rect 9042 29374 9044 29426
rect 8988 28868 9044 29374
rect 8988 28802 9044 28812
rect 8876 27970 8932 27982
rect 8876 27918 8878 27970
rect 8930 27918 8932 27970
rect 8764 27858 8820 27870
rect 8764 27806 8766 27858
rect 8818 27806 8820 27858
rect 8764 27076 8820 27806
rect 8876 27188 8932 27918
rect 9212 27972 9268 27982
rect 8876 27122 8932 27132
rect 9100 27858 9156 27870
rect 9100 27806 9102 27858
rect 9154 27806 9156 27858
rect 8764 27010 8820 27020
rect 8876 26516 8932 26526
rect 8876 26422 8932 26460
rect 9100 25844 9156 27806
rect 9100 25778 9156 25788
rect 9212 26850 9268 27916
rect 9212 26798 9214 26850
rect 9266 26798 9268 26850
rect 9212 25730 9268 26798
rect 9212 25678 9214 25730
rect 9266 25678 9268 25730
rect 9212 25666 9268 25678
rect 8988 25620 9044 25630
rect 8988 25526 9044 25564
rect 9324 25508 9380 30716
rect 9884 29988 9940 29998
rect 9884 29650 9940 29932
rect 9884 29598 9886 29650
rect 9938 29598 9940 29650
rect 9884 29586 9940 29598
rect 9772 29428 9828 29438
rect 9772 29334 9828 29372
rect 9884 29202 9940 29214
rect 9884 29150 9886 29202
rect 9938 29150 9940 29202
rect 9884 28532 9940 29150
rect 9884 28466 9940 28476
rect 9660 27972 9716 27982
rect 9660 27858 9716 27916
rect 9660 27806 9662 27858
rect 9714 27806 9716 27858
rect 9660 27794 9716 27806
rect 10108 27858 10164 32396
rect 10668 30994 10724 32510
rect 10780 32564 10836 34190
rect 10892 32788 10948 34972
rect 11116 34914 11172 35252
rect 12796 35028 12852 35038
rect 12460 34972 12796 35028
rect 11116 34862 11118 34914
rect 11170 34862 11172 34914
rect 11116 34850 11172 34862
rect 11452 34916 11508 34926
rect 11900 34916 11956 34926
rect 11452 34914 11956 34916
rect 11452 34862 11454 34914
rect 11506 34862 11902 34914
rect 11954 34862 11956 34914
rect 11452 34860 11956 34862
rect 11452 34850 11508 34860
rect 11900 34850 11956 34860
rect 12460 34914 12516 34972
rect 12796 34934 12852 34972
rect 12460 34862 12462 34914
rect 12514 34862 12516 34914
rect 12460 34850 12516 34862
rect 12908 34804 12964 35756
rect 12572 34748 12964 34804
rect 11116 34690 11172 34702
rect 11116 34638 11118 34690
rect 11170 34638 11172 34690
rect 10892 32786 11060 32788
rect 10892 32734 10894 32786
rect 10946 32734 11060 32786
rect 10892 32732 11060 32734
rect 10892 32722 10948 32732
rect 10780 32498 10836 32508
rect 11004 32004 11060 32732
rect 11116 32676 11172 34638
rect 11788 34692 11844 34702
rect 12012 34692 12068 34702
rect 11788 34598 11844 34636
rect 11900 34636 12012 34692
rect 11452 33458 11508 33470
rect 11452 33406 11454 33458
rect 11506 33406 11508 33458
rect 11452 32788 11508 33406
rect 11116 32610 11172 32620
rect 11228 32732 11508 32788
rect 11116 32004 11172 32014
rect 11004 32002 11172 32004
rect 11004 31950 11118 32002
rect 11170 31950 11172 32002
rect 11004 31948 11172 31950
rect 11116 31938 11172 31948
rect 10668 30942 10670 30994
rect 10722 30942 10724 30994
rect 10668 30884 10724 30942
rect 11228 30884 11284 32732
rect 11452 32562 11508 32574
rect 11452 32510 11454 32562
rect 11506 32510 11508 32562
rect 11452 32452 11508 32510
rect 11508 32396 11732 32452
rect 11452 32386 11508 32396
rect 11340 32002 11396 32014
rect 11340 31950 11342 32002
rect 11394 31950 11396 32002
rect 11340 31890 11396 31950
rect 11340 31838 11342 31890
rect 11394 31838 11396 31890
rect 11340 31826 11396 31838
rect 11676 31890 11732 32396
rect 11676 31838 11678 31890
rect 11730 31838 11732 31890
rect 11676 31826 11732 31838
rect 10668 30828 11284 30884
rect 10556 30772 10612 30782
rect 10556 30678 10612 30716
rect 10220 30100 10276 30110
rect 10220 30006 10276 30044
rect 10668 30100 10724 30110
rect 10668 30006 10724 30044
rect 11116 30100 11172 30110
rect 11116 30006 11172 30044
rect 10556 29988 10612 29998
rect 10556 29538 10612 29932
rect 11004 29986 11060 29998
rect 11004 29934 11006 29986
rect 11058 29934 11060 29986
rect 10668 29652 10724 29662
rect 10668 29558 10724 29596
rect 10556 29486 10558 29538
rect 10610 29486 10612 29538
rect 10556 29474 10612 29486
rect 10332 29428 10388 29438
rect 10332 29334 10388 29372
rect 11004 29426 11060 29934
rect 11228 29538 11284 30828
rect 11452 30882 11508 30894
rect 11452 30830 11454 30882
rect 11506 30830 11508 30882
rect 11452 30660 11508 30830
rect 11452 29988 11508 30604
rect 11452 29922 11508 29932
rect 11788 30210 11844 30222
rect 11788 30158 11790 30210
rect 11842 30158 11844 30210
rect 11788 30100 11844 30158
rect 11228 29486 11230 29538
rect 11282 29486 11284 29538
rect 11228 29474 11284 29486
rect 11004 29374 11006 29426
rect 11058 29374 11060 29426
rect 11004 29362 11060 29374
rect 11788 29426 11844 30044
rect 11900 29652 11956 34636
rect 12012 34598 12068 34636
rect 12012 33236 12068 33246
rect 12012 30882 12068 33180
rect 12236 32676 12292 32686
rect 12236 32582 12292 32620
rect 12012 30830 12014 30882
rect 12066 30830 12068 30882
rect 12012 29764 12068 30830
rect 12124 30100 12180 30110
rect 12124 30006 12180 30044
rect 12236 29988 12292 29998
rect 12236 29894 12292 29932
rect 12348 29986 12404 29998
rect 12348 29934 12350 29986
rect 12402 29934 12404 29986
rect 12348 29876 12404 29934
rect 12348 29810 12404 29820
rect 12012 29708 12292 29764
rect 11900 29596 12180 29652
rect 11788 29374 11790 29426
rect 11842 29374 11844 29426
rect 10780 29204 10836 29214
rect 10668 29202 10836 29204
rect 10668 29150 10782 29202
rect 10834 29150 10836 29202
rect 10668 29148 10836 29150
rect 10668 28868 10724 29148
rect 10780 29138 10836 29148
rect 10108 27806 10110 27858
rect 10162 27806 10164 27858
rect 9660 27634 9716 27646
rect 9660 27582 9662 27634
rect 9714 27582 9716 27634
rect 9660 27300 9716 27582
rect 9660 27244 9940 27300
rect 9660 26852 9716 26862
rect 9660 26758 9716 26796
rect 9212 25452 9380 25508
rect 9436 25730 9492 25742
rect 9436 25678 9438 25730
rect 9490 25678 9492 25730
rect 8764 25396 8820 25406
rect 8764 24500 8820 25340
rect 9212 24948 9268 25452
rect 9212 24882 9268 24892
rect 9324 25284 9380 25294
rect 9436 25284 9492 25678
rect 9772 25284 9828 25294
rect 9324 25282 9828 25284
rect 9324 25230 9326 25282
rect 9378 25230 9774 25282
rect 9826 25230 9828 25282
rect 9324 25228 9828 25230
rect 8876 24836 8932 24846
rect 8876 24742 8932 24780
rect 8988 24722 9044 24734
rect 8988 24670 8990 24722
rect 9042 24670 9044 24722
rect 8876 24500 8932 24510
rect 8764 24498 8932 24500
rect 8764 24446 8878 24498
rect 8930 24446 8932 24498
rect 8764 24444 8932 24446
rect 8876 24434 8932 24444
rect 8988 24164 9044 24670
rect 8876 24108 9044 24164
rect 9100 24388 9156 24398
rect 9324 24388 9380 25228
rect 9772 25218 9828 25228
rect 9548 24724 9604 24734
rect 9548 24630 9604 24668
rect 9772 24722 9828 24734
rect 9772 24670 9774 24722
rect 9826 24670 9828 24722
rect 9660 24612 9716 24622
rect 9660 24518 9716 24556
rect 9156 24332 9380 24388
rect 8876 24052 8932 24108
rect 8876 23986 8932 23996
rect 8764 23938 8820 23950
rect 8764 23886 8766 23938
rect 8818 23886 8820 23938
rect 8764 23828 8820 23886
rect 8988 23940 9044 23950
rect 9100 23940 9156 24332
rect 8988 23938 9156 23940
rect 8988 23886 8990 23938
rect 9042 23886 9156 23938
rect 8988 23884 9156 23886
rect 8988 23874 9044 23884
rect 8764 23772 8932 23828
rect 8876 23716 8932 23772
rect 9212 23826 9268 23838
rect 9212 23774 9214 23826
rect 9266 23774 9268 23826
rect 8876 23660 9156 23716
rect 9100 23492 9156 23660
rect 8316 23436 8596 23492
rect 8652 23436 9044 23492
rect 8540 23378 8596 23436
rect 8540 23326 8542 23378
rect 8594 23326 8596 23378
rect 8540 23314 8596 23326
rect 8764 23268 8820 23278
rect 8652 23266 8820 23268
rect 8652 23214 8766 23266
rect 8818 23214 8820 23266
rect 8652 23212 8820 23214
rect 8316 23156 8372 23166
rect 8316 23042 8372 23100
rect 8316 22990 8318 23042
rect 8370 22990 8372 23042
rect 8316 22596 8372 22990
rect 8316 22530 8372 22540
rect 8204 22318 8206 22370
rect 8258 22318 8260 22370
rect 8204 22306 8260 22318
rect 7980 22146 8036 22158
rect 7980 22094 7982 22146
rect 8034 22094 8036 22146
rect 7980 21812 8036 22094
rect 8652 21924 8708 23212
rect 8764 23202 8820 23212
rect 8876 23156 8932 23166
rect 8876 23062 8932 23100
rect 7980 21746 8036 21756
rect 8204 21868 8708 21924
rect 7980 21588 8036 21598
rect 7980 19458 8036 21532
rect 8204 21026 8260 21868
rect 8204 20974 8206 21026
rect 8258 20974 8260 21026
rect 8204 20962 8260 20974
rect 8764 21028 8820 21038
rect 8988 21028 9044 23436
rect 9100 23156 9156 23436
rect 9212 23268 9268 23774
rect 9772 23828 9828 24670
rect 9884 24276 9940 27244
rect 10108 27188 10164 27806
rect 10220 27860 10276 27870
rect 10220 27298 10276 27804
rect 10220 27246 10222 27298
rect 10274 27246 10276 27298
rect 10220 27234 10276 27246
rect 10332 27412 10388 27422
rect 10332 27298 10388 27356
rect 10332 27246 10334 27298
rect 10386 27246 10388 27298
rect 10332 27234 10388 27246
rect 10556 27300 10612 27310
rect 10556 27206 10612 27244
rect 10668 27298 10724 28812
rect 11004 29092 11060 29102
rect 10668 27246 10670 27298
rect 10722 27246 10724 27298
rect 10108 27122 10164 27132
rect 10668 26908 10724 27246
rect 10444 26852 10724 26908
rect 10780 28756 10836 28766
rect 10780 28082 10836 28700
rect 10780 28030 10782 28082
rect 10834 28030 10836 28082
rect 10780 26908 10836 28030
rect 11004 28530 11060 29036
rect 11788 28756 11844 29374
rect 11788 28690 11844 28700
rect 11900 29314 11956 29326
rect 11900 29262 11902 29314
rect 11954 29262 11956 29314
rect 11004 28478 11006 28530
rect 11058 28478 11060 28530
rect 10780 26852 10948 26908
rect 10220 25844 10276 25854
rect 10108 25284 10164 25294
rect 10108 25190 10164 25228
rect 10108 24724 10164 24734
rect 10220 24724 10276 25788
rect 10444 25730 10500 26852
rect 10444 25678 10446 25730
rect 10498 25678 10500 25730
rect 10332 25508 10388 25518
rect 10332 25414 10388 25452
rect 10444 25284 10500 25678
rect 10892 26178 10948 26852
rect 10892 26126 10894 26178
rect 10946 26126 10948 26178
rect 10892 25620 10948 26126
rect 10108 24722 10276 24724
rect 10108 24670 10110 24722
rect 10162 24670 10276 24722
rect 10108 24668 10276 24670
rect 10332 25228 10500 25284
rect 10668 25564 10948 25620
rect 10668 25394 10724 25564
rect 10668 25342 10670 25394
rect 10722 25342 10724 25394
rect 10108 24658 10164 24668
rect 9884 23938 9940 24220
rect 9884 23886 9886 23938
rect 9938 23886 9940 23938
rect 9884 23874 9940 23886
rect 10108 23940 10164 23950
rect 9772 23762 9828 23772
rect 10108 23378 10164 23884
rect 10332 23492 10388 25228
rect 10668 25172 10724 25342
rect 10556 24834 10612 24846
rect 10556 24782 10558 24834
rect 10610 24782 10612 24834
rect 10332 23436 10500 23492
rect 10108 23326 10110 23378
rect 10162 23326 10164 23378
rect 10108 23314 10164 23326
rect 9212 23202 9268 23212
rect 9100 23090 9156 23100
rect 10332 23154 10388 23166
rect 10332 23102 10334 23154
rect 10386 23102 10388 23154
rect 9772 23042 9828 23054
rect 9772 22990 9774 23042
rect 9826 22990 9828 23042
rect 9772 22596 9828 22990
rect 9772 22484 9828 22540
rect 10220 22484 10276 22494
rect 9772 22482 10276 22484
rect 9772 22430 9774 22482
rect 9826 22430 10222 22482
rect 10274 22430 10276 22482
rect 9772 22428 10276 22430
rect 9772 22418 9828 22428
rect 10220 22418 10276 22428
rect 9548 21812 9604 21822
rect 9548 21718 9604 21756
rect 10332 21700 10388 23102
rect 10444 23156 10500 23436
rect 10444 23062 10500 23100
rect 10332 21634 10388 21644
rect 9772 21588 9828 21598
rect 9772 21494 9828 21532
rect 8764 21026 9044 21028
rect 8764 20974 8766 21026
rect 8818 20974 9044 21026
rect 8764 20972 9044 20974
rect 8764 20962 8820 20972
rect 9324 20916 9380 20926
rect 8988 20860 9324 20916
rect 7980 19406 7982 19458
rect 8034 19406 8036 19458
rect 7980 19394 8036 19406
rect 8092 20690 8148 20702
rect 8092 20638 8094 20690
rect 8146 20638 8148 20690
rect 7420 19234 7476 19246
rect 7420 19182 7422 19234
rect 7474 19182 7476 19234
rect 7420 18674 7476 19182
rect 7420 18622 7422 18674
rect 7474 18622 7476 18674
rect 7420 18610 7476 18622
rect 7644 19234 7700 19246
rect 7644 19182 7646 19234
rect 7698 19182 7700 19234
rect 7196 18564 7252 18574
rect 7196 18450 7252 18508
rect 7196 18398 7198 18450
rect 7250 18398 7252 18450
rect 7196 18004 7252 18398
rect 7196 17938 7252 17948
rect 7308 18452 7364 18462
rect 7532 18452 7588 18462
rect 7364 18450 7588 18452
rect 7364 18398 7534 18450
rect 7586 18398 7588 18450
rect 7364 18396 7588 18398
rect 7308 17780 7364 18396
rect 7532 18386 7588 18396
rect 7420 17892 7476 17902
rect 7644 17892 7700 19182
rect 8092 18676 8148 20638
rect 8876 20690 8932 20702
rect 8876 20638 8878 20690
rect 8930 20638 8932 20690
rect 8204 20580 8260 20590
rect 8204 20578 8372 20580
rect 8204 20526 8206 20578
rect 8258 20526 8372 20578
rect 8204 20524 8372 20526
rect 8204 20514 8260 20524
rect 8316 19236 8372 20524
rect 8876 19346 8932 20638
rect 8988 20018 9044 20860
rect 9324 20822 9380 20860
rect 8988 19966 8990 20018
rect 9042 19966 9044 20018
rect 8988 19954 9044 19966
rect 9660 20580 9716 20590
rect 9660 19906 9716 20524
rect 9660 19854 9662 19906
rect 9714 19854 9716 19906
rect 9660 19842 9716 19854
rect 8876 19294 8878 19346
rect 8930 19294 8932 19346
rect 8876 19282 8932 19294
rect 8428 19236 8484 19246
rect 8316 19234 8484 19236
rect 8316 19182 8430 19234
rect 8482 19182 8484 19234
rect 8316 19180 8484 19182
rect 8092 18610 8148 18620
rect 8204 18788 8260 18798
rect 7756 18562 7812 18574
rect 7980 18564 8036 18574
rect 7756 18510 7758 18562
rect 7810 18510 7812 18562
rect 7756 18340 7812 18510
rect 7756 18274 7812 18284
rect 7868 18508 7980 18564
rect 7420 17890 7700 17892
rect 7420 17838 7422 17890
rect 7474 17838 7700 17890
rect 7420 17836 7700 17838
rect 7420 17826 7476 17836
rect 7196 17724 7364 17780
rect 7868 17780 7924 18508
rect 7980 18498 8036 18508
rect 8092 18452 8148 18462
rect 8092 18226 8148 18396
rect 8204 18450 8260 18732
rect 8204 18398 8206 18450
rect 8258 18398 8260 18450
rect 8204 18386 8260 18398
rect 8092 18174 8094 18226
rect 8146 18174 8148 18226
rect 7196 17108 7252 17724
rect 7532 17668 7588 17678
rect 7532 17574 7588 17612
rect 7868 17666 7924 17724
rect 7868 17614 7870 17666
rect 7922 17614 7924 17666
rect 7868 17602 7924 17614
rect 7980 18004 8036 18014
rect 7308 17554 7364 17566
rect 7308 17502 7310 17554
rect 7362 17502 7364 17554
rect 7308 17444 7364 17502
rect 7308 17378 7364 17388
rect 7756 17444 7812 17454
rect 7980 17444 8036 17948
rect 8092 17556 8148 18174
rect 8316 18340 8372 18350
rect 8316 17892 8372 18284
rect 8428 18228 8484 19180
rect 8764 19010 8820 19022
rect 8764 18958 8766 19010
rect 8818 18958 8820 19010
rect 8652 18788 8708 18798
rect 8764 18788 8820 18958
rect 8708 18732 8820 18788
rect 8988 19010 9044 19022
rect 8988 18958 8990 19010
rect 9042 18958 9044 19010
rect 8652 18674 8708 18732
rect 8652 18622 8654 18674
rect 8706 18622 8708 18674
rect 8652 18610 8708 18622
rect 8540 18562 8596 18574
rect 8540 18510 8542 18562
rect 8594 18510 8596 18562
rect 8540 18452 8596 18510
rect 8540 18386 8596 18396
rect 8652 18228 8708 18238
rect 8428 18226 8708 18228
rect 8428 18174 8654 18226
rect 8706 18174 8708 18226
rect 8428 18172 8708 18174
rect 8652 18162 8708 18172
rect 8876 17892 8932 17902
rect 8988 17892 9044 18958
rect 9436 18676 9492 18686
rect 9436 18450 9492 18620
rect 9660 18564 9716 18574
rect 9660 18470 9716 18508
rect 9436 18398 9438 18450
rect 9490 18398 9492 18450
rect 9436 18386 9492 18398
rect 9772 18450 9828 18462
rect 9772 18398 9774 18450
rect 9826 18398 9828 18450
rect 9436 18004 9492 18014
rect 8316 17836 8484 17892
rect 8316 17668 8372 17678
rect 8092 17490 8148 17500
rect 8204 17666 8372 17668
rect 8204 17614 8318 17666
rect 8370 17614 8372 17666
rect 8204 17612 8372 17614
rect 7756 17442 8036 17444
rect 7756 17390 7758 17442
rect 7810 17390 8036 17442
rect 7756 17388 8036 17390
rect 7756 17378 7812 17388
rect 7756 17220 7812 17230
rect 7756 17108 7812 17164
rect 7196 17106 7812 17108
rect 7196 17054 7198 17106
rect 7250 17054 7758 17106
rect 7810 17054 7812 17106
rect 7196 17052 7812 17054
rect 7196 17042 7252 17052
rect 7756 17042 7812 17052
rect 7980 17106 8036 17388
rect 8204 17220 8260 17612
rect 8316 17602 8372 17612
rect 8204 17154 8260 17164
rect 8428 17556 8484 17836
rect 8876 17890 9044 17892
rect 8876 17838 8878 17890
rect 8930 17838 9044 17890
rect 8876 17836 9044 17838
rect 9324 17890 9380 17902
rect 9324 17838 9326 17890
rect 9378 17838 9380 17890
rect 8876 17826 8932 17836
rect 7980 17054 7982 17106
rect 8034 17054 8036 17106
rect 7980 17042 8036 17054
rect 8092 17108 8148 17118
rect 7532 16884 7588 16894
rect 7532 16790 7588 16828
rect 8092 16770 8148 17052
rect 8428 16884 8484 17500
rect 8540 17668 8596 17678
rect 8540 16996 8596 17612
rect 9324 17668 9380 17838
rect 9324 17602 9380 17612
rect 9212 17556 9268 17566
rect 9212 17462 9268 17500
rect 9324 17444 9380 17454
rect 9436 17444 9492 17948
rect 9324 17442 9492 17444
rect 9324 17390 9326 17442
rect 9378 17390 9492 17442
rect 9324 17388 9492 17390
rect 9324 17378 9380 17388
rect 9772 17108 9828 18398
rect 9772 17042 9828 17052
rect 8540 16930 8596 16940
rect 8428 16818 8484 16828
rect 8092 16718 8094 16770
rect 8146 16718 8148 16770
rect 8092 16706 8148 16718
rect 10556 16772 10612 24782
rect 10668 24276 10724 25116
rect 10780 25396 10836 25406
rect 10780 24722 10836 25340
rect 10780 24670 10782 24722
rect 10834 24670 10836 24722
rect 10780 24658 10836 24670
rect 10892 25394 10948 25406
rect 10892 25342 10894 25394
rect 10946 25342 10948 25394
rect 10892 24500 10948 25342
rect 10892 24434 10948 24444
rect 10668 24220 10948 24276
rect 10668 23154 10724 24220
rect 10668 23102 10670 23154
rect 10722 23102 10724 23154
rect 10668 22596 10724 23102
rect 10668 22530 10724 22540
rect 10780 24050 10836 24062
rect 10780 23998 10782 24050
rect 10834 23998 10836 24050
rect 10780 18564 10836 23998
rect 10892 23938 10948 24220
rect 10892 23886 10894 23938
rect 10946 23886 10948 23938
rect 10892 23874 10948 23886
rect 10892 23154 10948 23166
rect 10892 23102 10894 23154
rect 10946 23102 10948 23154
rect 10892 22596 10948 23102
rect 10892 22530 10948 22540
rect 10892 22370 10948 22382
rect 10892 22318 10894 22370
rect 10946 22318 10948 22370
rect 10892 21700 10948 22318
rect 10892 21634 10948 21644
rect 11004 20916 11060 28478
rect 11116 28532 11172 28542
rect 11116 27858 11172 28476
rect 11116 27806 11118 27858
rect 11170 27806 11172 27858
rect 11116 27794 11172 27806
rect 11900 27972 11956 29262
rect 11788 27412 11844 27422
rect 11340 27188 11396 27198
rect 11340 27094 11396 27132
rect 11676 26964 11732 26974
rect 11676 25620 11732 26908
rect 11788 26850 11844 27356
rect 11900 27300 11956 27916
rect 11900 27234 11956 27244
rect 12012 27746 12068 27758
rect 12012 27694 12014 27746
rect 12066 27694 12068 27746
rect 11788 26798 11790 26850
rect 11842 26798 11844 26850
rect 11788 26786 11844 26798
rect 11340 25506 11396 25518
rect 11340 25454 11342 25506
rect 11394 25454 11396 25506
rect 11228 25396 11284 25406
rect 11228 25302 11284 25340
rect 11340 25172 11396 25454
rect 11676 25506 11732 25564
rect 11676 25454 11678 25506
rect 11730 25454 11732 25506
rect 11676 25442 11732 25454
rect 11340 25106 11396 25116
rect 11900 25172 11956 25182
rect 11900 24722 11956 25116
rect 11900 24670 11902 24722
rect 11954 24670 11956 24722
rect 11900 24658 11956 24670
rect 11228 24164 11284 24174
rect 11228 23154 11284 24108
rect 11676 23826 11732 23838
rect 11676 23774 11678 23826
rect 11730 23774 11732 23826
rect 11676 23604 11732 23774
rect 11676 23538 11732 23548
rect 11228 23102 11230 23154
rect 11282 23102 11284 23154
rect 11228 23090 11284 23102
rect 11676 22596 11732 22606
rect 11228 22484 11284 22494
rect 11004 20850 11060 20860
rect 11116 22146 11172 22158
rect 11116 22094 11118 22146
rect 11170 22094 11172 22146
rect 10780 18508 10948 18564
rect 10780 18338 10836 18350
rect 10780 18286 10782 18338
rect 10834 18286 10836 18338
rect 10780 17892 10836 18286
rect 10780 17826 10836 17836
rect 10556 16706 10612 16716
rect 10668 16100 10724 16110
rect 10668 15426 10724 16044
rect 10668 15374 10670 15426
rect 10722 15374 10724 15426
rect 9772 15314 9828 15326
rect 9772 15262 9774 15314
rect 9826 15262 9828 15314
rect 9772 15204 9828 15262
rect 10556 15316 10612 15354
rect 10556 15250 10612 15260
rect 9772 15138 9828 15148
rect 9996 15202 10052 15214
rect 9996 15150 9998 15202
rect 10050 15150 10052 15202
rect 9996 14644 10052 15150
rect 10668 15148 10724 15374
rect 10556 15092 10724 15148
rect 10444 14980 10500 14990
rect 9996 14642 10276 14644
rect 9996 14590 9998 14642
rect 10050 14590 10276 14642
rect 9996 14588 10276 14590
rect 9996 14578 10052 14588
rect 9884 14532 9940 14542
rect 9884 14438 9940 14476
rect 7420 14420 7476 14430
rect 6524 14028 6692 14084
rect 7084 14028 7252 14084
rect 6412 13234 6468 13244
rect 6524 13860 6580 13870
rect 5740 13186 6020 13188
rect 5740 13134 5966 13186
rect 6018 13134 6020 13186
rect 5740 13132 6020 13134
rect 5740 12180 5796 13132
rect 5964 13122 6020 13132
rect 6188 13132 6356 13188
rect 5628 11954 5684 11966
rect 5628 11902 5630 11954
rect 5682 11902 5684 11954
rect 5628 11620 5684 11902
rect 5628 11554 5684 11564
rect 5516 11396 5572 11452
rect 5740 11506 5796 12124
rect 5852 12964 5908 12974
rect 5852 12178 5908 12908
rect 6076 12964 6132 12974
rect 6076 12870 6132 12908
rect 5964 12740 6020 12750
rect 6188 12740 6244 13132
rect 6524 13076 6580 13804
rect 6300 13020 6580 13076
rect 6300 12962 6356 13020
rect 6300 12910 6302 12962
rect 6354 12910 6356 12962
rect 6300 12898 6356 12910
rect 6636 12740 6692 14028
rect 7196 13860 7252 14028
rect 6860 13802 6916 13814
rect 6860 13750 6862 13802
rect 6914 13750 6916 13802
rect 5964 12738 6244 12740
rect 5964 12686 5966 12738
rect 6018 12686 6244 12738
rect 5964 12684 6244 12686
rect 6524 12684 6692 12740
rect 6748 13636 6804 13646
rect 6860 13636 6916 13750
rect 6804 13580 6916 13636
rect 7084 13804 7252 13860
rect 5964 12674 6020 12684
rect 6188 12516 6244 12526
rect 6412 12516 6468 12526
rect 5852 12126 5854 12178
rect 5906 12126 5908 12178
rect 5852 12114 5908 12126
rect 5964 12402 6020 12414
rect 5964 12350 5966 12402
rect 6018 12350 6020 12402
rect 5964 12180 6020 12350
rect 6076 12180 6132 12190
rect 5964 12124 6076 12180
rect 6076 12114 6132 12124
rect 5740 11454 5742 11506
rect 5794 11454 5796 11506
rect 5740 11442 5796 11454
rect 5852 11956 5908 11966
rect 5516 11394 5684 11396
rect 5516 11342 5518 11394
rect 5570 11342 5684 11394
rect 5516 11340 5684 11342
rect 5516 11330 5572 11340
rect 5628 11060 5684 11340
rect 5852 11394 5908 11900
rect 5852 11342 5854 11394
rect 5906 11342 5908 11394
rect 5852 11284 5908 11342
rect 6188 11396 6244 12460
rect 6188 11302 6244 11340
rect 6300 12460 6412 12516
rect 5852 11218 5908 11228
rect 5628 11004 6020 11060
rect 5964 10834 6020 11004
rect 5964 10782 5966 10834
rect 6018 10782 6020 10834
rect 5964 10770 6020 10782
rect 5292 10546 5348 10556
rect 6076 10612 6132 10622
rect 6076 10518 6132 10556
rect 3500 9426 3556 9436
rect 4620 9884 5012 9940
rect 2156 6916 2212 7532
rect 2380 7476 2436 7486
rect 1596 6860 1764 6916
rect 1820 6860 2212 6916
rect 2268 7474 2436 7476
rect 2268 7422 2382 7474
rect 2434 7422 2436 7474
rect 2268 7420 2436 7422
rect 2268 6916 2324 7420
rect 2380 7410 2436 7420
rect 1596 6468 1652 6860
rect 1708 6692 1764 6702
rect 1708 6598 1764 6636
rect 1820 6468 1876 6860
rect 2268 6850 2324 6860
rect 2044 6692 2100 6702
rect 2268 6692 2324 6702
rect 2100 6690 2324 6692
rect 2100 6638 2270 6690
rect 2322 6638 2324 6690
rect 2100 6636 2324 6638
rect 2044 6626 2100 6636
rect 2268 6626 2324 6636
rect 1596 6412 1764 6468
rect 1708 5122 1764 6412
rect 1820 6374 1876 6412
rect 2044 6468 2100 6478
rect 2268 6468 2324 6478
rect 2044 6466 2212 6468
rect 2044 6414 2046 6466
rect 2098 6414 2212 6466
rect 2044 6412 2212 6414
rect 2044 6402 2100 6412
rect 1708 5070 1710 5122
rect 1762 5070 1764 5122
rect 1708 3554 1764 5070
rect 2156 5124 2212 6412
rect 2268 6130 2324 6412
rect 2268 6078 2270 6130
rect 2322 6078 2324 6130
rect 2268 6066 2324 6078
rect 2492 5236 2548 9212
rect 2716 9174 2772 9212
rect 2828 9212 3220 9268
rect 3388 9268 3444 9278
rect 4620 9268 4676 9884
rect 3388 9266 4676 9268
rect 3388 9214 3390 9266
rect 3442 9214 4622 9266
rect 4674 9214 4676 9266
rect 3388 9212 4676 9214
rect 2604 9044 2660 9054
rect 2828 9044 2884 9212
rect 3388 9202 3444 9212
rect 2604 9042 2884 9044
rect 2604 8990 2606 9042
rect 2658 8990 2884 9042
rect 2604 8988 2884 8990
rect 2604 8978 2660 8988
rect 2716 8708 2772 8718
rect 2604 8036 2660 8046
rect 2604 7698 2660 7980
rect 2604 7646 2606 7698
rect 2658 7646 2660 7698
rect 2604 7364 2660 7646
rect 2716 7586 2772 8652
rect 2828 8428 2884 8988
rect 2940 9044 2996 9054
rect 3164 9044 3220 9054
rect 2940 9042 3220 9044
rect 2940 8990 2942 9042
rect 2994 8990 3166 9042
rect 3218 8990 3220 9042
rect 2940 8988 3220 8990
rect 2940 8978 2996 8988
rect 2828 8372 3108 8428
rect 2716 7534 2718 7586
rect 2770 7534 2772 7586
rect 2716 7522 2772 7534
rect 3052 7474 3108 8372
rect 3052 7422 3054 7474
rect 3106 7422 3108 7474
rect 3052 7410 3108 7422
rect 2604 7308 2996 7364
rect 2940 7252 2996 7308
rect 3052 7252 3108 7262
rect 2940 7196 3052 7252
rect 2940 6690 2996 6702
rect 2940 6638 2942 6690
rect 2994 6638 2996 6690
rect 2940 6580 2996 6638
rect 2940 6514 2996 6524
rect 3052 6130 3108 7196
rect 3164 6802 3220 8988
rect 3612 9044 3668 9054
rect 3276 8930 3332 8942
rect 3276 8878 3278 8930
rect 3330 8878 3332 8930
rect 3276 8708 3332 8878
rect 3276 8642 3332 8652
rect 3276 7588 3332 7598
rect 3276 7586 3444 7588
rect 3276 7534 3278 7586
rect 3330 7534 3444 7586
rect 3276 7532 3444 7534
rect 3276 7522 3332 7532
rect 3164 6750 3166 6802
rect 3218 6750 3220 6802
rect 3164 6738 3220 6750
rect 3388 6580 3444 7532
rect 3388 6514 3444 6524
rect 3612 7474 3668 8988
rect 3836 9042 3892 9054
rect 3836 8990 3838 9042
rect 3890 8990 3892 9042
rect 3836 8932 3892 8990
rect 4172 8932 4228 8942
rect 3836 8930 4228 8932
rect 3836 8878 4174 8930
rect 4226 8878 4228 8930
rect 3836 8876 4228 8878
rect 4172 8260 4228 8876
rect 4172 8194 4228 8204
rect 3612 7422 3614 7474
rect 3666 7422 3668 7474
rect 3052 6078 3054 6130
rect 3106 6078 3108 6130
rect 3052 6066 3108 6078
rect 2492 5180 2660 5236
rect 2156 5068 2548 5124
rect 2492 5010 2548 5068
rect 2492 4958 2494 5010
rect 2546 4958 2548 5010
rect 2492 4946 2548 4958
rect 2492 3668 2548 3678
rect 2604 3668 2660 5180
rect 2492 3666 2660 3668
rect 2492 3614 2494 3666
rect 2546 3614 2660 3666
rect 2492 3612 2660 3614
rect 3612 3668 3668 7422
rect 3836 6692 3892 6702
rect 4284 6692 4340 9212
rect 4620 9202 4676 9212
rect 5628 9156 5684 9166
rect 5852 9156 5908 9166
rect 6300 9156 6356 12460
rect 6412 12450 6468 12460
rect 6524 12180 6580 12684
rect 6748 12292 6804 13580
rect 6972 13524 7028 13534
rect 6972 13430 7028 13468
rect 6748 12226 6804 12236
rect 6860 13076 6916 13086
rect 6524 12114 6580 12124
rect 6860 12178 6916 13020
rect 6860 12126 6862 12178
rect 6914 12126 6916 12178
rect 6860 11844 6916 12126
rect 6860 11778 6916 11788
rect 6524 11620 6580 11630
rect 6524 11526 6580 11564
rect 6860 11508 6916 11518
rect 6860 11414 6916 11452
rect 6636 11394 6692 11406
rect 6636 11342 6638 11394
rect 6690 11342 6692 11394
rect 6636 11284 6692 11342
rect 6636 11218 6692 11228
rect 6972 11396 7028 11406
rect 6972 10724 7028 11340
rect 6972 10658 7028 10668
rect 6860 10612 6916 10622
rect 5628 9154 5852 9156
rect 5628 9102 5630 9154
rect 5682 9102 5852 9154
rect 5628 9100 5852 9102
rect 5628 9090 5684 9100
rect 5852 9062 5908 9100
rect 6188 9100 6356 9156
rect 6748 10164 6804 10174
rect 6748 9938 6804 10108
rect 6748 9886 6750 9938
rect 6802 9886 6804 9938
rect 5964 9044 6020 9054
rect 5964 8950 6020 8988
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4508 8372 4564 8382
rect 4508 8278 4564 8316
rect 4956 8260 5012 8270
rect 4508 7476 4564 7486
rect 4844 7476 4900 7486
rect 4508 7382 4564 7420
rect 4620 7474 4900 7476
rect 4620 7422 4846 7474
rect 4898 7422 4900 7474
rect 4620 7420 4900 7422
rect 4620 7250 4676 7420
rect 4844 7410 4900 7420
rect 4620 7198 4622 7250
rect 4674 7198 4676 7250
rect 4620 7186 4676 7198
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4396 6692 4452 6702
rect 4284 6690 4452 6692
rect 4284 6638 4398 6690
rect 4450 6638 4452 6690
rect 4284 6636 4452 6638
rect 3836 6598 3892 6636
rect 4396 6626 4452 6636
rect 4956 6690 5012 8204
rect 5852 8260 5908 8270
rect 5852 8166 5908 8204
rect 5404 7252 5460 7262
rect 5404 7158 5460 7196
rect 4956 6638 4958 6690
rect 5010 6638 5012 6690
rect 4508 6580 4564 6590
rect 3948 6468 4004 6478
rect 3948 6374 4004 6412
rect 4172 6466 4228 6478
rect 4172 6414 4174 6466
rect 4226 6414 4228 6466
rect 2492 3602 2548 3612
rect 3612 3602 3668 3612
rect 1708 3502 1710 3554
rect 1762 3502 1764 3554
rect 1708 3332 1764 3502
rect 1708 3266 1764 3276
rect 3388 3332 3444 3342
rect 3388 2770 3444 3276
rect 4172 2882 4228 6414
rect 4284 6468 4340 6478
rect 4508 6468 4564 6524
rect 4508 6412 4900 6468
rect 4284 6132 4340 6412
rect 4396 6132 4452 6142
rect 4284 6130 4452 6132
rect 4284 6078 4398 6130
rect 4450 6078 4452 6130
rect 4284 6076 4452 6078
rect 4396 6066 4452 6076
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4620 5236 4676 5246
rect 4844 5236 4900 6412
rect 4956 6356 5012 6638
rect 5068 6580 5124 6590
rect 5068 6486 5124 6524
rect 5964 6580 6020 6590
rect 5964 6486 6020 6524
rect 4956 6300 5460 6356
rect 5404 6130 5460 6300
rect 5404 6078 5406 6130
rect 5458 6078 5460 6130
rect 5404 6066 5460 6078
rect 4620 5234 4900 5236
rect 4620 5182 4622 5234
rect 4674 5182 4900 5234
rect 4620 5180 4900 5182
rect 4620 5170 4676 5180
rect 6076 5012 6132 5022
rect 5068 4898 5124 4910
rect 5068 4846 5070 4898
rect 5122 4846 5124 4898
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 4620 3668 4676 3678
rect 4620 3574 4676 3612
rect 5068 3666 5124 4846
rect 6076 4898 6132 4956
rect 6076 4846 6078 4898
rect 6130 4846 6132 4898
rect 6076 4834 6132 4846
rect 5068 3614 5070 3666
rect 5122 3614 5124 3666
rect 5068 3388 5124 3614
rect 6188 3388 6244 9100
rect 6524 9044 6580 9054
rect 6524 8950 6580 8988
rect 6412 8258 6468 8270
rect 6412 8206 6414 8258
rect 6466 8206 6468 8258
rect 6412 7476 6468 8206
rect 6748 8260 6804 9886
rect 6860 8818 6916 10556
rect 7084 9156 7140 13804
rect 7308 12850 7364 12862
rect 7308 12798 7310 12850
rect 7362 12798 7364 12850
rect 7308 12292 7364 12798
rect 7308 12226 7364 12236
rect 7196 12066 7252 12078
rect 7196 12014 7198 12066
rect 7250 12014 7252 12066
rect 7196 11956 7252 12014
rect 7196 11890 7252 11900
rect 7420 10612 7476 14364
rect 10220 13858 10276 14588
rect 10444 14532 10500 14924
rect 10444 13970 10500 14476
rect 10556 14196 10612 15092
rect 10556 14130 10612 14140
rect 10444 13918 10446 13970
rect 10498 13918 10500 13970
rect 10444 13906 10500 13918
rect 10220 13806 10222 13858
rect 10274 13806 10276 13858
rect 10220 13794 10276 13806
rect 9660 13636 9716 13646
rect 9660 13542 9716 13580
rect 10332 13634 10388 13646
rect 10332 13582 10334 13634
rect 10386 13582 10388 13634
rect 9548 13522 9604 13534
rect 9548 13470 9550 13522
rect 9602 13470 9604 13522
rect 8652 12964 8708 12974
rect 8652 12870 8708 12908
rect 9324 12962 9380 12974
rect 9324 12910 9326 12962
rect 9378 12910 9380 12962
rect 7868 12738 7924 12750
rect 7868 12686 7870 12738
rect 7922 12686 7924 12738
rect 7420 10546 7476 10556
rect 7756 11732 7812 11742
rect 7756 11506 7812 11676
rect 7756 11454 7758 11506
rect 7810 11454 7812 11506
rect 7756 10164 7812 11454
rect 7868 11508 7924 12686
rect 8316 12738 8372 12750
rect 8316 12686 8318 12738
rect 8370 12686 8372 12738
rect 8316 12516 8372 12686
rect 9324 12628 9380 12910
rect 9548 12964 9604 13470
rect 10332 13076 10388 13582
rect 10892 13188 10948 18508
rect 11004 18452 11060 18462
rect 11004 18358 11060 18396
rect 11116 16996 11172 22094
rect 11228 21810 11284 22428
rect 11676 22370 11732 22540
rect 11676 22318 11678 22370
rect 11730 22318 11732 22370
rect 11676 22306 11732 22318
rect 11900 22484 11956 22494
rect 11900 22370 11956 22428
rect 11900 22318 11902 22370
rect 11954 22318 11956 22370
rect 11228 21758 11230 21810
rect 11282 21758 11284 21810
rect 11228 21746 11284 21758
rect 11564 21700 11620 21710
rect 11564 21606 11620 21644
rect 11900 21474 11956 22318
rect 11900 21422 11902 21474
rect 11954 21422 11956 21474
rect 11900 21410 11956 21422
rect 11788 19908 11844 19918
rect 11564 19906 11844 19908
rect 11564 19854 11790 19906
rect 11842 19854 11844 19906
rect 11564 19852 11844 19854
rect 11340 19234 11396 19246
rect 11340 19182 11342 19234
rect 11394 19182 11396 19234
rect 11340 18674 11396 19182
rect 11564 19122 11620 19852
rect 11788 19842 11844 19852
rect 11564 19070 11566 19122
rect 11618 19070 11620 19122
rect 11564 19058 11620 19070
rect 11340 18622 11342 18674
rect 11394 18622 11396 18674
rect 11340 18610 11396 18622
rect 11788 18452 11844 18462
rect 11788 18358 11844 18396
rect 11116 16940 11508 16996
rect 11004 16212 11060 16222
rect 11004 15316 11060 16156
rect 11116 16100 11172 16940
rect 11452 16770 11508 16940
rect 11900 16884 11956 16894
rect 12012 16884 12068 27694
rect 12124 26964 12180 29596
rect 12236 29426 12292 29708
rect 12236 29374 12238 29426
rect 12290 29374 12292 29426
rect 12236 29362 12292 29374
rect 12124 26898 12180 26908
rect 12572 26908 12628 34748
rect 12908 30772 12964 30782
rect 12796 29986 12852 29998
rect 12796 29934 12798 29986
rect 12850 29934 12852 29986
rect 12796 29876 12852 29934
rect 12796 29426 12852 29820
rect 12796 29374 12798 29426
rect 12850 29374 12852 29426
rect 12684 28756 12740 28766
rect 12684 28662 12740 28700
rect 12796 28644 12852 29374
rect 12796 28578 12852 28588
rect 12908 27860 12964 30716
rect 13020 29092 13076 29102
rect 13132 29092 13188 36988
rect 13580 35252 13636 35262
rect 13580 34692 13636 35196
rect 13580 34598 13636 34636
rect 13468 31666 13524 31678
rect 13468 31614 13470 31666
rect 13522 31614 13524 31666
rect 13468 30434 13524 31614
rect 13468 30382 13470 30434
rect 13522 30382 13524 30434
rect 13468 30370 13524 30382
rect 13244 29988 13300 29998
rect 13300 29932 13412 29988
rect 13244 29922 13300 29932
rect 13356 29538 13412 29932
rect 13356 29486 13358 29538
rect 13410 29486 13412 29538
rect 13356 29474 13412 29486
rect 13244 29428 13300 29438
rect 13244 29334 13300 29372
rect 13076 29036 13188 29092
rect 13020 29026 13076 29036
rect 13356 28756 13412 28766
rect 13356 28644 13412 28700
rect 13580 28644 13636 28654
rect 13356 28588 13524 28644
rect 13356 27860 13412 27870
rect 12908 27858 13412 27860
rect 12908 27806 13358 27858
rect 13410 27806 13412 27858
rect 12908 27804 13412 27806
rect 13356 27794 13412 27804
rect 13468 27746 13524 28588
rect 13580 28550 13636 28588
rect 13468 27694 13470 27746
rect 13522 27694 13524 27746
rect 13468 27682 13524 27694
rect 13692 26908 13748 38668
rect 14028 33572 14084 40348
rect 14476 40292 14532 41916
rect 14476 40226 14532 40236
rect 14588 38668 14644 51660
rect 14700 51492 14756 51502
rect 14700 51490 14868 51492
rect 14700 51438 14702 51490
rect 14754 51438 14868 51490
rect 14700 51436 14868 51438
rect 14700 51426 14756 51436
rect 14812 49924 14868 51436
rect 14924 50596 14980 50606
rect 14924 50370 14980 50540
rect 15260 50428 15316 60620
rect 15596 60452 15652 63084
rect 15596 59330 15652 60396
rect 16492 60898 16548 67900
rect 16828 67842 16884 67900
rect 16828 67790 16830 67842
rect 16882 67790 16884 67842
rect 16828 67778 16884 67790
rect 17388 65380 17444 73948
rect 17500 73938 17556 73948
rect 18620 73938 18676 73948
rect 19404 73554 19460 73948
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 19404 73502 19406 73554
rect 19458 73502 19460 73554
rect 19404 73490 19460 73502
rect 19628 73332 19684 73342
rect 19516 73330 19684 73332
rect 19516 73278 19630 73330
rect 19682 73278 19684 73330
rect 19516 73276 19684 73278
rect 18956 73218 19012 73230
rect 18956 73166 18958 73218
rect 19010 73166 19012 73218
rect 18956 73108 19012 73166
rect 19180 73108 19236 73118
rect 19292 73108 19348 73118
rect 18956 73052 19180 73108
rect 19236 73106 19348 73108
rect 19236 73054 19294 73106
rect 19346 73054 19348 73106
rect 19236 73052 19348 73054
rect 17724 71652 17780 71662
rect 17724 70644 17780 71596
rect 17724 70194 17780 70588
rect 17724 70142 17726 70194
rect 17778 70142 17780 70194
rect 17724 70130 17780 70142
rect 19180 71204 19236 73052
rect 19292 73042 19348 73052
rect 18396 70084 18452 70094
rect 18396 70082 18788 70084
rect 18396 70030 18398 70082
rect 18450 70030 18788 70082
rect 18396 70028 18788 70030
rect 18396 70018 18452 70028
rect 18732 69410 18788 70028
rect 18732 69358 18734 69410
rect 18786 69358 18788 69410
rect 18732 69346 18788 69358
rect 18508 69300 18564 69310
rect 18508 69206 18564 69244
rect 19068 69300 19124 69310
rect 19068 69206 19124 69244
rect 18956 69186 19012 69198
rect 18956 69134 18958 69186
rect 19010 69134 19012 69186
rect 18956 68852 19012 69134
rect 18956 68786 19012 68796
rect 17500 67732 17556 67742
rect 17500 67730 18004 67732
rect 17500 67678 17502 67730
rect 17554 67678 18004 67730
rect 17500 67676 18004 67678
rect 17500 67666 17556 67676
rect 17948 67282 18004 67676
rect 17948 67230 17950 67282
rect 18002 67230 18004 67282
rect 17948 67218 18004 67230
rect 18284 67060 18340 67070
rect 18284 66966 18340 67004
rect 17948 65490 18004 65502
rect 17948 65438 17950 65490
rect 18002 65438 18004 65490
rect 17612 65380 17668 65390
rect 17948 65380 18004 65438
rect 17388 65378 18004 65380
rect 17388 65326 17614 65378
rect 17666 65326 18004 65378
rect 17388 65324 18004 65326
rect 18732 65380 18788 65390
rect 16828 63924 16884 63934
rect 17388 63924 17444 63934
rect 17612 63924 17668 65324
rect 18732 65286 18788 65324
rect 16828 63922 17668 63924
rect 16828 63870 16830 63922
rect 16882 63870 17390 63922
rect 17442 63870 17668 63922
rect 16828 63868 17668 63870
rect 18508 64594 18564 64606
rect 18508 64542 18510 64594
rect 18562 64542 18564 64594
rect 16828 63140 16884 63868
rect 17388 63858 17444 63868
rect 16828 63074 16884 63084
rect 18172 63810 18228 63822
rect 18172 63758 18174 63810
rect 18226 63758 18228 63810
rect 17724 62468 17780 62478
rect 17724 62374 17780 62412
rect 17948 62466 18004 62478
rect 17948 62414 17950 62466
rect 18002 62414 18004 62466
rect 17948 62244 18004 62414
rect 17948 62178 18004 62188
rect 18060 62244 18116 62254
rect 18172 62244 18228 63758
rect 18508 63250 18564 64542
rect 18508 63198 18510 63250
rect 18562 63198 18564 63250
rect 18508 63186 18564 63198
rect 18620 64482 18676 64494
rect 18620 64430 18622 64482
rect 18674 64430 18676 64482
rect 18620 62804 18676 64430
rect 19180 63364 19236 71148
rect 19516 68068 19572 73276
rect 19628 73266 19684 73276
rect 20636 73108 20692 75628
rect 20748 75590 20804 75628
rect 21644 75684 21700 75694
rect 21644 75590 21700 75628
rect 22428 75684 22484 75694
rect 22764 75684 22820 75694
rect 22484 75682 22820 75684
rect 22484 75630 22766 75682
rect 22818 75630 22820 75682
rect 22484 75628 22820 75630
rect 22428 75590 22484 75628
rect 22764 75618 22820 75628
rect 23100 75684 23156 75694
rect 23436 75684 23492 75694
rect 23100 75682 23492 75684
rect 23100 75630 23102 75682
rect 23154 75630 23438 75682
rect 23490 75630 23492 75682
rect 23100 75628 23492 75630
rect 23100 75618 23156 75628
rect 21420 75458 21476 75470
rect 21420 75406 21422 75458
rect 21474 75406 21476 75458
rect 20748 74228 20804 74238
rect 21308 74228 21364 74238
rect 20748 74226 21364 74228
rect 20748 74174 20750 74226
rect 20802 74174 21310 74226
rect 21362 74174 21364 74226
rect 20748 74172 21364 74174
rect 20748 74162 20804 74172
rect 21308 74162 21364 74172
rect 21420 74004 21476 75406
rect 21420 74002 21588 74004
rect 21420 73950 21422 74002
rect 21474 73950 21588 74002
rect 21420 73948 21588 73950
rect 21420 73938 21476 73948
rect 20636 73042 20692 73052
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 20300 71764 20356 71774
rect 20748 71764 20804 71774
rect 20300 71762 20916 71764
rect 20300 71710 20302 71762
rect 20354 71710 20750 71762
rect 20802 71710 20916 71762
rect 20300 71708 20916 71710
rect 20300 71652 20356 71708
rect 20748 71698 20804 71708
rect 20300 71586 20356 71596
rect 20748 71204 20804 71214
rect 20748 71090 20804 71148
rect 20748 71038 20750 71090
rect 20802 71038 20804 71090
rect 20748 71026 20804 71038
rect 20860 70644 20916 71708
rect 21420 71650 21476 71662
rect 21420 71598 21422 71650
rect 21474 71598 21476 71650
rect 21420 71090 21476 71598
rect 21420 71038 21422 71090
rect 21474 71038 21476 71090
rect 21420 71026 21476 71038
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20860 70578 20916 70588
rect 21420 70754 21476 70766
rect 21420 70702 21422 70754
rect 21474 70702 21476 70754
rect 19836 70522 20100 70532
rect 20524 70084 20580 70094
rect 20860 70084 20916 70094
rect 20524 70082 20916 70084
rect 20524 70030 20526 70082
rect 20578 70030 20862 70082
rect 20914 70030 20916 70082
rect 20524 70028 20916 70030
rect 20524 70018 20580 70028
rect 20860 70018 20916 70028
rect 20972 69970 21028 69982
rect 20972 69918 20974 69970
rect 21026 69918 21028 69970
rect 20972 69412 21028 69918
rect 21420 69412 21476 70702
rect 20972 69410 21476 69412
rect 20972 69358 21422 69410
rect 21474 69358 21476 69410
rect 20972 69356 21476 69358
rect 21420 69346 21476 69356
rect 21532 69412 21588 73948
rect 21644 71204 21700 71214
rect 21644 71110 21700 71148
rect 22876 70978 22932 70990
rect 22876 70926 22878 70978
rect 22930 70926 22932 70978
rect 22428 70754 22484 70766
rect 22428 70702 22430 70754
rect 22482 70702 22484 70754
rect 22428 70644 22484 70702
rect 22428 70578 22484 70588
rect 22876 70644 22932 70926
rect 22876 70578 22932 70588
rect 23100 70194 23156 70206
rect 23100 70142 23102 70194
rect 23154 70142 23156 70194
rect 21532 69346 21588 69356
rect 21868 69410 21924 69422
rect 21868 69358 21870 69410
rect 21922 69358 21924 69410
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 19740 68852 19796 68862
rect 19796 68796 20132 68852
rect 19740 68758 19796 68796
rect 20076 68628 20132 68796
rect 20300 68628 20356 68638
rect 20076 68626 20356 68628
rect 20076 68574 20302 68626
rect 20354 68574 20356 68626
rect 20076 68572 20356 68574
rect 20300 68562 20356 68572
rect 20860 68628 20916 68638
rect 20860 68534 20916 68572
rect 21420 68626 21476 68638
rect 21420 68574 21422 68626
rect 21474 68574 21476 68626
rect 19516 68002 19572 68012
rect 19628 68514 19684 68526
rect 19628 68462 19630 68514
rect 19682 68462 19684 68514
rect 19628 67954 19684 68462
rect 20300 68068 20356 68078
rect 20300 67974 20356 68012
rect 21420 68068 21476 68574
rect 21868 68628 21924 69358
rect 22540 69412 22596 69422
rect 22540 69318 22596 69356
rect 23100 69410 23156 70142
rect 23436 70194 23492 75628
rect 24220 75684 24276 75694
rect 24220 75590 24276 75628
rect 24556 75682 24612 75740
rect 26796 75796 26852 76300
rect 27804 75906 27860 77086
rect 30940 77138 31220 77140
rect 30940 77086 31166 77138
rect 31218 77086 31220 77138
rect 30940 77084 31220 77086
rect 28140 77028 28196 77038
rect 27916 77026 28196 77028
rect 27916 76974 28142 77026
rect 28194 76974 28196 77026
rect 27916 76972 28196 76974
rect 27916 76578 27972 76972
rect 28140 76962 28196 76972
rect 30940 76690 30996 77084
rect 31164 77074 31220 77084
rect 30940 76638 30942 76690
rect 30994 76638 30996 76690
rect 30940 76626 30996 76638
rect 27916 76526 27918 76578
rect 27970 76526 27972 76578
rect 27916 76514 27972 76526
rect 30604 76466 30660 76478
rect 30604 76414 30606 76466
rect 30658 76414 30660 76466
rect 30044 76356 30100 76366
rect 27804 75854 27806 75906
rect 27858 75854 27860 75906
rect 27804 75842 27860 75854
rect 29932 76354 30100 76356
rect 29932 76302 30046 76354
rect 30098 76302 30100 76354
rect 29932 76300 30100 76302
rect 26796 75730 26852 75740
rect 27468 75796 27524 75806
rect 28140 75796 28196 75806
rect 27468 75794 27636 75796
rect 27468 75742 27470 75794
rect 27522 75742 27636 75794
rect 27468 75740 27636 75742
rect 27468 75730 27524 75740
rect 24556 75630 24558 75682
rect 24610 75630 24612 75682
rect 24108 74900 24164 74910
rect 23548 72322 23604 72334
rect 23548 72270 23550 72322
rect 23602 72270 23604 72322
rect 23548 72100 23604 72270
rect 24108 72100 24164 74844
rect 24220 74788 24276 74798
rect 24556 74788 24612 75630
rect 25228 75684 25284 75694
rect 25228 75348 25284 75628
rect 25340 75572 25396 75582
rect 25340 75570 25620 75572
rect 25340 75518 25342 75570
rect 25394 75518 25620 75570
rect 25340 75516 25620 75518
rect 25340 75506 25396 75516
rect 25228 75292 25396 75348
rect 25340 75012 25396 75292
rect 25564 75122 25620 75516
rect 25564 75070 25566 75122
rect 25618 75070 25620 75122
rect 25564 75058 25620 75070
rect 27580 75460 27636 75740
rect 28140 75702 28196 75740
rect 29372 75796 29428 75806
rect 29260 75684 29316 75694
rect 29372 75684 29428 75740
rect 29260 75682 29428 75684
rect 29260 75630 29262 75682
rect 29314 75630 29428 75682
rect 29260 75628 29428 75630
rect 29260 75618 29316 75628
rect 28364 75570 28420 75582
rect 28364 75518 28366 75570
rect 28418 75518 28420 75570
rect 28364 75460 28420 75518
rect 27580 75404 28420 75460
rect 25340 75010 25508 75012
rect 25340 74958 25342 75010
rect 25394 74958 25508 75010
rect 25340 74956 25508 74958
rect 25340 74946 25396 74956
rect 25228 74900 25284 74910
rect 25228 74806 25284 74844
rect 24220 74786 24612 74788
rect 24220 74734 24222 74786
rect 24274 74734 24612 74786
rect 24220 74732 24612 74734
rect 24220 73220 24276 74732
rect 24220 73154 24276 73164
rect 25228 73220 25284 73230
rect 23548 72044 24164 72100
rect 23772 71762 23828 71774
rect 23772 71710 23774 71762
rect 23826 71710 23828 71762
rect 23660 71652 23716 71662
rect 23548 71623 23660 71652
rect 23548 71571 23550 71623
rect 23602 71596 23660 71623
rect 23602 71571 23604 71596
rect 23660 71586 23716 71596
rect 23548 71559 23604 71571
rect 23548 71092 23604 71102
rect 23772 71092 23828 71710
rect 23548 71090 23828 71092
rect 23548 71038 23550 71090
rect 23602 71038 23828 71090
rect 23548 71036 23828 71038
rect 23548 71026 23604 71036
rect 23436 70142 23438 70194
rect 23490 70142 23492 70194
rect 23436 70130 23492 70142
rect 23324 70082 23380 70094
rect 23324 70030 23326 70082
rect 23378 70030 23380 70082
rect 23324 69524 23380 70030
rect 23436 69524 23492 69534
rect 23324 69522 23492 69524
rect 23324 69470 23438 69522
rect 23490 69470 23492 69522
rect 23324 69468 23492 69470
rect 23100 69358 23102 69410
rect 23154 69358 23156 69410
rect 22316 69298 22372 69310
rect 22316 69246 22318 69298
rect 22370 69246 22372 69298
rect 21868 68562 21924 68572
rect 21980 68852 22036 68862
rect 21980 68626 22036 68796
rect 21980 68574 21982 68626
rect 22034 68574 22036 68626
rect 21980 68562 22036 68574
rect 21868 68404 21924 68414
rect 21868 68310 21924 68348
rect 21420 68002 21476 68012
rect 19628 67902 19630 67954
rect 19682 67902 19684 67954
rect 19628 67890 19684 67902
rect 20412 67732 20468 67742
rect 21420 67732 21476 67742
rect 20412 67730 21476 67732
rect 20412 67678 20414 67730
rect 20466 67678 21422 67730
rect 21474 67678 21476 67730
rect 20412 67676 21476 67678
rect 20412 67666 20468 67676
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 19068 63362 19236 63364
rect 19068 63310 19182 63362
rect 19234 63310 19236 63362
rect 19068 63308 19236 63310
rect 18956 63252 19012 63262
rect 18956 63158 19012 63196
rect 18060 62242 18228 62244
rect 18060 62190 18062 62242
rect 18114 62190 18228 62242
rect 18060 62188 18228 62190
rect 18396 62748 18676 62804
rect 18844 63138 18900 63150
rect 18844 63086 18846 63138
rect 18898 63086 18900 63138
rect 18396 62244 18452 62748
rect 18508 62468 18564 62478
rect 18508 62374 18564 62412
rect 18508 62244 18564 62254
rect 18396 62188 18508 62244
rect 18060 62178 18116 62188
rect 17836 61570 17892 61582
rect 17836 61518 17838 61570
rect 17890 61518 17892 61570
rect 16492 60846 16494 60898
rect 16546 60846 16548 60898
rect 15708 59892 15764 59902
rect 15708 59798 15764 59836
rect 16492 59444 16548 60846
rect 17500 61348 17556 61358
rect 17836 61348 17892 61518
rect 17500 61346 17892 61348
rect 17500 61294 17502 61346
rect 17554 61294 17892 61346
rect 17500 61292 17892 61294
rect 17500 60452 17556 61292
rect 17500 60386 17556 60396
rect 18284 60452 18340 60462
rect 17836 60116 17892 60126
rect 17836 60114 18004 60116
rect 17836 60062 17838 60114
rect 17890 60062 18004 60114
rect 17836 60060 18004 60062
rect 17836 60050 17892 60060
rect 16940 59444 16996 59454
rect 16492 59442 16996 59444
rect 16492 59390 16942 59442
rect 16994 59390 16996 59442
rect 16492 59388 16996 59390
rect 15596 59278 15598 59330
rect 15650 59278 15652 59330
rect 15596 59108 15652 59278
rect 15596 58434 15652 59052
rect 16268 59332 16324 59342
rect 16268 58546 16324 59276
rect 16380 59332 16436 59342
rect 16492 59332 16548 59388
rect 16940 59378 16996 59388
rect 16380 59330 16548 59332
rect 16380 59278 16382 59330
rect 16434 59278 16548 59330
rect 16380 59276 16548 59278
rect 17388 59332 17444 59342
rect 16380 59266 16436 59276
rect 17388 59238 17444 59276
rect 17612 59220 17668 59230
rect 16268 58494 16270 58546
rect 16322 58494 16324 58546
rect 16268 58482 16324 58494
rect 17500 59218 17668 59220
rect 17500 59166 17614 59218
rect 17666 59166 17668 59218
rect 17500 59164 17668 59166
rect 15596 58382 15598 58434
rect 15650 58382 15652 58434
rect 15596 58370 15652 58382
rect 17388 57876 17444 57886
rect 17500 57876 17556 59164
rect 17612 59154 17668 59164
rect 17388 57874 17556 57876
rect 17388 57822 17390 57874
rect 17442 57822 17556 57874
rect 17388 57820 17556 57822
rect 17388 57810 17444 57820
rect 17948 57762 18004 60060
rect 18284 60114 18340 60396
rect 18284 60062 18286 60114
rect 18338 60062 18340 60114
rect 18060 59892 18116 59902
rect 18060 59442 18116 59836
rect 18060 59390 18062 59442
rect 18114 59390 18116 59442
rect 18060 59378 18116 59390
rect 18284 59108 18340 60062
rect 18508 59556 18564 62188
rect 18620 61460 18676 61470
rect 18620 61366 18676 61404
rect 18508 59490 18564 59500
rect 18844 59444 18900 63086
rect 18956 62468 19012 62478
rect 19068 62468 19124 63308
rect 19180 63298 19236 63308
rect 20300 63810 20356 63822
rect 20300 63758 20302 63810
rect 20354 63758 20356 63810
rect 19628 63140 19684 63150
rect 19628 63046 19684 63084
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 19628 62468 19684 62478
rect 19012 62412 19348 62468
rect 18956 62374 19012 62412
rect 19292 62188 19348 62412
rect 19628 62374 19684 62412
rect 20300 62468 20356 63758
rect 20300 62402 20356 62412
rect 20412 62916 20468 62926
rect 19292 62132 19460 62188
rect 19404 60674 19460 62132
rect 19740 62132 19796 62142
rect 19740 62130 20244 62132
rect 19740 62078 19742 62130
rect 19794 62078 20244 62130
rect 19740 62076 20244 62078
rect 19740 62066 19796 62076
rect 19516 61460 19572 61470
rect 19572 61404 19684 61460
rect 19516 61394 19572 61404
rect 19628 61012 19684 61404
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 19852 61012 19908 61022
rect 19628 61010 19908 61012
rect 19628 60958 19854 61010
rect 19906 60958 19908 61010
rect 19628 60956 19908 60958
rect 19852 60946 19908 60956
rect 19404 60622 19406 60674
rect 19458 60622 19460 60674
rect 19404 60564 19460 60622
rect 19964 60898 20020 60910
rect 19964 60846 19966 60898
rect 20018 60846 20020 60898
rect 19740 60564 19796 60574
rect 19404 60562 19796 60564
rect 19404 60510 19742 60562
rect 19794 60510 19796 60562
rect 19404 60508 19796 60510
rect 19740 60004 19796 60508
rect 19740 59938 19796 59948
rect 19964 59780 20020 60846
rect 19628 59724 20020 59780
rect 18620 59388 18900 59444
rect 19516 59556 19572 59566
rect 18396 59220 18452 59230
rect 18396 59126 18452 59164
rect 18284 59042 18340 59052
rect 18396 58546 18452 58558
rect 18396 58494 18398 58546
rect 18450 58494 18452 58546
rect 17948 57710 17950 57762
rect 18002 57710 18004 57762
rect 17948 57652 18004 57710
rect 17948 57586 18004 57596
rect 18284 58324 18340 58334
rect 18284 57650 18340 58268
rect 18284 57598 18286 57650
rect 18338 57598 18340 57650
rect 17724 57426 17780 57438
rect 17724 57374 17726 57426
rect 17778 57374 17780 57426
rect 17052 56868 17108 56878
rect 17052 55522 17108 56812
rect 17724 56644 17780 57374
rect 18284 57204 18340 57598
rect 18284 57138 18340 57148
rect 18396 58212 18452 58494
rect 17724 56578 17780 56588
rect 18172 56644 18228 56654
rect 18172 56550 18228 56588
rect 17052 55470 17054 55522
rect 17106 55470 17108 55522
rect 17052 55458 17108 55470
rect 18060 55412 18116 55422
rect 18396 55412 18452 58156
rect 18508 57652 18564 57662
rect 18508 57558 18564 57596
rect 18620 56868 18676 59388
rect 18844 59108 18900 59118
rect 18844 59014 18900 59052
rect 19292 59108 19348 59118
rect 18844 58324 18900 58334
rect 18844 58230 18900 58268
rect 19292 58322 19348 59052
rect 19292 58270 19294 58322
rect 19346 58270 19348 58322
rect 19292 58258 19348 58270
rect 19068 58212 19124 58222
rect 19068 58118 19124 58156
rect 19404 58210 19460 58222
rect 19404 58158 19406 58210
rect 19458 58158 19460 58210
rect 18620 56802 18676 56812
rect 18732 57762 18788 57774
rect 18732 57710 18734 57762
rect 18786 57710 18788 57762
rect 18060 55410 18452 55412
rect 18060 55358 18062 55410
rect 18114 55358 18452 55410
rect 18060 55356 18452 55358
rect 18508 56644 18564 56654
rect 18060 55346 18116 55356
rect 17836 55298 17892 55310
rect 17836 55246 17838 55298
rect 17890 55246 17892 55298
rect 16940 55188 16996 55198
rect 16604 55186 16996 55188
rect 16604 55134 16942 55186
rect 16994 55134 16996 55186
rect 16604 55132 16996 55134
rect 16604 54402 16660 55132
rect 16940 55122 16996 55132
rect 17500 55076 17556 55086
rect 17836 55076 17892 55246
rect 17500 55074 17668 55076
rect 17500 55022 17502 55074
rect 17554 55022 17668 55074
rect 17500 55020 17668 55022
rect 17500 55010 17556 55020
rect 17388 54628 17444 54638
rect 16604 54350 16606 54402
rect 16658 54350 16660 54402
rect 16604 54338 16660 54350
rect 17052 54626 17444 54628
rect 17052 54574 17390 54626
rect 17442 54574 17444 54626
rect 17052 54572 17444 54574
rect 16380 54292 16436 54302
rect 15932 53732 15988 53742
rect 16380 53732 16436 54236
rect 17052 53842 17108 54572
rect 17388 54562 17444 54572
rect 17612 54514 17668 55020
rect 17836 55010 17892 55020
rect 18508 55076 18564 56588
rect 18508 54982 18564 55020
rect 18732 56642 18788 57710
rect 18956 57650 19012 57662
rect 18956 57598 18958 57650
rect 19010 57598 19012 57650
rect 18844 57540 18900 57550
rect 18956 57540 19012 57598
rect 18844 57538 19012 57540
rect 18844 57486 18846 57538
rect 18898 57486 19012 57538
rect 18844 57484 19012 57486
rect 18844 57474 18900 57484
rect 18732 56590 18734 56642
rect 18786 56590 18788 56642
rect 18732 54740 18788 56590
rect 18732 54674 18788 54684
rect 18844 57204 18900 57214
rect 17612 54462 17614 54514
rect 17666 54462 17668 54514
rect 17612 54450 17668 54462
rect 18172 54402 18228 54414
rect 18172 54350 18174 54402
rect 18226 54350 18228 54402
rect 18172 54292 18228 54350
rect 18844 54404 18900 57148
rect 19404 56866 19460 58158
rect 19404 56814 19406 56866
rect 19458 56814 19460 56866
rect 19404 56802 19460 56814
rect 19516 56756 19572 59500
rect 19628 59332 19684 59724
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 19628 59276 19796 59332
rect 19628 59108 19684 59118
rect 19628 59014 19684 59052
rect 19740 58212 19796 59276
rect 19852 58324 19908 58334
rect 19852 58230 19908 58268
rect 19628 58156 19796 58212
rect 19628 57764 19684 58156
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 19852 57764 19908 57774
rect 19628 57708 19796 57764
rect 19740 57092 19796 57708
rect 19740 57026 19796 57036
rect 19852 57090 19908 57708
rect 19852 57038 19854 57090
rect 19906 57038 19908 57090
rect 19852 57026 19908 57038
rect 19964 57650 20020 57662
rect 19964 57598 19966 57650
rect 20018 57598 20020 57650
rect 19740 56866 19796 56878
rect 19740 56814 19742 56866
rect 19794 56814 19796 56866
rect 19740 56756 19796 56814
rect 19852 56868 19908 56878
rect 19964 56868 20020 57598
rect 19908 56812 20020 56868
rect 20076 57426 20132 57438
rect 20076 57374 20078 57426
rect 20130 57374 20132 57426
rect 19852 56802 19908 56812
rect 19516 56700 19796 56756
rect 20076 56756 20132 57374
rect 20076 56690 20132 56700
rect 19068 56644 19124 56654
rect 18844 54402 19012 54404
rect 18844 54350 18846 54402
rect 18898 54350 19012 54402
rect 18844 54348 19012 54350
rect 18844 54338 18900 54348
rect 18172 54226 18228 54236
rect 17052 53790 17054 53842
rect 17106 53790 17108 53842
rect 17052 53778 17108 53790
rect 15932 53730 16436 53732
rect 15932 53678 15934 53730
rect 15986 53678 16382 53730
rect 16434 53678 16436 53730
rect 15932 53676 16436 53678
rect 15932 53666 15988 53676
rect 16380 53666 16436 53676
rect 18956 53732 19012 54348
rect 15372 53618 15428 53630
rect 15372 53566 15374 53618
rect 15426 53566 15428 53618
rect 15372 52836 15428 53566
rect 15372 52770 15428 52780
rect 18284 53620 18340 53630
rect 17948 51492 18004 51502
rect 15820 50708 15876 50718
rect 15820 50614 15876 50652
rect 17948 50706 18004 51436
rect 17948 50654 17950 50706
rect 18002 50654 18004 50706
rect 17948 50642 18004 50654
rect 16156 50596 16212 50606
rect 15260 50372 15428 50428
rect 14924 50318 14926 50370
rect 14978 50318 14980 50370
rect 14924 50148 14980 50318
rect 14924 50092 15092 50148
rect 14924 49924 14980 49934
rect 14812 49922 14980 49924
rect 14812 49870 14926 49922
rect 14978 49870 14980 49922
rect 14812 49868 14980 49870
rect 14924 49858 14980 49868
rect 14924 49700 14980 49710
rect 14924 49138 14980 49644
rect 14924 49086 14926 49138
rect 14978 49086 14980 49138
rect 14700 49026 14756 49038
rect 14700 48974 14702 49026
rect 14754 48974 14756 49026
rect 14700 48580 14756 48974
rect 14924 48916 14980 49086
rect 14924 48850 14980 48860
rect 14756 48524 14980 48580
rect 14700 48514 14756 48524
rect 14924 48468 14980 48524
rect 15036 48468 15092 50092
rect 15148 48468 15204 48478
rect 14924 48466 15204 48468
rect 14924 48414 15150 48466
rect 15202 48414 15204 48466
rect 14924 48412 15204 48414
rect 15148 48402 15204 48412
rect 15372 47068 15428 50372
rect 15484 50372 15540 50382
rect 15484 50370 15652 50372
rect 15484 50318 15486 50370
rect 15538 50318 15652 50370
rect 15484 50316 15652 50318
rect 15484 50306 15540 50316
rect 15596 49810 15652 50316
rect 15596 49758 15598 49810
rect 15650 49758 15652 49810
rect 15596 49700 15652 49758
rect 15484 49028 15540 49038
rect 15596 49028 15652 49644
rect 16156 49700 16212 50540
rect 17724 50484 17780 50494
rect 16156 49606 16212 49644
rect 16604 49812 16660 49822
rect 15484 49026 15652 49028
rect 15484 48974 15486 49026
rect 15538 48974 15652 49026
rect 15484 48972 15652 48974
rect 15484 48804 15540 48972
rect 16268 48916 16324 48926
rect 16268 48914 16436 48916
rect 16268 48862 16270 48914
rect 16322 48862 16436 48914
rect 16268 48860 16436 48862
rect 16268 48850 16324 48860
rect 15484 48738 15540 48748
rect 16156 48468 16212 48478
rect 16212 48412 16324 48468
rect 16156 48374 16212 48412
rect 15372 47012 15540 47068
rect 15372 46564 15428 46574
rect 15372 46470 15428 46508
rect 15484 46340 15540 47012
rect 15372 46284 15540 46340
rect 16156 46676 16212 46686
rect 14924 45892 14980 45902
rect 14924 45778 14980 45836
rect 14924 45726 14926 45778
rect 14978 45726 14980 45778
rect 14924 45714 14980 45726
rect 15148 44098 15204 44110
rect 15148 44046 15150 44098
rect 15202 44046 15204 44098
rect 15148 43708 15204 44046
rect 14700 43652 15204 43708
rect 14700 43650 14756 43652
rect 14700 43598 14702 43650
rect 14754 43598 14756 43650
rect 14700 43586 14756 43598
rect 14812 43540 14868 43550
rect 14812 42194 14868 43484
rect 14812 42142 14814 42194
rect 14866 42142 14868 42194
rect 14812 39620 14868 42142
rect 15372 41972 15428 46284
rect 16156 45890 16212 46620
rect 16156 45838 16158 45890
rect 16210 45838 16212 45890
rect 15708 45668 15764 45678
rect 15708 45574 15764 45612
rect 16156 45668 16212 45838
rect 16156 45602 16212 45612
rect 16268 44436 16324 48412
rect 16380 48466 16436 48860
rect 16380 48414 16382 48466
rect 16434 48414 16436 48466
rect 16380 48402 16436 48414
rect 16604 48354 16660 49756
rect 17612 48804 17668 48814
rect 16604 48302 16606 48354
rect 16658 48302 16660 48354
rect 16380 47570 16436 47582
rect 16380 47518 16382 47570
rect 16434 47518 16436 47570
rect 16380 45780 16436 47518
rect 16604 46676 16660 48302
rect 16716 48468 16772 48478
rect 16716 48354 16772 48412
rect 16716 48302 16718 48354
rect 16770 48302 16772 48354
rect 16716 48290 16772 48302
rect 16828 47236 16884 47246
rect 16828 46676 16884 47180
rect 17612 46898 17668 48748
rect 17612 46846 17614 46898
rect 17666 46846 17668 46898
rect 17612 46834 17668 46846
rect 16604 46620 16772 46676
rect 16604 45780 16660 45790
rect 16380 45724 16604 45780
rect 16156 44380 16268 44436
rect 15484 44212 15540 44222
rect 16044 44212 16100 44222
rect 15484 44210 16100 44212
rect 15484 44158 15486 44210
rect 15538 44158 16046 44210
rect 16098 44158 16100 44210
rect 15484 44156 16100 44158
rect 15484 44146 15540 44156
rect 16044 44146 16100 44156
rect 16156 43876 16212 44380
rect 16268 44370 16324 44380
rect 16492 44994 16548 45006
rect 16492 44942 16494 44994
rect 16546 44942 16548 44994
rect 15372 41906 15428 41916
rect 15932 43820 16212 43876
rect 16380 44322 16436 44334
rect 16380 44270 16382 44322
rect 16434 44270 16436 44322
rect 16380 44100 16436 44270
rect 15932 41298 15988 43820
rect 15932 41246 15934 41298
rect 15986 41246 15988 41298
rect 15932 41234 15988 41246
rect 16044 43652 16100 43662
rect 16380 43652 16436 44044
rect 16100 43596 16436 43652
rect 15372 40404 15428 40414
rect 15260 40402 15428 40404
rect 15260 40350 15374 40402
rect 15426 40350 15428 40402
rect 15260 40348 15428 40350
rect 14812 39554 14868 39564
rect 14924 40292 14980 40302
rect 14700 39508 14756 39518
rect 14700 39414 14756 39452
rect 14476 38612 14644 38668
rect 14700 38722 14756 38734
rect 14700 38670 14702 38722
rect 14754 38670 14756 38722
rect 14364 37156 14420 37166
rect 14252 34914 14308 34926
rect 14252 34862 14254 34914
rect 14306 34862 14308 34914
rect 14028 33570 14196 33572
rect 14028 33518 14030 33570
rect 14082 33518 14196 33570
rect 14028 33516 14196 33518
rect 14028 33506 14084 33516
rect 13804 33236 13860 33246
rect 13804 33142 13860 33180
rect 14140 31948 14196 33516
rect 14252 32452 14308 34862
rect 14364 34130 14420 37100
rect 14364 34078 14366 34130
rect 14418 34078 14420 34130
rect 14364 34066 14420 34078
rect 14364 33572 14420 33582
rect 14476 33572 14532 38612
rect 14700 38052 14756 38670
rect 14700 37986 14756 37996
rect 14700 36932 14756 36942
rect 14700 36484 14756 36876
rect 14700 36390 14756 36428
rect 14364 33570 14532 33572
rect 14364 33518 14366 33570
rect 14418 33518 14532 33570
rect 14364 33516 14532 33518
rect 14364 33506 14420 33516
rect 14364 32452 14420 32462
rect 14252 32450 14420 32452
rect 14252 32398 14366 32450
rect 14418 32398 14420 32450
rect 14252 32396 14420 32398
rect 14364 32386 14420 32396
rect 14700 32452 14756 32462
rect 14140 31892 14644 31948
rect 13804 31556 13860 31566
rect 13804 31554 14196 31556
rect 13804 31502 13806 31554
rect 13858 31502 14196 31554
rect 13804 31500 14196 31502
rect 13804 31490 13860 31500
rect 14140 31106 14196 31500
rect 14140 31054 14142 31106
rect 14194 31054 14196 31106
rect 14140 31042 14196 31054
rect 14476 30322 14532 31892
rect 14588 31890 14644 31892
rect 14588 31838 14590 31890
rect 14642 31838 14644 31890
rect 14588 31826 14644 31838
rect 14476 30270 14478 30322
rect 14530 30270 14532 30322
rect 13804 30212 13860 30222
rect 13804 30118 13860 30156
rect 14476 30212 14532 30270
rect 14028 30100 14084 30110
rect 13916 30044 14028 30100
rect 13916 29314 13972 30044
rect 14028 30006 14084 30044
rect 13916 29262 13918 29314
rect 13970 29262 13972 29314
rect 13916 29250 13972 29262
rect 14476 28868 14532 30156
rect 14140 27972 14196 27982
rect 14140 27878 14196 27916
rect 12572 26852 12964 26908
rect 13692 26852 13860 26908
rect 12572 25620 12628 25630
rect 12572 25526 12628 25564
rect 12796 24834 12852 24846
rect 12796 24782 12798 24834
rect 12850 24782 12852 24834
rect 12796 24500 12852 24782
rect 12796 24434 12852 24444
rect 12908 23940 12964 26852
rect 13244 24948 13300 24958
rect 13244 24722 13300 24892
rect 13244 24670 13246 24722
rect 13298 24670 13300 24722
rect 13244 24658 13300 24670
rect 13468 24164 13524 24174
rect 13468 24050 13524 24108
rect 13468 23998 13470 24050
rect 13522 23998 13524 24050
rect 13468 23986 13524 23998
rect 13804 24052 13860 26852
rect 14028 26066 14084 26078
rect 14028 26014 14030 26066
rect 14082 26014 14084 26066
rect 14028 25284 14084 26014
rect 14476 25732 14532 28812
rect 14700 27188 14756 32396
rect 14812 32450 14868 32462
rect 14812 32398 14814 32450
rect 14866 32398 14868 32450
rect 14812 30996 14868 32398
rect 14812 30902 14868 30940
rect 14812 27188 14868 27198
rect 14700 27186 14868 27188
rect 14700 27134 14814 27186
rect 14866 27134 14868 27186
rect 14700 27132 14868 27134
rect 14700 26908 14756 27132
rect 14812 27122 14868 27132
rect 14588 26852 14756 26908
rect 14588 26402 14644 26852
rect 14588 26350 14590 26402
rect 14642 26350 14644 26402
rect 14588 26338 14644 26350
rect 14476 25676 14644 25732
rect 14476 25506 14532 25518
rect 14476 25454 14478 25506
rect 14530 25454 14532 25506
rect 14476 25284 14532 25454
rect 14028 25282 14532 25284
rect 14028 25230 14030 25282
rect 14082 25230 14532 25282
rect 14028 25228 14532 25230
rect 14028 25218 14084 25228
rect 14476 24948 14532 25228
rect 14476 24882 14532 24892
rect 13916 24610 13972 24622
rect 13916 24558 13918 24610
rect 13970 24558 13972 24610
rect 13916 24164 13972 24558
rect 13916 24098 13972 24108
rect 12796 23884 12964 23940
rect 13580 23938 13636 23950
rect 13580 23886 13582 23938
rect 13634 23886 13636 23938
rect 12572 23716 12628 23726
rect 12124 23268 12180 23278
rect 12124 23154 12180 23212
rect 12124 23102 12126 23154
rect 12178 23102 12180 23154
rect 12124 22820 12180 23102
rect 12124 22754 12180 22764
rect 12572 23154 12628 23660
rect 12572 23102 12574 23154
rect 12626 23102 12628 23154
rect 12572 22484 12628 23102
rect 12572 22418 12628 22428
rect 12796 21812 12852 23884
rect 12908 23716 12964 23726
rect 12908 23622 12964 23660
rect 13580 23716 13636 23886
rect 13804 23938 13860 23996
rect 13804 23886 13806 23938
rect 13858 23886 13860 23938
rect 13804 23874 13860 23886
rect 13580 23650 13636 23660
rect 12124 21810 12852 21812
rect 12124 21758 12798 21810
rect 12850 21758 12852 21810
rect 12124 21756 12852 21758
rect 12124 21586 12180 21756
rect 12796 21746 12852 21756
rect 13132 23042 13188 23054
rect 13132 22990 13134 23042
rect 13186 22990 13188 23042
rect 12124 21534 12126 21586
rect 12178 21534 12180 21586
rect 12124 21522 12180 21534
rect 12572 20020 12628 20030
rect 13020 20020 13076 20030
rect 12628 19964 12852 20020
rect 12572 19926 12628 19964
rect 12796 19346 12852 19964
rect 13020 19926 13076 19964
rect 12796 19294 12798 19346
rect 12850 19294 12852 19346
rect 12796 19282 12852 19294
rect 11900 16882 12068 16884
rect 11900 16830 11902 16882
rect 11954 16830 12068 16882
rect 11900 16828 12068 16830
rect 11900 16818 11956 16828
rect 11452 16718 11454 16770
rect 11506 16718 11508 16770
rect 11452 16706 11508 16718
rect 11564 16658 11620 16670
rect 11564 16606 11566 16658
rect 11618 16606 11620 16658
rect 11564 16212 11620 16606
rect 11564 16146 11620 16156
rect 11172 16044 11396 16100
rect 11116 16006 11172 16044
rect 11340 15540 11396 16044
rect 11788 15988 11844 15998
rect 11116 15316 11172 15326
rect 11004 15260 11116 15316
rect 11116 13636 11172 15260
rect 11340 15314 11396 15484
rect 11340 15262 11342 15314
rect 11394 15262 11396 15314
rect 11340 15250 11396 15262
rect 11676 15986 11844 15988
rect 11676 15934 11790 15986
rect 11842 15934 11844 15986
rect 11676 15932 11844 15934
rect 11452 15204 11508 15214
rect 11452 14868 11508 15148
rect 11676 15148 11732 15932
rect 11788 15922 11844 15932
rect 12012 15314 12068 16828
rect 12012 15262 12014 15314
rect 12066 15262 12068 15314
rect 11676 15092 11844 15148
rect 11340 14812 11508 14868
rect 11228 14196 11284 14206
rect 11228 13858 11284 14140
rect 11228 13806 11230 13858
rect 11282 13806 11284 13858
rect 11228 13794 11284 13806
rect 11116 13570 11172 13580
rect 9548 12898 9604 12908
rect 10108 13020 10388 13076
rect 10556 13132 10948 13188
rect 10108 12962 10164 13020
rect 10108 12910 10110 12962
rect 10162 12910 10164 12962
rect 10108 12898 10164 12910
rect 10444 12964 10500 12974
rect 10444 12870 10500 12908
rect 9436 12852 9492 12862
rect 9436 12758 9492 12796
rect 9996 12852 10052 12862
rect 9884 12738 9940 12750
rect 9884 12686 9886 12738
rect 9938 12686 9940 12738
rect 9884 12628 9940 12686
rect 9324 12572 9940 12628
rect 8092 12460 8372 12516
rect 8092 12178 8148 12460
rect 9548 12290 9604 12302
rect 9548 12238 9550 12290
rect 9602 12238 9604 12290
rect 8092 12126 8094 12178
rect 8146 12126 8148 12178
rect 8092 12114 8148 12126
rect 8988 12178 9044 12190
rect 8988 12126 8990 12178
rect 9042 12126 9044 12178
rect 8540 11956 8596 11966
rect 8092 11732 8148 11742
rect 8092 11618 8148 11676
rect 8092 11566 8094 11618
rect 8146 11566 8148 11618
rect 8092 11554 8148 11566
rect 7868 11442 7924 11452
rect 8316 11396 8372 11406
rect 8316 11302 8372 11340
rect 8540 11394 8596 11900
rect 8652 11508 8708 11518
rect 8652 11414 8708 11452
rect 8540 11342 8542 11394
rect 8594 11342 8596 11394
rect 8540 11330 8596 11342
rect 8764 11284 8820 11294
rect 8764 11190 8820 11228
rect 7756 10098 7812 10108
rect 7084 9090 7140 9100
rect 6860 8766 6862 8818
rect 6914 8766 6916 8818
rect 6860 8754 6916 8766
rect 7420 9044 7476 9054
rect 6748 8194 6804 8204
rect 7196 8260 7252 8270
rect 7084 8146 7140 8158
rect 7084 8094 7086 8146
rect 7138 8094 7140 8146
rect 6524 7588 6580 7598
rect 6524 7494 6580 7532
rect 6412 6692 6468 7420
rect 6636 7476 6692 7486
rect 6636 7382 6692 7420
rect 6748 7476 6804 7486
rect 7084 7476 7140 8094
rect 7196 8146 7252 8204
rect 7420 8258 7476 8988
rect 7420 8206 7422 8258
rect 7474 8206 7476 8258
rect 7420 8194 7476 8206
rect 7868 9042 7924 9054
rect 7868 8990 7870 9042
rect 7922 8990 7924 9042
rect 7196 8094 7198 8146
rect 7250 8094 7252 8146
rect 7196 8082 7252 8094
rect 7868 7812 7924 8990
rect 8204 9044 8260 9054
rect 8204 8950 8260 8988
rect 8428 8370 8484 8382
rect 8428 8318 8430 8370
rect 8482 8318 8484 8370
rect 7868 7746 7924 7756
rect 7980 8258 8036 8270
rect 7980 8206 7982 8258
rect 8034 8206 8036 8258
rect 7196 7700 7252 7710
rect 7196 7606 7252 7644
rect 7756 7588 7812 7598
rect 7532 7476 7588 7486
rect 6748 7474 7588 7476
rect 6748 7422 6750 7474
rect 6802 7422 7534 7474
rect 7586 7422 7588 7474
rect 6748 7420 7588 7422
rect 6748 7410 6804 7420
rect 6524 6692 6580 6702
rect 6412 6690 6580 6692
rect 6412 6638 6526 6690
rect 6578 6638 6580 6690
rect 6412 6636 6580 6638
rect 6412 5124 6468 5134
rect 6412 5030 6468 5068
rect 6524 3556 6580 6636
rect 7308 6468 7364 6478
rect 7308 6374 7364 6412
rect 6636 5908 6692 5918
rect 7420 5908 7476 7420
rect 7532 7410 7588 7420
rect 7756 6580 7812 7532
rect 7980 7362 8036 8206
rect 8428 7700 8484 8318
rect 8428 7634 8484 7644
rect 8428 7476 8484 7486
rect 7980 7310 7982 7362
rect 8034 7310 8036 7362
rect 7980 7298 8036 7310
rect 8316 7364 8372 7374
rect 7980 6692 8036 6702
rect 8316 6692 8372 7308
rect 7980 6690 8372 6692
rect 7980 6638 7982 6690
rect 8034 6638 8318 6690
rect 8370 6638 8372 6690
rect 7980 6636 8372 6638
rect 7980 6626 8036 6636
rect 7756 6514 7812 6524
rect 7532 6132 7588 6142
rect 7532 6038 7588 6076
rect 8092 6132 8148 6142
rect 7644 5908 7700 5918
rect 7420 5852 7588 5908
rect 6636 5122 6692 5852
rect 7420 5684 7476 5694
rect 6636 5070 6638 5122
rect 6690 5070 6692 5122
rect 6636 5058 6692 5070
rect 6860 5682 7476 5684
rect 6860 5630 7422 5682
rect 7474 5630 7476 5682
rect 6860 5628 7476 5630
rect 6636 3556 6692 3566
rect 6524 3554 6692 3556
rect 6524 3502 6638 3554
rect 6690 3502 6692 3554
rect 6524 3500 6692 3502
rect 4956 3332 5124 3388
rect 5852 3332 6244 3388
rect 4956 3266 5012 3276
rect 5852 2996 5908 3332
rect 5852 2930 5908 2940
rect 6412 2996 6468 3006
rect 6636 2996 6692 3500
rect 6860 3554 6916 5628
rect 7420 5618 7476 5628
rect 7420 5236 7476 5246
rect 7196 4676 7252 4686
rect 7196 4338 7252 4620
rect 7196 4286 7198 4338
rect 7250 4286 7252 4338
rect 7196 4274 7252 4286
rect 7420 4338 7476 5180
rect 7532 5122 7588 5852
rect 7532 5070 7534 5122
rect 7586 5070 7588 5122
rect 7532 4900 7588 5070
rect 7532 4834 7588 4844
rect 7420 4286 7422 4338
rect 7474 4286 7476 4338
rect 7420 4274 7476 4286
rect 7644 4116 7700 5852
rect 7756 5906 7812 5918
rect 7756 5854 7758 5906
rect 7810 5854 7812 5906
rect 7756 4564 7812 5854
rect 7980 5908 8036 5918
rect 7980 5814 8036 5852
rect 7756 4498 7812 4508
rect 6860 3502 6862 3554
rect 6914 3502 6916 3554
rect 6860 3490 6916 3502
rect 7308 4060 7700 4116
rect 6972 3442 7028 3454
rect 6972 3390 6974 3442
rect 7026 3390 7028 3442
rect 6412 2994 6692 2996
rect 6412 2942 6414 2994
rect 6466 2942 6692 2994
rect 6412 2940 6692 2942
rect 6748 3332 6804 3342
rect 6412 2930 6468 2940
rect 4172 2830 4174 2882
rect 4226 2830 4228 2882
rect 4172 2818 4228 2830
rect 3388 2718 3390 2770
rect 3442 2718 3444 2770
rect 3388 2706 3444 2718
rect 4476 2380 4740 2390
rect 4532 2324 4580 2380
rect 4636 2324 4684 2380
rect 4476 2314 4740 2324
rect 6748 2100 6804 3276
rect 6860 2996 6916 3006
rect 6972 2996 7028 3390
rect 6860 2994 7028 2996
rect 6860 2942 6862 2994
rect 6914 2942 7028 2994
rect 6860 2940 7028 2942
rect 6860 2930 6916 2940
rect 7308 2548 7364 4060
rect 7420 3780 7476 3790
rect 7420 3686 7476 3724
rect 8092 3556 8148 6076
rect 8204 4676 8260 6636
rect 8316 6626 8372 6636
rect 8428 6244 8484 7420
rect 8316 6188 8484 6244
rect 8540 6580 8596 6590
rect 8316 6130 8372 6188
rect 8316 6078 8318 6130
rect 8370 6078 8372 6130
rect 8316 6066 8372 6078
rect 8204 4610 8260 4620
rect 8316 5124 8372 5134
rect 8540 5124 8596 6524
rect 8876 6020 8932 6030
rect 8372 5122 8596 5124
rect 8372 5070 8542 5122
rect 8594 5070 8596 5122
rect 8372 5068 8596 5070
rect 8204 3556 8260 3566
rect 7532 3554 8260 3556
rect 7532 3502 8206 3554
rect 8258 3502 8260 3554
rect 7532 3500 8260 3502
rect 7532 2770 7588 3500
rect 8204 3490 8260 3500
rect 7532 2718 7534 2770
rect 7586 2718 7588 2770
rect 7532 2706 7588 2718
rect 7756 2772 7812 2782
rect 8316 2772 8372 5068
rect 8540 5058 8596 5068
rect 8652 5682 8708 5694
rect 8652 5630 8654 5682
rect 8706 5630 8708 5682
rect 8428 4452 8484 4462
rect 8652 4452 8708 5630
rect 8876 5236 8932 5964
rect 8876 5170 8932 5180
rect 8988 5010 9044 12126
rect 9324 11732 9380 11742
rect 9548 11732 9604 12238
rect 9380 11676 9604 11732
rect 9324 11506 9380 11676
rect 9324 11454 9326 11506
rect 9378 11454 9380 11506
rect 9324 11442 9380 11454
rect 9884 10948 9940 12572
rect 9996 12738 10052 12796
rect 9996 12686 9998 12738
rect 10050 12686 10052 12738
rect 9996 12178 10052 12686
rect 9996 12126 9998 12178
rect 10050 12126 10052 12178
rect 9996 12114 10052 12126
rect 10220 12066 10276 12078
rect 10220 12014 10222 12066
rect 10274 12014 10276 12066
rect 10220 11284 10276 12014
rect 10220 11218 10276 11228
rect 10556 11060 10612 13132
rect 11340 12962 11396 14812
rect 11340 12910 11342 12962
rect 11394 12910 11396 12962
rect 9660 10892 9940 10948
rect 10220 11004 10612 11060
rect 10668 12404 10724 12414
rect 9548 9940 9604 9950
rect 9548 9846 9604 9884
rect 9100 7812 9156 7822
rect 9100 6468 9156 7756
rect 9100 5122 9156 6412
rect 9324 7700 9380 7710
rect 9324 6578 9380 7644
rect 9548 7700 9604 7710
rect 9660 7700 9716 10892
rect 10220 10612 10276 11004
rect 10668 10948 10724 12348
rect 11340 12404 11396 12910
rect 11340 12338 11396 12348
rect 11452 14642 11508 14654
rect 11452 14590 11454 14642
rect 11506 14590 11508 14642
rect 11340 11508 11396 11518
rect 11340 11414 11396 11452
rect 11452 11396 11508 14590
rect 11564 13634 11620 13646
rect 11564 13582 11566 13634
rect 11618 13582 11620 13634
rect 11564 12292 11620 13582
rect 11676 13524 11732 13534
rect 11676 13074 11732 13468
rect 11676 13022 11678 13074
rect 11730 13022 11732 13074
rect 11676 13010 11732 13022
rect 11788 12628 11844 15092
rect 11900 15092 11956 15102
rect 11900 14998 11956 15036
rect 11900 14530 11956 14542
rect 11900 14478 11902 14530
rect 11954 14478 11956 14530
rect 11900 13634 11956 14478
rect 12012 14532 12068 15262
rect 12012 14466 12068 14476
rect 12460 18452 12516 18462
rect 12460 14308 12516 18396
rect 12796 16772 12852 16782
rect 12572 15540 12628 15550
rect 12572 14754 12628 15484
rect 12796 15538 12852 16716
rect 12796 15486 12798 15538
rect 12850 15486 12852 15538
rect 12796 15316 12852 15486
rect 12796 15250 12852 15260
rect 12572 14702 12574 14754
rect 12626 14702 12628 14754
rect 12572 14690 12628 14702
rect 13020 15092 13076 15102
rect 12796 14532 12852 14542
rect 12796 14418 12852 14476
rect 12796 14366 12798 14418
rect 12850 14366 12852 14418
rect 12796 14354 12852 14366
rect 12684 14308 12740 14318
rect 12460 14242 12516 14252
rect 12572 14306 12740 14308
rect 12572 14254 12686 14306
rect 12738 14254 12740 14306
rect 12572 14252 12740 14254
rect 11900 13582 11902 13634
rect 11954 13582 11956 13634
rect 11900 13524 11956 13582
rect 11900 13458 11956 13468
rect 12236 13860 12292 13870
rect 12236 12964 12292 13804
rect 12572 13746 12628 14252
rect 12684 14242 12740 14252
rect 13020 13970 13076 15036
rect 13020 13918 13022 13970
rect 13074 13918 13076 13970
rect 13020 13906 13076 13918
rect 12572 13694 12574 13746
rect 12626 13694 12628 13746
rect 12460 13188 12516 13198
rect 12572 13188 12628 13694
rect 12908 13746 12964 13758
rect 12908 13694 12910 13746
rect 12962 13694 12964 13746
rect 12908 13524 12964 13694
rect 12908 13458 12964 13468
rect 13020 13522 13076 13534
rect 13020 13470 13022 13522
rect 13074 13470 13076 13522
rect 12460 13186 12628 13188
rect 12460 13134 12462 13186
rect 12514 13134 12628 13186
rect 12460 13132 12628 13134
rect 12460 13122 12516 13132
rect 12236 12962 12964 12964
rect 12236 12910 12238 12962
rect 12290 12910 12964 12962
rect 12236 12908 12964 12910
rect 12236 12898 12292 12908
rect 11788 12562 11844 12572
rect 11900 12850 11956 12862
rect 11900 12798 11902 12850
rect 11954 12798 11956 12850
rect 11564 12178 11620 12236
rect 11564 12126 11566 12178
rect 11618 12126 11620 12178
rect 11564 12114 11620 12126
rect 11676 12066 11732 12078
rect 11676 12014 11678 12066
rect 11730 12014 11732 12066
rect 11564 11956 11620 11966
rect 11676 11956 11732 12014
rect 11620 11900 11732 11956
rect 11564 11890 11620 11900
rect 11900 11732 11956 12798
rect 12796 12738 12852 12750
rect 12796 12686 12798 12738
rect 12850 12686 12852 12738
rect 12236 12628 12292 12638
rect 12124 12516 12180 12526
rect 12012 12066 12068 12078
rect 12012 12014 12014 12066
rect 12066 12014 12068 12066
rect 12012 11844 12068 12014
rect 12012 11778 12068 11788
rect 11900 11666 11956 11676
rect 12124 11508 12180 12460
rect 11900 11452 12180 11508
rect 11452 11394 11732 11396
rect 11452 11342 11454 11394
rect 11506 11342 11732 11394
rect 11452 11340 11732 11342
rect 11452 11330 11508 11340
rect 10892 11284 10948 11294
rect 10780 11170 10836 11182
rect 10780 11118 10782 11170
rect 10834 11118 10836 11170
rect 10780 10948 10836 11118
rect 10332 10892 10836 10948
rect 10332 10834 10388 10892
rect 10332 10782 10334 10834
rect 10386 10782 10388 10834
rect 10332 10770 10388 10782
rect 10668 10724 10724 10734
rect 10220 10556 10388 10612
rect 10332 9940 10388 10556
rect 10220 9884 10388 9940
rect 10108 9826 10164 9838
rect 10108 9774 10110 9826
rect 10162 9774 10164 9826
rect 10108 9604 10164 9774
rect 10108 9538 10164 9548
rect 10108 9156 10164 9166
rect 9772 8258 9828 8270
rect 9772 8206 9774 8258
rect 9826 8206 9828 8258
rect 9772 7812 9828 8206
rect 9772 7746 9828 7756
rect 9548 7698 9716 7700
rect 9548 7646 9550 7698
rect 9602 7646 9716 7698
rect 9548 7644 9716 7646
rect 9548 7634 9604 7644
rect 9772 7586 9828 7598
rect 9772 7534 9774 7586
rect 9826 7534 9828 7586
rect 9772 6916 9828 7534
rect 9884 7588 9940 7598
rect 9884 7494 9940 7532
rect 9772 6860 10052 6916
rect 9996 6692 10052 6860
rect 9996 6626 10052 6636
rect 10108 6804 10164 9100
rect 10220 7364 10276 9884
rect 10556 9826 10612 9838
rect 10556 9774 10558 9826
rect 10610 9774 10612 9826
rect 10444 9602 10500 9614
rect 10444 9550 10446 9602
rect 10498 9550 10500 9602
rect 10444 9042 10500 9550
rect 10444 8990 10446 9042
rect 10498 8990 10500 9042
rect 10444 7700 10500 8990
rect 10556 8932 10612 9774
rect 10556 8866 10612 8876
rect 10668 8482 10724 10668
rect 10780 10610 10836 10892
rect 10780 10558 10782 10610
rect 10834 10558 10836 10610
rect 10780 9604 10836 10558
rect 10780 9538 10836 9548
rect 10668 8430 10670 8482
rect 10722 8430 10724 8482
rect 10668 8418 10724 8430
rect 10892 8258 10948 11228
rect 11228 11282 11284 11294
rect 11228 11230 11230 11282
rect 11282 11230 11284 11282
rect 11228 10386 11284 11230
rect 11228 10334 11230 10386
rect 11282 10334 11284 10386
rect 11228 9828 11284 10334
rect 11564 9828 11620 9838
rect 11228 9772 11564 9828
rect 11004 9044 11060 9054
rect 11004 8950 11060 8988
rect 10892 8206 10894 8258
rect 10946 8206 10948 8258
rect 10892 8194 10948 8206
rect 11452 8930 11508 8942
rect 11452 8878 11454 8930
rect 11506 8878 11508 8930
rect 11452 7924 11508 8878
rect 10444 7634 10500 7644
rect 11340 7868 11508 7924
rect 11340 7588 11396 7868
rect 11564 7588 11620 9772
rect 11676 9716 11732 11340
rect 11900 10164 11956 11452
rect 12236 11394 12292 12572
rect 12572 12292 12628 12302
rect 12460 12236 12572 12292
rect 12236 11342 12238 11394
rect 12290 11342 12292 11394
rect 12236 11330 12292 11342
rect 12348 11732 12404 11742
rect 12124 10610 12180 10622
rect 12124 10558 12126 10610
rect 12178 10558 12180 10610
rect 11900 10108 12068 10164
rect 11900 9940 11956 9950
rect 11900 9826 11956 9884
rect 11900 9774 11902 9826
rect 11954 9774 11956 9826
rect 11900 9762 11956 9774
rect 11676 9660 11844 9716
rect 11676 8932 11732 8942
rect 11676 8370 11732 8876
rect 11676 8318 11678 8370
rect 11730 8318 11732 8370
rect 11676 8306 11732 8318
rect 11676 7588 11732 7598
rect 11564 7586 11732 7588
rect 11564 7534 11678 7586
rect 11730 7534 11732 7586
rect 11564 7532 11732 7534
rect 10220 7298 10276 7308
rect 10332 7474 10388 7486
rect 10332 7422 10334 7474
rect 10386 7422 10388 7474
rect 9324 6526 9326 6578
rect 9378 6526 9380 6578
rect 9324 5908 9380 6526
rect 9548 6580 9604 6590
rect 9548 6486 9604 6524
rect 9324 5842 9380 5852
rect 9436 6466 9492 6478
rect 9436 6414 9438 6466
rect 9490 6414 9492 6466
rect 9100 5070 9102 5122
rect 9154 5070 9156 5122
rect 9100 5058 9156 5070
rect 9436 5124 9492 6414
rect 9884 5908 9940 5918
rect 9884 5814 9940 5852
rect 10108 5906 10164 6748
rect 10220 6802 10276 6814
rect 10220 6750 10222 6802
rect 10274 6750 10276 6802
rect 10220 6020 10276 6750
rect 10220 5954 10276 5964
rect 10108 5854 10110 5906
rect 10162 5854 10164 5906
rect 10108 5842 10164 5854
rect 10332 5348 10388 7422
rect 10668 7474 10724 7486
rect 10668 7422 10670 7474
rect 10722 7422 10724 7474
rect 10668 5908 10724 7422
rect 10892 7476 10948 7486
rect 10892 7474 11172 7476
rect 10892 7422 10894 7474
rect 10946 7422 11172 7474
rect 10892 7420 11172 7422
rect 10892 7410 10948 7420
rect 10780 7362 10836 7374
rect 10780 7310 10782 7362
rect 10834 7310 10836 7362
rect 10780 6132 10836 7310
rect 10892 6692 10948 6702
rect 10892 6598 10948 6636
rect 10780 6076 11060 6132
rect 10780 5908 10836 5918
rect 10668 5906 10836 5908
rect 10668 5854 10782 5906
rect 10834 5854 10836 5906
rect 10668 5852 10836 5854
rect 10444 5684 10500 5694
rect 10444 5682 10612 5684
rect 10444 5630 10446 5682
rect 10498 5630 10612 5682
rect 10444 5628 10612 5630
rect 10444 5618 10500 5628
rect 10332 5282 10388 5292
rect 9436 5068 10164 5124
rect 8988 4958 8990 5010
rect 9042 4958 9044 5010
rect 8988 4946 9044 4958
rect 8428 4450 8708 4452
rect 8428 4398 8430 4450
rect 8482 4398 8708 4450
rect 8428 4396 8708 4398
rect 8764 4900 8820 4910
rect 8428 3780 8484 4396
rect 8428 3714 8484 3724
rect 8764 3666 8820 4844
rect 9660 4676 9716 4686
rect 8876 4564 8932 4574
rect 8876 4116 8932 4508
rect 9660 4562 9716 4620
rect 9660 4510 9662 4562
rect 9714 4510 9716 4562
rect 9660 4498 9716 4510
rect 8876 4050 8932 4060
rect 8764 3614 8766 3666
rect 8818 3614 8820 3666
rect 8764 3602 8820 3614
rect 7756 2770 8372 2772
rect 7756 2718 7758 2770
rect 7810 2718 8372 2770
rect 7756 2716 8372 2718
rect 10108 2770 10164 5068
rect 10332 5012 10388 5022
rect 10332 4918 10388 4956
rect 10332 4564 10388 4574
rect 10332 4470 10388 4508
rect 10444 4452 10500 4462
rect 10444 4358 10500 4396
rect 10556 4340 10612 5628
rect 10668 4564 10724 5852
rect 10780 5842 10836 5852
rect 10892 5908 10948 5918
rect 10668 4498 10724 4508
rect 10780 4340 10836 4350
rect 10556 4338 10836 4340
rect 10556 4286 10782 4338
rect 10834 4286 10836 4338
rect 10556 4284 10836 4286
rect 10780 4274 10836 4284
rect 10332 4114 10388 4126
rect 10332 4062 10334 4114
rect 10386 4062 10388 4114
rect 10332 3388 10388 4062
rect 10444 4116 10500 4126
rect 10892 4116 10948 5852
rect 11004 4562 11060 6076
rect 11116 5796 11172 7420
rect 11340 6690 11396 7532
rect 11676 7252 11732 7532
rect 11788 7474 11844 9660
rect 12012 9042 12068 10108
rect 12124 9716 12180 10558
rect 12124 9650 12180 9660
rect 12012 8990 12014 9042
rect 12066 8990 12068 9042
rect 12012 8484 12068 8990
rect 12348 9042 12404 11676
rect 12460 9826 12516 12236
rect 12572 12198 12628 12236
rect 12572 11508 12628 11518
rect 12628 11452 12740 11508
rect 12572 11442 12628 11452
rect 12460 9774 12462 9826
rect 12514 9774 12516 9826
rect 12460 9762 12516 9774
rect 12572 10612 12628 10622
rect 12572 9714 12628 10556
rect 12572 9662 12574 9714
rect 12626 9662 12628 9714
rect 12572 9650 12628 9662
rect 12348 8990 12350 9042
rect 12402 8990 12404 9042
rect 12348 8978 12404 8990
rect 12684 9042 12740 11452
rect 12796 9716 12852 12686
rect 12908 12178 12964 12908
rect 12908 12126 12910 12178
rect 12962 12126 12964 12178
rect 12908 11508 12964 12126
rect 12908 11170 12964 11452
rect 12908 11118 12910 11170
rect 12962 11118 12964 11170
rect 12908 9940 12964 11118
rect 12908 9874 12964 9884
rect 12796 9650 12852 9660
rect 12684 8990 12686 9042
rect 12738 8990 12740 9042
rect 12684 8978 12740 8990
rect 12012 8418 12068 8428
rect 12908 8484 12964 8494
rect 12908 8372 12964 8428
rect 11788 7422 11790 7474
rect 11842 7422 11844 7474
rect 11788 7410 11844 7422
rect 12684 8370 12964 8372
rect 12684 8318 12910 8370
rect 12962 8318 12964 8370
rect 12684 8316 12964 8318
rect 12684 7476 12740 8316
rect 12908 8306 12964 8316
rect 12460 7362 12516 7374
rect 12460 7310 12462 7362
rect 12514 7310 12516 7362
rect 11676 7196 11844 7252
rect 11340 6638 11342 6690
rect 11394 6638 11396 6690
rect 11340 6626 11396 6638
rect 11788 6356 11844 7196
rect 12236 6804 12292 6814
rect 12236 6690 12292 6748
rect 12236 6638 12238 6690
rect 12290 6638 12292 6690
rect 12236 6626 12292 6638
rect 11788 6290 11844 6300
rect 11116 5730 11172 5740
rect 11228 6132 11284 6142
rect 12460 6132 12516 7310
rect 12684 6804 12740 7420
rect 11228 6018 11284 6076
rect 11228 5966 11230 6018
rect 11282 5966 11284 6018
rect 11228 5122 11284 5966
rect 11228 5070 11230 5122
rect 11282 5070 11284 5122
rect 11228 5058 11284 5070
rect 12124 6076 12516 6132
rect 12012 4898 12068 4910
rect 12012 4846 12014 4898
rect 12066 4846 12068 4898
rect 11004 4510 11006 4562
rect 11058 4510 11060 4562
rect 11004 4498 11060 4510
rect 11116 4562 11172 4574
rect 11116 4510 11118 4562
rect 11170 4510 11172 4562
rect 10444 3554 10500 4060
rect 10444 3502 10446 3554
rect 10498 3502 10500 3554
rect 10444 3490 10500 3502
rect 10668 4060 10948 4116
rect 10332 3332 10612 3388
rect 10108 2718 10110 2770
rect 10162 2718 10164 2770
rect 7756 2706 7812 2716
rect 10108 2706 10164 2718
rect 10556 2770 10612 3332
rect 10556 2718 10558 2770
rect 10610 2718 10612 2770
rect 10556 2706 10612 2718
rect 10332 2658 10388 2670
rect 10332 2606 10334 2658
rect 10386 2606 10388 2658
rect 7308 2454 7364 2492
rect 10108 2548 10164 2558
rect 10332 2548 10388 2606
rect 10668 2548 10724 4060
rect 10892 3668 10948 3678
rect 11116 3668 11172 4510
rect 11788 4564 11844 4574
rect 12012 4564 12068 4846
rect 11844 4508 12068 4564
rect 11788 4450 11844 4508
rect 11788 4398 11790 4450
rect 11842 4398 11844 4450
rect 11788 4386 11844 4398
rect 11340 3780 11396 3790
rect 11340 3686 11396 3724
rect 10892 3666 11172 3668
rect 10892 3614 10894 3666
rect 10946 3614 11172 3666
rect 10892 3612 11172 3614
rect 10892 3602 10948 3612
rect 11900 3554 11956 3566
rect 11900 3502 11902 3554
rect 11954 3502 11956 3554
rect 11900 3332 11956 3502
rect 12012 3554 12068 4508
rect 12124 4452 12180 6076
rect 12460 6020 12516 6076
rect 12460 5954 12516 5964
rect 12572 6468 12628 6478
rect 12124 4338 12180 4396
rect 12124 4286 12126 4338
rect 12178 4286 12180 4338
rect 12124 4274 12180 4286
rect 12236 5906 12292 5918
rect 12236 5854 12238 5906
rect 12290 5854 12292 5906
rect 12236 5124 12292 5854
rect 12460 5348 12516 5358
rect 12236 3666 12292 5068
rect 12348 5236 12404 5246
rect 12348 5122 12404 5180
rect 12348 5070 12350 5122
rect 12402 5070 12404 5122
rect 12348 5058 12404 5070
rect 12236 3614 12238 3666
rect 12290 3614 12292 3666
rect 12236 3602 12292 3614
rect 12460 4564 12516 5292
rect 12572 5122 12628 6412
rect 12572 5070 12574 5122
rect 12626 5070 12628 5122
rect 12572 5058 12628 5070
rect 12572 4564 12628 4574
rect 12460 4562 12628 4564
rect 12460 4510 12574 4562
rect 12626 4510 12628 4562
rect 12460 4508 12628 4510
rect 12012 3502 12014 3554
rect 12066 3502 12068 3554
rect 12012 3490 12068 3502
rect 12460 3388 12516 4508
rect 12572 4498 12628 4508
rect 12684 4452 12740 6748
rect 13020 6580 13076 13470
rect 13132 12516 13188 22990
rect 14476 23042 14532 23054
rect 14476 22990 14478 23042
rect 14530 22990 14532 23042
rect 13692 21476 13748 21486
rect 13468 21140 13524 21150
rect 13468 20802 13524 21084
rect 13692 21026 13748 21420
rect 14252 21476 14308 21486
rect 14252 21382 14308 21420
rect 14476 21476 14532 22990
rect 14476 21410 14532 21420
rect 13692 20974 13694 21026
rect 13746 20974 13748 21026
rect 13692 20962 13748 20974
rect 14588 21028 14644 25676
rect 14700 24052 14756 24062
rect 14700 23940 14756 23996
rect 14812 23940 14868 23950
rect 14700 23938 14868 23940
rect 14700 23886 14814 23938
rect 14866 23886 14868 23938
rect 14700 23884 14868 23886
rect 14812 23874 14868 23884
rect 14700 23380 14756 23390
rect 14700 22930 14756 23324
rect 14700 22878 14702 22930
rect 14754 22878 14756 22930
rect 14700 21588 14756 22878
rect 14700 21522 14756 21532
rect 14588 20972 14756 21028
rect 13468 20750 13470 20802
rect 13522 20750 13524 20802
rect 13468 20580 13524 20750
rect 14028 20804 14084 20814
rect 14588 20804 14644 20814
rect 14028 20802 14644 20804
rect 14028 20750 14030 20802
rect 14082 20750 14590 20802
rect 14642 20750 14644 20802
rect 14028 20748 14644 20750
rect 14028 20738 14084 20748
rect 14588 20738 14644 20748
rect 14364 20580 14420 20590
rect 13468 20514 13524 20524
rect 13692 20578 14420 20580
rect 13692 20526 14366 20578
rect 14418 20526 14420 20578
rect 13692 20524 14420 20526
rect 13692 20130 13748 20524
rect 14364 20514 14420 20524
rect 13692 20078 13694 20130
rect 13746 20078 13748 20130
rect 13692 20066 13748 20078
rect 14588 18452 14644 18462
rect 14700 18452 14756 20972
rect 14644 18396 14756 18452
rect 14812 18676 14868 18686
rect 14588 18386 14644 18396
rect 13580 17444 13636 17454
rect 13580 16098 13636 17388
rect 14700 17444 14756 17454
rect 14700 17350 14756 17388
rect 14476 16994 14532 17006
rect 14476 16942 14478 16994
rect 14530 16942 14532 16994
rect 13580 16046 13582 16098
rect 13634 16046 13636 16098
rect 13580 15148 13636 16046
rect 14140 16884 14196 16894
rect 13580 15092 13972 15148
rect 13468 14532 13524 14542
rect 13468 13858 13524 14476
rect 13468 13806 13470 13858
rect 13522 13806 13524 13858
rect 13468 13794 13524 13806
rect 13580 14306 13636 14318
rect 13580 14254 13582 14306
rect 13634 14254 13636 14306
rect 13580 13860 13636 14254
rect 13580 13794 13636 13804
rect 13916 13746 13972 15092
rect 13916 13694 13918 13746
rect 13970 13694 13972 13746
rect 13580 13522 13636 13534
rect 13580 13470 13582 13522
rect 13634 13470 13636 13522
rect 13580 12516 13636 13470
rect 13916 13524 13972 13694
rect 13916 13458 13972 13468
rect 14028 14644 14084 14654
rect 14028 13076 14084 14588
rect 14140 13860 14196 16828
rect 14252 16212 14308 16222
rect 14476 16212 14532 16942
rect 14812 16994 14868 18620
rect 14812 16942 14814 16994
rect 14866 16942 14868 16994
rect 14812 16930 14868 16942
rect 14252 16210 14532 16212
rect 14252 16158 14254 16210
rect 14306 16158 14532 16210
rect 14252 16156 14532 16158
rect 14252 16146 14308 16156
rect 14924 14644 14980 40236
rect 15260 38724 15316 40348
rect 15372 40338 15428 40348
rect 15372 39508 15428 39518
rect 15372 39058 15428 39452
rect 15372 39006 15374 39058
rect 15426 39006 15428 39058
rect 15372 38994 15428 39006
rect 15036 38668 15316 38724
rect 15708 38834 15764 38846
rect 15708 38782 15710 38834
rect 15762 38782 15764 38834
rect 15708 38668 15764 38782
rect 15036 37156 15092 38668
rect 15708 38612 15988 38668
rect 15932 38610 15988 38612
rect 15932 38558 15934 38610
rect 15986 38558 15988 38610
rect 15932 38546 15988 38558
rect 15372 38052 15428 38062
rect 15372 37958 15428 37996
rect 15036 37090 15092 37100
rect 16044 36708 16100 43596
rect 16492 43428 16548 44942
rect 16604 44434 16660 45724
rect 16604 44382 16606 44434
rect 16658 44382 16660 44434
rect 16604 44370 16660 44382
rect 16604 43428 16660 43438
rect 16492 43372 16604 43428
rect 16604 43362 16660 43372
rect 16156 42866 16212 42878
rect 16156 42814 16158 42866
rect 16210 42814 16212 42866
rect 16156 42532 16212 42814
rect 16156 42466 16212 42476
rect 16604 42196 16660 42206
rect 16716 42196 16772 46620
rect 16828 46610 16884 46620
rect 17500 46452 17556 46462
rect 16828 46450 17556 46452
rect 16828 46398 17502 46450
rect 17554 46398 17556 46450
rect 16828 46396 17556 46398
rect 16828 46002 16884 46396
rect 17500 46386 17556 46396
rect 16828 45950 16830 46002
rect 16882 45950 16884 46002
rect 16828 45938 16884 45950
rect 17052 45668 17108 45678
rect 17052 44098 17108 45612
rect 17052 44046 17054 44098
rect 17106 44046 17108 44098
rect 17052 43764 17108 44046
rect 17500 44100 17556 44110
rect 17500 44006 17556 44044
rect 17052 43698 17108 43708
rect 16828 43426 16884 43438
rect 16828 43374 16830 43426
rect 16882 43374 16884 43426
rect 16828 42644 16884 43374
rect 17612 43428 17668 43438
rect 17612 42866 17668 43372
rect 17612 42814 17614 42866
rect 17666 42814 17668 42866
rect 17612 42802 17668 42814
rect 16828 42578 16884 42588
rect 17500 42644 17556 42654
rect 16604 42194 16772 42196
rect 16604 42142 16606 42194
rect 16658 42142 16772 42194
rect 16604 42140 16772 42142
rect 17164 42530 17220 42542
rect 17164 42478 17166 42530
rect 17218 42478 17220 42530
rect 16604 42130 16660 42140
rect 16156 41972 16212 41982
rect 16156 40404 16212 41916
rect 16492 41858 16548 41870
rect 16492 41806 16494 41858
rect 16546 41806 16548 41858
rect 16492 40516 16548 41806
rect 17164 41860 17220 42478
rect 17500 42082 17556 42588
rect 17500 42030 17502 42082
rect 17554 42030 17556 42082
rect 17500 42018 17556 42030
rect 17724 41972 17780 50428
rect 18060 48132 18116 48142
rect 18060 47236 18116 48076
rect 18060 47170 18116 47180
rect 18284 46562 18340 53564
rect 18732 50596 18788 50606
rect 18732 50502 18788 50540
rect 18956 49364 19012 53676
rect 19068 53620 19124 56588
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 19516 55298 19572 55310
rect 19516 55246 19518 55298
rect 19570 55246 19572 55298
rect 19516 54738 19572 55246
rect 20188 55300 20244 62076
rect 20412 61012 20468 62860
rect 20412 60946 20468 60956
rect 20300 58324 20356 58334
rect 20300 58230 20356 58268
rect 20524 57988 20580 67676
rect 21420 67666 21476 67676
rect 22316 66500 22372 69246
rect 23100 68852 23156 69358
rect 23324 68852 23380 68862
rect 23100 68796 23324 68852
rect 22428 68740 22484 68750
rect 22428 68626 22484 68684
rect 22428 68574 22430 68626
rect 22482 68574 22484 68626
rect 22428 67620 22484 68574
rect 23100 68628 23156 68638
rect 23100 68534 23156 68572
rect 22988 68404 23044 68414
rect 22428 67554 22484 67564
rect 22876 67620 22932 67630
rect 22876 67526 22932 67564
rect 22316 66444 22596 66500
rect 21756 66276 21812 66286
rect 20860 66274 21812 66276
rect 20860 66222 21758 66274
rect 21810 66222 21812 66274
rect 20860 66220 21812 66222
rect 20860 65378 20916 66220
rect 21756 66210 21812 66220
rect 22316 66274 22372 66286
rect 22316 66222 22318 66274
rect 22370 66222 22372 66274
rect 21420 66052 21476 66062
rect 21308 65996 21420 66052
rect 20860 65326 20862 65378
rect 20914 65326 20916 65378
rect 20860 65314 20916 65326
rect 21196 65492 21252 65502
rect 21308 65492 21364 65996
rect 21420 65958 21476 65996
rect 21868 66050 21924 66062
rect 21868 65998 21870 66050
rect 21922 65998 21924 66050
rect 21196 65490 21364 65492
rect 21196 65438 21198 65490
rect 21250 65438 21364 65490
rect 21196 65436 21364 65438
rect 20748 64484 20804 64494
rect 21196 64484 21252 65436
rect 21420 65380 21476 65390
rect 21420 64930 21476 65324
rect 21420 64878 21422 64930
rect 21474 64878 21476 64930
rect 21420 64866 21476 64878
rect 21756 64594 21812 64606
rect 21756 64542 21758 64594
rect 21810 64542 21812 64594
rect 20748 64482 21252 64484
rect 20748 64430 20750 64482
rect 20802 64430 21252 64482
rect 20748 64428 21252 64430
rect 21532 64482 21588 64494
rect 21532 64430 21534 64482
rect 21586 64430 21588 64482
rect 20748 62916 20804 64428
rect 21532 63924 21588 64430
rect 21756 64148 21812 64542
rect 21868 64484 21924 65998
rect 22316 66052 22372 66222
rect 22316 65986 22372 65996
rect 21980 65378 22036 65390
rect 21980 65326 21982 65378
rect 22034 65326 22036 65378
rect 21980 64932 22036 65326
rect 22092 64932 22148 64942
rect 21980 64930 22148 64932
rect 21980 64878 22094 64930
rect 22146 64878 22148 64930
rect 21980 64876 22148 64878
rect 22092 64866 22148 64876
rect 22428 64594 22484 64606
rect 22428 64542 22430 64594
rect 22482 64542 22484 64594
rect 22204 64484 22260 64494
rect 21868 64482 22260 64484
rect 21868 64430 22206 64482
rect 22258 64430 22260 64482
rect 21868 64428 22260 64430
rect 21980 64148 22036 64158
rect 21756 64092 21980 64148
rect 21980 64054 22036 64092
rect 21532 63858 21588 63868
rect 22092 63924 22148 63934
rect 20748 62850 20804 62860
rect 20748 61684 20804 61694
rect 21644 61684 21700 61694
rect 20748 61682 21700 61684
rect 20748 61630 20750 61682
rect 20802 61630 21646 61682
rect 21698 61630 21700 61682
rect 20748 61628 21700 61630
rect 20748 61618 20804 61628
rect 21644 61618 21700 61628
rect 20972 61348 21028 61358
rect 21756 61348 21812 61358
rect 20636 61012 20692 61022
rect 20972 61012 21028 61292
rect 20692 60956 21028 61012
rect 20636 60918 20692 60956
rect 20972 60786 21028 60956
rect 20972 60734 20974 60786
rect 21026 60734 21028 60786
rect 20972 60722 21028 60734
rect 21644 61346 21812 61348
rect 21644 61294 21758 61346
rect 21810 61294 21812 61346
rect 21644 61292 21812 61294
rect 21644 60116 21700 61292
rect 21756 61282 21812 61292
rect 21756 60674 21812 60686
rect 21756 60622 21758 60674
rect 21810 60622 21812 60674
rect 21756 60340 21812 60622
rect 21756 60284 22036 60340
rect 21644 60060 21812 60116
rect 21420 60004 21476 60014
rect 20524 57932 21140 57988
rect 20860 57762 20916 57774
rect 20860 57710 20862 57762
rect 20914 57710 20916 57762
rect 20300 57650 20356 57662
rect 20300 57598 20302 57650
rect 20354 57598 20356 57650
rect 20300 56866 20356 57598
rect 20300 56814 20302 56866
rect 20354 56814 20356 56866
rect 20300 55300 20356 56814
rect 20636 55300 20692 55310
rect 20300 55298 20692 55300
rect 20300 55246 20638 55298
rect 20690 55246 20692 55298
rect 20300 55244 20692 55246
rect 20188 55206 20244 55244
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19516 54686 19518 54738
rect 19570 54686 19572 54738
rect 19516 54674 19572 54686
rect 19628 54740 19684 54750
rect 19684 54684 20020 54740
rect 19628 54646 19684 54684
rect 19180 54572 19460 54628
rect 19180 53844 19236 54572
rect 19404 54516 19460 54572
rect 19852 54516 19908 54526
rect 19404 54514 19908 54516
rect 19404 54462 19854 54514
rect 19906 54462 19908 54514
rect 19404 54460 19908 54462
rect 19852 54450 19908 54460
rect 19292 54404 19348 54414
rect 19292 54402 19572 54404
rect 19292 54350 19294 54402
rect 19346 54350 19572 54402
rect 19292 54348 19572 54350
rect 19292 54338 19348 54348
rect 19516 54292 19572 54348
rect 19180 53842 19460 53844
rect 19180 53790 19182 53842
rect 19234 53790 19460 53842
rect 19180 53788 19460 53790
rect 19180 53778 19236 53788
rect 19068 53564 19348 53620
rect 19068 52836 19124 52846
rect 19068 52834 19236 52836
rect 19068 52782 19070 52834
rect 19122 52782 19236 52834
rect 19068 52780 19236 52782
rect 19068 52770 19124 52780
rect 18956 49298 19012 49308
rect 19180 52724 19236 52780
rect 18396 49140 18452 49150
rect 18732 49140 18788 49150
rect 18396 49138 18788 49140
rect 18396 49086 18398 49138
rect 18450 49086 18734 49138
rect 18786 49086 18788 49138
rect 18396 49084 18788 49086
rect 18396 49074 18452 49084
rect 18732 49074 18788 49084
rect 18732 48916 18788 48926
rect 18732 48356 18788 48860
rect 18844 48804 18900 48814
rect 18844 48710 18900 48748
rect 18844 48356 18900 48366
rect 18732 48354 18900 48356
rect 18732 48302 18846 48354
rect 18898 48302 18900 48354
rect 18732 48300 18900 48302
rect 18844 48290 18900 48300
rect 18620 48244 18676 48254
rect 18620 48150 18676 48188
rect 18956 48242 19012 48254
rect 18956 48190 18958 48242
rect 19010 48190 19012 48242
rect 18508 47236 18564 47246
rect 18844 47236 18900 47246
rect 18508 47234 18844 47236
rect 18508 47182 18510 47234
rect 18562 47182 18844 47234
rect 18508 47180 18844 47182
rect 18508 47170 18564 47180
rect 18844 47170 18900 47180
rect 18284 46510 18286 46562
rect 18338 46510 18340 46562
rect 17836 46452 17892 46462
rect 18284 46452 18340 46510
rect 18844 46564 18900 46574
rect 18956 46564 19012 48190
rect 18900 46508 19012 46564
rect 18844 46470 18900 46508
rect 17836 46450 18340 46452
rect 17836 46398 17838 46450
rect 17890 46398 18340 46450
rect 17836 46396 18340 46398
rect 17836 46386 17892 46396
rect 17836 43764 17892 43774
rect 17836 43670 17892 43708
rect 17724 41878 17780 41916
rect 17164 41794 17220 41804
rect 17948 41298 18004 46396
rect 19180 46228 19236 52668
rect 19292 49922 19348 53564
rect 19404 52946 19460 53788
rect 19404 52894 19406 52946
rect 19458 52894 19460 52946
rect 19404 52882 19460 52894
rect 19516 51380 19572 54236
rect 19964 53508 20020 54684
rect 20076 54514 20132 54526
rect 20076 54462 20078 54514
rect 20130 54462 20132 54514
rect 20076 53732 20132 54462
rect 20524 54514 20580 54526
rect 20524 54462 20526 54514
rect 20578 54462 20580 54514
rect 20524 54292 20580 54462
rect 20524 54226 20580 54236
rect 20636 53844 20692 55244
rect 20748 55188 20804 55198
rect 20748 55094 20804 55132
rect 20636 53778 20692 53788
rect 20076 53666 20132 53676
rect 20300 53508 20356 53518
rect 19964 53506 20468 53508
rect 19964 53454 20302 53506
rect 20354 53454 20468 53506
rect 19964 53452 20468 53454
rect 20300 53442 20356 53452
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 20412 53060 20468 53452
rect 20524 53060 20580 53070
rect 20412 53004 20524 53060
rect 20524 52994 20580 53004
rect 20636 53058 20692 53070
rect 20636 53006 20638 53058
rect 20690 53006 20692 53058
rect 19964 52948 20020 52958
rect 20300 52948 20356 52958
rect 19964 52946 20356 52948
rect 19964 52894 19966 52946
rect 20018 52894 20302 52946
rect 20354 52894 20356 52946
rect 19964 52892 20356 52894
rect 19964 52882 20020 52892
rect 20300 52882 20356 52892
rect 19628 52724 19684 52734
rect 19628 52630 19684 52668
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 20636 51490 20692 53006
rect 20636 51438 20638 51490
rect 20690 51438 20692 51490
rect 20636 51426 20692 51438
rect 19852 51380 19908 51390
rect 19516 51378 19908 51380
rect 19516 51326 19518 51378
rect 19570 51326 19854 51378
rect 19906 51326 19908 51378
rect 19516 51324 19908 51326
rect 19516 51314 19572 51324
rect 19852 50596 19908 51324
rect 19852 50530 19908 50540
rect 20860 50428 20916 57710
rect 20972 55970 21028 55982
rect 20972 55918 20974 55970
rect 21026 55918 21028 55970
rect 20972 55858 21028 55918
rect 20972 55806 20974 55858
rect 21026 55806 21028 55858
rect 20972 55794 21028 55806
rect 21084 50428 21140 57932
rect 21308 56754 21364 56766
rect 21308 56702 21310 56754
rect 21362 56702 21364 56754
rect 21308 56644 21364 56702
rect 21308 56578 21364 56588
rect 21420 55860 21476 59948
rect 21644 59890 21700 59902
rect 21644 59838 21646 59890
rect 21698 59838 21700 59890
rect 21644 59444 21700 59838
rect 21756 59780 21812 60060
rect 21980 60002 22036 60284
rect 21980 59950 21982 60002
rect 22034 59950 22036 60002
rect 21980 59938 22036 59950
rect 21756 59686 21812 59724
rect 22092 59444 22148 63868
rect 21644 59378 21700 59388
rect 21868 59388 22148 59444
rect 21868 56082 21924 59388
rect 21980 59218 22036 59230
rect 21980 59166 21982 59218
rect 22034 59166 22036 59218
rect 21980 59108 22036 59166
rect 22204 59220 22260 64428
rect 22428 64484 22484 64542
rect 22428 64148 22484 64428
rect 22428 64082 22484 64092
rect 22316 62468 22372 62478
rect 22316 59778 22372 62412
rect 22316 59726 22318 59778
rect 22370 59726 22372 59778
rect 22316 59444 22372 59726
rect 22316 59378 22372 59388
rect 22428 59220 22484 59230
rect 22204 59218 22484 59220
rect 22204 59166 22430 59218
rect 22482 59166 22484 59218
rect 22204 59164 22484 59166
rect 22428 59154 22484 59164
rect 21980 58436 22036 59052
rect 22092 59106 22148 59118
rect 22092 59054 22094 59106
rect 22146 59054 22148 59106
rect 22092 58884 22148 59054
rect 22204 58884 22260 58894
rect 22092 58828 22204 58884
rect 22540 58828 22596 66444
rect 22876 64484 22932 64494
rect 22876 64390 22932 64428
rect 22876 64036 22932 64046
rect 22876 63942 22932 63980
rect 22764 63924 22820 63934
rect 22764 63830 22820 63868
rect 22988 62188 23044 68348
rect 23324 67954 23380 68796
rect 23436 68740 23492 69468
rect 23660 69300 23716 69310
rect 23884 69300 23940 72044
rect 23996 71874 24052 71886
rect 23996 71822 23998 71874
rect 24050 71822 24052 71874
rect 23996 71540 24052 71822
rect 24108 71874 24164 72044
rect 24108 71822 24110 71874
rect 24162 71822 24164 71874
rect 24108 71810 24164 71822
rect 24556 71652 24612 71662
rect 24556 71558 24612 71596
rect 24444 71540 24500 71550
rect 23996 71538 24500 71540
rect 23996 71486 24446 71538
rect 24498 71486 24500 71538
rect 23996 71484 24500 71486
rect 24108 70644 24164 70654
rect 23716 69244 23940 69300
rect 23996 70194 24052 70206
rect 23996 70142 23998 70194
rect 24050 70142 24052 70194
rect 23996 70084 24052 70142
rect 23548 68740 23604 68750
rect 23436 68684 23548 68740
rect 23548 68674 23604 68684
rect 23324 67902 23326 67954
rect 23378 67902 23380 67954
rect 23324 67890 23380 67902
rect 23100 66164 23156 66174
rect 23100 66162 23492 66164
rect 23100 66110 23102 66162
rect 23154 66110 23492 66162
rect 23100 66108 23492 66110
rect 23100 66098 23156 66108
rect 23436 64820 23492 66108
rect 23548 64820 23604 64830
rect 23436 64818 23604 64820
rect 23436 64766 23550 64818
rect 23602 64766 23604 64818
rect 23436 64764 23604 64766
rect 23548 64754 23604 64764
rect 23324 64594 23380 64606
rect 23324 64542 23326 64594
rect 23378 64542 23380 64594
rect 23324 64484 23380 64542
rect 23324 64418 23380 64428
rect 23548 64596 23604 64606
rect 23548 64482 23604 64540
rect 23548 64430 23550 64482
rect 23602 64430 23604 64482
rect 23324 62468 23380 62478
rect 23324 62374 23380 62412
rect 23548 62188 23604 64430
rect 23660 62468 23716 69244
rect 23772 68852 23828 68862
rect 23772 68758 23828 68796
rect 23996 68628 24052 70028
rect 23996 68562 24052 68572
rect 24108 69186 24164 70588
rect 24444 70082 24500 71484
rect 24444 70030 24446 70082
rect 24498 70030 24500 70082
rect 24444 70018 24500 70030
rect 24220 69972 24276 69982
rect 24220 69970 24388 69972
rect 24220 69918 24222 69970
rect 24274 69918 24388 69970
rect 24220 69916 24388 69918
rect 24220 69906 24276 69916
rect 24108 69134 24110 69186
rect 24162 69134 24164 69186
rect 24108 68516 24164 69134
rect 24108 68450 24164 68460
rect 24220 68628 24276 68638
rect 24220 68514 24276 68572
rect 24220 68462 24222 68514
rect 24274 68462 24276 68514
rect 24220 68402 24276 68462
rect 24220 68350 24222 68402
rect 24274 68350 24276 68402
rect 24220 68338 24276 68350
rect 24332 67228 24388 69916
rect 25004 69410 25060 69422
rect 25004 69358 25006 69410
rect 25058 69358 25060 69410
rect 24556 69186 24612 69198
rect 24556 69134 24558 69186
rect 24610 69134 24612 69186
rect 24556 68402 24612 69134
rect 24668 68740 24724 68750
rect 24668 68646 24724 68684
rect 25004 68516 25060 69358
rect 25004 68450 25060 68460
rect 24556 68350 24558 68402
rect 24610 68350 24612 68402
rect 24556 68338 24612 68350
rect 24780 68402 24836 68414
rect 24780 68350 24782 68402
rect 24834 68350 24836 68402
rect 23996 67172 24388 67228
rect 23660 62374 23716 62412
rect 23772 62468 23828 62478
rect 23772 62466 23940 62468
rect 23772 62414 23774 62466
rect 23826 62414 23940 62466
rect 23772 62412 23940 62414
rect 23772 62402 23828 62412
rect 22988 62132 23156 62188
rect 23548 62132 23716 62188
rect 22988 61570 23044 61582
rect 22988 61518 22990 61570
rect 23042 61518 23044 61570
rect 22652 61348 22708 61358
rect 22652 61254 22708 61292
rect 22988 61348 23044 61518
rect 22988 61282 23044 61292
rect 22876 59780 22932 59790
rect 22876 59218 22932 59724
rect 23100 59556 23156 62132
rect 22876 59166 22878 59218
rect 22930 59166 22932 59218
rect 22876 59154 22932 59166
rect 22988 59500 23156 59556
rect 22204 58818 22260 58828
rect 21980 57876 22036 58380
rect 22428 58772 22596 58828
rect 22652 59108 22708 59118
rect 21980 57820 22372 57876
rect 22316 56868 22372 57820
rect 22428 57650 22484 58772
rect 22428 57598 22430 57650
rect 22482 57598 22484 57650
rect 22428 57586 22484 57598
rect 22540 57538 22596 57550
rect 22540 57486 22542 57538
rect 22594 57486 22596 57538
rect 22316 56812 22484 56868
rect 22316 56642 22372 56654
rect 22316 56590 22318 56642
rect 22370 56590 22372 56642
rect 22316 56308 22372 56590
rect 21868 56030 21870 56082
rect 21922 56030 21924 56082
rect 21868 56018 21924 56030
rect 21980 56252 22372 56308
rect 21420 55858 21588 55860
rect 21420 55806 21422 55858
rect 21474 55806 21588 55858
rect 21420 55804 21588 55806
rect 21420 55794 21476 55804
rect 21308 55410 21364 55422
rect 21308 55358 21310 55410
rect 21362 55358 21364 55410
rect 21308 54626 21364 55358
rect 21420 55300 21476 55310
rect 21420 55186 21476 55244
rect 21420 55134 21422 55186
rect 21474 55134 21476 55186
rect 21420 55122 21476 55134
rect 21532 55188 21588 55804
rect 21644 55188 21700 55198
rect 21532 55186 21700 55188
rect 21532 55134 21646 55186
rect 21698 55134 21700 55186
rect 21532 55132 21700 55134
rect 21308 54574 21310 54626
rect 21362 54574 21364 54626
rect 21308 54562 21364 54574
rect 21644 53620 21700 55132
rect 21644 53554 21700 53564
rect 20748 50372 20916 50428
rect 20972 50372 21140 50428
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19292 49870 19294 49922
rect 19346 49870 19348 49922
rect 19292 49858 19348 49870
rect 19628 49812 19684 49822
rect 19628 49718 19684 49756
rect 20636 49810 20692 49822
rect 20636 49758 20638 49810
rect 20690 49758 20692 49810
rect 20076 49700 20132 49710
rect 20076 49698 20244 49700
rect 20076 49646 20078 49698
rect 20130 49646 20244 49698
rect 20076 49644 20244 49646
rect 20076 49634 20132 49644
rect 19516 49364 19572 49374
rect 19572 49308 19684 49364
rect 19516 49298 19572 49308
rect 19516 49026 19572 49038
rect 19516 48974 19518 49026
rect 19570 48974 19572 49026
rect 19516 48018 19572 48974
rect 19516 47966 19518 48018
rect 19570 47966 19572 48018
rect 19516 47954 19572 47966
rect 19516 47234 19572 47246
rect 19516 47182 19518 47234
rect 19570 47182 19572 47234
rect 19516 46900 19572 47182
rect 19516 46834 19572 46844
rect 19404 46674 19460 46686
rect 19404 46622 19406 46674
rect 19458 46622 19460 46674
rect 18732 46172 19236 46228
rect 19292 46564 19348 46574
rect 18620 44436 18676 44446
rect 18620 44342 18676 44380
rect 18284 43764 18340 43774
rect 18284 43538 18340 43708
rect 18284 43486 18286 43538
rect 18338 43486 18340 43538
rect 18284 43474 18340 43486
rect 18060 42532 18116 42542
rect 18060 42438 18116 42476
rect 18508 42530 18564 42542
rect 18508 42478 18510 42530
rect 18562 42478 18564 42530
rect 18508 42420 18564 42478
rect 18396 42364 18564 42420
rect 18396 41970 18452 42364
rect 18732 42308 18788 46172
rect 18956 46002 19012 46014
rect 18956 45950 18958 46002
rect 19010 45950 19012 46002
rect 18956 45220 19012 45950
rect 19292 45890 19348 46508
rect 19292 45838 19294 45890
rect 19346 45838 19348 45890
rect 19292 45668 19348 45838
rect 19292 45602 19348 45612
rect 19180 45332 19236 45342
rect 19404 45332 19460 46622
rect 19516 45780 19572 45790
rect 19516 45686 19572 45724
rect 19180 45330 19460 45332
rect 19180 45278 19182 45330
rect 19234 45278 19460 45330
rect 19180 45276 19460 45278
rect 19068 45220 19124 45230
rect 18956 45218 19124 45220
rect 18956 45166 19070 45218
rect 19122 45166 19124 45218
rect 18956 45164 19124 45166
rect 19068 45154 19124 45164
rect 19180 44996 19236 45276
rect 19628 45220 19684 49308
rect 20188 49138 20244 49644
rect 20636 49698 20692 49758
rect 20636 49646 20638 49698
rect 20690 49646 20692 49698
rect 20636 49634 20692 49646
rect 20188 49086 20190 49138
rect 20242 49086 20244 49138
rect 20076 49026 20132 49038
rect 20076 48974 20078 49026
rect 20130 48974 20132 49026
rect 20076 48804 20132 48974
rect 20076 48738 20132 48748
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20188 48468 20244 49086
rect 20076 48412 20244 48468
rect 20300 49028 20356 49038
rect 19740 48242 19796 48254
rect 19740 48190 19742 48242
rect 19794 48190 19796 48242
rect 19740 47236 19796 48190
rect 19964 47236 20020 47274
rect 19740 47180 19964 47236
rect 20076 47236 20132 48412
rect 20300 48244 20356 48972
rect 20748 48914 20804 50372
rect 20748 48862 20750 48914
rect 20802 48862 20804 48914
rect 20748 48850 20804 48862
rect 20300 47572 20356 48188
rect 20636 48242 20692 48254
rect 20636 48190 20638 48242
rect 20690 48190 20692 48242
rect 20636 48132 20692 48190
rect 20636 48066 20692 48076
rect 20300 47516 20580 47572
rect 20412 47236 20468 47246
rect 20076 47180 20244 47236
rect 19964 47170 20020 47180
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20188 46788 20244 47180
rect 19964 46732 20244 46788
rect 20300 47234 20468 47236
rect 20300 47182 20414 47234
rect 20466 47182 20468 47234
rect 20300 47180 20468 47182
rect 19852 46564 19908 46574
rect 19964 46564 20020 46732
rect 20300 46676 20356 47180
rect 20412 47170 20468 47180
rect 19852 46562 20020 46564
rect 19852 46510 19854 46562
rect 19906 46510 20020 46562
rect 19852 46508 20020 46510
rect 20076 46564 20132 46574
rect 19852 45780 19908 46508
rect 20076 46470 20132 46508
rect 19852 45714 19908 45724
rect 20188 46116 20244 46126
rect 20188 45890 20244 46060
rect 20188 45838 20190 45890
rect 20242 45838 20244 45890
rect 20188 45668 20244 45838
rect 20300 45892 20356 46620
rect 20412 46674 20468 46686
rect 20412 46622 20414 46674
rect 20466 46622 20468 46674
rect 20412 46114 20468 46622
rect 20412 46062 20414 46114
rect 20466 46062 20468 46114
rect 20412 46050 20468 46062
rect 20524 45892 20580 47516
rect 20636 47012 20692 47022
rect 20636 46116 20692 46956
rect 20636 46050 20692 46060
rect 20748 45892 20804 45902
rect 20524 45890 20804 45892
rect 20524 45838 20750 45890
rect 20802 45838 20804 45890
rect 20524 45836 20804 45838
rect 20300 45826 20356 45836
rect 20188 45612 20356 45668
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19068 44940 19236 44996
rect 19516 45164 19684 45220
rect 19068 44210 19124 44940
rect 19068 44158 19070 44210
rect 19122 44158 19124 44210
rect 19068 44146 19124 44158
rect 19180 44436 19236 44446
rect 19180 44322 19236 44380
rect 19180 44270 19182 44322
rect 19234 44270 19236 44322
rect 18844 44098 18900 44110
rect 18844 44046 18846 44098
rect 18898 44046 18900 44098
rect 18844 43652 18900 44046
rect 18956 43652 19012 43662
rect 18844 43650 19012 43652
rect 18844 43598 18958 43650
rect 19010 43598 19012 43650
rect 18844 43596 19012 43598
rect 18956 43586 19012 43596
rect 18956 43428 19012 43438
rect 18956 42868 19012 43372
rect 19180 43204 19236 44270
rect 19180 43138 19236 43148
rect 18396 41918 18398 41970
rect 18450 41918 18452 41970
rect 18060 41748 18116 41758
rect 18060 41654 18116 41692
rect 17948 41246 17950 41298
rect 18002 41246 18004 41298
rect 17948 41234 18004 41246
rect 18396 40628 18452 41918
rect 18396 40562 18452 40572
rect 18508 42252 18788 42308
rect 18844 42866 19012 42868
rect 18844 42814 18958 42866
rect 19010 42814 19012 42866
rect 18844 42812 19012 42814
rect 17500 40516 17556 40526
rect 16492 40460 16772 40516
rect 16156 40338 16212 40348
rect 16716 39732 16772 40460
rect 17500 40422 17556 40460
rect 18172 40404 18228 40414
rect 16828 39732 16884 39742
rect 16716 39730 16884 39732
rect 16716 39678 16830 39730
rect 16882 39678 16884 39730
rect 16716 39676 16884 39678
rect 16828 39666 16884 39676
rect 17948 39732 18004 39742
rect 17948 39638 18004 39676
rect 16268 39620 16324 39630
rect 16268 39058 16324 39564
rect 16268 39006 16270 39058
rect 16322 39006 16324 39058
rect 16268 38994 16324 39006
rect 17276 39618 17332 39630
rect 17276 39566 17278 39618
rect 17330 39566 17332 39618
rect 16604 38836 16660 38846
rect 16604 38668 16660 38780
rect 16156 38610 16212 38622
rect 16156 38558 16158 38610
rect 16210 38558 16212 38610
rect 16156 37490 16212 38558
rect 16156 37438 16158 37490
rect 16210 37438 16212 37490
rect 16156 37426 16212 37438
rect 16268 38612 16660 38668
rect 15820 36652 16100 36708
rect 15708 36596 15764 36606
rect 15820 36596 15876 36652
rect 15708 36594 15876 36596
rect 15708 36542 15710 36594
rect 15762 36542 15876 36594
rect 15708 36540 15876 36542
rect 15260 35588 15316 35598
rect 15148 33348 15204 33358
rect 15260 33348 15316 35532
rect 15708 34244 15764 36540
rect 15932 36484 15988 36494
rect 15932 35586 15988 36428
rect 15932 35534 15934 35586
rect 15986 35534 15988 35586
rect 15932 35028 15988 35534
rect 15932 34468 15988 34972
rect 15932 34402 15988 34412
rect 15708 34178 15764 34188
rect 15932 34132 15988 34142
rect 16268 34132 16324 38612
rect 16828 37380 16884 37390
rect 16716 37156 16772 37166
rect 16716 37062 16772 37100
rect 16492 37044 16548 37054
rect 16492 36950 16548 36988
rect 16828 37044 16884 37324
rect 17276 37156 17332 39566
rect 17948 38836 18004 38846
rect 17948 37490 18004 38780
rect 18172 38668 18228 40348
rect 17948 37438 17950 37490
rect 18002 37438 18004 37490
rect 17948 37426 18004 37438
rect 18060 38612 18228 38668
rect 17500 37156 17556 37166
rect 17276 37154 17556 37156
rect 17276 37102 17502 37154
rect 17554 37102 17556 37154
rect 17276 37100 17556 37102
rect 16380 35588 16436 35598
rect 16380 35494 16436 35532
rect 16828 35586 16884 36988
rect 17500 36484 17556 37100
rect 17836 36484 17892 36494
rect 17500 36482 17892 36484
rect 17500 36430 17838 36482
rect 17890 36430 17892 36482
rect 17500 36428 17892 36430
rect 17388 36370 17444 36382
rect 17388 36318 17390 36370
rect 17442 36318 17444 36370
rect 16828 35534 16830 35586
rect 16882 35534 16884 35586
rect 15932 34130 16324 34132
rect 15932 34078 15934 34130
rect 15986 34078 16324 34130
rect 15932 34076 16324 34078
rect 15820 33908 15876 33918
rect 15820 33458 15876 33852
rect 15820 33406 15822 33458
rect 15874 33406 15876 33458
rect 15820 33394 15876 33406
rect 15148 33346 15316 33348
rect 15148 33294 15150 33346
rect 15202 33294 15316 33346
rect 15148 33292 15316 33294
rect 15148 33282 15204 33292
rect 15260 30996 15316 33292
rect 15260 30884 15316 30940
rect 15484 32564 15540 32574
rect 15484 32450 15540 32508
rect 15820 32564 15876 32574
rect 15932 32564 15988 34076
rect 16380 34020 16436 34030
rect 16380 33684 16436 33964
rect 16380 33618 16436 33628
rect 15876 32508 15988 32564
rect 15820 32498 15876 32508
rect 15484 32398 15486 32450
rect 15538 32398 15540 32450
rect 15372 30884 15428 30894
rect 15260 30882 15428 30884
rect 15260 30830 15374 30882
rect 15426 30830 15428 30882
rect 15260 30828 15428 30830
rect 15148 30324 15204 30334
rect 15260 30324 15316 30828
rect 15372 30818 15428 30828
rect 15148 30322 15316 30324
rect 15148 30270 15150 30322
rect 15202 30270 15316 30322
rect 15148 30268 15316 30270
rect 15148 30258 15204 30268
rect 15260 30212 15316 30268
rect 15260 30146 15316 30156
rect 15260 27746 15316 27758
rect 15260 27694 15262 27746
rect 15314 27694 15316 27746
rect 15260 26964 15316 27694
rect 15484 27188 15540 32398
rect 16828 32004 16884 35534
rect 17052 36258 17108 36270
rect 17052 36206 17054 36258
rect 17106 36206 17108 36258
rect 17052 33908 17108 36206
rect 17388 35140 17444 36318
rect 17836 35588 17892 36428
rect 18060 35700 18116 38612
rect 18396 38162 18452 38174
rect 18396 38110 18398 38162
rect 18450 38110 18452 38162
rect 18172 35812 18228 35822
rect 18172 35718 18228 35756
rect 18060 35634 18116 35644
rect 17836 35522 17892 35532
rect 18396 35588 18452 38110
rect 18396 35522 18452 35532
rect 18508 35364 18564 42252
rect 18844 42196 18900 42812
rect 18956 42802 19012 42812
rect 19292 42756 19348 42766
rect 19292 42662 19348 42700
rect 19404 42644 19460 42654
rect 19404 42550 19460 42588
rect 18620 42140 18900 42196
rect 19068 42532 19124 42542
rect 18620 42082 18676 42140
rect 18620 42030 18622 42082
rect 18674 42030 18676 42082
rect 18620 42018 18676 42030
rect 18732 41970 18788 41982
rect 18732 41918 18734 41970
rect 18786 41918 18788 41970
rect 18732 41860 18788 41918
rect 19068 41972 19124 42476
rect 19404 41972 19460 41982
rect 19516 41972 19572 45164
rect 19628 44994 19684 45006
rect 19628 44942 19630 44994
rect 19682 44942 19684 44994
rect 19628 44772 19684 44942
rect 20300 44772 20356 45612
rect 20748 45220 20804 45836
rect 20972 45332 21028 50372
rect 21084 49700 21140 49710
rect 21084 49606 21140 49644
rect 21532 49698 21588 49710
rect 21532 49646 21534 49698
rect 21586 49646 21588 49698
rect 21196 49586 21252 49598
rect 21196 49534 21198 49586
rect 21250 49534 21252 49586
rect 21196 49250 21252 49534
rect 21196 49198 21198 49250
rect 21250 49198 21252 49250
rect 21196 49186 21252 49198
rect 21308 49028 21364 49066
rect 21308 48962 21364 48972
rect 21308 48804 21364 48814
rect 21532 48804 21588 49646
rect 21364 48748 21588 48804
rect 21756 49700 21812 49710
rect 21756 49028 21812 49644
rect 21868 49028 21924 49038
rect 21756 49026 21924 49028
rect 21756 48974 21870 49026
rect 21922 48974 21924 49026
rect 21756 48972 21924 48974
rect 21308 47236 21364 48748
rect 21420 48132 21476 48142
rect 21420 48038 21476 48076
rect 21420 47236 21476 47246
rect 21308 47234 21476 47236
rect 21308 47182 21422 47234
rect 21474 47182 21476 47234
rect 21308 47180 21476 47182
rect 21420 46788 21476 47180
rect 21308 46676 21364 46686
rect 20972 45276 21140 45332
rect 20748 45154 20804 45164
rect 20972 45108 21028 45118
rect 19628 44716 20356 44772
rect 20860 45106 21028 45108
rect 20860 45054 20974 45106
rect 21026 45054 21028 45106
rect 20860 45052 21028 45054
rect 19628 43428 19684 44716
rect 20636 44098 20692 44110
rect 20636 44046 20638 44098
rect 20690 44046 20692 44098
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20636 43540 20692 44046
rect 19628 43362 19684 43372
rect 20076 43428 20132 43438
rect 20076 42756 20132 43372
rect 20076 42754 20244 42756
rect 20076 42702 20078 42754
rect 20130 42702 20244 42754
rect 20076 42700 20244 42702
rect 20076 42690 20132 42700
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 20188 42084 20244 42700
rect 19068 41970 19348 41972
rect 19068 41918 19070 41970
rect 19122 41918 19348 41970
rect 19068 41916 19348 41918
rect 19068 41906 19124 41916
rect 18732 41636 18788 41804
rect 19180 41748 19236 41758
rect 18732 41580 18900 41636
rect 18732 40516 18788 40526
rect 18732 40422 18788 40460
rect 18844 40404 18900 41580
rect 19068 41186 19124 41198
rect 19068 41134 19070 41186
rect 19122 41134 19124 41186
rect 18844 40338 18900 40348
rect 18956 40514 19012 40526
rect 18956 40462 18958 40514
rect 19010 40462 19012 40514
rect 18956 39732 19012 40462
rect 18956 39666 19012 39676
rect 19068 38836 19124 41134
rect 19180 40402 19236 41692
rect 19292 40516 19348 41916
rect 19404 41970 19572 41972
rect 19404 41918 19406 41970
rect 19458 41918 19572 41970
rect 19404 41916 19572 41918
rect 19404 41906 19460 41916
rect 19292 40450 19348 40460
rect 19180 40350 19182 40402
rect 19234 40350 19236 40402
rect 19180 40338 19236 40350
rect 19068 38770 19124 38780
rect 19180 40180 19236 40190
rect 19180 38722 19236 40124
rect 19180 38670 19182 38722
rect 19234 38670 19236 38722
rect 19068 37380 19124 37390
rect 18620 37378 19124 37380
rect 18620 37326 19070 37378
rect 19122 37326 19124 37378
rect 18620 37324 19124 37326
rect 18620 36594 18676 37324
rect 19068 37314 19124 37324
rect 19180 37380 19236 38670
rect 19180 37314 19236 37324
rect 19292 38948 19348 38958
rect 18732 37154 18788 37166
rect 18732 37102 18734 37154
rect 18786 37102 18788 37154
rect 18732 36932 18788 37102
rect 18956 36932 19012 36942
rect 18732 36876 18956 36932
rect 18956 36866 19012 36876
rect 18620 36542 18622 36594
rect 18674 36542 18676 36594
rect 18620 36530 18676 36542
rect 19068 36820 19124 36830
rect 17388 35074 17444 35084
rect 18396 35308 18564 35364
rect 17948 35028 18004 35038
rect 17948 34934 18004 34972
rect 17052 33842 17108 33852
rect 17612 34130 17668 34142
rect 17612 34078 17614 34130
rect 17666 34078 17668 34130
rect 17612 33684 17668 34078
rect 17612 33618 17668 33628
rect 18396 33906 18452 35308
rect 18508 35140 18564 35150
rect 18508 35046 18564 35084
rect 19068 35026 19124 36764
rect 19292 35028 19348 38892
rect 19516 38668 19572 41916
rect 20076 42028 20244 42084
rect 19964 41858 20020 41870
rect 19964 41806 19966 41858
rect 20018 41806 20020 41858
rect 19964 41300 20020 41806
rect 19964 41206 20020 41244
rect 20076 40964 20132 42028
rect 20636 41860 20692 43484
rect 20860 42978 20916 45052
rect 20972 45042 21028 45052
rect 21084 44548 21140 45276
rect 20860 42926 20862 42978
rect 20914 42926 20916 42978
rect 20860 42914 20916 42926
rect 20972 44492 21140 44548
rect 20748 42754 20804 42766
rect 20748 42702 20750 42754
rect 20802 42702 20804 42754
rect 20748 42532 20804 42702
rect 20860 42532 20916 42542
rect 20748 42476 20860 42532
rect 20636 41794 20692 41804
rect 20748 41636 20804 41646
rect 20748 41298 20804 41580
rect 20748 41246 20750 41298
rect 20802 41246 20804 41298
rect 20748 41234 20804 41246
rect 20076 40908 20244 40964
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19964 40404 20020 40414
rect 19964 40310 20020 40348
rect 20188 39844 20244 40908
rect 20524 40516 20580 40526
rect 20524 40422 20580 40460
rect 20188 39788 20468 39844
rect 20076 39732 20132 39742
rect 20076 39730 20244 39732
rect 20076 39678 20078 39730
rect 20130 39678 20244 39730
rect 20076 39676 20244 39678
rect 20076 39666 20132 39676
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20188 39060 20244 39676
rect 20412 39172 20468 39788
rect 20860 39620 20916 42476
rect 20524 39396 20580 39406
rect 20524 39394 20692 39396
rect 20524 39342 20526 39394
rect 20578 39342 20692 39394
rect 20524 39340 20692 39342
rect 20524 39330 20580 39340
rect 20412 39060 20468 39116
rect 20524 39060 20580 39070
rect 20412 39058 20580 39060
rect 20412 39006 20526 39058
rect 20578 39006 20580 39058
rect 20412 39004 20580 39006
rect 19964 38948 20020 38958
rect 19516 38612 19796 38668
rect 19628 37828 19684 37838
rect 19404 37826 19684 37828
rect 19404 37774 19630 37826
rect 19682 37774 19684 37826
rect 19404 37772 19684 37774
rect 19740 37828 19796 38612
rect 19964 38274 20020 38892
rect 19964 38222 19966 38274
rect 20018 38222 20020 38274
rect 19964 38210 20020 38222
rect 20188 38162 20244 39004
rect 20524 38994 20580 39004
rect 20636 38612 20692 39340
rect 20860 38946 20916 39564
rect 20860 38894 20862 38946
rect 20914 38894 20916 38946
rect 20860 38882 20916 38894
rect 20636 38546 20692 38556
rect 20188 38110 20190 38162
rect 20242 38110 20244 38162
rect 20188 38098 20244 38110
rect 20972 38052 21028 44492
rect 21308 44436 21364 46620
rect 21420 45668 21476 46732
rect 21532 47124 21588 47134
rect 21532 46786 21588 47068
rect 21756 47012 21812 48972
rect 21868 48962 21924 48972
rect 21532 46734 21534 46786
rect 21586 46734 21588 46786
rect 21532 46676 21588 46734
rect 21532 46610 21588 46620
rect 21644 46900 21700 46910
rect 21644 46674 21700 46844
rect 21644 46622 21646 46674
rect 21698 46622 21700 46674
rect 21476 45612 21588 45668
rect 21420 45574 21476 45612
rect 21420 44436 21476 44446
rect 21308 44434 21476 44436
rect 21308 44382 21422 44434
rect 21474 44382 21476 44434
rect 21308 44380 21476 44382
rect 21308 43652 21364 44380
rect 21420 44370 21476 44380
rect 21308 43586 21364 43596
rect 21420 43540 21476 43550
rect 21420 43446 21476 43484
rect 21084 43428 21140 43438
rect 21084 43426 21364 43428
rect 21084 43374 21086 43426
rect 21138 43374 21364 43426
rect 21084 43372 21364 43374
rect 21084 43362 21140 43372
rect 21308 42866 21364 43372
rect 21308 42814 21310 42866
rect 21362 42814 21364 42866
rect 21308 42802 21364 42814
rect 21532 42756 21588 45612
rect 21644 43540 21700 46622
rect 21756 46676 21812 46956
rect 21868 46676 21924 46686
rect 21756 46620 21868 46676
rect 21868 46610 21924 46620
rect 21644 43474 21700 43484
rect 21756 45780 21812 45790
rect 21756 44994 21812 45724
rect 21868 45666 21924 45678
rect 21868 45614 21870 45666
rect 21922 45614 21924 45666
rect 21868 45220 21924 45614
rect 21868 45154 21924 45164
rect 21756 44942 21758 44994
rect 21810 44942 21812 44994
rect 21756 43426 21812 44942
rect 21980 44772 22036 56252
rect 22316 56084 22372 56094
rect 22428 56084 22484 56812
rect 22316 56082 22484 56084
rect 22316 56030 22318 56082
rect 22370 56030 22484 56082
rect 22316 56028 22484 56030
rect 22316 56018 22372 56028
rect 22428 55410 22484 56028
rect 22428 55358 22430 55410
rect 22482 55358 22484 55410
rect 22428 55346 22484 55358
rect 22540 53956 22596 57486
rect 22316 53900 22596 53956
rect 22204 52164 22260 52174
rect 22092 48132 22148 48142
rect 22092 47346 22148 48076
rect 22092 47294 22094 47346
rect 22146 47294 22148 47346
rect 22092 47282 22148 47294
rect 22204 45218 22260 52108
rect 22316 47236 22372 53900
rect 22652 52948 22708 59052
rect 22764 59106 22820 59118
rect 22764 59054 22766 59106
rect 22818 59054 22820 59106
rect 22764 57650 22820 59054
rect 22764 57598 22766 57650
rect 22818 57598 22820 57650
rect 22764 57586 22820 57598
rect 22988 56866 23044 59500
rect 23212 59444 23268 59454
rect 22988 56814 22990 56866
rect 23042 56814 23044 56866
rect 22988 56802 23044 56814
rect 23100 57092 23156 57102
rect 22764 56082 22820 56094
rect 22764 56030 22766 56082
rect 22818 56030 22820 56082
rect 22764 55972 22820 56030
rect 22764 55906 22820 55916
rect 23100 55970 23156 57036
rect 23100 55918 23102 55970
rect 23154 55918 23156 55970
rect 22764 55188 22820 55198
rect 22764 55186 23044 55188
rect 22764 55134 22766 55186
rect 22818 55134 23044 55186
rect 22764 55132 23044 55134
rect 22764 55122 22820 55132
rect 22764 53732 22820 53742
rect 22764 53172 22820 53676
rect 22764 53078 22820 53116
rect 22540 52892 22708 52948
rect 22540 51044 22596 52892
rect 22652 52722 22708 52734
rect 22652 52670 22654 52722
rect 22706 52670 22708 52722
rect 22652 52386 22708 52670
rect 22652 52334 22654 52386
rect 22706 52334 22708 52386
rect 22652 52322 22708 52334
rect 22764 52052 22820 52062
rect 22764 51958 22820 51996
rect 22764 51380 22820 51390
rect 22764 51266 22820 51324
rect 22764 51214 22766 51266
rect 22818 51214 22820 51266
rect 22764 51202 22820 51214
rect 22652 51044 22708 51054
rect 22540 50988 22652 51044
rect 22652 50978 22708 50988
rect 22988 50932 23044 55132
rect 23100 52722 23156 55918
rect 23212 54516 23268 59388
rect 23436 59218 23492 59230
rect 23436 59166 23438 59218
rect 23490 59166 23492 59218
rect 23436 58436 23492 59166
rect 23548 58436 23604 58446
rect 23436 58434 23604 58436
rect 23436 58382 23550 58434
rect 23602 58382 23604 58434
rect 23436 58380 23604 58382
rect 23324 57764 23380 57774
rect 23324 57670 23380 57708
rect 23548 57204 23604 58380
rect 23660 58324 23716 62132
rect 23772 62130 23828 62142
rect 23772 62078 23774 62130
rect 23826 62078 23828 62130
rect 23772 61682 23828 62078
rect 23772 61630 23774 61682
rect 23826 61630 23828 61682
rect 23772 61618 23828 61630
rect 23884 61124 23940 62412
rect 23996 62188 24052 67172
rect 24108 65380 24164 65390
rect 24444 65380 24500 65390
rect 24108 65378 24500 65380
rect 24108 65326 24110 65378
rect 24162 65326 24446 65378
rect 24498 65326 24500 65378
rect 24108 65324 24500 65326
rect 24108 65314 24164 65324
rect 24444 65314 24500 65324
rect 24556 65266 24612 65278
rect 24556 65214 24558 65266
rect 24610 65214 24612 65266
rect 24220 64596 24276 64606
rect 24556 64596 24612 65214
rect 24276 64540 24612 64596
rect 24220 64530 24276 64540
rect 24108 64484 24164 64494
rect 24108 63924 24164 64428
rect 24108 63858 24164 63868
rect 23996 62132 24500 62188
rect 23772 61068 23940 61124
rect 23772 60226 23828 61068
rect 23772 60174 23774 60226
rect 23826 60174 23828 60226
rect 23772 58546 23828 60174
rect 23884 60674 23940 60686
rect 23884 60622 23886 60674
rect 23938 60622 23940 60674
rect 23884 60114 23940 60622
rect 23884 60062 23886 60114
rect 23938 60062 23940 60114
rect 23884 60050 23940 60062
rect 24332 60562 24388 60574
rect 24332 60510 24334 60562
rect 24386 60510 24388 60562
rect 24332 60004 24388 60510
rect 24332 59910 24388 59948
rect 23772 58494 23774 58546
rect 23826 58494 23828 58546
rect 23772 58482 23828 58494
rect 24332 59106 24388 59118
rect 24332 59054 24334 59106
rect 24386 59054 24388 59106
rect 24332 58884 24388 59054
rect 24332 58548 24388 58828
rect 24332 58482 24388 58492
rect 24220 58436 24276 58446
rect 23884 58434 24276 58436
rect 23884 58382 24222 58434
rect 24274 58382 24276 58434
rect 23884 58380 24276 58382
rect 23884 58324 23940 58380
rect 24220 58370 24276 58380
rect 23660 58268 23940 58324
rect 23436 57148 23548 57204
rect 23324 56866 23380 56878
rect 23324 56814 23326 56866
rect 23378 56814 23380 56866
rect 23324 55858 23380 56814
rect 23436 56082 23492 57148
rect 23548 57138 23604 57148
rect 23884 56756 23940 56766
rect 23884 56662 23940 56700
rect 23436 56030 23438 56082
rect 23490 56030 23492 56082
rect 23436 56018 23492 56030
rect 23324 55806 23326 55858
rect 23378 55806 23380 55858
rect 23324 55794 23380 55806
rect 24332 55300 24388 55310
rect 24444 55300 24500 62132
rect 24780 61236 24836 68350
rect 25228 67228 25284 73164
rect 25340 70308 25396 70318
rect 25340 68850 25396 70252
rect 25452 70194 25508 74956
rect 25900 74900 25956 74910
rect 25900 74806 25956 74844
rect 27580 74786 27636 75404
rect 27580 74734 27582 74786
rect 27634 74734 27636 74786
rect 27580 73948 27636 74734
rect 27244 73892 27636 73948
rect 29372 73948 29428 75628
rect 29932 75684 29988 76300
rect 30044 76290 30100 76300
rect 30492 75908 30548 75918
rect 30604 75908 30660 76414
rect 30492 75906 30660 75908
rect 30492 75854 30494 75906
rect 30546 75854 30660 75906
rect 30492 75852 30660 75854
rect 31276 76244 31332 77196
rect 33516 76578 33572 77308
rect 33516 76526 33518 76578
rect 33570 76526 33572 76578
rect 33516 76514 33572 76526
rect 33740 77026 33796 77038
rect 33740 76974 33742 77026
rect 33794 76974 33796 77026
rect 33740 76468 33796 76974
rect 33964 76468 34020 76478
rect 33740 76466 34020 76468
rect 33740 76414 33966 76466
rect 34018 76414 34020 76466
rect 33740 76412 34020 76414
rect 30492 75842 30548 75852
rect 30156 75796 30212 75806
rect 30156 75702 30212 75740
rect 30940 75796 30996 75806
rect 30940 75702 30996 75740
rect 29932 75590 29988 75628
rect 30828 75684 30884 75694
rect 29820 74900 29876 74910
rect 29372 73892 29540 73948
rect 25900 73330 25956 73342
rect 25900 73278 25902 73330
rect 25954 73278 25956 73330
rect 25564 73220 25620 73230
rect 25900 73220 25956 73278
rect 25620 73164 25956 73220
rect 26684 73220 26740 73230
rect 25564 73126 25620 73164
rect 26684 73126 26740 73164
rect 25564 71650 25620 71662
rect 25564 71598 25566 71650
rect 25618 71598 25620 71650
rect 25564 71092 25620 71598
rect 26124 71652 26180 71662
rect 26180 71596 26404 71652
rect 26124 71558 26180 71596
rect 25676 71538 25732 71550
rect 25676 71486 25678 71538
rect 25730 71486 25732 71538
rect 25676 71316 25732 71486
rect 25676 71260 26180 71316
rect 25676 71092 25732 71102
rect 26012 71092 26068 71102
rect 25564 71090 25732 71092
rect 25564 71038 25678 71090
rect 25730 71038 25732 71090
rect 25564 71036 25732 71038
rect 25676 71026 25732 71036
rect 25788 71090 26068 71092
rect 25788 71038 26014 71090
rect 26066 71038 26068 71090
rect 25788 71036 26068 71038
rect 25788 70420 25844 71036
rect 26012 71026 26068 71036
rect 25452 70142 25454 70194
rect 25506 70142 25508 70194
rect 25452 70130 25508 70142
rect 25676 70364 25844 70420
rect 26124 70754 26180 71260
rect 26348 71204 26404 71596
rect 26348 71110 26404 71148
rect 26124 70702 26126 70754
rect 26178 70702 26180 70754
rect 25676 69522 25732 70364
rect 26012 70308 26068 70318
rect 25676 69470 25678 69522
rect 25730 69470 25732 69522
rect 25676 69458 25732 69470
rect 25788 70196 25844 70206
rect 25340 68798 25342 68850
rect 25394 68798 25396 68850
rect 25340 68740 25396 68798
rect 25340 68674 25396 68684
rect 25788 68852 25844 70140
rect 26012 70082 26068 70252
rect 26124 70196 26180 70702
rect 26908 70754 26964 70766
rect 26908 70702 26910 70754
rect 26962 70702 26964 70754
rect 26908 70532 26964 70702
rect 26908 70466 26964 70476
rect 26572 70196 26628 70206
rect 26124 70194 26628 70196
rect 26124 70142 26574 70194
rect 26626 70142 26628 70194
rect 26124 70140 26628 70142
rect 26572 70130 26628 70140
rect 26908 70194 26964 70206
rect 26908 70142 26910 70194
rect 26962 70142 26964 70194
rect 26012 70030 26014 70082
rect 26066 70030 26068 70082
rect 26012 70018 26068 70030
rect 26908 70084 26964 70142
rect 26908 70018 26964 70028
rect 25788 68514 25844 68796
rect 25788 68462 25790 68514
rect 25842 68462 25844 68514
rect 25228 67172 25396 67228
rect 25340 66946 25396 67172
rect 25340 66894 25342 66946
rect 25394 66894 25396 66946
rect 25228 66386 25284 66398
rect 25228 66334 25230 66386
rect 25282 66334 25284 66386
rect 25228 65604 25284 66334
rect 25340 66276 25396 66894
rect 25676 66276 25732 66286
rect 25340 66274 25732 66276
rect 25340 66222 25678 66274
rect 25730 66222 25732 66274
rect 25340 66220 25732 66222
rect 25340 65604 25396 65614
rect 25228 65602 25396 65604
rect 25228 65550 25342 65602
rect 25394 65550 25396 65602
rect 25228 65548 25396 65550
rect 25340 65538 25396 65548
rect 25452 65268 25508 65278
rect 25452 65266 25620 65268
rect 25452 65214 25454 65266
rect 25506 65214 25620 65266
rect 25452 65212 25620 65214
rect 25452 65202 25508 65212
rect 25340 65044 25396 65054
rect 25340 64484 25396 64988
rect 25228 64482 25396 64484
rect 25228 64430 25342 64482
rect 25394 64430 25396 64482
rect 25228 64428 25396 64430
rect 25004 61348 25060 61358
rect 25228 61348 25284 64428
rect 25340 64418 25396 64428
rect 24780 61170 24836 61180
rect 24892 61292 25004 61348
rect 25060 61292 25284 61348
rect 24556 61012 24612 61022
rect 24556 60918 24612 60956
rect 24668 60676 24724 60686
rect 24668 60582 24724 60620
rect 24892 60116 24948 61292
rect 25004 61282 25060 61292
rect 25228 60786 25284 61292
rect 25228 60734 25230 60786
rect 25282 60734 25284 60786
rect 25228 60722 25284 60734
rect 25340 63924 25396 63934
rect 24892 60022 24948 60060
rect 25004 60004 25060 60014
rect 24780 59106 24836 59118
rect 24780 59054 24782 59106
rect 24834 59054 24836 59106
rect 24780 58884 24836 59054
rect 24556 58828 24836 58884
rect 24556 58436 24612 58828
rect 24556 58342 24612 58380
rect 24668 58658 24724 58670
rect 24668 58606 24670 58658
rect 24722 58606 24724 58658
rect 24332 55298 24500 55300
rect 24332 55246 24334 55298
rect 24386 55246 24500 55298
rect 24332 55244 24500 55246
rect 24556 57540 24612 57550
rect 24556 55972 24612 57484
rect 24332 55234 24388 55244
rect 24220 55074 24276 55086
rect 24220 55022 24222 55074
rect 24274 55022 24276 55074
rect 23212 54450 23268 54460
rect 23324 54628 23380 54638
rect 23324 53730 23380 54572
rect 24108 54628 24164 54638
rect 24108 54534 24164 54572
rect 23436 54404 23492 54414
rect 23996 54404 24052 54414
rect 23436 54402 24052 54404
rect 23436 54350 23438 54402
rect 23490 54350 23998 54402
rect 24050 54350 24052 54402
rect 23436 54348 24052 54350
rect 23436 54338 23492 54348
rect 23996 54338 24052 54348
rect 24220 53956 24276 55022
rect 23884 53900 24276 53956
rect 24556 54402 24612 55916
rect 24668 55748 24724 58606
rect 24780 58548 24836 58558
rect 24780 57540 24836 58492
rect 25004 58100 25060 59948
rect 25004 58034 25060 58044
rect 25340 57764 25396 63868
rect 25452 59106 25508 59118
rect 25452 59054 25454 59106
rect 25506 59054 25508 59106
rect 25452 57876 25508 59054
rect 25564 58324 25620 65212
rect 25676 65044 25732 66220
rect 25788 65268 25844 68462
rect 26796 69970 26852 69982
rect 26796 69918 26798 69970
rect 26850 69918 26852 69970
rect 26348 66162 26404 66174
rect 26348 66110 26350 66162
rect 26402 66110 26404 66162
rect 26348 65716 26404 66110
rect 26460 65716 26516 65726
rect 26348 65714 26516 65716
rect 26348 65662 26462 65714
rect 26514 65662 26516 65714
rect 26348 65660 26516 65662
rect 26460 65650 26516 65660
rect 26684 65492 26740 65502
rect 25788 65202 25844 65212
rect 26460 65490 26740 65492
rect 26460 65438 26686 65490
rect 26738 65438 26740 65490
rect 26460 65436 26740 65438
rect 25676 64978 25732 64988
rect 25676 64818 25732 64830
rect 25676 64766 25678 64818
rect 25730 64766 25732 64818
rect 25676 64036 25732 64766
rect 25676 63970 25732 63980
rect 25900 61684 25956 61694
rect 26236 61684 26292 61694
rect 25900 61682 26292 61684
rect 25900 61630 25902 61682
rect 25954 61630 26238 61682
rect 26290 61630 26292 61682
rect 25900 61628 26292 61630
rect 25900 61618 25956 61628
rect 26236 61618 26292 61628
rect 26348 61348 26404 61358
rect 25900 61236 25956 61246
rect 25676 58548 25732 58558
rect 25676 58454 25732 58492
rect 25564 58258 25620 58268
rect 25900 58212 25956 61180
rect 26348 61012 26404 61292
rect 26348 60946 26404 60956
rect 26012 60676 26068 60686
rect 26012 60582 26068 60620
rect 26460 60226 26516 65436
rect 26684 65426 26740 65436
rect 26460 60174 26462 60226
rect 26514 60174 26516 60226
rect 26460 60162 26516 60174
rect 26572 65268 26628 65278
rect 26012 60116 26068 60126
rect 26012 59444 26068 60060
rect 26124 59780 26180 59790
rect 26348 59780 26404 59790
rect 26124 59778 26348 59780
rect 26124 59726 26126 59778
rect 26178 59726 26348 59778
rect 26124 59724 26348 59726
rect 26124 59714 26180 59724
rect 26348 59714 26404 59724
rect 26012 59442 26404 59444
rect 26012 59390 26014 59442
rect 26066 59390 26404 59442
rect 26012 59388 26404 59390
rect 26012 59378 26068 59388
rect 26348 59218 26404 59388
rect 26348 59166 26350 59218
rect 26402 59166 26404 59218
rect 26348 59154 26404 59166
rect 26572 58828 26628 65212
rect 26796 62188 26852 69918
rect 26908 68516 26964 68526
rect 26908 68422 26964 68460
rect 27244 68068 27300 73892
rect 28812 73218 28868 73230
rect 28812 73166 28814 73218
rect 28866 73166 28868 73218
rect 26460 58772 26628 58828
rect 26684 62132 26852 62188
rect 27132 68012 27300 68068
rect 27356 72324 27412 72334
rect 27356 68626 27412 72268
rect 28028 70196 28084 70206
rect 28028 70102 28084 70140
rect 28364 70084 28420 70094
rect 28364 69990 28420 70028
rect 28700 69970 28756 69982
rect 28700 69918 28702 69970
rect 28754 69918 28756 69970
rect 27804 69524 27860 69534
rect 27804 69522 27972 69524
rect 27804 69470 27806 69522
rect 27858 69470 27972 69522
rect 27804 69468 27972 69470
rect 27804 69458 27860 69468
rect 27356 68574 27358 68626
rect 27410 68574 27412 68626
rect 27356 68516 27412 68574
rect 27132 62188 27188 68012
rect 27356 67620 27412 68460
rect 27356 67554 27412 67564
rect 27468 67060 27524 67070
rect 27468 66966 27524 67004
rect 27244 66946 27300 66958
rect 27244 66894 27246 66946
rect 27298 66894 27300 66946
rect 27244 66836 27300 66894
rect 27244 66780 27524 66836
rect 27468 66724 27524 66780
rect 27804 66834 27860 66846
rect 27804 66782 27806 66834
rect 27858 66782 27860 66834
rect 27804 66724 27860 66782
rect 27468 66668 27860 66724
rect 27804 65492 27860 66668
rect 27916 65828 27972 69468
rect 28588 69412 28644 69422
rect 28700 69412 28756 69918
rect 28588 69410 28756 69412
rect 28588 69358 28590 69410
rect 28642 69358 28756 69410
rect 28588 69356 28756 69358
rect 28588 69346 28644 69356
rect 28252 69188 28308 69198
rect 28028 69186 28308 69188
rect 28028 69134 28254 69186
rect 28306 69134 28308 69186
rect 28028 69132 28308 69134
rect 28028 68738 28084 69132
rect 28252 69122 28308 69132
rect 28028 68686 28030 68738
rect 28082 68686 28084 68738
rect 28028 68674 28084 68686
rect 28028 66948 28084 66958
rect 28588 66948 28644 66958
rect 28028 66946 28644 66948
rect 28028 66894 28030 66946
rect 28082 66894 28590 66946
rect 28642 66894 28644 66946
rect 28028 66892 28644 66894
rect 28028 66882 28084 66892
rect 28476 66386 28532 66892
rect 28588 66882 28644 66892
rect 28476 66334 28478 66386
rect 28530 66334 28532 66386
rect 27916 65772 28084 65828
rect 27804 65426 27860 65436
rect 27804 64594 27860 64606
rect 27804 64542 27806 64594
rect 27858 64542 27860 64594
rect 27804 64148 27860 64542
rect 27916 64148 27972 64158
rect 27804 64146 27972 64148
rect 27804 64094 27918 64146
rect 27970 64094 27972 64146
rect 27804 64092 27972 64094
rect 27916 64082 27972 64092
rect 27132 62132 27748 62188
rect 26124 58436 26180 58446
rect 26124 58342 26180 58380
rect 25900 58156 26180 58212
rect 25452 57820 25732 57876
rect 24780 57474 24836 57484
rect 25228 57708 25396 57764
rect 25228 57092 25284 57708
rect 25452 57652 25508 57662
rect 25564 57652 25620 57662
rect 25452 57650 25564 57652
rect 25452 57598 25454 57650
rect 25506 57598 25564 57650
rect 25452 57596 25564 57598
rect 25452 57586 25508 57596
rect 25340 57540 25396 57550
rect 25340 57446 25396 57484
rect 25452 57092 25508 57102
rect 25228 57036 25452 57092
rect 25452 56998 25508 57036
rect 25564 56756 25620 57596
rect 25676 57650 25732 57820
rect 25676 57598 25678 57650
rect 25730 57598 25732 57650
rect 25676 56980 25732 57598
rect 25676 56914 25732 56924
rect 25788 56980 25844 56990
rect 25788 56978 26068 56980
rect 25788 56926 25790 56978
rect 25842 56926 26068 56978
rect 25788 56924 26068 56926
rect 25788 56914 25844 56924
rect 25676 56756 25732 56766
rect 25564 56754 25732 56756
rect 25564 56702 25678 56754
rect 25730 56702 25732 56754
rect 25564 56700 25732 56702
rect 25676 56690 25732 56700
rect 26012 56194 26068 56924
rect 26012 56142 26014 56194
rect 26066 56142 26068 56194
rect 26012 56130 26068 56142
rect 25228 56082 25284 56094
rect 25228 56030 25230 56082
rect 25282 56030 25284 56082
rect 24780 55972 24836 55982
rect 25228 55972 25284 56030
rect 24780 55970 25284 55972
rect 24780 55918 24782 55970
rect 24834 55918 25284 55970
rect 24780 55916 25284 55918
rect 24780 55906 24836 55916
rect 24668 55692 24836 55748
rect 24780 55298 24836 55692
rect 24780 55246 24782 55298
rect 24834 55246 24836 55298
rect 24780 55234 24836 55246
rect 24556 54350 24558 54402
rect 24610 54350 24612 54402
rect 23436 53844 23492 53854
rect 23436 53750 23492 53788
rect 23324 53678 23326 53730
rect 23378 53678 23380 53730
rect 23324 53666 23380 53678
rect 23212 53620 23268 53630
rect 23212 53526 23268 53564
rect 23324 53508 23380 53518
rect 23212 53060 23268 53070
rect 23212 52966 23268 53004
rect 23100 52670 23102 52722
rect 23154 52670 23156 52722
rect 23100 52658 23156 52670
rect 23212 52724 23268 52734
rect 23324 52724 23380 53452
rect 23436 53172 23492 53182
rect 23436 52946 23492 53116
rect 23772 52948 23828 52958
rect 23436 52894 23438 52946
rect 23490 52894 23492 52946
rect 23436 52882 23492 52894
rect 23660 52946 23828 52948
rect 23660 52894 23774 52946
rect 23826 52894 23828 52946
rect 23660 52892 23828 52894
rect 23268 52668 23380 52724
rect 23212 52276 23268 52668
rect 23212 52274 23492 52276
rect 23212 52222 23214 52274
rect 23266 52222 23492 52274
rect 23212 52220 23492 52222
rect 23212 52210 23268 52220
rect 23436 51378 23492 52220
rect 23436 51326 23438 51378
rect 23490 51326 23492 51378
rect 23436 51314 23492 51326
rect 23548 52052 23604 52062
rect 23100 51156 23156 51166
rect 23100 51154 23380 51156
rect 23100 51102 23102 51154
rect 23154 51102 23380 51154
rect 23100 51100 23380 51102
rect 23100 51090 23156 51100
rect 22764 50876 23044 50932
rect 22652 50708 22708 50718
rect 22540 50596 22596 50606
rect 22540 50502 22596 50540
rect 22540 49026 22596 49038
rect 22540 48974 22542 49026
rect 22594 48974 22596 49026
rect 22540 48804 22596 48974
rect 22652 48914 22708 50652
rect 22652 48862 22654 48914
rect 22706 48862 22708 48914
rect 22652 48850 22708 48862
rect 22540 48738 22596 48748
rect 22428 47348 22484 47358
rect 22428 47346 22708 47348
rect 22428 47294 22430 47346
rect 22482 47294 22708 47346
rect 22428 47292 22708 47294
rect 22428 47282 22484 47292
rect 22316 47170 22372 47180
rect 22316 46788 22372 46798
rect 22316 46694 22372 46732
rect 22652 46114 22708 47292
rect 22764 46564 22820 50876
rect 22988 50596 23044 50606
rect 22988 50502 23044 50540
rect 23324 49922 23380 51100
rect 23324 49870 23326 49922
rect 23378 49870 23380 49922
rect 23324 49858 23380 49870
rect 23436 51044 23492 51054
rect 23100 49698 23156 49710
rect 23100 49646 23102 49698
rect 23154 49646 23156 49698
rect 22876 49028 22932 49038
rect 23100 49028 23156 49646
rect 22932 48972 23156 49028
rect 22876 48962 22932 48972
rect 22764 46498 22820 46508
rect 23100 48804 23156 48814
rect 22652 46062 22654 46114
rect 22706 46062 22708 46114
rect 22652 46050 22708 46062
rect 22316 45892 22372 45902
rect 22316 45798 22372 45836
rect 22988 45892 23044 45902
rect 23100 45892 23156 48748
rect 23324 48804 23380 48814
rect 23324 48710 23380 48748
rect 23436 46564 23492 50988
rect 23548 48130 23604 51996
rect 23660 51380 23716 52892
rect 23772 52882 23828 52892
rect 23660 51286 23716 51324
rect 23660 50482 23716 50494
rect 23660 50430 23662 50482
rect 23714 50430 23716 50482
rect 23660 50034 23716 50430
rect 23884 50428 23940 53900
rect 24108 53730 24164 53742
rect 24108 53678 24110 53730
rect 24162 53678 24164 53730
rect 23660 49982 23662 50034
rect 23714 49982 23716 50034
rect 23660 49970 23716 49982
rect 23772 50372 23940 50428
rect 23996 53172 24052 53182
rect 23548 48078 23550 48130
rect 23602 48078 23604 48130
rect 23548 48066 23604 48078
rect 23548 47460 23604 47470
rect 23548 46900 23604 47404
rect 23548 46834 23604 46844
rect 23436 46470 23492 46508
rect 23044 45836 23156 45892
rect 22988 45798 23044 45836
rect 22204 45166 22206 45218
rect 22258 45166 22260 45218
rect 22204 45154 22260 45166
rect 22316 45220 22372 45230
rect 21980 44706 22036 44716
rect 22092 45106 22148 45118
rect 22092 45054 22094 45106
rect 22146 45054 22148 45106
rect 21756 43374 21758 43426
rect 21810 43374 21812 43426
rect 21756 43362 21812 43374
rect 21980 44546 22036 44558
rect 21980 44494 21982 44546
rect 22034 44494 22036 44546
rect 21980 44434 22036 44494
rect 21980 44382 21982 44434
rect 22034 44382 22036 44434
rect 21420 42530 21476 42542
rect 21420 42478 21422 42530
rect 21474 42478 21476 42530
rect 21420 42196 21476 42478
rect 21420 42130 21476 42140
rect 21532 42420 21588 42700
rect 21868 42530 21924 42542
rect 21868 42478 21870 42530
rect 21922 42478 21924 42530
rect 21868 42420 21924 42478
rect 21532 42364 21924 42420
rect 21420 41636 21476 41646
rect 21420 41186 21476 41580
rect 21420 41134 21422 41186
rect 21474 41134 21476 41186
rect 21420 41122 21476 41134
rect 21420 39394 21476 39406
rect 21420 39342 21422 39394
rect 21474 39342 21476 39394
rect 21308 39172 21364 39182
rect 21084 39060 21140 39070
rect 21084 38966 21140 39004
rect 21308 39058 21364 39116
rect 21308 39006 21310 39058
rect 21362 39006 21364 39058
rect 21308 38994 21364 39006
rect 21420 38948 21476 39342
rect 21420 38882 21476 38892
rect 21532 38834 21588 42364
rect 21980 41972 22036 44382
rect 22092 42196 22148 45054
rect 22316 43876 22372 45164
rect 22988 45106 23044 45118
rect 22988 45054 22990 45106
rect 23042 45054 23044 45106
rect 22988 44996 23044 45054
rect 22988 44930 23044 44940
rect 22540 44546 22596 44558
rect 22540 44494 22542 44546
rect 22594 44494 22596 44546
rect 22316 42532 22372 43820
rect 22428 44100 22484 44110
rect 22428 43764 22484 44044
rect 22428 43698 22484 43708
rect 22540 43652 22596 44494
rect 22764 44322 22820 44334
rect 22764 44270 22766 44322
rect 22818 44270 22820 44322
rect 22764 44100 22820 44270
rect 22764 44034 22820 44044
rect 23100 43988 23156 45836
rect 23660 45892 23716 45902
rect 23660 45798 23716 45836
rect 23212 45778 23268 45790
rect 23212 45726 23214 45778
rect 23266 45726 23268 45778
rect 23212 44660 23268 45726
rect 23324 45220 23380 45230
rect 23324 45218 23604 45220
rect 23324 45166 23326 45218
rect 23378 45166 23604 45218
rect 23324 45164 23604 45166
rect 23324 45154 23380 45164
rect 23212 44594 23268 44604
rect 23548 44434 23604 45164
rect 23660 44996 23716 45006
rect 23660 44902 23716 44940
rect 23548 44382 23550 44434
rect 23602 44382 23604 44434
rect 23548 44370 23604 44382
rect 23212 43988 23268 43998
rect 23100 43932 23212 43988
rect 22876 43652 22932 43662
rect 22540 43650 22932 43652
rect 22540 43598 22878 43650
rect 22930 43598 22932 43650
rect 22540 43596 22932 43598
rect 22876 43586 22932 43596
rect 22316 42438 22372 42476
rect 22092 42130 22148 42140
rect 23100 41972 23156 41982
rect 21756 41970 22036 41972
rect 21756 41918 21982 41970
rect 22034 41918 22036 41970
rect 21756 41916 22036 41918
rect 21756 41300 21812 41916
rect 21980 41906 22036 41916
rect 22092 41970 23156 41972
rect 22092 41918 23102 41970
rect 23154 41918 23156 41970
rect 22092 41916 23156 41918
rect 21756 40402 21812 41244
rect 22092 41298 22148 41916
rect 23100 41906 23156 41916
rect 22652 41748 22708 41758
rect 22652 41654 22708 41692
rect 22092 41246 22094 41298
rect 22146 41246 22148 41298
rect 22092 41234 22148 41246
rect 21756 40350 21758 40402
rect 21810 40350 21812 40402
rect 21532 38782 21534 38834
rect 21586 38782 21588 38834
rect 21532 38612 21588 38782
rect 21644 38836 21700 38846
rect 21644 38742 21700 38780
rect 21756 38668 21812 40350
rect 21868 40292 21924 40302
rect 21868 40290 22036 40292
rect 21868 40238 21870 40290
rect 21922 40238 22036 40290
rect 21868 40236 22036 40238
rect 21868 40226 21924 40236
rect 21980 39620 22036 40236
rect 23212 40180 23268 43932
rect 23548 43652 23604 43662
rect 23548 43538 23604 43596
rect 23548 43486 23550 43538
rect 23602 43486 23604 43538
rect 23548 43474 23604 43486
rect 23436 43204 23492 43214
rect 23436 42308 23492 43148
rect 23324 42196 23380 42206
rect 23324 42102 23380 42140
rect 23436 42084 23492 42252
rect 23436 42082 23716 42084
rect 23436 42030 23438 42082
rect 23490 42030 23716 42082
rect 23436 42028 23716 42030
rect 23436 42018 23492 42028
rect 23660 41746 23716 42028
rect 23660 41694 23662 41746
rect 23714 41694 23716 41746
rect 23660 41188 23716 41694
rect 23772 41412 23828 50372
rect 23996 50036 24052 53116
rect 24108 53170 24164 53678
rect 24108 53118 24110 53170
rect 24162 53118 24164 53170
rect 24108 53106 24164 53118
rect 24444 53618 24500 53630
rect 24444 53566 24446 53618
rect 24498 53566 24500 53618
rect 24444 52164 24500 53566
rect 24444 52098 24500 52108
rect 24108 50036 24164 50046
rect 23996 50034 24164 50036
rect 23996 49982 24110 50034
rect 24162 49982 24164 50034
rect 23996 49980 24164 49982
rect 24108 48916 24164 49980
rect 24444 49026 24500 49038
rect 24444 48974 24446 49026
rect 24498 48974 24500 49026
rect 24164 48860 24276 48916
rect 24108 48850 24164 48860
rect 23884 48802 23940 48814
rect 23884 48750 23886 48802
rect 23938 48750 23940 48802
rect 23884 48356 23940 48750
rect 24220 48468 24276 48860
rect 23884 47460 23940 48300
rect 23884 47394 23940 47404
rect 23996 48466 24276 48468
rect 23996 48414 24222 48466
rect 24274 48414 24276 48466
rect 23996 48412 24276 48414
rect 23996 47570 24052 48412
rect 24220 48402 24276 48412
rect 24444 48804 24500 48974
rect 23996 47518 23998 47570
rect 24050 47518 24052 47570
rect 23996 47068 24052 47518
rect 24444 47460 24500 48748
rect 24444 47366 24500 47404
rect 23884 47012 24052 47068
rect 23884 42084 23940 47012
rect 23996 46788 24052 46798
rect 23996 46674 24052 46732
rect 23996 46622 23998 46674
rect 24050 46622 24052 46674
rect 23996 46610 24052 46622
rect 24220 44996 24276 45006
rect 24108 44940 24220 44996
rect 23996 44882 24052 44894
rect 23996 44830 23998 44882
rect 24050 44830 24052 44882
rect 23996 43988 24052 44830
rect 23996 43922 24052 43932
rect 23884 42018 23940 42028
rect 23996 43650 24052 43662
rect 23996 43598 23998 43650
rect 24050 43598 24052 43650
rect 23996 43428 24052 43598
rect 23884 41858 23940 41870
rect 23884 41806 23886 41858
rect 23938 41806 23940 41858
rect 23884 41746 23940 41806
rect 23884 41694 23886 41746
rect 23938 41694 23940 41746
rect 23884 41682 23940 41694
rect 23884 41412 23940 41422
rect 23772 41356 23884 41412
rect 23884 41346 23940 41356
rect 23660 41132 23940 41188
rect 23212 40114 23268 40124
rect 21980 39058 22036 39564
rect 23436 39620 23492 39630
rect 23436 39526 23492 39564
rect 23548 39508 23604 39518
rect 23548 39414 23604 39452
rect 23660 39396 23716 39406
rect 23660 39302 23716 39340
rect 21980 39006 21982 39058
rect 22034 39006 22036 39058
rect 21980 38994 22036 39006
rect 20524 37996 21028 38052
rect 21308 38050 21364 38062
rect 21308 37998 21310 38050
rect 21362 37998 21364 38050
rect 19740 37772 20244 37828
rect 19404 37378 19460 37772
rect 19628 37762 19684 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 37492 20244 37772
rect 19404 37326 19406 37378
rect 19458 37326 19460 37378
rect 19404 37314 19460 37326
rect 20076 37436 20244 37492
rect 19740 37266 19796 37278
rect 19740 37214 19742 37266
rect 19794 37214 19796 37266
rect 19740 36932 19796 37214
rect 19740 36260 19796 36876
rect 19628 36204 19796 36260
rect 20076 36260 20132 37436
rect 19516 35028 19572 35038
rect 19068 34974 19070 35026
rect 19122 34974 19124 35026
rect 19068 34962 19124 34974
rect 19180 35026 19572 35028
rect 19180 34974 19518 35026
rect 19570 34974 19572 35026
rect 19180 34972 19572 34974
rect 18844 34914 18900 34926
rect 18844 34862 18846 34914
rect 18898 34862 18900 34914
rect 18844 34804 18900 34862
rect 19180 34804 19236 34972
rect 18844 34748 19236 34804
rect 18396 33854 18398 33906
rect 18450 33854 18452 33906
rect 18396 33796 18452 33854
rect 17948 33460 18004 33470
rect 16828 31938 16884 31948
rect 17164 33458 18004 33460
rect 17164 33406 17950 33458
rect 18002 33406 18004 33458
rect 17164 33404 18004 33406
rect 16940 31554 16996 31566
rect 16940 31502 16942 31554
rect 16994 31502 16996 31554
rect 16268 30324 16324 30334
rect 15596 30212 15652 30222
rect 15596 30118 15652 30156
rect 16268 30210 16324 30268
rect 16940 30324 16996 31502
rect 16940 30258 16996 30268
rect 16268 30158 16270 30210
rect 16322 30158 16324 30210
rect 16268 30146 16324 30158
rect 17052 30212 17108 30222
rect 16044 29540 16100 29550
rect 16044 29446 16100 29484
rect 16604 29428 16660 29438
rect 16268 28868 16324 28878
rect 16268 28774 16324 28812
rect 16604 28866 16660 29372
rect 16604 28814 16606 28866
rect 16658 28814 16660 28866
rect 16604 28802 16660 28814
rect 16828 29426 16884 29438
rect 16828 29374 16830 29426
rect 16882 29374 16884 29426
rect 16828 28868 16884 29374
rect 17052 28868 17108 30156
rect 16828 28812 17108 28868
rect 16044 28530 16100 28542
rect 16044 28478 16046 28530
rect 16098 28478 16100 28530
rect 15596 28084 15652 28094
rect 15596 27858 15652 28028
rect 15596 27806 15598 27858
rect 15650 27806 15652 27858
rect 15596 27412 15652 27806
rect 15596 27346 15652 27356
rect 15484 27132 15652 27188
rect 15260 26908 15428 26964
rect 15372 26852 15540 26908
rect 15148 26402 15204 26414
rect 15148 26350 15150 26402
rect 15202 26350 15204 26402
rect 15148 25618 15204 26350
rect 15372 26292 15428 26302
rect 15148 25566 15150 25618
rect 15202 25566 15204 25618
rect 15148 25554 15204 25566
rect 15260 26290 15428 26292
rect 15260 26238 15374 26290
rect 15426 26238 15428 26290
rect 15260 26236 15428 26238
rect 15148 24164 15204 24174
rect 15260 24164 15316 26236
rect 15372 26226 15428 26236
rect 15484 24164 15540 26852
rect 15148 24162 15316 24164
rect 15148 24110 15150 24162
rect 15202 24110 15316 24162
rect 15148 24108 15316 24110
rect 15372 24108 15540 24164
rect 15148 24098 15204 24108
rect 15372 23940 15428 24108
rect 15148 23884 15428 23940
rect 15484 23940 15540 23950
rect 15036 23828 15092 23838
rect 15036 23378 15092 23772
rect 15036 23326 15038 23378
rect 15090 23326 15092 23378
rect 15036 23314 15092 23326
rect 15148 17892 15204 23884
rect 15484 23380 15540 23884
rect 15596 23548 15652 27132
rect 16044 26628 16100 28478
rect 16268 28084 16324 28094
rect 16268 27990 16324 28028
rect 16828 28082 16884 28812
rect 17052 28754 17108 28812
rect 17052 28702 17054 28754
rect 17106 28702 17108 28754
rect 17052 28690 17108 28702
rect 16828 28030 16830 28082
rect 16882 28030 16884 28082
rect 16828 28018 16884 28030
rect 16940 28644 16996 28654
rect 16044 26562 16100 26572
rect 16492 24948 16548 24958
rect 16492 24854 16548 24892
rect 15708 24612 15764 24622
rect 15708 24050 15764 24556
rect 16044 24612 16100 24622
rect 16044 24518 16100 24556
rect 15708 23998 15710 24050
rect 15762 23998 15764 24050
rect 15708 23986 15764 23998
rect 16044 24164 16100 24174
rect 16044 23826 16100 24108
rect 16828 24050 16884 24062
rect 16828 23998 16830 24050
rect 16882 23998 16884 24050
rect 16716 23940 16772 23950
rect 16828 23940 16884 23998
rect 16772 23884 16884 23940
rect 16716 23874 16772 23884
rect 16044 23774 16046 23826
rect 16098 23774 16100 23826
rect 16044 23762 16100 23774
rect 16380 23828 16436 23838
rect 16940 23828 16996 28588
rect 16380 23734 16436 23772
rect 16828 23772 16996 23828
rect 17052 26068 17108 26078
rect 15596 23492 15764 23548
rect 15484 23286 15540 23324
rect 15036 17836 15204 17892
rect 15260 20804 15316 20814
rect 15596 20804 15652 20814
rect 15260 20802 15652 20804
rect 15260 20750 15262 20802
rect 15314 20750 15598 20802
rect 15650 20750 15652 20802
rect 15260 20748 15652 20750
rect 15036 17108 15092 17836
rect 15148 17668 15204 17678
rect 15260 17668 15316 20748
rect 15596 20738 15652 20748
rect 15148 17666 15316 17668
rect 15148 17614 15150 17666
rect 15202 17614 15316 17666
rect 15148 17612 15316 17614
rect 15596 20020 15652 20030
rect 15148 17444 15204 17612
rect 15148 17378 15204 17388
rect 15260 17108 15316 17118
rect 15036 17106 15316 17108
rect 15036 17054 15262 17106
rect 15314 17054 15316 17106
rect 15036 17052 15316 17054
rect 15036 16884 15092 17052
rect 15260 17042 15316 17052
rect 15036 16818 15092 16828
rect 14924 14530 14980 14588
rect 14924 14478 14926 14530
rect 14978 14478 14980 14530
rect 14924 14466 14980 14478
rect 14140 13794 14196 13804
rect 14588 14308 14644 14318
rect 14028 13010 14084 13020
rect 14252 12962 14308 12974
rect 14252 12910 14254 12962
rect 14306 12910 14308 12962
rect 13804 12740 13860 12750
rect 14252 12740 14308 12910
rect 13804 12738 14308 12740
rect 13804 12686 13806 12738
rect 13858 12686 14308 12738
rect 13804 12684 14308 12686
rect 13804 12674 13860 12684
rect 13580 12460 14084 12516
rect 13132 12450 13188 12460
rect 14028 12180 14084 12460
rect 14252 12404 14308 12684
rect 14252 12338 14308 12348
rect 14140 12180 14196 12190
rect 14028 12178 14196 12180
rect 14028 12126 14142 12178
rect 14194 12126 14196 12178
rect 14028 12124 14196 12126
rect 14140 12114 14196 12124
rect 13692 12066 13748 12078
rect 13692 12014 13694 12066
rect 13746 12014 13748 12066
rect 13468 11282 13524 11294
rect 13468 11230 13470 11282
rect 13522 11230 13524 11282
rect 13468 10612 13524 11230
rect 13468 10546 13524 10556
rect 13580 11172 13636 11182
rect 13692 11172 13748 12014
rect 14476 11732 14532 11742
rect 14364 11620 14420 11630
rect 14140 11508 14196 11518
rect 14140 11414 14196 11452
rect 13580 11170 13748 11172
rect 13580 11118 13582 11170
rect 13634 11118 13748 11170
rect 13580 11116 13748 11118
rect 13804 11170 13860 11182
rect 13804 11118 13806 11170
rect 13858 11118 13860 11170
rect 13580 10610 13636 11116
rect 13580 10558 13582 10610
rect 13634 10558 13636 10610
rect 13356 10498 13412 10510
rect 13356 10446 13358 10498
rect 13410 10446 13412 10498
rect 13356 8932 13412 10446
rect 13580 9826 13636 10558
rect 13580 9774 13582 9826
rect 13634 9774 13636 9826
rect 13580 9762 13636 9774
rect 13356 8866 13412 8876
rect 13356 6692 13412 6702
rect 13356 6598 13412 6636
rect 13468 6690 13524 6702
rect 13468 6638 13470 6690
rect 13522 6638 13524 6690
rect 12796 6524 13020 6580
rect 12796 5122 12852 6524
rect 13020 6514 13076 6524
rect 13468 6132 13524 6638
rect 13804 6692 13860 11118
rect 14252 10612 14308 10622
rect 14252 9940 14308 10556
rect 13916 9884 14308 9940
rect 13916 8372 13972 9884
rect 13916 8278 13972 8316
rect 14028 9716 14084 9726
rect 13804 6626 13860 6636
rect 13692 6580 13748 6590
rect 13692 6486 13748 6524
rect 13804 6356 13860 6366
rect 13468 6076 13748 6132
rect 13132 6020 13188 6030
rect 13132 5926 13188 5964
rect 13692 5908 13748 6076
rect 13804 6018 13860 6300
rect 13804 5966 13806 6018
rect 13858 5966 13860 6018
rect 13804 5954 13860 5966
rect 13692 5796 13748 5852
rect 14028 5906 14084 9660
rect 14364 9042 14420 11564
rect 14364 8990 14366 9042
rect 14418 8990 14420 9042
rect 14364 8978 14420 8990
rect 14476 11394 14532 11676
rect 14476 11342 14478 11394
rect 14530 11342 14532 11394
rect 14364 8260 14420 8270
rect 14476 8260 14532 11342
rect 14588 10724 14644 14252
rect 14700 13636 14756 13646
rect 14700 13634 15092 13636
rect 14700 13582 14702 13634
rect 14754 13582 15092 13634
rect 14700 13580 15092 13582
rect 14700 13570 14756 13580
rect 14700 13412 14756 13422
rect 14700 13074 14756 13356
rect 14700 13022 14702 13074
rect 14754 13022 14756 13074
rect 14700 13010 14756 13022
rect 15036 12850 15092 13580
rect 15372 13524 15428 13534
rect 15372 12962 15428 13468
rect 15372 12910 15374 12962
rect 15426 12910 15428 12962
rect 15372 12898 15428 12910
rect 15036 12798 15038 12850
rect 15090 12798 15092 12850
rect 15036 12786 15092 12798
rect 15260 12404 15316 12414
rect 15260 12178 15316 12348
rect 15260 12126 15262 12178
rect 15314 12126 15316 12178
rect 15260 12114 15316 12126
rect 15596 12402 15652 19964
rect 15708 12964 15764 23492
rect 16828 22372 16884 23772
rect 16940 23604 16996 23614
rect 16940 22594 16996 23548
rect 16940 22542 16942 22594
rect 16994 22542 16996 22594
rect 16940 22530 16996 22542
rect 16828 22306 16884 22316
rect 16380 21700 16436 21710
rect 15820 21476 15876 21486
rect 15820 19906 15876 21420
rect 16380 20914 16436 21644
rect 16380 20862 16382 20914
rect 16434 20862 16436 20914
rect 16380 20850 16436 20862
rect 16380 20020 16436 20030
rect 16380 19926 16436 19964
rect 15820 19854 15822 19906
rect 15874 19854 15876 19906
rect 15820 19842 15876 19854
rect 15932 18562 15988 18574
rect 15932 18510 15934 18562
rect 15986 18510 15988 18562
rect 15820 17780 15876 17790
rect 15932 17780 15988 18510
rect 16156 18452 16212 18462
rect 15820 17778 15988 17780
rect 15820 17726 15822 17778
rect 15874 17726 15988 17778
rect 15820 17724 15988 17726
rect 16044 18450 16212 18452
rect 16044 18398 16158 18450
rect 16210 18398 16212 18450
rect 16044 18396 16212 18398
rect 15820 17714 15876 17724
rect 15932 17108 15988 17118
rect 16044 17108 16100 18396
rect 16156 18386 16212 18396
rect 15932 17106 16100 17108
rect 15932 17054 15934 17106
rect 15986 17054 16100 17106
rect 15932 17052 16100 17054
rect 16604 17444 16660 17454
rect 15932 17042 15988 17052
rect 16268 16772 16324 16782
rect 16268 16678 16324 16716
rect 16492 16770 16548 16782
rect 16492 16718 16494 16770
rect 16546 16718 16548 16770
rect 16380 16212 16436 16222
rect 16492 16212 16548 16718
rect 16380 16210 16548 16212
rect 16380 16158 16382 16210
rect 16434 16158 16548 16210
rect 16380 16156 16548 16158
rect 16380 16100 16436 16156
rect 16380 16034 16436 16044
rect 16604 15538 16660 17388
rect 17052 16772 17108 26012
rect 16828 16716 17052 16772
rect 16828 16210 16884 16716
rect 17052 16706 17108 16716
rect 16828 16158 16830 16210
rect 16882 16158 16884 16210
rect 16828 16146 16884 16158
rect 17164 16212 17220 33404
rect 17948 33394 18004 33404
rect 17948 32562 18004 32574
rect 17948 32510 17950 32562
rect 18002 32510 18004 32562
rect 17500 32450 17556 32462
rect 17500 32398 17502 32450
rect 17554 32398 17556 32450
rect 17500 32228 17556 32398
rect 17500 32162 17556 32172
rect 17948 32228 18004 32510
rect 17948 32162 18004 32172
rect 18172 32004 18228 32014
rect 17276 31666 17332 31678
rect 17276 31614 17278 31666
rect 17330 31614 17332 31666
rect 17276 31556 17332 31614
rect 17948 31556 18004 31566
rect 17276 31554 18004 31556
rect 17276 31502 17950 31554
rect 18002 31502 18004 31554
rect 17276 31500 18004 31502
rect 17948 31490 18004 31500
rect 17388 29540 17444 29550
rect 17388 29446 17444 29484
rect 17612 29428 17668 29438
rect 17612 29334 17668 29372
rect 17500 28868 17556 28878
rect 17500 28754 17556 28812
rect 17500 28702 17502 28754
rect 17554 28702 17556 28754
rect 17500 28690 17556 28702
rect 17612 27858 17668 27870
rect 17612 27806 17614 27858
rect 17666 27806 17668 27858
rect 17612 26852 17668 27806
rect 18060 26962 18116 26974
rect 18060 26910 18062 26962
rect 18114 26910 18116 26962
rect 18060 26908 18116 26910
rect 17276 26628 17332 26638
rect 17276 25620 17332 26572
rect 17276 25526 17332 25564
rect 17612 25508 17668 26796
rect 17724 26852 18116 26908
rect 17724 26514 17780 26852
rect 17724 26462 17726 26514
rect 17778 26462 17780 26514
rect 17724 26450 17780 26462
rect 18172 26292 18228 31948
rect 18284 31892 18340 31902
rect 18284 31798 18340 31836
rect 18396 31668 18452 33740
rect 18508 34020 18564 34030
rect 18508 31890 18564 33964
rect 19068 34018 19124 34030
rect 19068 33966 19070 34018
rect 19122 33966 19124 34018
rect 19068 33684 19124 33966
rect 19068 33618 19124 33628
rect 19292 33908 19348 33918
rect 18620 32452 18676 32462
rect 18620 32450 19236 32452
rect 18620 32398 18622 32450
rect 18674 32398 19236 32450
rect 18620 32396 19236 32398
rect 18620 32386 18676 32396
rect 18508 31838 18510 31890
rect 18562 31838 18564 31890
rect 18508 31826 18564 31838
rect 18732 32228 18788 32238
rect 18396 31612 18676 31668
rect 18396 30324 18452 30334
rect 18284 30322 18452 30324
rect 18284 30270 18398 30322
rect 18450 30270 18452 30322
rect 18284 30268 18452 30270
rect 18284 26404 18340 30268
rect 18396 30258 18452 30268
rect 18396 27746 18452 27758
rect 18396 27694 18398 27746
rect 18450 27694 18452 27746
rect 18396 26962 18452 27694
rect 18396 26910 18398 26962
rect 18450 26910 18452 26962
rect 18396 26898 18452 26910
rect 18284 26348 18452 26404
rect 18060 26236 18228 26292
rect 18060 26068 18116 26236
rect 18284 26180 18340 26190
rect 18060 25974 18116 26012
rect 18172 26178 18340 26180
rect 18172 26126 18286 26178
rect 18338 26126 18340 26178
rect 18172 26124 18340 26126
rect 17724 25508 17780 25518
rect 17500 25506 17780 25508
rect 17500 25454 17726 25506
rect 17778 25454 17780 25506
rect 17500 25452 17780 25454
rect 17500 24948 17556 25452
rect 17724 25442 17780 25452
rect 17500 24854 17556 24892
rect 17948 23156 18004 23166
rect 17724 23044 17780 23054
rect 17276 23042 17780 23044
rect 17276 22990 17726 23042
rect 17778 22990 17780 23042
rect 17276 22988 17780 22990
rect 17276 20188 17332 22988
rect 17724 22978 17780 22988
rect 17836 22932 17892 22942
rect 17836 22596 17892 22876
rect 17724 22540 17892 22596
rect 17500 22482 17556 22494
rect 17500 22430 17502 22482
rect 17554 22430 17556 22482
rect 17388 21700 17444 21710
rect 17388 21606 17444 21644
rect 17500 21140 17556 22430
rect 17612 22372 17668 22382
rect 17612 22278 17668 22316
rect 17724 21698 17780 22540
rect 17724 21646 17726 21698
rect 17778 21646 17780 21698
rect 17724 21634 17780 21646
rect 17500 21074 17556 21084
rect 17276 20132 17556 20188
rect 17500 17556 17556 20132
rect 17724 18676 17780 18686
rect 17724 18582 17780 18620
rect 17948 18228 18004 23100
rect 18060 18452 18116 18462
rect 18060 18358 18116 18396
rect 17164 16156 17444 16212
rect 16604 15486 16606 15538
rect 16658 15486 16660 15538
rect 15932 14642 15988 14654
rect 15932 14590 15934 14642
rect 15986 14590 15988 14642
rect 15708 12908 15876 12964
rect 15596 12350 15598 12402
rect 15650 12350 15652 12402
rect 15596 11732 15652 12350
rect 15596 11666 15652 11676
rect 15708 12738 15764 12750
rect 15708 12686 15710 12738
rect 15762 12686 15764 12738
rect 15260 11508 15316 11518
rect 15708 11508 15764 12686
rect 15260 11506 15764 11508
rect 15260 11454 15262 11506
rect 15314 11454 15764 11506
rect 15260 11452 15764 11454
rect 15260 11442 15316 11452
rect 14588 10658 14644 10668
rect 15820 10612 15876 12908
rect 15932 12404 15988 14590
rect 16604 14308 16660 15486
rect 17276 15986 17332 15998
rect 17276 15934 17278 15986
rect 17330 15934 17332 15986
rect 17276 14644 17332 15934
rect 16604 14242 16660 14252
rect 16828 14588 17332 14644
rect 16828 13636 16884 14588
rect 17388 14532 17444 16156
rect 17276 14476 17388 14532
rect 16828 13634 17108 13636
rect 16828 13582 16830 13634
rect 16882 13582 17108 13634
rect 16828 13580 17108 13582
rect 16828 13570 16884 13580
rect 16940 13188 16996 13198
rect 16828 13132 16940 13188
rect 16828 13074 16884 13132
rect 16940 13122 16996 13132
rect 16828 13022 16830 13074
rect 16882 13022 16884 13074
rect 16044 12852 16100 12862
rect 16492 12852 16548 12862
rect 16044 12850 16548 12852
rect 16044 12798 16046 12850
rect 16098 12798 16494 12850
rect 16546 12798 16548 12850
rect 16044 12796 16548 12798
rect 16044 12786 16100 12796
rect 16492 12786 16548 12796
rect 15932 12338 15988 12348
rect 16828 12402 16884 13022
rect 17052 13074 17108 13580
rect 17052 13022 17054 13074
rect 17106 13022 17108 13074
rect 17052 13010 17108 13022
rect 16828 12350 16830 12402
rect 16882 12350 16884 12402
rect 15820 10546 15876 10556
rect 16604 10724 16660 10734
rect 16604 10498 16660 10668
rect 16604 10446 16606 10498
rect 16658 10446 16660 10498
rect 16604 10434 16660 10446
rect 15260 9940 15316 9950
rect 16828 9940 16884 12350
rect 17276 9940 17332 14476
rect 17388 14466 17444 14476
rect 17388 14308 17444 14318
rect 17388 14214 17444 14252
rect 17388 13524 17444 13534
rect 17388 13430 17444 13468
rect 17388 11508 17444 11518
rect 17500 11508 17556 17500
rect 17724 18172 17948 18228
rect 17724 13748 17780 18172
rect 17948 18162 18004 18172
rect 17948 17780 18004 17790
rect 18172 17780 18228 26124
rect 18284 26114 18340 26124
rect 18284 24722 18340 24734
rect 18284 24670 18286 24722
rect 18338 24670 18340 24722
rect 18284 23378 18340 24670
rect 18284 23326 18286 23378
rect 18338 23326 18340 23378
rect 18284 23314 18340 23326
rect 18396 20188 18452 26348
rect 18508 25394 18564 25406
rect 18508 25342 18510 25394
rect 18562 25342 18564 25394
rect 18508 24946 18564 25342
rect 18508 24894 18510 24946
rect 18562 24894 18564 24946
rect 18508 24882 18564 24894
rect 18508 24052 18564 24062
rect 18620 24052 18676 31612
rect 18732 30882 18788 32172
rect 19180 31666 19236 32396
rect 19292 32228 19348 33852
rect 19292 32162 19348 32172
rect 19516 33348 19572 34972
rect 19628 35028 19684 36204
rect 20076 36194 20132 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19964 35698 20020 35710
rect 19964 35646 19966 35698
rect 20018 35646 20020 35698
rect 19964 35588 20020 35646
rect 19964 35522 20020 35532
rect 20412 35588 20468 35598
rect 20412 35494 20468 35532
rect 19628 34244 19684 34972
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19628 34178 19684 34188
rect 19516 31892 19572 33292
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20524 32452 20580 37996
rect 20748 37828 20804 37838
rect 21308 37828 21364 37998
rect 20636 37826 21364 37828
rect 20636 37774 20750 37826
rect 20802 37774 21364 37826
rect 20636 37772 21364 37774
rect 20636 33908 20692 37772
rect 20748 37762 20804 37772
rect 21196 37492 21252 37502
rect 21196 37398 21252 37436
rect 21532 37492 21588 38556
rect 21532 37426 21588 37436
rect 21644 38612 21812 38668
rect 23884 38668 23940 41132
rect 23996 39508 24052 43372
rect 23996 39442 24052 39452
rect 24108 38668 24164 44940
rect 24220 44902 24276 44940
rect 24220 41300 24276 41310
rect 24556 41300 24612 54350
rect 24668 52836 24724 52846
rect 24892 52836 24948 55916
rect 25340 55188 25396 55198
rect 25340 55094 25396 55132
rect 25340 54628 25396 54638
rect 25340 54534 25396 54572
rect 25228 54516 25284 54526
rect 25228 54422 25284 54460
rect 25564 54516 25620 54526
rect 25900 54516 25956 54526
rect 25564 54514 25844 54516
rect 25564 54462 25566 54514
rect 25618 54462 25844 54514
rect 25564 54460 25844 54462
rect 25564 54450 25620 54460
rect 25676 53844 25732 53854
rect 25340 53506 25396 53518
rect 25340 53454 25342 53506
rect 25394 53454 25396 53506
rect 25228 52946 25284 52958
rect 25228 52894 25230 52946
rect 25282 52894 25284 52946
rect 25228 52836 25284 52894
rect 24668 52834 25284 52836
rect 24668 52782 24670 52834
rect 24722 52782 25284 52834
rect 24668 52780 25284 52782
rect 24668 50596 24724 52780
rect 25340 51940 25396 53454
rect 24668 50530 24724 50540
rect 25116 51884 25396 51940
rect 25004 48914 25060 48926
rect 25004 48862 25006 48914
rect 25058 48862 25060 48914
rect 24668 48132 24724 48142
rect 24668 47124 24724 48076
rect 25004 48132 25060 48862
rect 25004 48066 25060 48076
rect 24668 47058 24724 47068
rect 25116 47068 25172 51884
rect 25340 50596 25396 50606
rect 25340 50036 25396 50540
rect 25676 50428 25732 53788
rect 25788 53060 25844 54460
rect 25900 54422 25956 54460
rect 26012 53732 26068 53742
rect 26012 53638 26068 53676
rect 26012 53060 26068 53070
rect 25788 53058 26068 53060
rect 25788 53006 26014 53058
rect 26066 53006 26068 53058
rect 25788 53004 26068 53006
rect 26012 52994 26068 53004
rect 25788 50708 25844 50718
rect 25788 50706 26068 50708
rect 25788 50654 25790 50706
rect 25842 50654 26068 50706
rect 25788 50652 26068 50654
rect 25788 50642 25844 50652
rect 25676 50372 25844 50428
rect 25340 50034 25732 50036
rect 25340 49982 25342 50034
rect 25394 49982 25732 50034
rect 25340 49980 25732 49982
rect 25340 49970 25396 49980
rect 25676 49810 25732 49980
rect 25676 49758 25678 49810
rect 25730 49758 25732 49810
rect 25676 49746 25732 49758
rect 25788 49138 25844 50372
rect 25788 49086 25790 49138
rect 25842 49086 25844 49138
rect 25788 49074 25844 49086
rect 25676 48916 25732 48926
rect 25676 48822 25732 48860
rect 25228 48356 25284 48366
rect 25228 48242 25284 48300
rect 25228 48190 25230 48242
rect 25282 48190 25284 48242
rect 25228 48178 25284 48190
rect 25900 48356 25956 48366
rect 25676 47348 25732 47358
rect 25116 47012 25396 47068
rect 24668 45108 24724 45118
rect 24668 44994 24724 45052
rect 24668 44942 24670 44994
rect 24722 44942 24724 44994
rect 24668 43876 24724 44942
rect 25340 44548 25396 47012
rect 25452 45108 25508 45118
rect 25452 45014 25508 45052
rect 25676 45108 25732 47292
rect 25900 46898 25956 48300
rect 25900 46846 25902 46898
rect 25954 46846 25956 46898
rect 25900 46676 25956 46846
rect 25900 46610 25956 46620
rect 26012 45108 26068 50652
rect 26124 48130 26180 58156
rect 26348 57426 26404 57438
rect 26348 57374 26350 57426
rect 26402 57374 26404 57426
rect 26236 57092 26292 57102
rect 26236 56978 26292 57036
rect 26236 56926 26238 56978
rect 26290 56926 26292 56978
rect 26236 54628 26292 56926
rect 26236 54562 26292 54572
rect 26348 53730 26404 57374
rect 26348 53678 26350 53730
rect 26402 53678 26404 53730
rect 26348 53666 26404 53678
rect 26460 52276 26516 58772
rect 26572 58436 26628 58446
rect 26572 57428 26628 58380
rect 26572 57362 26628 57372
rect 26684 53732 26740 62132
rect 26908 61348 26964 61358
rect 26796 60002 26852 60014
rect 26796 59950 26798 60002
rect 26850 59950 26852 60002
rect 26796 59780 26852 59950
rect 26796 58436 26852 59724
rect 26796 58370 26852 58380
rect 26684 53666 26740 53676
rect 26796 57650 26852 57662
rect 26796 57598 26798 57650
rect 26850 57598 26852 57650
rect 26796 57204 26852 57598
rect 26908 57538 26964 61292
rect 27580 60004 27636 60014
rect 27468 60002 27636 60004
rect 27468 59950 27582 60002
rect 27634 59950 27636 60002
rect 27468 59948 27636 59950
rect 26908 57486 26910 57538
rect 26962 57486 26964 57538
rect 26908 57474 26964 57486
rect 27020 59892 27076 59902
rect 26796 53508 26852 57148
rect 27020 56980 27076 59836
rect 27356 59780 27412 59790
rect 27132 59778 27412 59780
rect 27132 59726 27358 59778
rect 27410 59726 27412 59778
rect 27132 59724 27412 59726
rect 27132 59330 27188 59724
rect 27356 59714 27412 59724
rect 27132 59278 27134 59330
rect 27186 59278 27188 59330
rect 27132 59266 27188 59278
rect 27468 58658 27524 59948
rect 27580 59938 27636 59948
rect 27468 58606 27470 58658
rect 27522 58606 27524 58658
rect 27468 58594 27524 58606
rect 27132 58436 27188 58446
rect 27132 57316 27188 58380
rect 27132 57250 27188 57260
rect 27020 56924 27188 56980
rect 26908 53620 26964 53630
rect 26908 53526 26964 53564
rect 26460 52210 26516 52220
rect 26684 53452 26852 53508
rect 26572 51492 26628 51502
rect 26572 51398 26628 51436
rect 26236 50484 26292 50522
rect 26236 50418 26292 50428
rect 26572 50372 26628 50382
rect 26460 50370 26628 50372
rect 26460 50318 26574 50370
rect 26626 50318 26628 50370
rect 26460 50316 26628 50318
rect 26460 49922 26516 50316
rect 26572 50306 26628 50316
rect 26460 49870 26462 49922
rect 26514 49870 26516 49922
rect 26460 49858 26516 49870
rect 26124 48078 26126 48130
rect 26178 48078 26180 48130
rect 26124 48066 26180 48078
rect 26684 47570 26740 53452
rect 26796 51378 26852 51390
rect 26796 51326 26798 51378
rect 26850 51326 26852 51378
rect 26796 49252 26852 51326
rect 27020 50596 27076 50606
rect 26908 50540 27020 50596
rect 26908 50482 26964 50540
rect 27020 50530 27076 50540
rect 26908 50430 26910 50482
rect 26962 50430 26964 50482
rect 26908 50418 26964 50430
rect 27132 50428 27188 56924
rect 27580 50820 27636 50830
rect 27580 50726 27636 50764
rect 27244 50706 27300 50718
rect 27244 50654 27246 50706
rect 27298 50654 27300 50706
rect 27244 50596 27300 50654
rect 27244 50530 27300 50540
rect 27692 50428 27748 62132
rect 27804 58436 27860 58446
rect 27804 58342 27860 58380
rect 28028 58322 28084 65772
rect 28252 63924 28308 63934
rect 28252 63830 28308 63868
rect 28364 62356 28420 62394
rect 28364 62290 28420 62300
rect 28476 62188 28532 66334
rect 28588 65044 28644 65054
rect 28588 64706 28644 64988
rect 28588 64654 28590 64706
rect 28642 64654 28644 64706
rect 28588 64642 28644 64654
rect 28700 63924 28756 63934
rect 28700 63830 28756 63868
rect 28364 62132 28532 62188
rect 28140 60674 28196 60686
rect 28140 60622 28142 60674
rect 28194 60622 28196 60674
rect 28140 59892 28196 60622
rect 28140 59826 28196 59836
rect 28028 58270 28030 58322
rect 28082 58270 28084 58322
rect 28028 58212 28084 58270
rect 28028 58146 28084 58156
rect 27916 57652 27972 57662
rect 27916 57558 27972 57596
rect 28140 55972 28196 55982
rect 27916 55970 28196 55972
rect 27916 55918 28142 55970
rect 28194 55918 28196 55970
rect 27916 55916 28196 55918
rect 27804 54402 27860 54414
rect 27804 54350 27806 54402
rect 27858 54350 27860 54402
rect 27804 53844 27860 54350
rect 27804 53778 27860 53788
rect 27804 50708 27860 50718
rect 27804 50614 27860 50652
rect 27916 50428 27972 55916
rect 28140 55906 28196 55916
rect 28028 54740 28084 54750
rect 28028 54626 28084 54684
rect 28028 54574 28030 54626
rect 28082 54574 28084 54626
rect 28028 54562 28084 54574
rect 28140 54516 28196 54526
rect 28140 53060 28196 54460
rect 28252 54290 28308 54302
rect 28252 54238 28254 54290
rect 28306 54238 28308 54290
rect 28252 53844 28308 54238
rect 28252 53778 28308 53788
rect 28140 53004 28308 53060
rect 28140 52836 28196 52846
rect 28140 52742 28196 52780
rect 28140 52052 28196 52062
rect 26796 49186 26852 49196
rect 27020 50372 27188 50428
rect 27580 50372 27748 50428
rect 27804 50372 27972 50428
rect 28028 51996 28140 52052
rect 28028 50820 28084 51996
rect 28140 51986 28196 51996
rect 26684 47518 26686 47570
rect 26738 47518 26740 47570
rect 26684 47506 26740 47518
rect 26796 48916 26852 48926
rect 26796 48354 26852 48860
rect 26796 48302 26798 48354
rect 26850 48302 26852 48354
rect 26124 47460 26180 47470
rect 26124 47366 26180 47404
rect 26572 47348 26628 47358
rect 26796 47348 26852 48302
rect 26572 47346 26852 47348
rect 26572 47294 26574 47346
rect 26626 47294 26852 47346
rect 26572 47292 26852 47294
rect 26572 47282 26628 47292
rect 26572 47124 26628 47134
rect 26572 46786 26628 47068
rect 26572 46734 26574 46786
rect 26626 46734 26628 46786
rect 26572 46722 26628 46734
rect 26236 46676 26292 46686
rect 26236 46340 26292 46620
rect 26236 46274 26292 46284
rect 26460 45666 26516 45678
rect 26460 45614 26462 45666
rect 26514 45614 26516 45666
rect 26460 45332 26516 45614
rect 26908 45332 26964 45342
rect 26460 45330 26964 45332
rect 26460 45278 26910 45330
rect 26962 45278 26964 45330
rect 26460 45276 26964 45278
rect 27020 45332 27076 50372
rect 27356 49026 27412 49038
rect 27356 48974 27358 49026
rect 27410 48974 27412 49026
rect 27356 47124 27412 48974
rect 27580 48580 27636 50372
rect 27692 49252 27748 49262
rect 27692 49158 27748 49196
rect 27356 47058 27412 47068
rect 27468 48524 27636 48580
rect 27244 45780 27300 45790
rect 27132 45332 27188 45342
rect 27020 45330 27188 45332
rect 27020 45278 27134 45330
rect 27186 45278 27188 45330
rect 27020 45276 27188 45278
rect 25676 45014 25732 45052
rect 25900 45052 26068 45108
rect 26684 45106 26740 45118
rect 26684 45054 26686 45106
rect 26738 45054 26740 45106
rect 25676 44660 25732 44670
rect 25340 44492 25508 44548
rect 24668 43810 24724 43820
rect 25340 43428 25396 43438
rect 25340 43334 25396 43372
rect 24668 41972 24724 41982
rect 25228 41972 25284 41982
rect 24668 41970 25284 41972
rect 24668 41918 24670 41970
rect 24722 41918 25230 41970
rect 25282 41918 25284 41970
rect 24668 41916 25284 41918
rect 24668 41636 24724 41916
rect 25228 41906 25284 41916
rect 24668 41570 24724 41580
rect 24220 41206 24276 41244
rect 24444 41244 24612 41300
rect 24220 39508 24276 39518
rect 24220 39414 24276 39452
rect 23884 38612 24052 38668
rect 24108 38612 24276 38668
rect 20748 36820 20804 36830
rect 20748 36594 20804 36764
rect 20748 36542 20750 36594
rect 20802 36542 20804 36594
rect 20748 36530 20804 36542
rect 21420 36260 21476 36270
rect 21420 36166 21476 36204
rect 21644 35588 21700 38612
rect 22092 37940 22148 37950
rect 21868 37938 22148 37940
rect 21868 37886 22094 37938
rect 22146 37886 22148 37938
rect 21868 37884 22148 37886
rect 21756 37156 21812 37166
rect 21756 37062 21812 37100
rect 21868 36260 21924 37884
rect 22092 37874 22148 37884
rect 21644 35522 21700 35532
rect 21756 36204 21924 36260
rect 22540 37828 22596 37838
rect 21420 34804 21476 34814
rect 20636 33842 20692 33852
rect 21308 34802 21476 34804
rect 21308 34750 21422 34802
rect 21474 34750 21476 34802
rect 21308 34748 21476 34750
rect 20748 33796 20804 33806
rect 20748 33458 20804 33740
rect 21308 33570 21364 34748
rect 21420 34738 21476 34748
rect 21756 34802 21812 36204
rect 21756 34750 21758 34802
rect 21810 34750 21812 34802
rect 21756 34738 21812 34750
rect 21420 34018 21476 34030
rect 21420 33966 21422 34018
rect 21474 33966 21476 34018
rect 21420 33908 21476 33966
rect 21756 34020 21812 34030
rect 21756 33926 21812 33964
rect 21420 33842 21476 33852
rect 21308 33518 21310 33570
rect 21362 33518 21364 33570
rect 21308 33506 21364 33518
rect 21644 33796 21700 33806
rect 21644 33570 21700 33740
rect 21644 33518 21646 33570
rect 21698 33518 21700 33570
rect 21644 33506 21700 33518
rect 20748 33406 20750 33458
rect 20802 33406 20804 33458
rect 20748 33394 20804 33406
rect 22540 33460 22596 37772
rect 23884 37156 23940 37166
rect 23772 37154 23940 37156
rect 23772 37102 23886 37154
rect 23938 37102 23940 37154
rect 23772 37100 23940 37102
rect 23772 36370 23828 37100
rect 23884 37090 23940 37100
rect 23772 36318 23774 36370
rect 23826 36318 23828 36370
rect 23772 36306 23828 36318
rect 23548 36260 23604 36270
rect 22540 33458 22708 33460
rect 22540 33406 22542 33458
rect 22594 33406 22708 33458
rect 22540 33404 22708 33406
rect 22540 33394 22596 33404
rect 21868 33346 21924 33358
rect 21868 33294 21870 33346
rect 21922 33294 21924 33346
rect 20748 32452 20804 32462
rect 20524 32450 20804 32452
rect 20524 32398 20750 32450
rect 20802 32398 20804 32450
rect 20524 32396 20804 32398
rect 20748 32386 20804 32396
rect 19404 31780 19460 31790
rect 19180 31614 19182 31666
rect 19234 31614 19236 31666
rect 19180 31602 19236 31614
rect 19292 31778 19460 31780
rect 19292 31726 19406 31778
rect 19458 31726 19460 31778
rect 19292 31724 19460 31726
rect 19292 31332 19348 31724
rect 19404 31714 19460 31724
rect 19068 31276 19348 31332
rect 19068 31218 19124 31276
rect 19068 31166 19070 31218
rect 19122 31166 19124 31218
rect 19068 31154 19124 31166
rect 19404 30996 19460 31006
rect 19516 30996 19572 31836
rect 19964 31892 20020 31902
rect 19964 31798 20020 31836
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19404 30994 19572 30996
rect 19404 30942 19406 30994
rect 19458 30942 19572 30994
rect 19404 30940 19572 30942
rect 19404 30930 19460 30940
rect 18732 30830 18734 30882
rect 18786 30830 18788 30882
rect 18732 30212 18788 30830
rect 19516 30660 19572 30940
rect 20076 30994 20132 31006
rect 20076 30942 20078 30994
rect 20130 30942 20132 30994
rect 19628 30884 19684 30894
rect 19628 30790 19684 30828
rect 19516 30604 19908 30660
rect 18732 30146 18788 30156
rect 19852 30322 19908 30604
rect 19852 30270 19854 30322
rect 19906 30270 19908 30322
rect 19852 30100 19908 30270
rect 20076 30212 20132 30942
rect 20748 30884 20804 30894
rect 20748 30882 21364 30884
rect 20748 30830 20750 30882
rect 20802 30830 21364 30882
rect 20748 30828 21364 30830
rect 20748 30818 20804 30828
rect 20076 30146 20132 30156
rect 19852 30034 19908 30044
rect 20636 30100 20692 30110
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20636 29540 20692 30044
rect 21308 30098 21364 30828
rect 21532 30212 21588 30222
rect 21308 30046 21310 30098
rect 21362 30046 21364 30098
rect 21308 30034 21364 30046
rect 21420 30210 21588 30212
rect 21420 30158 21534 30210
rect 21586 30158 21588 30210
rect 21420 30156 21588 30158
rect 21420 29764 21476 30156
rect 21532 30146 21588 30156
rect 20972 29708 21476 29764
rect 20972 29650 21028 29708
rect 20972 29598 20974 29650
rect 21026 29598 21028 29650
rect 20972 29586 21028 29598
rect 20636 29426 20692 29484
rect 21420 29540 21476 29550
rect 21420 29446 21476 29484
rect 20636 29374 20638 29426
rect 20690 29374 20692 29426
rect 20636 29362 20692 29374
rect 20412 29314 20468 29326
rect 20412 29262 20414 29314
rect 20466 29262 20468 29314
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19404 27076 19460 27086
rect 18732 26178 18788 26190
rect 18732 26126 18734 26178
rect 18786 26126 18788 26178
rect 18732 26068 18788 26126
rect 18732 26002 18788 26012
rect 18508 24050 18676 24052
rect 18508 23998 18510 24050
rect 18562 23998 18676 24050
rect 18508 23996 18676 23998
rect 18508 23156 18564 23996
rect 18508 23090 18564 23100
rect 18956 23268 19012 23278
rect 18620 22932 18676 22942
rect 18956 22932 19012 23212
rect 18620 22838 18676 22876
rect 18844 22930 19012 22932
rect 18844 22878 18958 22930
rect 19010 22878 19012 22930
rect 18844 22876 19012 22878
rect 18508 22820 18564 22830
rect 18508 21362 18564 22764
rect 18620 21476 18676 21486
rect 18620 21382 18676 21420
rect 18508 21310 18510 21362
rect 18562 21310 18564 21362
rect 18508 21298 18564 21310
rect 18284 20132 18452 20188
rect 18508 20914 18564 20926
rect 18508 20862 18510 20914
rect 18562 20862 18564 20914
rect 18284 18340 18340 20132
rect 18284 18246 18340 18284
rect 17948 17778 18228 17780
rect 17948 17726 17950 17778
rect 18002 17726 18228 17778
rect 17948 17724 18228 17726
rect 17948 17668 18004 17724
rect 17948 17602 18004 17612
rect 18508 17332 18564 20862
rect 18844 20188 18900 22876
rect 18956 22866 19012 22876
rect 19180 23042 19236 23054
rect 19180 22990 19182 23042
rect 19234 22990 19236 23042
rect 19180 22708 19236 22990
rect 19404 23044 19460 27020
rect 20412 26908 20468 29262
rect 20524 27748 20580 27758
rect 20524 27654 20580 27692
rect 21868 27748 21924 33294
rect 22652 33124 22708 33404
rect 22764 33348 22820 33358
rect 22764 33254 22820 33292
rect 23436 33234 23492 33246
rect 23436 33182 23438 33234
rect 23490 33182 23492 33234
rect 23100 33124 23156 33134
rect 23436 33124 23492 33182
rect 22652 33068 22932 33124
rect 22876 30882 22932 33068
rect 23100 33122 23492 33124
rect 23100 33070 23102 33122
rect 23154 33070 23492 33122
rect 23100 33068 23492 33070
rect 23100 33058 23156 33068
rect 23548 32452 23604 36204
rect 23884 34020 23940 34030
rect 23772 34018 23940 34020
rect 23772 33966 23886 34018
rect 23938 33966 23940 34018
rect 23772 33964 23940 33966
rect 23772 33234 23828 33964
rect 23884 33954 23940 33964
rect 23772 33182 23774 33234
rect 23826 33182 23828 33234
rect 23772 33170 23828 33182
rect 23548 32386 23604 32396
rect 22876 30830 22878 30882
rect 22930 30830 22932 30882
rect 22876 30818 22932 30830
rect 22316 30212 22372 30222
rect 21308 27076 21364 27114
rect 20860 27020 21140 27076
rect 20860 26908 20916 27020
rect 20412 26852 20916 26908
rect 21084 26908 21140 27020
rect 21308 27010 21364 27020
rect 21420 26962 21476 26974
rect 21420 26910 21422 26962
rect 21474 26910 21476 26962
rect 21420 26908 21476 26910
rect 21868 26964 21924 27692
rect 21980 29316 22036 29326
rect 22316 29316 22372 30156
rect 23100 30100 23156 30110
rect 23100 30098 23380 30100
rect 23100 30046 23102 30098
rect 23154 30046 23380 30098
rect 23100 30044 23380 30046
rect 23100 30034 23156 30044
rect 21980 29314 22372 29316
rect 21980 29262 21982 29314
rect 22034 29262 22372 29314
rect 21980 29260 22372 29262
rect 21980 27188 22036 29260
rect 23324 28530 23380 30044
rect 23884 29540 23940 29550
rect 23324 28478 23326 28530
rect 23378 28478 23380 28530
rect 23324 28466 23380 28478
rect 23436 28756 23492 28766
rect 23212 28420 23268 28430
rect 22316 28308 22372 28318
rect 22204 27748 22260 27758
rect 22316 27748 22372 28252
rect 22764 27972 22820 27982
rect 22764 27878 22820 27916
rect 22204 27746 22372 27748
rect 22204 27694 22206 27746
rect 22258 27694 22372 27746
rect 22204 27692 22372 27694
rect 22204 27682 22260 27692
rect 21980 27122 22036 27132
rect 22204 27074 22260 27086
rect 22204 27022 22206 27074
rect 22258 27022 22260 27074
rect 22204 26964 22260 27022
rect 22316 27076 22372 27692
rect 22316 27010 22372 27020
rect 23212 27186 23268 28364
rect 23436 27858 23492 28700
rect 23436 27806 23438 27858
rect 23490 27806 23492 27858
rect 23436 27794 23492 27806
rect 23548 28642 23604 28654
rect 23548 28590 23550 28642
rect 23602 28590 23604 28642
rect 23548 27298 23604 28590
rect 23548 27246 23550 27298
rect 23602 27246 23604 27298
rect 23548 27234 23604 27246
rect 23884 27298 23940 29484
rect 23996 28532 24052 38612
rect 24220 38162 24276 38612
rect 24220 38110 24222 38162
rect 24274 38110 24276 38162
rect 24220 38098 24276 38110
rect 24444 37268 24500 41244
rect 24668 41188 24724 41198
rect 25228 41188 25284 41198
rect 24668 41186 25284 41188
rect 24668 41134 24670 41186
rect 24722 41134 25230 41186
rect 25282 41134 25284 41186
rect 24668 41132 25284 41134
rect 24668 41122 24724 41132
rect 25228 41122 25284 41132
rect 24892 40964 24948 40974
rect 24892 40870 24948 40908
rect 24668 40740 24724 40750
rect 24668 40626 24724 40684
rect 24668 40574 24670 40626
rect 24722 40574 24724 40626
rect 24668 40562 24724 40574
rect 24780 39396 24836 39406
rect 24780 39060 24836 39340
rect 24444 37202 24500 37212
rect 24668 37266 24724 37278
rect 24668 37214 24670 37266
rect 24722 37214 24724 37266
rect 24108 36372 24164 36382
rect 24556 36372 24612 36382
rect 24108 36370 24612 36372
rect 24108 36318 24110 36370
rect 24162 36318 24558 36370
rect 24610 36318 24612 36370
rect 24108 36316 24612 36318
rect 24108 36306 24164 36316
rect 24556 36306 24612 36316
rect 24668 36260 24724 37214
rect 24668 36194 24724 36204
rect 24556 34130 24612 34142
rect 24556 34078 24558 34130
rect 24610 34078 24612 34130
rect 24556 33908 24612 34078
rect 24556 33842 24612 33852
rect 24220 33348 24276 33358
rect 24220 33254 24276 33292
rect 24668 32452 24724 32462
rect 24668 32358 24724 32396
rect 24556 31556 24612 31566
rect 24444 29764 24500 29774
rect 24444 28756 24500 29708
rect 24444 28662 24500 28700
rect 24556 28532 24612 31500
rect 23996 28466 24052 28476
rect 24444 28476 24612 28532
rect 23884 27246 23886 27298
rect 23938 27246 23940 27298
rect 23212 27134 23214 27186
rect 23266 27134 23268 27186
rect 21868 26908 22260 26964
rect 22540 26964 22596 27002
rect 20972 26852 21028 26862
rect 21084 26852 21476 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20636 25618 20692 26852
rect 20972 26180 21028 26796
rect 22428 26850 22484 26862
rect 22428 26798 22430 26850
rect 22482 26798 22484 26850
rect 20972 26086 21028 26124
rect 21420 26290 21476 26302
rect 21420 26238 21422 26290
rect 21474 26238 21476 26290
rect 21420 26180 21476 26238
rect 21420 26114 21476 26124
rect 22092 26180 22148 26190
rect 22092 26178 22372 26180
rect 22092 26126 22094 26178
rect 22146 26126 22372 26178
rect 22092 26124 22372 26126
rect 22092 26114 22148 26124
rect 20636 25566 20638 25618
rect 20690 25566 20692 25618
rect 20636 25554 20692 25566
rect 22092 25620 22148 25630
rect 21980 25396 22036 25406
rect 21756 25394 22036 25396
rect 21756 25342 21982 25394
rect 22034 25342 22036 25394
rect 21756 25340 22036 25342
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20972 24722 21028 24734
rect 20972 24670 20974 24722
rect 21026 24670 21028 24722
rect 19740 24612 19796 24622
rect 19740 24518 19796 24556
rect 20188 24500 20244 24510
rect 20188 24406 20244 24444
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19628 23268 19684 23278
rect 19628 23174 19684 23212
rect 19404 22988 19684 23044
rect 19180 22642 19236 22652
rect 18956 22370 19012 22382
rect 18956 22318 18958 22370
rect 19010 22318 19012 22370
rect 18956 20692 19012 22318
rect 19516 22372 19572 22382
rect 19516 21586 19572 22316
rect 19516 21534 19518 21586
rect 19570 21534 19572 21586
rect 19516 21522 19572 21534
rect 18956 20626 19012 20636
rect 18732 20132 18900 20188
rect 19516 20244 19572 20254
rect 18732 18452 18788 20132
rect 19068 20020 19124 20030
rect 19292 20020 19348 20030
rect 19124 20018 19348 20020
rect 19124 19966 19294 20018
rect 19346 19966 19348 20018
rect 19124 19964 19348 19966
rect 19068 19926 19124 19964
rect 19292 19954 19348 19964
rect 18732 18358 18788 18396
rect 18956 18340 19012 18350
rect 18844 17892 18900 17902
rect 18844 17666 18900 17836
rect 18844 17614 18846 17666
rect 18898 17614 18900 17666
rect 18732 17556 18788 17566
rect 18732 17462 18788 17500
rect 18396 17276 18564 17332
rect 18396 16996 18452 17276
rect 18172 16994 18452 16996
rect 18172 16942 18398 16994
rect 18450 16942 18452 16994
rect 18172 16940 18452 16942
rect 17836 16884 17892 16894
rect 17836 16098 17892 16828
rect 18172 16660 18228 16940
rect 18396 16930 18452 16940
rect 18620 16884 18676 16894
rect 18844 16884 18900 17614
rect 17836 16046 17838 16098
rect 17890 16046 17892 16098
rect 17836 16034 17892 16046
rect 17948 16604 18228 16660
rect 18508 16828 18620 16884
rect 18676 16828 18900 16884
rect 18956 16882 19012 18284
rect 19180 17668 19236 17678
rect 19516 17668 19572 20188
rect 19628 18564 19684 22988
rect 20972 23042 21028 24670
rect 21756 24162 21812 25340
rect 21980 25330 22036 25340
rect 22092 24164 22148 25564
rect 22316 25394 22372 26124
rect 22316 25342 22318 25394
rect 22370 25342 22372 25394
rect 22316 25330 22372 25342
rect 22428 25060 22484 26798
rect 21756 24110 21758 24162
rect 21810 24110 21812 24162
rect 21756 24098 21812 24110
rect 21980 24108 22148 24164
rect 22204 25004 22484 25060
rect 20972 22990 20974 23042
rect 21026 22990 21028 23042
rect 20524 22484 20580 22494
rect 19964 22370 20020 22382
rect 19964 22318 19966 22370
rect 20018 22318 20020 22370
rect 19964 22148 20020 22318
rect 20524 22370 20580 22428
rect 20524 22318 20526 22370
rect 20578 22318 20580 22370
rect 20524 22306 20580 22318
rect 20972 22372 21028 22990
rect 21420 22484 21476 22494
rect 21420 22390 21476 22428
rect 21980 22482 22036 24108
rect 22092 23940 22148 23950
rect 22092 23846 22148 23884
rect 22204 23266 22260 25004
rect 22316 24724 22372 24734
rect 22316 24630 22372 24668
rect 22204 23214 22206 23266
rect 22258 23214 22260 23266
rect 22204 23202 22260 23214
rect 22316 23826 22372 23838
rect 22316 23774 22318 23826
rect 22370 23774 22372 23826
rect 22204 22596 22260 22606
rect 22204 22502 22260 22540
rect 21980 22430 21982 22482
rect 22034 22430 22036 22482
rect 21980 22418 22036 22430
rect 20972 22306 21028 22316
rect 19964 22092 20244 22148
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20188 21812 20244 22092
rect 20188 21756 20356 21812
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20300 20188 20356 21756
rect 20860 21588 20916 21598
rect 20860 21494 20916 21532
rect 21644 21474 21700 21486
rect 21644 21422 21646 21474
rect 21698 21422 21700 21474
rect 21644 20244 21700 21422
rect 20300 20132 20580 20188
rect 21644 20178 21700 20188
rect 22204 20692 22260 20702
rect 22316 20692 22372 23774
rect 22428 21586 22484 21598
rect 22428 21534 22430 21586
rect 22482 21534 22484 21586
rect 22428 21476 22484 21534
rect 22428 21410 22484 21420
rect 22540 20916 22596 26908
rect 23212 26964 23268 27134
rect 23212 26898 23268 26908
rect 23884 26852 23940 27246
rect 24108 27860 24164 27870
rect 23212 26292 23268 26302
rect 22988 24722 23044 24734
rect 22988 24670 22990 24722
rect 23042 24670 23044 24722
rect 22988 24612 23044 24670
rect 22988 24546 23044 24556
rect 23100 24610 23156 24622
rect 23100 24558 23102 24610
rect 23154 24558 23156 24610
rect 23100 24164 23156 24558
rect 22204 20690 22372 20692
rect 22204 20638 22206 20690
rect 22258 20638 22372 20690
rect 22204 20636 22372 20638
rect 22428 20860 22596 20916
rect 22652 24108 23156 24164
rect 20076 19908 20132 19918
rect 20076 19906 20356 19908
rect 20076 19854 20078 19906
rect 20130 19854 20356 19906
rect 20076 19852 20356 19854
rect 20076 19842 20132 19852
rect 19964 19122 20020 19134
rect 19964 19070 19966 19122
rect 20018 19070 20020 19122
rect 19964 19012 20020 19070
rect 20300 19122 20356 19852
rect 20300 19070 20302 19122
rect 20354 19070 20356 19122
rect 20300 19058 20356 19070
rect 19964 18956 20244 19012
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20188 18676 20244 18956
rect 20076 18620 20244 18676
rect 19628 18508 20020 18564
rect 19628 17892 19684 18508
rect 19964 18450 20020 18508
rect 19964 18398 19966 18450
rect 20018 18398 20020 18450
rect 19964 18386 20020 18398
rect 19628 17826 19684 17836
rect 20076 17890 20132 18620
rect 20076 17838 20078 17890
rect 20130 17838 20132 17890
rect 20076 17826 20132 17838
rect 20412 18338 20468 18350
rect 20412 18286 20414 18338
rect 20466 18286 20468 18338
rect 20412 18228 20468 18286
rect 19516 17612 19684 17668
rect 19180 17574 19236 17612
rect 19404 17442 19460 17454
rect 19404 17390 19406 17442
rect 19458 17390 19460 17442
rect 18956 16830 18958 16882
rect 19010 16830 19012 16882
rect 17724 13746 17892 13748
rect 17724 13694 17726 13746
rect 17778 13694 17892 13746
rect 17724 13692 17892 13694
rect 17724 13188 17780 13692
rect 17836 13524 17892 13692
rect 17948 13746 18004 16604
rect 18172 16100 18228 16110
rect 18172 16006 18228 16044
rect 18396 15874 18452 15886
rect 18396 15822 18398 15874
rect 18450 15822 18452 15874
rect 18060 14532 18116 14542
rect 18060 14418 18116 14476
rect 18060 14366 18062 14418
rect 18114 14366 18116 14418
rect 18060 14354 18116 14366
rect 18396 13972 18452 15822
rect 18508 15540 18564 16828
rect 18620 16790 18676 16828
rect 18956 16818 19012 16830
rect 19180 17106 19236 17118
rect 19180 17054 19182 17106
rect 19234 17054 19236 17106
rect 19180 16772 19236 17054
rect 19180 16706 19236 16716
rect 19292 17108 19348 17118
rect 19292 16212 19348 17052
rect 19068 16210 19348 16212
rect 19068 16158 19294 16210
rect 19346 16158 19348 16210
rect 19068 16156 19348 16158
rect 18620 15876 18676 15886
rect 19068 15876 19124 16156
rect 19292 16146 19348 16156
rect 18620 15874 19124 15876
rect 18620 15822 18622 15874
rect 18674 15822 19124 15874
rect 18620 15820 19124 15822
rect 18620 15810 18676 15820
rect 18620 15540 18676 15550
rect 18508 15538 18676 15540
rect 18508 15486 18622 15538
rect 18674 15486 18676 15538
rect 18508 15484 18676 15486
rect 18620 15474 18676 15484
rect 19068 15538 19124 15820
rect 19068 15486 19070 15538
rect 19122 15486 19124 15538
rect 19068 15474 19124 15486
rect 19404 15428 19460 17390
rect 19516 17442 19572 17454
rect 19516 17390 19518 17442
rect 19570 17390 19572 17442
rect 19516 17108 19572 17390
rect 19516 17042 19572 17052
rect 19404 15362 19460 15372
rect 19068 14532 19124 14542
rect 18956 14476 19068 14532
rect 18844 14420 18900 14430
rect 18396 13906 18452 13916
rect 18508 14364 18844 14420
rect 17948 13694 17950 13746
rect 18002 13694 18004 13746
rect 17948 13682 18004 13694
rect 18396 13634 18452 13646
rect 18396 13582 18398 13634
rect 18450 13582 18452 13634
rect 18396 13524 18452 13582
rect 17836 13468 18452 13524
rect 17724 13122 17780 13132
rect 17612 12964 17668 12974
rect 17612 12962 18452 12964
rect 17612 12910 17614 12962
rect 17666 12910 18452 12962
rect 17612 12908 18452 12910
rect 17612 12898 17668 12908
rect 17388 11506 17556 11508
rect 17388 11454 17390 11506
rect 17442 11454 17556 11506
rect 17388 11452 17556 11454
rect 17612 12404 17668 12414
rect 17388 11442 17444 11452
rect 17612 10834 17668 12348
rect 17612 10782 17614 10834
rect 17666 10782 17668 10834
rect 17612 10770 17668 10782
rect 17724 12290 17780 12302
rect 17724 12238 17726 12290
rect 17778 12238 17780 12290
rect 15260 9846 15316 9884
rect 16604 9938 16884 9940
rect 16604 9886 16830 9938
rect 16882 9886 16884 9938
rect 16604 9884 16884 9886
rect 14924 9602 14980 9614
rect 14924 9550 14926 9602
rect 14978 9550 14980 9602
rect 14924 9044 14980 9550
rect 14364 8258 14532 8260
rect 14364 8206 14366 8258
rect 14418 8206 14532 8258
rect 14364 8204 14532 8206
rect 14588 8372 14644 8382
rect 14364 8194 14420 8204
rect 14364 7476 14420 7486
rect 14364 7382 14420 7420
rect 14252 6692 14308 6702
rect 14252 6578 14308 6636
rect 14252 6526 14254 6578
rect 14306 6526 14308 6578
rect 14252 6514 14308 6526
rect 14588 6244 14644 8316
rect 14924 7474 14980 8988
rect 15372 9604 15428 9614
rect 15372 9044 15428 9548
rect 16604 9044 16660 9884
rect 16828 9874 16884 9884
rect 16940 9938 17332 9940
rect 16940 9886 17278 9938
rect 17330 9886 17332 9938
rect 16940 9884 17332 9886
rect 15372 9042 15540 9044
rect 15372 8990 15374 9042
rect 15426 8990 15540 9042
rect 15372 8988 15540 8990
rect 15372 8978 15428 8988
rect 15148 8932 15204 8942
rect 15148 8838 15204 8876
rect 15372 8818 15428 8830
rect 15372 8766 15374 8818
rect 15426 8766 15428 8818
rect 15036 8148 15092 8158
rect 15036 8146 15316 8148
rect 15036 8094 15038 8146
rect 15090 8094 15316 8146
rect 15036 8092 15316 8094
rect 15036 8082 15092 8092
rect 15148 7812 15204 7822
rect 14924 7422 14926 7474
rect 14978 7422 14980 7474
rect 14924 7410 14980 7422
rect 15036 7756 15148 7812
rect 14588 6178 14644 6188
rect 14476 6020 14532 6030
rect 15036 6020 15092 7756
rect 15148 7746 15204 7756
rect 15260 7698 15316 8092
rect 15372 7812 15428 8766
rect 15372 7746 15428 7756
rect 15260 7646 15262 7698
rect 15314 7646 15316 7698
rect 15260 7634 15316 7646
rect 15484 7476 15540 8988
rect 16604 8950 16660 8988
rect 16828 9044 16884 9054
rect 16940 9044 16996 9884
rect 17276 9874 17332 9884
rect 17724 9268 17780 12238
rect 16828 9042 16996 9044
rect 16828 8990 16830 9042
rect 16882 8990 16996 9042
rect 16828 8988 16996 8990
rect 17388 9212 17780 9268
rect 17836 11732 17892 11742
rect 17836 11506 17892 11676
rect 17836 11454 17838 11506
rect 17890 11454 17892 11506
rect 16828 8978 16884 8988
rect 16268 8818 16324 8830
rect 16268 8766 16270 8818
rect 16322 8766 16324 8818
rect 16268 8428 16324 8766
rect 17388 8428 17444 9212
rect 17500 9042 17556 9054
rect 17500 8990 17502 9042
rect 17554 8990 17556 9042
rect 17500 8932 17556 8990
rect 17836 8932 17892 11454
rect 18284 9714 18340 9726
rect 18284 9662 18286 9714
rect 18338 9662 18340 9714
rect 17948 9604 18004 9614
rect 17948 9602 18228 9604
rect 17948 9550 17950 9602
rect 18002 9550 18228 9602
rect 17948 9548 18228 9550
rect 17948 9538 18004 9548
rect 18172 9154 18228 9548
rect 18172 9102 18174 9154
rect 18226 9102 18228 9154
rect 18172 9090 18228 9102
rect 17500 8876 17892 8932
rect 15596 8372 16324 8428
rect 17164 8372 17780 8428
rect 15596 7586 15652 8372
rect 17164 8370 17220 8372
rect 17164 8318 17166 8370
rect 17218 8318 17220 8370
rect 17164 8306 17220 8318
rect 17724 8370 17780 8372
rect 17724 8318 17726 8370
rect 17778 8318 17780 8370
rect 17724 8306 17780 8318
rect 15596 7534 15598 7586
rect 15650 7534 15652 7586
rect 15596 7522 15652 7534
rect 15148 7420 15540 7476
rect 16044 7476 16100 7486
rect 15148 6690 15204 7420
rect 16044 7382 16100 7420
rect 15148 6638 15150 6690
rect 15202 6638 15204 6690
rect 15148 6626 15204 6638
rect 17500 7364 17556 7374
rect 17836 7364 17892 8876
rect 17948 9044 18004 9054
rect 17948 8482 18004 8988
rect 17948 8430 17950 8482
rect 18002 8430 18004 8482
rect 17948 8372 18004 8430
rect 18284 8482 18340 9662
rect 18284 8430 18286 8482
rect 18338 8430 18340 8482
rect 18284 8418 18340 8430
rect 17948 8306 18004 8316
rect 17948 7364 18004 7374
rect 17500 7362 18004 7364
rect 17500 7310 17502 7362
rect 17554 7310 17950 7362
rect 18002 7310 18004 7362
rect 17500 7308 18004 7310
rect 17500 6580 17556 7308
rect 17948 7298 18004 7308
rect 15484 6244 15540 6254
rect 15484 6132 15540 6188
rect 15484 6130 15764 6132
rect 15484 6078 15486 6130
rect 15538 6078 15764 6130
rect 15484 6076 15764 6078
rect 15484 6066 15540 6076
rect 14476 5926 14532 5964
rect 14812 6018 15092 6020
rect 14812 5966 15038 6018
rect 15090 5966 15092 6018
rect 14812 5964 15092 5966
rect 14028 5854 14030 5906
rect 14082 5854 14084 5906
rect 14028 5842 14084 5854
rect 14700 5908 14756 5918
rect 14700 5814 14756 5852
rect 13804 5796 13860 5806
rect 13692 5794 13860 5796
rect 13692 5742 13806 5794
rect 13858 5742 13860 5794
rect 13692 5740 13860 5742
rect 12796 5070 12798 5122
rect 12850 5070 12852 5122
rect 12796 5058 12852 5070
rect 13468 5234 13524 5246
rect 13468 5182 13470 5234
rect 13522 5182 13524 5234
rect 13468 5124 13524 5182
rect 13468 5058 13524 5068
rect 13804 5236 13860 5740
rect 14812 5684 14868 5964
rect 15036 5954 15092 5964
rect 14924 5796 14980 5806
rect 14924 5702 14980 5740
rect 13804 5010 13860 5180
rect 14140 5628 14868 5684
rect 14140 5122 14196 5628
rect 14812 5348 14868 5358
rect 14700 5124 14756 5134
rect 14140 5070 14142 5122
rect 14194 5070 14196 5122
rect 14140 5058 14196 5070
rect 14588 5122 14756 5124
rect 14588 5070 14702 5122
rect 14754 5070 14756 5122
rect 14588 5068 14756 5070
rect 13804 4958 13806 5010
rect 13858 4958 13860 5010
rect 13804 4946 13860 4958
rect 14476 4900 14532 4910
rect 13916 4898 14532 4900
rect 13916 4846 14478 4898
rect 14530 4846 14532 4898
rect 13916 4844 14532 4846
rect 12684 4450 13076 4452
rect 12684 4398 12686 4450
rect 12738 4398 13076 4450
rect 12684 4396 13076 4398
rect 12684 4386 12740 4396
rect 13020 3666 13076 4396
rect 13916 4450 13972 4844
rect 14476 4834 14532 4844
rect 13916 4398 13918 4450
rect 13970 4398 13972 4450
rect 13916 4386 13972 4398
rect 13244 4340 13300 4350
rect 14588 4340 14644 5068
rect 14700 5058 14756 5068
rect 13244 4246 13300 4284
rect 14140 4284 14644 4340
rect 14140 3778 14196 4284
rect 14140 3726 14142 3778
rect 14194 3726 14196 3778
rect 14140 3714 14196 3726
rect 14700 4228 14756 4238
rect 13020 3614 13022 3666
rect 13074 3614 13076 3666
rect 13020 3602 13076 3614
rect 14700 3666 14756 4172
rect 14700 3614 14702 3666
rect 14754 3614 14756 3666
rect 14700 3602 14756 3614
rect 13916 3556 13972 3566
rect 14476 3556 14532 3566
rect 13916 3554 14532 3556
rect 13916 3502 13918 3554
rect 13970 3502 14478 3554
rect 14530 3502 14532 3554
rect 13916 3500 14532 3502
rect 13916 3490 13972 3500
rect 14476 3444 14532 3500
rect 14812 3444 14868 5292
rect 15708 5348 15764 6076
rect 15708 5254 15764 5292
rect 15484 5236 15540 5246
rect 15484 5142 15540 5180
rect 15820 5236 15876 5246
rect 15148 4900 15204 4910
rect 15148 4340 15204 4844
rect 15148 3554 15204 4284
rect 15820 4228 15876 5180
rect 16044 4900 16100 4910
rect 16492 4900 16548 4910
rect 16044 4898 16436 4900
rect 16044 4846 16046 4898
rect 16098 4846 16436 4898
rect 16044 4844 16436 4846
rect 16044 4834 16100 4844
rect 16380 4676 16436 4844
rect 16492 4806 16548 4844
rect 17052 4900 17108 4910
rect 17052 4806 17108 4844
rect 17500 4900 17556 6524
rect 18284 6468 18340 6478
rect 17724 6018 17780 6030
rect 18284 6020 18340 6412
rect 18396 6130 18452 12908
rect 18508 12290 18564 14364
rect 18844 14326 18900 14364
rect 18956 13972 19012 14476
rect 19068 14438 19124 14476
rect 18508 12238 18510 12290
rect 18562 12238 18564 12290
rect 18508 11618 18564 12238
rect 18620 13916 19012 13972
rect 19180 14418 19236 14430
rect 19180 14366 19182 14418
rect 19234 14366 19236 14418
rect 18620 12180 18676 13916
rect 19180 13860 19236 14366
rect 19516 13860 19572 13870
rect 19180 13804 19516 13860
rect 19516 13794 19572 13804
rect 18844 13746 18900 13758
rect 18844 13694 18846 13746
rect 18898 13694 18900 13746
rect 18844 13076 18900 13694
rect 19516 13076 19572 13086
rect 19628 13076 19684 17612
rect 20412 17666 20468 18172
rect 20412 17614 20414 17666
rect 20466 17614 20468 17666
rect 20412 17332 20468 17614
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20412 17266 20468 17276
rect 19836 17210 20100 17220
rect 20188 17108 20244 17118
rect 20188 17014 20244 17052
rect 20412 16212 20468 16222
rect 19740 16098 19796 16110
rect 19740 16046 19742 16098
rect 19794 16046 19796 16098
rect 19740 15876 19796 16046
rect 20188 16100 20244 16110
rect 19964 15986 20020 15998
rect 19964 15934 19966 15986
rect 20018 15934 20020 15986
rect 19964 15876 20020 15934
rect 20188 15876 20244 16044
rect 19964 15820 20244 15876
rect 19740 15810 19796 15820
rect 20188 15764 20244 15820
rect 20412 15986 20468 16156
rect 20412 15934 20414 15986
rect 20466 15934 20468 15986
rect 19836 15708 20100 15718
rect 20188 15708 20356 15764
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20188 15540 20244 15550
rect 19740 14644 19796 14654
rect 19740 14550 19796 14588
rect 20188 14644 20244 15484
rect 20188 14550 20244 14588
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 18844 13020 19348 13076
rect 18956 12850 19012 12862
rect 18956 12798 18958 12850
rect 19010 12798 19012 12850
rect 18844 12292 18900 12302
rect 18956 12292 19012 12798
rect 18844 12290 19012 12292
rect 18844 12238 18846 12290
rect 18898 12238 19012 12290
rect 18844 12236 19012 12238
rect 18844 12226 18900 12236
rect 18620 12086 18676 12124
rect 19068 12178 19124 12190
rect 19068 12126 19070 12178
rect 19122 12126 19124 12178
rect 19068 12068 19124 12126
rect 18508 11566 18510 11618
rect 18562 11566 18564 11618
rect 18508 11554 18564 11566
rect 18732 11732 18788 11742
rect 18732 11506 18788 11676
rect 19068 11732 19124 12012
rect 19068 11666 19124 11676
rect 19180 12180 19236 12190
rect 18732 11454 18734 11506
rect 18786 11454 18788 11506
rect 18732 11442 18788 11454
rect 19180 11506 19236 12124
rect 19180 11454 19182 11506
rect 19234 11454 19236 11506
rect 19180 11060 19236 11454
rect 19068 11004 19236 11060
rect 18844 8372 18900 8382
rect 18844 8278 18900 8316
rect 19068 6692 19124 11004
rect 19292 8428 19348 13020
rect 19516 13074 19684 13076
rect 19516 13022 19518 13074
rect 19570 13022 19684 13074
rect 19516 13020 19684 13022
rect 19852 13972 19908 13982
rect 19516 13010 19572 13020
rect 19852 12850 19908 13916
rect 20076 13972 20132 13982
rect 20076 12962 20132 13916
rect 20188 13860 20244 13870
rect 20188 13766 20244 13804
rect 20076 12910 20078 12962
rect 20130 12910 20132 12962
rect 20076 12898 20132 12910
rect 19852 12798 19854 12850
rect 19906 12798 19908 12850
rect 19852 12786 19908 12798
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19852 12068 19908 12078
rect 19852 12066 20132 12068
rect 19852 12014 19854 12066
rect 19906 12014 20132 12066
rect 19852 12012 20132 12014
rect 19852 12002 19908 12012
rect 20076 11788 20132 12012
rect 20076 11732 20244 11788
rect 19740 11618 19796 11630
rect 19740 11566 19742 11618
rect 19794 11566 19796 11618
rect 19740 11506 19796 11566
rect 19740 11454 19742 11506
rect 19794 11454 19796 11506
rect 19740 11442 19796 11454
rect 20188 11282 20244 11732
rect 20188 11230 20190 11282
rect 20242 11230 20244 11282
rect 20188 11218 20244 11230
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20300 8930 20356 15708
rect 20412 14754 20468 15934
rect 20412 14702 20414 14754
rect 20466 14702 20468 14754
rect 20412 14420 20468 14702
rect 20412 14354 20468 14364
rect 20524 13634 20580 20132
rect 22204 19906 22260 20636
rect 22428 20580 22484 20860
rect 22204 19854 22206 19906
rect 22258 19854 22260 19906
rect 22204 19842 22260 19854
rect 22316 20524 22484 20580
rect 22540 20690 22596 20702
rect 22540 20638 22542 20690
rect 22594 20638 22596 20690
rect 22540 20580 22596 20638
rect 20636 17666 20692 17678
rect 20636 17614 20638 17666
rect 20690 17614 20692 17666
rect 20636 16100 20692 17614
rect 21308 17666 21364 17678
rect 21308 17614 21310 17666
rect 21362 17614 21364 17666
rect 21308 17556 21364 17614
rect 22092 17556 22148 17566
rect 20972 16996 21028 17006
rect 21308 16996 21364 17500
rect 21644 17554 22148 17556
rect 21644 17502 22094 17554
rect 22146 17502 22148 17554
rect 21644 17500 22148 17502
rect 21644 17106 21700 17500
rect 22092 17490 22148 17500
rect 21644 17054 21646 17106
rect 21698 17054 21700 17106
rect 21644 17042 21700 17054
rect 22092 17332 22148 17342
rect 20972 16994 21364 16996
rect 20972 16942 20974 16994
rect 21026 16942 21364 16994
rect 20972 16940 21364 16942
rect 20972 16930 21028 16940
rect 21308 16884 21364 16940
rect 21308 16818 21364 16828
rect 21420 16884 21476 16894
rect 21420 16882 21588 16884
rect 21420 16830 21422 16882
rect 21474 16830 21588 16882
rect 21420 16828 21588 16830
rect 21420 16818 21476 16828
rect 20636 16034 20692 16044
rect 21084 16772 21140 16782
rect 20636 15874 20692 15886
rect 20636 15822 20638 15874
rect 20690 15822 20692 15874
rect 20636 15428 20692 15822
rect 20748 15428 20804 15438
rect 20636 15426 20804 15428
rect 20636 15374 20750 15426
rect 20802 15374 20804 15426
rect 20636 15372 20804 15374
rect 20748 15362 20804 15372
rect 20860 15314 20916 15326
rect 20860 15262 20862 15314
rect 20914 15262 20916 15314
rect 20636 14754 20692 14766
rect 20636 14702 20638 14754
rect 20690 14702 20692 14754
rect 20636 14642 20692 14702
rect 20636 14590 20638 14642
rect 20690 14590 20692 14642
rect 20636 14578 20692 14590
rect 20524 13582 20526 13634
rect 20578 13582 20580 13634
rect 20524 13570 20580 13582
rect 20860 11844 20916 15262
rect 21084 13858 21140 16716
rect 21532 16322 21588 16828
rect 22092 16770 22148 17276
rect 22316 17108 22372 20524
rect 22540 20514 22596 20524
rect 22316 17042 22372 17052
rect 22540 20020 22596 20030
rect 22092 16718 22094 16770
rect 22146 16718 22148 16770
rect 21532 16270 21534 16322
rect 21586 16270 21588 16322
rect 21532 16258 21588 16270
rect 21868 16324 21924 16334
rect 22092 16324 22148 16718
rect 21868 16322 22148 16324
rect 21868 16270 21870 16322
rect 21922 16270 22148 16322
rect 21868 16268 22148 16270
rect 21868 16258 21924 16268
rect 22540 16210 22596 19964
rect 22540 16158 22542 16210
rect 22594 16158 22596 16210
rect 22092 16098 22148 16110
rect 22092 16046 22094 16098
rect 22146 16046 22148 16098
rect 21868 15428 21924 15438
rect 21868 15334 21924 15372
rect 22092 14532 22148 16046
rect 22540 15876 22596 16158
rect 22540 15810 22596 15820
rect 22652 15652 22708 24108
rect 22764 23940 22820 23950
rect 22764 23714 22820 23884
rect 22764 23662 22766 23714
rect 22818 23662 22820 23714
rect 22764 23604 22820 23662
rect 23212 23604 23268 26236
rect 23884 26292 23940 26796
rect 23884 26226 23940 26236
rect 23996 27188 24052 27198
rect 23996 26180 24052 27132
rect 24108 27186 24164 27804
rect 24108 27134 24110 27186
rect 24162 27134 24164 27186
rect 24108 26908 24164 27134
rect 24332 27858 24388 27870
rect 24332 27806 24334 27858
rect 24386 27806 24388 27858
rect 24108 26852 24276 26908
rect 23436 25508 23492 25518
rect 23884 25508 23940 25518
rect 23996 25508 24052 26124
rect 24220 26178 24276 26852
rect 24220 26126 24222 26178
rect 24274 26126 24276 26178
rect 24220 26114 24276 26126
rect 23436 25506 24052 25508
rect 23436 25454 23438 25506
rect 23490 25454 23886 25506
rect 23938 25454 24052 25506
rect 23436 25452 24052 25454
rect 23436 25442 23492 25452
rect 23884 25442 23940 25452
rect 22764 23548 23268 23604
rect 22988 23266 23044 23278
rect 22988 23214 22990 23266
rect 23042 23214 23044 23266
rect 22764 23154 22820 23166
rect 22764 23102 22766 23154
rect 22818 23102 22820 23154
rect 22764 21028 22820 23102
rect 22764 20962 22820 20972
rect 22988 20916 23044 23214
rect 23100 22372 23156 22382
rect 23100 22278 23156 22316
rect 23100 20916 23156 20926
rect 22988 20914 23156 20916
rect 22988 20862 23102 20914
rect 23154 20862 23156 20914
rect 22988 20860 23156 20862
rect 23100 20850 23156 20860
rect 22876 20804 22932 20814
rect 22764 20802 22932 20804
rect 22764 20750 22878 20802
rect 22930 20750 22932 20802
rect 22764 20748 22932 20750
rect 22764 20188 22820 20748
rect 22876 20738 22932 20748
rect 22764 20122 22820 20132
rect 22876 20580 22932 20590
rect 22876 20242 22932 20524
rect 22876 20190 22878 20242
rect 22930 20190 22932 20242
rect 22876 20020 22932 20190
rect 23212 20188 23268 23548
rect 23884 22372 23940 22382
rect 23772 22370 23940 22372
rect 23772 22318 23886 22370
rect 23938 22318 23940 22370
rect 23772 22316 23940 22318
rect 23436 21476 23492 21486
rect 23436 20356 23492 21420
rect 23772 21252 23828 22316
rect 23884 22306 23940 22316
rect 23996 21812 24052 25452
rect 24332 24052 24388 27806
rect 24332 23986 24388 23996
rect 24332 23828 24388 23838
rect 24332 22372 24388 23772
rect 24220 21812 24276 21822
rect 24332 21812 24388 22316
rect 24052 21756 24164 21812
rect 23996 21746 24052 21756
rect 23884 21588 23940 21598
rect 23884 21476 23940 21532
rect 23884 21474 24052 21476
rect 23884 21422 23886 21474
rect 23938 21422 24052 21474
rect 23884 21420 24052 21422
rect 23884 21410 23940 21420
rect 23660 21196 23828 21252
rect 23436 20290 23492 20300
rect 23548 20804 23604 20814
rect 23212 20132 23380 20188
rect 23212 20020 23268 20030
rect 22764 19964 22932 20020
rect 22988 20018 23268 20020
rect 22988 19966 23214 20018
rect 23266 19966 23268 20018
rect 22988 19964 23268 19966
rect 22764 16212 22820 19964
rect 22876 19460 22932 19470
rect 22988 19460 23044 19964
rect 23212 19954 23268 19964
rect 22876 19458 23044 19460
rect 22876 19406 22878 19458
rect 22930 19406 23044 19458
rect 22876 19404 23044 19406
rect 22876 19394 22932 19404
rect 23212 19236 23268 19246
rect 23324 19236 23380 20132
rect 23548 20130 23604 20748
rect 23548 20078 23550 20130
rect 23602 20078 23604 20130
rect 23548 20066 23604 20078
rect 23100 19180 23212 19236
rect 23268 19180 23380 19236
rect 23100 18564 23156 19180
rect 23212 19142 23268 19180
rect 23436 19122 23492 19134
rect 23436 19070 23438 19122
rect 23490 19070 23492 19122
rect 23100 18498 23156 18508
rect 23212 18676 23268 18686
rect 22988 16212 23044 16222
rect 22820 16210 23044 16212
rect 22820 16158 22990 16210
rect 23042 16158 23044 16210
rect 22820 16156 23044 16158
rect 22764 16118 22820 16156
rect 22988 16146 23044 16156
rect 22428 15596 22708 15652
rect 22428 15202 22484 15596
rect 22540 15316 22596 15326
rect 22540 15314 22708 15316
rect 22540 15262 22542 15314
rect 22594 15262 22708 15314
rect 22540 15260 22708 15262
rect 22540 15250 22596 15260
rect 22428 15150 22430 15202
rect 22482 15150 22484 15202
rect 22428 15138 22484 15150
rect 22540 14644 22596 14654
rect 22428 14532 22484 14542
rect 22092 14530 22484 14532
rect 22092 14478 22430 14530
rect 22482 14478 22484 14530
rect 22092 14476 22484 14478
rect 21084 13806 21086 13858
rect 21138 13806 21140 13858
rect 21084 13794 21140 13806
rect 21756 13746 21812 13758
rect 22316 13748 22372 13758
rect 21756 13694 21758 13746
rect 21810 13694 21812 13746
rect 21756 13188 21812 13694
rect 21756 13122 21812 13132
rect 21980 13746 22372 13748
rect 21980 13694 22318 13746
rect 22370 13694 22372 13746
rect 21980 13692 22372 13694
rect 21868 12962 21924 12974
rect 21868 12910 21870 12962
rect 21922 12910 21924 12962
rect 21420 12740 21476 12750
rect 21868 12740 21924 12910
rect 21420 12738 21924 12740
rect 21420 12686 21422 12738
rect 21474 12686 21924 12738
rect 21420 12684 21924 12686
rect 21420 12180 21476 12684
rect 21868 12516 21924 12684
rect 21868 12450 21924 12460
rect 21420 12114 21476 12124
rect 21868 12180 21924 12190
rect 20300 8878 20302 8930
rect 20354 8878 20356 8930
rect 20300 8866 20356 8878
rect 20412 11788 20916 11844
rect 20188 8596 20244 8606
rect 20188 8484 20244 8540
rect 18620 6468 18676 6478
rect 19068 6468 19124 6636
rect 18620 6374 18676 6412
rect 18844 6466 19124 6468
rect 18844 6414 19070 6466
rect 19122 6414 19124 6466
rect 18844 6412 19124 6414
rect 18396 6078 18398 6130
rect 18450 6078 18452 6130
rect 18396 6066 18452 6078
rect 17724 5966 17726 6018
rect 17778 5966 17780 6018
rect 17724 5236 17780 5966
rect 17724 5170 17780 5180
rect 17836 6018 18340 6020
rect 17836 5966 18286 6018
rect 18338 5966 18340 6018
rect 17836 5964 18340 5966
rect 17724 5012 17780 5022
rect 17836 5012 17892 5964
rect 18284 5954 18340 5964
rect 18620 5908 18676 5918
rect 18844 5908 18900 6412
rect 19068 6402 19124 6412
rect 19180 8372 19348 8428
rect 20076 8428 20244 8484
rect 20076 8372 20132 8428
rect 19068 6132 19124 6142
rect 18676 5852 18900 5908
rect 18956 6130 19124 6132
rect 18956 6078 19070 6130
rect 19122 6078 19124 6130
rect 18956 6076 19124 6078
rect 18620 5814 18676 5852
rect 18732 5348 18788 5358
rect 17724 5010 17892 5012
rect 17724 4958 17726 5010
rect 17778 4958 17892 5010
rect 17724 4956 17892 4958
rect 18396 5010 18452 5022
rect 18396 4958 18398 5010
rect 18450 4958 18452 5010
rect 17724 4946 17780 4956
rect 16380 4620 16660 4676
rect 16380 4452 16436 4462
rect 16156 4450 16436 4452
rect 16156 4398 16382 4450
rect 16434 4398 16436 4450
rect 16156 4396 16436 4398
rect 16044 4228 16100 4238
rect 15820 4226 16100 4228
rect 15820 4174 16046 4226
rect 16098 4174 16100 4226
rect 15820 4172 16100 4174
rect 16044 4162 16100 4172
rect 15932 3668 15988 3678
rect 16156 3668 16212 4396
rect 16380 4386 16436 4396
rect 16604 4338 16660 4620
rect 16604 4286 16606 4338
rect 16658 4286 16660 4338
rect 16604 4274 16660 4286
rect 17500 4340 17556 4844
rect 18060 4898 18116 4910
rect 18060 4846 18062 4898
rect 18114 4846 18116 4898
rect 18060 4452 18116 4846
rect 18396 4564 18452 4958
rect 18396 4498 18452 4508
rect 18172 4452 18228 4462
rect 18060 4450 18228 4452
rect 18060 4398 18174 4450
rect 18226 4398 18228 4450
rect 18060 4396 18228 4398
rect 18172 4386 18228 4396
rect 17500 4246 17556 4284
rect 18284 4340 18340 4350
rect 15932 3666 16212 3668
rect 15932 3614 15934 3666
rect 15986 3614 16212 3666
rect 15932 3612 16212 3614
rect 18060 3668 18116 3678
rect 15932 3602 15988 3612
rect 18060 3574 18116 3612
rect 15148 3502 15150 3554
rect 15202 3502 15204 3554
rect 15148 3490 15204 3502
rect 14476 3388 14868 3444
rect 12124 3332 12516 3388
rect 11900 3276 12180 3332
rect 18284 2996 18340 4284
rect 18732 3666 18788 5292
rect 18732 3614 18734 3666
rect 18786 3614 18788 3666
rect 18732 3444 18788 3614
rect 18956 3668 19012 6076
rect 19068 6066 19124 6076
rect 19068 5010 19124 5022
rect 19068 4958 19070 5010
rect 19122 4958 19124 5010
rect 19068 4228 19124 4958
rect 19180 4900 19236 8372
rect 20076 8306 20132 8316
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19740 7474 19796 7486
rect 19740 7422 19742 7474
rect 19794 7422 19796 7474
rect 19404 7364 19460 7374
rect 19740 7364 19796 7422
rect 19404 7362 19796 7364
rect 19404 7310 19406 7362
rect 19458 7310 19796 7362
rect 19404 7308 19796 7310
rect 19404 6580 19460 7308
rect 20300 6692 20356 6702
rect 20300 6598 20356 6636
rect 19404 6514 19460 6524
rect 19516 6468 19572 6478
rect 19292 6130 19348 6142
rect 19292 6078 19294 6130
rect 19346 6078 19348 6130
rect 19292 6018 19348 6078
rect 19292 5966 19294 6018
rect 19346 5966 19348 6018
rect 19292 5954 19348 5966
rect 19516 6020 19572 6412
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20412 6244 20468 11788
rect 21868 11506 21924 12124
rect 21868 11454 21870 11506
rect 21922 11454 21924 11506
rect 21868 11442 21924 11454
rect 21980 12066 22036 13692
rect 22316 13682 22372 13692
rect 22428 12852 22484 14476
rect 22540 14418 22596 14588
rect 22540 14366 22542 14418
rect 22594 14366 22596 14418
rect 22540 13970 22596 14366
rect 22652 14306 22708 15260
rect 22652 14254 22654 14306
rect 22706 14254 22708 14306
rect 22652 14242 22708 14254
rect 23212 14644 23268 18620
rect 23436 18452 23492 19070
rect 23548 18452 23604 18462
rect 23436 18396 23548 18452
rect 23548 18358 23604 18396
rect 23660 17108 23716 21196
rect 23772 21028 23828 21038
rect 23772 18676 23828 20972
rect 23884 20916 23940 20926
rect 23884 20822 23940 20860
rect 23996 20580 24052 21420
rect 24108 20916 24164 21756
rect 24220 21810 24388 21812
rect 24220 21758 24222 21810
rect 24274 21758 24388 21810
rect 24220 21756 24388 21758
rect 24220 21746 24276 21756
rect 24108 20802 24164 20860
rect 24108 20750 24110 20802
rect 24162 20750 24164 20802
rect 24108 20738 24164 20750
rect 23996 20514 24052 20524
rect 23996 20020 24052 20030
rect 23996 19926 24052 19964
rect 24332 19348 24388 19358
rect 24444 19348 24500 28476
rect 24668 27972 24724 27982
rect 24668 27746 24724 27916
rect 24668 27694 24670 27746
rect 24722 27694 24724 27746
rect 24668 27188 24724 27694
rect 24668 27122 24724 27132
rect 24556 27074 24612 27086
rect 24556 27022 24558 27074
rect 24610 27022 24612 27074
rect 24556 26852 24612 27022
rect 24780 26908 24836 39004
rect 25452 38500 25508 44492
rect 25676 44434 25732 44604
rect 25676 44382 25678 44434
rect 25730 44382 25732 44434
rect 25676 44370 25732 44382
rect 25676 42980 25732 42990
rect 25452 38434 25508 38444
rect 25564 42978 25732 42980
rect 25564 42926 25678 42978
rect 25730 42926 25732 42978
rect 25564 42924 25732 42926
rect 25564 41410 25620 42924
rect 25676 42914 25732 42924
rect 25564 41358 25566 41410
rect 25618 41358 25620 41410
rect 25564 37380 25620 41358
rect 25788 41300 25844 41310
rect 25788 39620 25844 41244
rect 25900 39844 25956 45052
rect 26684 44996 26740 45054
rect 26684 44930 26740 44940
rect 26012 44882 26068 44894
rect 26012 44830 26014 44882
rect 26066 44830 26068 44882
rect 26012 44212 26068 44830
rect 26236 44660 26292 44670
rect 26124 44212 26180 44222
rect 26012 44156 26124 44212
rect 26124 44118 26180 44156
rect 26236 44210 26292 44604
rect 26236 44158 26238 44210
rect 26290 44158 26292 44210
rect 26236 44146 26292 44158
rect 26684 44212 26740 44222
rect 26460 44100 26516 44110
rect 26460 44006 26516 44044
rect 26684 44100 26740 44156
rect 26796 44100 26852 45276
rect 26908 45266 26964 45276
rect 27132 45266 27188 45276
rect 27132 44996 27188 45006
rect 26684 44098 26852 44100
rect 26684 44046 26798 44098
rect 26850 44046 26852 44098
rect 26684 44044 26852 44046
rect 26572 42978 26628 42990
rect 26572 42926 26574 42978
rect 26626 42926 26628 42978
rect 26572 42866 26628 42926
rect 26572 42814 26574 42866
rect 26626 42814 26628 42866
rect 26572 42802 26628 42814
rect 26012 42530 26068 42542
rect 26012 42478 26014 42530
rect 26066 42478 26068 42530
rect 26012 42196 26068 42478
rect 26012 42130 26068 42140
rect 26012 41858 26068 41870
rect 26012 41806 26014 41858
rect 26066 41806 26068 41858
rect 26012 40964 26068 41806
rect 26348 40964 26404 40974
rect 26012 40898 26068 40908
rect 26124 40962 26404 40964
rect 26124 40910 26350 40962
rect 26402 40910 26404 40962
rect 26124 40908 26404 40910
rect 25900 39788 26068 39844
rect 25900 39620 25956 39630
rect 25788 39618 25956 39620
rect 25788 39566 25902 39618
rect 25954 39566 25956 39618
rect 25788 39564 25956 39566
rect 25900 39554 25956 39564
rect 26012 39284 26068 39788
rect 26124 39620 26180 40908
rect 26348 40898 26404 40908
rect 26460 40852 26516 40862
rect 26460 40514 26516 40796
rect 26460 40462 26462 40514
rect 26514 40462 26516 40514
rect 26460 40450 26516 40462
rect 26124 39526 26180 39564
rect 26236 39508 26292 39518
rect 26236 39414 26292 39452
rect 26348 39394 26404 39406
rect 26348 39342 26350 39394
rect 26402 39342 26404 39394
rect 26348 39284 26404 39342
rect 25452 37324 25564 37380
rect 25340 37156 25396 37166
rect 25452 37156 25508 37324
rect 25564 37286 25620 37324
rect 25676 39228 26404 39284
rect 26460 39394 26516 39406
rect 26460 39342 26462 39394
rect 26514 39342 26516 39394
rect 25340 37154 25508 37156
rect 25340 37102 25342 37154
rect 25394 37102 25508 37154
rect 25340 37100 25508 37102
rect 25564 37156 25620 37166
rect 25340 37044 25396 37100
rect 25116 36988 25396 37044
rect 24892 36708 24948 36718
rect 25116 36708 25172 36988
rect 24892 36706 25172 36708
rect 24892 36654 24894 36706
rect 24946 36654 25172 36706
rect 24892 36652 25172 36654
rect 24892 36642 24948 36652
rect 25116 36482 25172 36494
rect 25116 36430 25118 36482
rect 25170 36430 25172 36482
rect 25116 36372 25172 36430
rect 25564 36482 25620 37100
rect 25564 36430 25566 36482
rect 25618 36430 25620 36482
rect 25564 36418 25620 36430
rect 25116 35588 25172 36316
rect 25564 35588 25620 35598
rect 25116 35586 25620 35588
rect 25116 35534 25566 35586
rect 25618 35534 25620 35586
rect 25116 35532 25620 35534
rect 25228 33906 25284 33918
rect 25228 33854 25230 33906
rect 25282 33854 25284 33906
rect 25004 33348 25060 33358
rect 24892 33124 24948 33134
rect 25004 33124 25060 33292
rect 25228 33346 25284 33854
rect 25228 33294 25230 33346
rect 25282 33294 25284 33346
rect 25228 33282 25284 33294
rect 24892 33122 25060 33124
rect 24892 33070 24894 33122
rect 24946 33070 25060 33122
rect 24892 33068 25060 33070
rect 24892 33058 24948 33068
rect 24556 26786 24612 26796
rect 24668 26852 24836 26908
rect 25004 32004 25060 33068
rect 25228 32562 25284 32574
rect 25228 32510 25230 32562
rect 25282 32510 25284 32562
rect 25228 32452 25284 32510
rect 25228 32386 25284 32396
rect 24556 26068 24612 26078
rect 24556 25618 24612 26012
rect 24556 25566 24558 25618
rect 24610 25566 24612 25618
rect 24556 25554 24612 25566
rect 24668 25396 24724 26852
rect 25004 26740 25060 31948
rect 25452 31332 25508 35532
rect 25564 35522 25620 35532
rect 25676 34244 25732 39228
rect 26460 39172 26516 39342
rect 26460 39106 26516 39116
rect 26460 38946 26516 38958
rect 26460 38894 26462 38946
rect 26514 38894 26516 38946
rect 26460 38836 26516 38894
rect 26460 38770 26516 38780
rect 26348 38722 26404 38734
rect 26348 38670 26350 38722
rect 26402 38670 26404 38722
rect 26348 38668 26404 38670
rect 26124 38612 26404 38668
rect 26124 37490 26180 38612
rect 26124 37438 26126 37490
rect 26178 37438 26180 37490
rect 26124 37426 26180 37438
rect 26572 37940 26628 37950
rect 26348 37378 26404 37390
rect 26348 37326 26350 37378
rect 26402 37326 26404 37378
rect 25900 37154 25956 37166
rect 25900 37102 25902 37154
rect 25954 37102 25956 37154
rect 25900 36932 25956 37102
rect 25788 36484 25844 36494
rect 25788 36390 25844 36428
rect 25900 36372 25956 36876
rect 26348 36932 26404 37326
rect 26348 36866 26404 36876
rect 26460 37266 26516 37278
rect 26460 37214 26462 37266
rect 26514 37214 26516 37266
rect 26460 36708 26516 37214
rect 26124 36596 26180 36606
rect 26124 36502 26180 36540
rect 26460 36484 26516 36652
rect 26460 36418 26516 36428
rect 25900 36306 25956 36316
rect 26124 36372 26180 36382
rect 26124 36278 26180 36316
rect 26572 36372 26628 37884
rect 26684 36484 26740 44044
rect 26796 44034 26852 44044
rect 27020 44884 27076 44894
rect 27020 43988 27076 44828
rect 27020 43922 27076 43932
rect 27020 43428 27076 43438
rect 26908 43372 27020 43428
rect 26796 41188 26852 41198
rect 26796 41094 26852 41132
rect 26908 41186 26964 43372
rect 27020 43362 27076 43372
rect 27132 42642 27188 44940
rect 27244 44994 27300 45724
rect 27356 45220 27412 45230
rect 27356 45106 27412 45164
rect 27356 45054 27358 45106
rect 27410 45054 27412 45106
rect 27356 45042 27412 45054
rect 27244 44942 27246 44994
rect 27298 44942 27300 44994
rect 27244 44930 27300 44942
rect 27356 44548 27412 44558
rect 27356 44434 27412 44492
rect 27356 44382 27358 44434
rect 27410 44382 27412 44434
rect 27356 43540 27412 44382
rect 27468 44436 27524 48524
rect 27580 48354 27636 48366
rect 27580 48302 27582 48354
rect 27634 48302 27636 48354
rect 27580 47348 27636 48302
rect 27580 47282 27636 47292
rect 27692 45668 27748 45678
rect 27692 44996 27748 45612
rect 27692 44902 27748 44940
rect 27804 44772 27860 50372
rect 28028 49252 28084 50764
rect 28252 51604 28308 53004
rect 28252 50708 28308 51548
rect 28252 50614 28308 50652
rect 28364 50428 28420 62132
rect 28476 58212 28532 58222
rect 28476 57204 28532 58156
rect 28476 57138 28532 57148
rect 28588 57538 28644 57550
rect 28588 57486 28590 57538
rect 28642 57486 28644 57538
rect 28588 54628 28644 57486
rect 28476 54572 28644 54628
rect 28476 54180 28532 54572
rect 28812 54516 28868 73166
rect 29148 73218 29204 73230
rect 29148 73166 29150 73218
rect 29202 73166 29204 73218
rect 29036 70196 29092 70206
rect 29036 70102 29092 70140
rect 29148 70084 29204 73166
rect 29260 72324 29316 72334
rect 29260 72230 29316 72268
rect 29484 71090 29540 73892
rect 29820 73892 29876 74844
rect 30828 74788 30884 75628
rect 31276 75682 31332 76188
rect 33180 76354 33236 76366
rect 33180 76302 33182 76354
rect 33234 76302 33236 76354
rect 33180 76244 33236 76302
rect 33180 76178 33236 76188
rect 33628 76242 33684 76254
rect 33628 76190 33630 76242
rect 33682 76190 33684 76242
rect 33628 76020 33684 76190
rect 33964 76244 34020 76412
rect 33964 76178 34020 76188
rect 34748 76354 34804 76366
rect 36876 76356 36932 76366
rect 34748 76302 34750 76354
rect 34802 76302 34804 76354
rect 33628 75964 34356 76020
rect 34188 75796 34244 75806
rect 33516 75794 34244 75796
rect 33516 75742 34190 75794
rect 34242 75742 34244 75794
rect 33516 75740 34244 75742
rect 34300 75796 34356 75964
rect 34300 75740 34692 75796
rect 31276 75630 31278 75682
rect 31330 75630 31332 75682
rect 31276 75618 31332 75630
rect 32060 75684 32116 75694
rect 32060 75590 32116 75628
rect 30940 74788 30996 74798
rect 30828 74786 30996 74788
rect 30828 74734 30942 74786
rect 30994 74734 30996 74786
rect 30828 74732 30996 74734
rect 30268 74002 30324 74014
rect 30268 73950 30270 74002
rect 30322 73950 30324 74002
rect 29932 73892 29988 73902
rect 30268 73892 30324 73950
rect 30380 74004 30436 74014
rect 30940 74004 30996 74732
rect 32508 74788 32564 74798
rect 32508 74694 32564 74732
rect 33404 74788 33460 74798
rect 33404 74694 33460 74732
rect 33516 74226 33572 75740
rect 34188 75730 34244 75740
rect 33628 75572 33684 75582
rect 33684 75516 33796 75572
rect 33628 75506 33684 75516
rect 33628 75012 33684 75022
rect 33628 74918 33684 74956
rect 33740 74786 33796 75516
rect 33740 74734 33742 74786
rect 33794 74734 33796 74786
rect 33740 74722 33796 74734
rect 34188 74788 34244 74798
rect 33516 74174 33518 74226
rect 33570 74174 33572 74226
rect 33516 74162 33572 74174
rect 33964 74674 34020 74686
rect 33964 74622 33966 74674
rect 34018 74622 34020 74674
rect 33404 74004 33460 74014
rect 30940 73948 31444 74004
rect 30380 73910 30436 73948
rect 29820 73890 30324 73892
rect 29820 73838 29934 73890
rect 29986 73838 30324 73890
rect 29820 73836 30324 73838
rect 30604 73890 30660 73902
rect 30604 73838 30606 73890
rect 30658 73838 30660 73890
rect 29820 72324 29876 73836
rect 29932 73826 29988 73836
rect 30604 73444 30660 73838
rect 31276 73444 31332 73454
rect 30604 73442 31332 73444
rect 30604 73390 31278 73442
rect 31330 73390 31332 73442
rect 30604 73388 31332 73390
rect 31276 73378 31332 73388
rect 30044 73220 30100 73230
rect 30044 72546 30100 73164
rect 30380 72548 30436 72558
rect 30044 72494 30046 72546
rect 30098 72494 30100 72546
rect 30044 72482 30100 72494
rect 30156 72546 30436 72548
rect 30156 72494 30382 72546
rect 30434 72494 30436 72546
rect 30156 72492 30436 72494
rect 30156 72324 30212 72492
rect 30380 72482 30436 72492
rect 30828 72548 30884 72558
rect 29820 72322 30212 72324
rect 29820 72270 29822 72322
rect 29874 72270 30212 72322
rect 29820 72268 30212 72270
rect 30268 72324 30324 72334
rect 29820 72258 29876 72268
rect 30268 72230 30324 72268
rect 29484 71038 29486 71090
rect 29538 71038 29540 71090
rect 29484 70196 29540 71038
rect 29484 70130 29540 70140
rect 29932 70196 29988 70206
rect 29932 70102 29988 70140
rect 29260 70084 29316 70094
rect 29148 70082 29316 70084
rect 29148 70030 29262 70082
rect 29314 70030 29316 70082
rect 29148 70028 29316 70030
rect 29260 69972 29316 70028
rect 29260 68404 29316 69916
rect 29708 70084 29764 70094
rect 29596 69410 29652 69422
rect 29596 69358 29598 69410
rect 29650 69358 29652 69410
rect 29596 69188 29652 69358
rect 29596 69122 29652 69132
rect 29708 68516 29764 70028
rect 30716 70082 30772 70094
rect 30716 70030 30718 70082
rect 30770 70030 30772 70082
rect 30268 69972 30324 69982
rect 30716 69972 30772 70030
rect 30268 69970 30660 69972
rect 30268 69918 30270 69970
rect 30322 69918 30660 69970
rect 30268 69916 30660 69918
rect 30268 69906 30324 69916
rect 30380 69298 30436 69310
rect 30380 69246 30382 69298
rect 30434 69246 30436 69298
rect 30380 68852 30436 69246
rect 30492 68852 30548 68862
rect 30380 68850 30548 68852
rect 30380 68798 30494 68850
rect 30546 68798 30548 68850
rect 30380 68796 30548 68798
rect 30492 68786 30548 68796
rect 30604 68628 30660 69916
rect 30716 69906 30772 69916
rect 30828 69188 30884 72492
rect 30828 69122 30884 69132
rect 31164 70196 31220 70206
rect 30716 68628 30772 68638
rect 30604 68626 30772 68628
rect 30604 68574 30718 68626
rect 30770 68574 30772 68626
rect 30604 68572 30772 68574
rect 30716 68562 30772 68572
rect 30156 68516 30212 68526
rect 29708 68514 30212 68516
rect 29708 68462 30158 68514
rect 30210 68462 30212 68514
rect 29708 68460 30212 68462
rect 29260 68348 29876 68404
rect 29372 64706 29428 64718
rect 29372 64654 29374 64706
rect 29426 64654 29428 64706
rect 29372 62356 29428 64654
rect 29372 62290 29428 62300
rect 29148 62242 29204 62254
rect 29148 62190 29150 62242
rect 29202 62190 29204 62242
rect 29148 62188 29204 62190
rect 29148 62132 29764 62188
rect 29708 61458 29764 62132
rect 29708 61406 29710 61458
rect 29762 61406 29764 61458
rect 29708 61394 29764 61406
rect 29148 59220 29204 59230
rect 29148 58658 29204 59164
rect 29148 58606 29150 58658
rect 29202 58606 29204 58658
rect 29148 58594 29204 58606
rect 29260 59106 29316 59118
rect 29260 59054 29262 59106
rect 29314 59054 29316 59106
rect 29260 58660 29316 59054
rect 29260 58604 29652 58660
rect 29484 58434 29540 58446
rect 29484 58382 29486 58434
rect 29538 58382 29540 58434
rect 29484 58212 29540 58382
rect 29596 58436 29652 58604
rect 29708 58436 29764 58446
rect 29596 58434 29764 58436
rect 29596 58382 29710 58434
rect 29762 58382 29764 58434
rect 29596 58380 29764 58382
rect 29484 57988 29540 58156
rect 29036 57932 29540 57988
rect 28812 54450 28868 54460
rect 28924 54514 28980 54526
rect 28924 54462 28926 54514
rect 28978 54462 28980 54514
rect 28588 54404 28644 54414
rect 28588 54310 28644 54348
rect 28924 54404 28980 54462
rect 28924 54338 28980 54348
rect 28476 54124 28756 54180
rect 28588 53732 28644 53742
rect 28588 53638 28644 53676
rect 28588 52948 28644 52958
rect 28588 52854 28644 52892
rect 28700 50428 28756 54124
rect 29036 53508 29092 57932
rect 29708 57428 29764 58380
rect 29484 57372 29764 57428
rect 29260 54626 29316 54638
rect 29260 54574 29262 54626
rect 29314 54574 29316 54626
rect 29036 53442 29092 53452
rect 29148 53618 29204 53630
rect 29148 53566 29150 53618
rect 29202 53566 29204 53618
rect 29148 52836 29204 53566
rect 29260 53058 29316 54574
rect 29372 53732 29428 53742
rect 29372 53638 29428 53676
rect 29484 53508 29540 57372
rect 29820 57316 29876 68348
rect 29260 53006 29262 53058
rect 29314 53006 29316 53058
rect 29260 52994 29316 53006
rect 29372 53452 29540 53508
rect 29596 57260 29876 57316
rect 28924 52276 28980 52286
rect 28924 50484 28980 52220
rect 28364 50372 28532 50428
rect 28700 50372 28868 50428
rect 28028 49158 28084 49196
rect 28252 49924 28308 49934
rect 28252 49138 28308 49868
rect 28252 49086 28254 49138
rect 28306 49086 28308 49138
rect 28252 49074 28308 49086
rect 28364 48244 28420 48254
rect 28364 48150 28420 48188
rect 27916 47458 27972 47470
rect 28140 47460 28196 47470
rect 27916 47406 27918 47458
rect 27970 47406 27972 47458
rect 27916 47124 27972 47406
rect 27916 45106 27972 47068
rect 27916 45054 27918 45106
rect 27970 45054 27972 45106
rect 27916 44884 27972 45054
rect 27916 44818 27972 44828
rect 28028 47404 28140 47460
rect 28028 45218 28084 47404
rect 28140 47394 28196 47404
rect 28140 46788 28196 46798
rect 28140 46694 28196 46732
rect 28028 45166 28030 45218
rect 28082 45166 28084 45218
rect 27580 44716 27860 44772
rect 27580 44548 27636 44716
rect 28028 44660 28084 45166
rect 28028 44594 28084 44604
rect 28140 45666 28196 45678
rect 28140 45614 28142 45666
rect 28194 45614 28196 45666
rect 28140 45444 28196 45614
rect 27580 44492 27972 44548
rect 27468 44370 27524 44380
rect 27356 43474 27412 43484
rect 27580 43988 27636 43998
rect 27244 43428 27300 43438
rect 27244 42754 27300 43372
rect 27244 42702 27246 42754
rect 27298 42702 27300 42754
rect 27244 42690 27300 42702
rect 27132 42590 27134 42642
rect 27186 42590 27188 42642
rect 27132 42084 27188 42590
rect 27356 42644 27412 42654
rect 27356 42642 27524 42644
rect 27356 42590 27358 42642
rect 27410 42590 27524 42642
rect 27356 42588 27524 42590
rect 27356 42578 27412 42588
rect 27132 42018 27188 42028
rect 26908 41134 26910 41186
rect 26962 41134 26964 41186
rect 26908 41122 26964 41134
rect 27020 41860 27076 41870
rect 27020 41074 27076 41804
rect 27468 41412 27524 42588
rect 27468 41318 27524 41356
rect 27580 41636 27636 43932
rect 27804 43876 27860 43886
rect 27804 42980 27860 43820
rect 27020 41022 27022 41074
rect 27074 41022 27076 41074
rect 26908 40740 26964 40750
rect 26908 40402 26964 40684
rect 26908 40350 26910 40402
rect 26962 40350 26964 40402
rect 26908 40338 26964 40350
rect 26908 39508 26964 39518
rect 26796 38946 26852 38958
rect 26796 38894 26798 38946
rect 26850 38894 26852 38946
rect 26796 38164 26852 38894
rect 26908 38834 26964 39452
rect 26908 38782 26910 38834
rect 26962 38782 26964 38834
rect 26908 38770 26964 38782
rect 27020 38668 27076 41022
rect 27580 41074 27636 41580
rect 27580 41022 27582 41074
rect 27634 41022 27636 41074
rect 27580 41010 27636 41022
rect 27692 42978 27860 42980
rect 27692 42926 27806 42978
rect 27858 42926 27860 42978
rect 27692 42924 27860 42926
rect 27468 40516 27524 40526
rect 27356 40404 27412 40414
rect 27356 40310 27412 40348
rect 27244 39620 27300 39630
rect 27244 39526 27300 39564
rect 27356 39508 27412 39518
rect 27468 39508 27524 40460
rect 27356 39506 27524 39508
rect 27356 39454 27358 39506
rect 27410 39454 27524 39506
rect 27356 39452 27524 39454
rect 27580 39508 27636 39518
rect 27356 39442 27412 39452
rect 27580 39414 27636 39452
rect 27356 38836 27412 38846
rect 27692 38836 27748 42924
rect 27804 42914 27860 42924
rect 27804 41412 27860 41422
rect 27804 40628 27860 41356
rect 27804 40562 27860 40572
rect 27356 38742 27412 38780
rect 27468 38780 27748 38836
rect 26796 38098 26852 38108
rect 26908 38612 27076 38668
rect 26908 36820 26964 38612
rect 27356 38500 27412 38510
rect 27132 38444 27356 38500
rect 27020 37492 27076 37502
rect 27020 37398 27076 37436
rect 26908 36764 27076 36820
rect 26908 36596 26964 36606
rect 26684 36428 26852 36484
rect 26012 36258 26068 36270
rect 26572 36260 26628 36316
rect 26684 36260 26740 36270
rect 26012 36206 26014 36258
rect 26066 36206 26068 36258
rect 25788 36148 25844 36158
rect 25788 35364 25844 36092
rect 25788 35026 25844 35308
rect 25788 34974 25790 35026
rect 25842 34974 25844 35026
rect 25788 34962 25844 34974
rect 25900 35588 25956 35598
rect 25788 34244 25844 34254
rect 25676 34242 25844 34244
rect 25676 34190 25790 34242
rect 25842 34190 25844 34242
rect 25676 34188 25844 34190
rect 25788 34178 25844 34188
rect 25564 33906 25620 33918
rect 25564 33854 25566 33906
rect 25618 33854 25620 33906
rect 25564 33348 25620 33854
rect 25900 33796 25956 35532
rect 26012 34020 26068 36206
rect 26460 36258 26740 36260
rect 26460 36206 26686 36258
rect 26738 36206 26740 36258
rect 26460 36204 26740 36206
rect 26236 36036 26292 36046
rect 26460 36036 26516 36204
rect 26684 36194 26740 36204
rect 26124 34356 26180 34366
rect 26236 34356 26292 35980
rect 26124 34354 26292 34356
rect 26124 34302 26126 34354
rect 26178 34302 26292 34354
rect 26124 34300 26292 34302
rect 26124 34290 26180 34300
rect 26012 33954 26068 33964
rect 25900 33740 26180 33796
rect 25564 33282 25620 33292
rect 25564 33124 25620 33134
rect 25564 33122 26068 33124
rect 25564 33070 25566 33122
rect 25618 33070 26068 33122
rect 25564 33068 26068 33070
rect 25564 33058 25620 33068
rect 26012 32674 26068 33068
rect 26124 33122 26180 33740
rect 26124 33070 26126 33122
rect 26178 33070 26180 33122
rect 26124 32900 26180 33070
rect 26124 32834 26180 32844
rect 26012 32622 26014 32674
rect 26066 32622 26068 32674
rect 26012 32610 26068 32622
rect 25900 32564 25956 32574
rect 25788 32508 25900 32564
rect 25676 31666 25732 31678
rect 25676 31614 25678 31666
rect 25730 31614 25732 31666
rect 25564 31332 25620 31342
rect 25452 31276 25564 31332
rect 25564 31266 25620 31276
rect 25228 30884 25284 30894
rect 25228 30324 25284 30828
rect 25676 30548 25732 31614
rect 25676 30482 25732 30492
rect 25788 30436 25844 32508
rect 25900 32498 25956 32508
rect 26236 32116 26292 34300
rect 26012 32060 26292 32116
rect 26348 35980 26516 36036
rect 25900 31556 25956 31566
rect 26012 31556 26068 32060
rect 26236 31892 26292 31902
rect 26236 31798 26292 31836
rect 26124 31780 26180 31790
rect 26124 31686 26180 31724
rect 26236 31556 26292 31566
rect 26012 31554 26292 31556
rect 26012 31502 26238 31554
rect 26290 31502 26292 31554
rect 26012 31500 26292 31502
rect 25900 31462 25956 31500
rect 26236 31490 26292 31500
rect 26348 30884 26404 35980
rect 26460 35364 26516 35374
rect 26460 34130 26516 35308
rect 26460 34078 26462 34130
rect 26514 34078 26516 34130
rect 26460 33460 26516 34078
rect 26684 34018 26740 34030
rect 26684 33966 26686 34018
rect 26738 33966 26740 34018
rect 26684 33908 26740 33966
rect 26572 33460 26628 33470
rect 26460 33404 26572 33460
rect 26572 33366 26628 33404
rect 26684 32116 26740 33852
rect 26796 32564 26852 36428
rect 26908 36482 26964 36540
rect 26908 36430 26910 36482
rect 26962 36430 26964 36482
rect 26908 36418 26964 36430
rect 27020 35812 27076 36764
rect 27020 35746 27076 35756
rect 27020 34690 27076 34702
rect 27020 34638 27022 34690
rect 27074 34638 27076 34690
rect 27020 34468 27076 34638
rect 27020 34402 27076 34412
rect 27132 34244 27188 38444
rect 27356 38434 27412 38444
rect 27244 38164 27300 38174
rect 27244 38070 27300 38108
rect 27468 38052 27524 38780
rect 27916 38668 27972 44492
rect 28028 44436 28084 44446
rect 28028 44342 28084 44380
rect 28028 43540 28084 43550
rect 28028 41412 28084 43484
rect 28140 42196 28196 45388
rect 28252 45332 28308 45342
rect 28252 45106 28308 45276
rect 28252 45054 28254 45106
rect 28306 45054 28308 45106
rect 28252 43428 28308 45054
rect 28364 45220 28420 45230
rect 28364 44996 28420 45164
rect 28364 44322 28420 44940
rect 28364 44270 28366 44322
rect 28418 44270 28420 44322
rect 28364 44258 28420 44270
rect 28476 44212 28532 50372
rect 28588 49924 28644 49934
rect 28588 49698 28644 49868
rect 28588 49646 28590 49698
rect 28642 49646 28644 49698
rect 28588 49634 28644 49646
rect 28588 48244 28644 48254
rect 28644 48188 28756 48244
rect 28588 48178 28644 48188
rect 28588 47460 28644 47470
rect 28588 47366 28644 47404
rect 28700 47068 28756 48188
rect 28588 47012 28756 47068
rect 28588 46898 28644 47012
rect 28588 46846 28590 46898
rect 28642 46846 28644 46898
rect 28588 46834 28644 46846
rect 28588 46004 28644 46014
rect 28588 45666 28644 45948
rect 28588 45614 28590 45666
rect 28642 45614 28644 45666
rect 28588 45108 28644 45614
rect 28812 45556 28868 50372
rect 28924 48356 28980 50428
rect 28924 48290 28980 48300
rect 29036 50260 29092 50270
rect 28812 45490 28868 45500
rect 28924 48132 28980 48142
rect 28924 45332 28980 48076
rect 29036 46900 29092 50204
rect 29148 47012 29204 52780
rect 29372 50482 29428 53452
rect 29484 50708 29540 50718
rect 29484 50614 29540 50652
rect 29372 50430 29374 50482
rect 29426 50430 29428 50482
rect 29372 50418 29428 50430
rect 29260 49252 29316 49262
rect 29260 49138 29316 49196
rect 29260 49086 29262 49138
rect 29314 49086 29316 49138
rect 29260 49074 29316 49086
rect 29596 48356 29652 57260
rect 29932 57092 29988 68460
rect 30156 68450 30212 68460
rect 30492 65602 30548 65614
rect 30492 65550 30494 65602
rect 30546 65550 30548 65602
rect 30156 64820 30212 64830
rect 30492 64820 30548 65550
rect 30156 64818 30548 64820
rect 30156 64766 30158 64818
rect 30210 64766 30548 64818
rect 30156 64764 30548 64766
rect 30604 65492 30660 65502
rect 30156 64754 30212 64764
rect 30604 64148 30660 65436
rect 30828 65492 30884 65502
rect 30828 65490 30996 65492
rect 30828 65438 30830 65490
rect 30882 65438 30996 65490
rect 30828 65436 30996 65438
rect 30828 65426 30884 65436
rect 30268 64092 30604 64148
rect 30044 62914 30100 62926
rect 30044 62862 30046 62914
rect 30098 62862 30100 62914
rect 30044 61570 30100 62862
rect 30044 61518 30046 61570
rect 30098 61518 30100 61570
rect 30044 61506 30100 61518
rect 29820 57036 29988 57092
rect 30044 58994 30100 59006
rect 30044 58942 30046 58994
rect 30098 58942 30100 58994
rect 29820 56980 29876 57036
rect 29708 56924 29876 56980
rect 29708 56308 29764 56924
rect 29820 56756 29876 56766
rect 30044 56756 30100 58942
rect 30268 58884 30324 64092
rect 30604 64054 30660 64092
rect 30940 64146 30996 65436
rect 30940 64094 30942 64146
rect 30994 64094 30996 64146
rect 30940 64082 30996 64094
rect 30156 58828 30324 58884
rect 30380 63420 30772 63476
rect 30380 63362 30436 63420
rect 30380 63310 30382 63362
rect 30434 63310 30436 63362
rect 30380 58994 30436 63310
rect 30604 63252 30660 63262
rect 30716 63252 30772 63420
rect 31052 63252 31108 63262
rect 31164 63252 31220 70140
rect 31276 64148 31332 64158
rect 31276 63922 31332 64092
rect 31276 63870 31278 63922
rect 31330 63870 31332 63922
rect 31276 63858 31332 63870
rect 30716 63250 31220 63252
rect 30716 63198 31054 63250
rect 31106 63198 31220 63250
rect 30716 63196 31220 63198
rect 30604 63158 30660 63196
rect 31052 63186 31108 63196
rect 31276 62242 31332 62254
rect 31276 62190 31278 62242
rect 31330 62190 31332 62242
rect 31276 62188 31332 62190
rect 30380 58942 30382 58994
rect 30434 58942 30436 58994
rect 30156 58212 30212 58828
rect 30156 58118 30212 58156
rect 30380 58100 30436 58942
rect 30604 62132 31332 62188
rect 30604 59330 30660 62132
rect 31388 60564 31444 73948
rect 33460 73948 33684 74004
rect 33964 73948 34020 74622
rect 34188 74004 34244 74732
rect 34300 74004 34356 74014
rect 34188 73948 34300 74004
rect 33404 73910 33460 73948
rect 33628 73892 33796 73948
rect 31948 73330 32004 73342
rect 31948 73278 31950 73330
rect 32002 73278 32004 73330
rect 31500 72434 31556 72446
rect 31500 72382 31502 72434
rect 31554 72382 31556 72434
rect 31500 71988 31556 72382
rect 31948 72436 32004 73278
rect 33180 73220 33236 73230
rect 33180 73218 33684 73220
rect 33180 73166 33182 73218
rect 33234 73166 33684 73218
rect 33180 73164 33684 73166
rect 33180 73154 33236 73164
rect 33068 73108 33124 73118
rect 31948 72370 32004 72380
rect 32956 73106 33124 73108
rect 32956 73054 33070 73106
rect 33122 73054 33124 73106
rect 32956 73052 33124 73054
rect 31500 71922 31556 71932
rect 32956 72324 33012 73052
rect 33068 73042 33124 73052
rect 33628 72658 33684 73164
rect 33628 72606 33630 72658
rect 33682 72606 33684 72658
rect 33628 72594 33684 72606
rect 32844 71764 32900 71774
rect 32508 71652 32564 71662
rect 32508 71558 32564 71596
rect 32844 70978 32900 71708
rect 32956 71090 33012 72268
rect 33180 71988 33236 71998
rect 33180 71894 33236 71932
rect 33404 71762 33460 71774
rect 33404 71710 33406 71762
rect 33458 71710 33460 71762
rect 33068 71652 33124 71662
rect 33068 71558 33124 71596
rect 33404 71652 33460 71710
rect 33404 71586 33460 71596
rect 32956 71038 32958 71090
rect 33010 71038 33012 71090
rect 32956 71026 33012 71038
rect 32844 70926 32846 70978
rect 32898 70926 32900 70978
rect 32844 70914 32900 70926
rect 33628 70980 33684 70990
rect 33740 70980 33796 73892
rect 33852 73892 34020 73948
rect 34300 73938 34356 73948
rect 34412 73948 34468 75740
rect 34524 75570 34580 75582
rect 34524 75518 34526 75570
rect 34578 75518 34580 75570
rect 34524 74788 34580 75518
rect 34636 75572 34692 75740
rect 34748 75794 34804 76302
rect 36428 76354 36932 76356
rect 36428 76302 36878 76354
rect 36930 76302 36932 76354
rect 36428 76300 36932 76302
rect 34748 75742 34750 75794
rect 34802 75742 34804 75794
rect 34748 75730 34804 75742
rect 34972 76244 35028 76254
rect 34748 75572 34804 75582
rect 34636 75570 34804 75572
rect 34636 75518 34750 75570
rect 34802 75518 34804 75570
rect 34636 75516 34804 75518
rect 34748 75506 34804 75516
rect 34972 75348 35028 76188
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 36428 75794 36484 76300
rect 36876 76290 36932 76300
rect 36428 75742 36430 75794
rect 36482 75742 36484 75794
rect 36428 75730 36484 75742
rect 35308 75684 35364 75694
rect 35196 75682 35364 75684
rect 35196 75630 35310 75682
rect 35362 75630 35364 75682
rect 35196 75628 35364 75630
rect 35196 75348 35252 75628
rect 35308 75618 35364 75628
rect 34972 75292 35252 75348
rect 36316 75458 36372 75470
rect 36316 75406 36318 75458
rect 36370 75406 36372 75458
rect 34972 75012 35028 75292
rect 35196 75012 35252 75022
rect 34524 74722 34580 74732
rect 34636 74956 35028 75012
rect 34636 74786 34692 74956
rect 34972 74898 35028 74956
rect 34972 74846 34974 74898
rect 35026 74846 35028 74898
rect 34972 74834 35028 74846
rect 35084 74956 35196 75012
rect 34636 74734 34638 74786
rect 34690 74734 34692 74786
rect 34636 74674 34692 74734
rect 34636 74622 34638 74674
rect 34690 74622 34692 74674
rect 34636 74610 34692 74622
rect 34412 73892 34580 73948
rect 33852 73218 33908 73892
rect 33852 73166 33854 73218
rect 33906 73166 33908 73218
rect 33852 72548 33908 73166
rect 33852 72482 33908 72492
rect 34300 72324 34356 72334
rect 34300 72322 34468 72324
rect 34300 72270 34302 72322
rect 34354 72270 34468 72322
rect 34300 72268 34468 72270
rect 34300 72258 34356 72268
rect 34412 71764 34468 72268
rect 34412 71698 34468 71708
rect 33628 70978 33796 70980
rect 33628 70926 33630 70978
rect 33682 70926 33796 70978
rect 33628 70924 33796 70926
rect 33852 71652 33908 71662
rect 34300 71652 34356 71662
rect 33852 71650 34356 71652
rect 33852 71598 33854 71650
rect 33906 71598 34302 71650
rect 34354 71598 34356 71650
rect 33852 71596 34356 71598
rect 33852 71090 33908 71596
rect 34300 71586 34356 71596
rect 33852 71038 33854 71090
rect 33906 71038 33908 71090
rect 33628 70914 33684 70924
rect 33292 70866 33348 70878
rect 33292 70814 33294 70866
rect 33346 70814 33348 70866
rect 31612 70084 31668 70094
rect 31612 69990 31668 70028
rect 32508 69522 32564 69534
rect 32508 69470 32510 69522
rect 32562 69470 32564 69522
rect 32396 69188 32452 69198
rect 31836 67842 31892 67854
rect 31836 67790 31838 67842
rect 31890 67790 31892 67842
rect 31500 67620 31556 67630
rect 31836 67620 31892 67790
rect 31556 67564 31892 67620
rect 31500 67526 31556 67564
rect 31500 63924 31556 63934
rect 31500 63830 31556 63868
rect 31164 60508 31444 60564
rect 30716 60116 30772 60126
rect 30716 60022 30772 60060
rect 30604 59278 30606 59330
rect 30658 59278 30660 59330
rect 30604 58324 30660 59278
rect 30940 59780 30996 59790
rect 30940 58434 30996 59724
rect 30940 58382 30942 58434
rect 30994 58382 30996 58434
rect 30940 58370 30996 58382
rect 31052 59106 31108 59118
rect 31052 59054 31054 59106
rect 31106 59054 31108 59106
rect 30604 58258 30660 58268
rect 31052 58100 31108 59054
rect 30380 58044 31108 58100
rect 29820 56754 30100 56756
rect 29820 56702 29822 56754
rect 29874 56702 30100 56754
rect 29820 56700 30100 56702
rect 30156 57540 30212 57550
rect 30156 56754 30212 57484
rect 30156 56702 30158 56754
rect 30210 56702 30212 56754
rect 29820 56690 29876 56700
rect 30156 56690 30212 56702
rect 30268 57204 30324 57214
rect 29708 56252 29988 56308
rect 29708 54740 29764 54750
rect 29708 54646 29764 54684
rect 29708 53956 29764 53966
rect 29708 53862 29764 53900
rect 29820 53732 29876 53742
rect 29708 53172 29764 53182
rect 29708 51940 29764 53116
rect 29820 52724 29876 53676
rect 29820 52052 29876 52668
rect 29820 51986 29876 51996
rect 29708 51604 29764 51884
rect 29820 51604 29876 51614
rect 29708 51602 29876 51604
rect 29708 51550 29822 51602
rect 29874 51550 29876 51602
rect 29708 51548 29876 51550
rect 29820 51538 29876 51548
rect 29708 50594 29764 50606
rect 29708 50542 29710 50594
rect 29762 50542 29764 50594
rect 29708 50036 29764 50542
rect 29708 49970 29764 49980
rect 29820 50484 29876 50494
rect 29708 49812 29764 49822
rect 29708 49718 29764 49756
rect 29820 49810 29876 50428
rect 29820 49758 29822 49810
rect 29874 49758 29876 49810
rect 29820 49746 29876 49758
rect 29820 49252 29876 49262
rect 29820 49158 29876 49196
rect 29596 48300 29764 48356
rect 29596 48130 29652 48142
rect 29596 48078 29598 48130
rect 29650 48078 29652 48130
rect 29596 47684 29652 48078
rect 29260 47628 29596 47684
rect 29260 47234 29316 47628
rect 29596 47570 29652 47628
rect 29596 47518 29598 47570
rect 29650 47518 29652 47570
rect 29596 47506 29652 47518
rect 29260 47182 29262 47234
rect 29314 47182 29316 47234
rect 29260 47124 29316 47182
rect 29484 47460 29540 47470
rect 29260 47068 29428 47124
rect 29148 46956 29316 47012
rect 29036 46844 29204 46900
rect 29036 46676 29092 46686
rect 29036 46562 29092 46620
rect 29036 46510 29038 46562
rect 29090 46510 29092 46562
rect 29036 45668 29092 46510
rect 29148 46002 29204 46844
rect 29148 45950 29150 46002
rect 29202 45950 29204 46002
rect 29148 45938 29204 45950
rect 29036 45602 29092 45612
rect 28924 45266 28980 45276
rect 29036 45444 29092 45454
rect 29036 45218 29092 45388
rect 29036 45166 29038 45218
rect 29090 45166 29092 45218
rect 29036 45154 29092 45166
rect 28924 45108 28980 45118
rect 28588 45106 28980 45108
rect 28588 45054 28926 45106
rect 28978 45054 28980 45106
rect 28588 45052 28980 45054
rect 28700 44882 28756 44894
rect 28700 44830 28702 44882
rect 28754 44830 28756 44882
rect 28700 44324 28756 44830
rect 28924 44660 28980 45052
rect 29148 44660 29204 44670
rect 28924 44604 29148 44660
rect 29148 44594 29204 44604
rect 29148 44324 29204 44334
rect 29260 44324 29316 46956
rect 29372 46004 29428 47068
rect 29372 45938 29428 45948
rect 29372 45780 29428 45790
rect 29372 45686 29428 45724
rect 29372 44996 29428 45006
rect 29372 44902 29428 44940
rect 28700 44268 29092 44324
rect 28476 44210 28644 44212
rect 28476 44158 28478 44210
rect 28530 44158 28644 44210
rect 28476 44156 28644 44158
rect 28476 44146 28532 44156
rect 28252 43362 28308 43372
rect 28364 44100 28420 44110
rect 28140 42130 28196 42140
rect 28252 42530 28308 42542
rect 28252 42478 28254 42530
rect 28306 42478 28308 42530
rect 28252 42084 28308 42478
rect 28252 42018 28308 42028
rect 28028 41346 28084 41356
rect 28140 41858 28196 41870
rect 28140 41806 28142 41858
rect 28194 41806 28196 41858
rect 28028 40740 28084 40750
rect 28028 39732 28084 40684
rect 28140 40516 28196 41806
rect 28252 41412 28308 41422
rect 28252 41298 28308 41356
rect 28252 41246 28254 41298
rect 28306 41246 28308 41298
rect 28252 41234 28308 41246
rect 28140 40450 28196 40460
rect 28252 40404 28308 40414
rect 28140 39732 28196 39742
rect 28028 39730 28196 39732
rect 28028 39678 28142 39730
rect 28194 39678 28196 39730
rect 28028 39676 28196 39678
rect 28140 39666 28196 39676
rect 28252 39172 28308 40348
rect 28140 39116 28308 39172
rect 28028 38836 28084 38846
rect 28028 38742 28084 38780
rect 27916 38612 28084 38668
rect 27804 38164 27860 38174
rect 27580 38052 27636 38062
rect 27468 38050 27636 38052
rect 27468 37998 27582 38050
rect 27634 37998 27636 38050
rect 27468 37996 27636 37998
rect 27580 37986 27636 37996
rect 27804 38050 27860 38108
rect 27804 37998 27806 38050
rect 27858 37998 27860 38050
rect 27804 37986 27860 37998
rect 27244 37940 27300 37950
rect 27244 37846 27300 37884
rect 27356 37828 27412 37838
rect 27356 37734 27412 37772
rect 27244 37716 27300 37726
rect 27244 37380 27300 37660
rect 27356 37380 27412 37390
rect 27244 37324 27356 37380
rect 27356 37286 27412 37324
rect 27580 37268 27636 37278
rect 27468 37044 27524 37054
rect 27244 36370 27300 36382
rect 27244 36318 27246 36370
rect 27298 36318 27300 36370
rect 27244 36260 27300 36318
rect 27468 36370 27524 36988
rect 27580 36706 27636 37212
rect 27916 37266 27972 37278
rect 27916 37214 27918 37266
rect 27970 37214 27972 37266
rect 27916 36820 27972 37214
rect 27916 36754 27972 36764
rect 27580 36654 27582 36706
rect 27634 36654 27636 36706
rect 27580 36642 27636 36654
rect 27804 36708 27860 36718
rect 27804 36614 27860 36652
rect 27468 36318 27470 36370
rect 27522 36318 27524 36370
rect 27468 36306 27524 36318
rect 27916 36370 27972 36382
rect 27916 36318 27918 36370
rect 27970 36318 27972 36370
rect 27356 36260 27412 36270
rect 27244 36204 27356 36260
rect 27356 36194 27412 36204
rect 27916 36036 27972 36318
rect 27916 35970 27972 35980
rect 26796 32498 26852 32508
rect 26908 34188 27188 34244
rect 27244 35252 27300 35262
rect 26348 30818 26404 30828
rect 26460 32060 26740 32116
rect 26460 30548 26516 32060
rect 26684 31892 26740 31902
rect 26684 31666 26740 31836
rect 26796 31780 26852 31790
rect 26908 31780 26964 34188
rect 26796 31778 26964 31780
rect 26796 31726 26798 31778
rect 26850 31726 26964 31778
rect 26796 31724 26964 31726
rect 27020 34020 27076 34030
rect 26796 31714 26852 31724
rect 26684 31614 26686 31666
rect 26738 31614 26740 31666
rect 26684 31602 26740 31614
rect 26572 31556 26628 31566
rect 26572 31218 26628 31500
rect 26572 31166 26574 31218
rect 26626 31166 26628 31218
rect 26572 31154 26628 31166
rect 26796 31332 26852 31342
rect 26684 30548 26740 30558
rect 26460 30492 26628 30548
rect 26236 30436 26292 30446
rect 25788 30380 26068 30436
rect 25228 30322 25956 30324
rect 25228 30270 25230 30322
rect 25282 30270 25956 30322
rect 25228 30268 25956 30270
rect 25228 30258 25284 30268
rect 25900 30210 25956 30268
rect 25900 30158 25902 30210
rect 25954 30158 25956 30210
rect 25900 30146 25956 30158
rect 25676 30098 25732 30110
rect 25676 30046 25678 30098
rect 25730 30046 25732 30098
rect 25676 29540 25732 30046
rect 26012 29652 26068 30380
rect 26236 30342 26292 30380
rect 26572 30322 26628 30492
rect 26572 30270 26574 30322
rect 26626 30270 26628 30322
rect 26572 30100 26628 30270
rect 25228 29484 25676 29540
rect 25116 28532 25172 28542
rect 25116 26908 25172 28476
rect 25228 27970 25284 29484
rect 25676 29474 25732 29484
rect 25788 29596 26068 29652
rect 26124 30044 26628 30100
rect 26124 29986 26180 30044
rect 26124 29934 26126 29986
rect 26178 29934 26180 29986
rect 25788 28420 25844 29596
rect 26012 29428 26068 29438
rect 26012 29334 26068 29372
rect 26124 28980 26180 29934
rect 26460 29652 26516 29662
rect 26460 29558 26516 29596
rect 26684 28980 26740 30492
rect 25788 28354 25844 28364
rect 25900 28924 26180 28980
rect 26572 28924 26740 28980
rect 25900 28754 25956 28924
rect 25900 28702 25902 28754
rect 25954 28702 25956 28754
rect 25900 28196 25956 28702
rect 25676 28140 25900 28196
rect 26572 28196 26628 28924
rect 26684 28756 26740 28766
rect 26684 28662 26740 28700
rect 26572 28140 26740 28196
rect 25676 28082 25732 28140
rect 25900 28102 25956 28140
rect 25676 28030 25678 28082
rect 25730 28030 25732 28082
rect 25676 28018 25732 28030
rect 25228 27918 25230 27970
rect 25282 27918 25284 27970
rect 25228 27748 25284 27918
rect 25788 27972 25844 27982
rect 26572 27972 26628 27982
rect 25788 27970 26628 27972
rect 25788 27918 25790 27970
rect 25842 27918 26574 27970
rect 26626 27918 26628 27970
rect 25788 27916 26628 27918
rect 25788 27906 25844 27916
rect 26572 27906 26628 27916
rect 25452 27860 25508 27870
rect 25452 27766 25508 27804
rect 25228 27682 25284 27692
rect 25900 27748 25956 27758
rect 26124 27748 26180 27758
rect 26684 27748 26740 28140
rect 25956 27746 26404 27748
rect 25956 27694 26126 27746
rect 26178 27694 26404 27746
rect 25956 27692 26404 27694
rect 25900 27682 25956 27692
rect 26124 27682 26180 27692
rect 25676 27524 25732 27534
rect 25340 27188 25396 27198
rect 25676 27188 25732 27468
rect 25340 27186 25732 27188
rect 25340 27134 25342 27186
rect 25394 27134 25678 27186
rect 25730 27134 25732 27186
rect 25340 27132 25732 27134
rect 25340 27122 25396 27132
rect 25676 27122 25732 27132
rect 26124 27188 26180 27198
rect 26124 27094 26180 27132
rect 25900 27074 25956 27086
rect 25900 27022 25902 27074
rect 25954 27022 25956 27074
rect 25564 26964 25620 26974
rect 25116 26852 25620 26908
rect 25004 26674 25060 26684
rect 24556 25340 24724 25396
rect 24556 23828 24612 25340
rect 24556 23762 24612 23772
rect 24668 24724 24724 24734
rect 24668 24610 24724 24668
rect 24668 24558 24670 24610
rect 24722 24558 24724 24610
rect 24668 23716 24724 24558
rect 25340 24052 25396 26852
rect 25452 26516 25508 26526
rect 25452 26422 25508 26460
rect 25564 26402 25620 26852
rect 25564 26350 25566 26402
rect 25618 26350 25620 26402
rect 25564 26338 25620 26350
rect 25452 26068 25508 26078
rect 25452 25974 25508 26012
rect 25452 24612 25508 24622
rect 25452 24518 25508 24556
rect 25228 24050 25396 24052
rect 25228 23998 25342 24050
rect 25394 23998 25396 24050
rect 25228 23996 25396 23998
rect 24892 23716 24948 23726
rect 24668 23650 24724 23660
rect 24780 23714 24948 23716
rect 24780 23662 24894 23714
rect 24946 23662 24948 23714
rect 24780 23660 24948 23662
rect 24668 23156 24724 23166
rect 24780 23156 24836 23660
rect 24892 23650 24948 23660
rect 25116 23156 25172 23166
rect 24668 23154 24836 23156
rect 24668 23102 24670 23154
rect 24722 23102 24836 23154
rect 24668 23100 24836 23102
rect 24892 23154 25172 23156
rect 24892 23102 25118 23154
rect 25170 23102 25172 23154
rect 24892 23100 25172 23102
rect 25228 23156 25284 23996
rect 25340 23986 25396 23996
rect 25340 23380 25396 23390
rect 25788 23380 25844 23390
rect 25900 23380 25956 27022
rect 26012 26964 26068 26974
rect 26012 26514 26068 26908
rect 26012 26462 26014 26514
rect 26066 26462 26068 26514
rect 26012 26450 26068 26462
rect 25340 23378 25956 23380
rect 25340 23326 25342 23378
rect 25394 23326 25790 23378
rect 25842 23326 25956 23378
rect 25340 23324 25956 23326
rect 26012 24052 26068 24062
rect 25340 23314 25396 23324
rect 25788 23314 25844 23324
rect 25452 23156 25508 23166
rect 25228 23154 25844 23156
rect 25228 23102 25454 23154
rect 25506 23102 25844 23154
rect 25228 23100 25844 23102
rect 24556 22932 24612 22942
rect 24556 22838 24612 22876
rect 24668 22372 24724 23100
rect 24108 19346 24500 19348
rect 24108 19294 24334 19346
rect 24386 19294 24500 19346
rect 24108 19292 24500 19294
rect 24556 22316 24724 22372
rect 23884 19236 23940 19246
rect 23884 19142 23940 19180
rect 23884 18676 23940 18686
rect 23772 18674 23940 18676
rect 23772 18622 23886 18674
rect 23938 18622 23940 18674
rect 23772 18620 23940 18622
rect 23884 18610 23940 18620
rect 23660 17042 23716 17052
rect 24108 18450 24164 19292
rect 24332 19282 24388 19292
rect 24556 18788 24612 22316
rect 24668 21812 24724 21822
rect 24668 21718 24724 21756
rect 24892 20914 24948 23100
rect 25116 23090 25172 23100
rect 25452 23090 25508 23100
rect 25340 22932 25396 22942
rect 25340 22482 25396 22876
rect 25340 22430 25342 22482
rect 25394 22430 25396 22482
rect 25340 22418 25396 22430
rect 25676 22932 25732 22942
rect 25228 21812 25284 21822
rect 25228 21586 25284 21756
rect 25228 21534 25230 21586
rect 25282 21534 25284 21586
rect 25228 21522 25284 21534
rect 24892 20862 24894 20914
rect 24946 20862 24948 20914
rect 24892 20850 24948 20862
rect 25676 20188 25732 22876
rect 25340 20132 25396 20142
rect 24332 18732 24612 18788
rect 24668 19236 24724 19246
rect 24108 18398 24110 18450
rect 24162 18398 24164 18450
rect 23996 15540 24052 15550
rect 24108 15540 24164 18398
rect 24220 18452 24276 18462
rect 24220 17778 24276 18396
rect 24220 17726 24222 17778
rect 24274 17726 24276 17778
rect 24220 17714 24276 17726
rect 23996 15538 24164 15540
rect 23996 15486 23998 15538
rect 24050 15486 24164 15538
rect 23996 15484 24164 15486
rect 22540 13918 22542 13970
rect 22594 13918 22596 13970
rect 22540 13906 22596 13918
rect 22652 13972 22708 13982
rect 22652 13878 22708 13916
rect 22988 13860 23044 13870
rect 22540 13524 22596 13534
rect 22540 13074 22596 13468
rect 22540 13022 22542 13074
rect 22594 13022 22596 13074
rect 22540 13010 22596 13022
rect 22428 12796 22596 12852
rect 21980 12014 21982 12066
rect 22034 12014 22036 12066
rect 21644 11394 21700 11406
rect 21644 11342 21646 11394
rect 21698 11342 21700 11394
rect 20524 11284 20580 11294
rect 21308 11284 21364 11294
rect 20524 11282 21364 11284
rect 20524 11230 20526 11282
rect 20578 11230 21310 11282
rect 21362 11230 21364 11282
rect 20524 11228 21364 11230
rect 20524 11218 20580 11228
rect 21308 11218 21364 11228
rect 21644 11172 21700 11342
rect 20972 10498 21028 10510
rect 20972 10446 20974 10498
rect 21026 10446 21028 10498
rect 20748 9604 20804 9614
rect 20972 9604 21028 10446
rect 21644 9826 21700 11116
rect 21868 9940 21924 9950
rect 21980 9940 22036 12014
rect 21868 9938 22036 9940
rect 21868 9886 21870 9938
rect 21922 9886 22036 9938
rect 21868 9884 22036 9886
rect 21868 9874 21924 9884
rect 21644 9774 21646 9826
rect 21698 9774 21700 9826
rect 21308 9604 21364 9614
rect 20748 9602 21028 9604
rect 20748 9550 20750 9602
rect 20802 9550 21028 9602
rect 20748 9548 21028 9550
rect 21196 9602 21364 9604
rect 21196 9550 21310 9602
rect 21362 9550 21364 9602
rect 21196 9548 21364 9550
rect 20748 8596 20804 9548
rect 20748 8530 20804 8540
rect 20860 9154 20916 9166
rect 20860 9102 20862 9154
rect 20914 9102 20916 9154
rect 20860 8428 20916 9102
rect 21196 9154 21252 9548
rect 21308 9538 21364 9548
rect 21196 9102 21198 9154
rect 21250 9102 21252 9154
rect 21196 9090 21252 9102
rect 21644 8596 21700 9774
rect 21868 8596 21924 8606
rect 21644 8540 21868 8596
rect 20524 8372 20916 8428
rect 21868 8372 21924 8540
rect 22428 8372 22484 8382
rect 20524 7586 20580 8372
rect 21868 8370 22484 8372
rect 21868 8318 21870 8370
rect 21922 8318 22430 8370
rect 22482 8318 22484 8370
rect 21868 8316 22484 8318
rect 21868 8306 21924 8316
rect 22428 8306 22484 8316
rect 20524 7534 20526 7586
rect 20578 7534 20580 7586
rect 20524 7522 20580 7534
rect 22092 8034 22148 8046
rect 22092 7982 22094 8034
rect 22146 7982 22148 8034
rect 21420 6692 21476 6702
rect 22092 6692 22148 7982
rect 22540 7364 22596 12796
rect 22652 12516 22708 12526
rect 22652 11508 22708 12460
rect 22652 9266 22708 11452
rect 22764 11172 22820 11182
rect 22764 11078 22820 11116
rect 22652 9214 22654 9266
rect 22706 9214 22708 9266
rect 22652 9202 22708 9214
rect 22988 8428 23044 13804
rect 23212 12292 23268 14588
rect 23324 15092 23380 15102
rect 23324 14532 23380 15036
rect 23996 15092 24052 15484
rect 23996 15026 24052 15036
rect 24332 14756 24388 18732
rect 24444 18562 24500 18574
rect 24444 18510 24446 18562
rect 24498 18510 24500 18562
rect 24444 17556 24500 18510
rect 24668 17892 24724 19180
rect 24780 19236 24836 19246
rect 24780 19234 25172 19236
rect 24780 19182 24782 19234
rect 24834 19182 25172 19234
rect 24780 19180 25172 19182
rect 24780 19170 24836 19180
rect 25004 19010 25060 19022
rect 25004 18958 25006 19010
rect 25058 18958 25060 19010
rect 25004 18452 25060 18958
rect 25004 18386 25060 18396
rect 24780 17892 24836 17902
rect 24668 17836 24780 17892
rect 24780 17798 24836 17836
rect 25116 17890 25172 19180
rect 25116 17838 25118 17890
rect 25170 17838 25172 17890
rect 25116 17826 25172 17838
rect 25228 18450 25284 18462
rect 25228 18398 25230 18450
rect 25282 18398 25284 18450
rect 24556 17556 24612 17566
rect 24444 17554 24612 17556
rect 24444 17502 24558 17554
rect 24610 17502 24612 17554
rect 24444 17500 24612 17502
rect 24332 14700 24500 14756
rect 24332 14532 24388 14542
rect 23324 14530 23492 14532
rect 23324 14478 23326 14530
rect 23378 14478 23492 14530
rect 23324 14476 23492 14478
rect 23324 14466 23380 14476
rect 23436 13972 23492 14476
rect 23660 14530 24388 14532
rect 23660 14478 24334 14530
rect 24386 14478 24388 14530
rect 23660 14476 24388 14478
rect 23324 13860 23380 13870
rect 23324 13766 23380 13804
rect 23436 13746 23492 13916
rect 23436 13694 23438 13746
rect 23490 13694 23492 13746
rect 23436 13682 23492 13694
rect 23548 14418 23604 14430
rect 23548 14366 23550 14418
rect 23602 14366 23604 14418
rect 23324 12292 23380 12302
rect 23212 12290 23380 12292
rect 23212 12238 23326 12290
rect 23378 12238 23380 12290
rect 23212 12236 23380 12238
rect 23100 12180 23156 12190
rect 23100 12086 23156 12124
rect 23324 11732 23380 12236
rect 23324 11666 23380 11676
rect 23100 11394 23156 11406
rect 23100 11342 23102 11394
rect 23154 11342 23156 11394
rect 23100 11172 23156 11342
rect 23324 11396 23380 11406
rect 23324 11302 23380 11340
rect 23548 11172 23604 14366
rect 23660 11618 23716 14476
rect 24332 14466 24388 14476
rect 24108 14306 24164 14318
rect 24108 14254 24110 14306
rect 24162 14254 24164 14306
rect 24108 13524 24164 14254
rect 24220 14308 24276 14318
rect 24220 13970 24276 14252
rect 24220 13918 24222 13970
rect 24274 13918 24276 13970
rect 24220 13906 24276 13918
rect 24108 13458 24164 13468
rect 23996 13188 24052 13198
rect 23996 12402 24052 13132
rect 24444 12516 24500 14700
rect 24556 13076 24612 17500
rect 25228 16996 25284 18398
rect 25116 16940 25284 16996
rect 24668 16884 24724 16894
rect 24668 16790 24724 16828
rect 25116 16884 25172 16940
rect 25116 16818 25172 16828
rect 25228 16772 25284 16782
rect 25340 16772 25396 20076
rect 25452 20132 25732 20188
rect 25452 19346 25508 20132
rect 25452 19294 25454 19346
rect 25506 19294 25508 19346
rect 25452 18676 25508 19294
rect 25452 18610 25508 18620
rect 25564 17442 25620 17454
rect 25564 17390 25566 17442
rect 25618 17390 25620 17442
rect 25564 16884 25620 17390
rect 25564 16818 25620 16828
rect 25228 16770 25396 16772
rect 25228 16718 25230 16770
rect 25282 16718 25396 16770
rect 25228 16716 25396 16718
rect 25228 16706 25284 16716
rect 25788 16212 25844 23100
rect 25900 23042 25956 23054
rect 25900 22990 25902 23042
rect 25954 22990 25956 23042
rect 25900 21476 25956 22990
rect 26012 22932 26068 23996
rect 26012 22866 26068 22876
rect 26124 22596 26180 22606
rect 26124 22370 26180 22540
rect 26124 22318 26126 22370
rect 26178 22318 26180 22370
rect 26124 22306 26180 22318
rect 25900 21410 25956 21420
rect 26012 21474 26068 21486
rect 26012 21422 26014 21474
rect 26066 21422 26068 21474
rect 26012 20804 26068 21422
rect 26012 20738 26068 20748
rect 26348 20020 26404 27692
rect 26348 19954 26404 19964
rect 26460 27692 26740 27748
rect 26460 25620 26516 27692
rect 26572 27300 26628 27310
rect 26572 27206 26628 27244
rect 26684 27188 26740 27198
rect 26684 26514 26740 27132
rect 26684 26462 26686 26514
rect 26738 26462 26740 26514
rect 26684 26450 26740 26462
rect 26684 25620 26740 25630
rect 26460 25618 26740 25620
rect 26460 25566 26686 25618
rect 26738 25566 26740 25618
rect 26460 25564 26740 25566
rect 26012 18452 26068 18462
rect 26012 18358 26068 18396
rect 26236 17892 26292 17902
rect 26236 17798 26292 17836
rect 26460 17778 26516 25564
rect 26684 25554 26740 25564
rect 26796 25396 26852 31276
rect 26908 29652 26964 29662
rect 27020 29652 27076 33964
rect 27132 34020 27188 34030
rect 27244 34020 27300 35196
rect 27468 34690 27524 34702
rect 27468 34638 27470 34690
rect 27522 34638 27524 34690
rect 27468 34244 27524 34638
rect 27916 34692 27972 34702
rect 27916 34598 27972 34636
rect 27468 34178 27524 34188
rect 27132 34018 27300 34020
rect 27132 33966 27134 34018
rect 27186 33966 27300 34018
rect 27132 33964 27300 33966
rect 27132 33908 27188 33964
rect 27132 33842 27188 33852
rect 27356 33236 27412 33246
rect 27356 33142 27412 33180
rect 27692 33122 27748 33134
rect 27692 33070 27694 33122
rect 27746 33070 27748 33122
rect 27356 32116 27412 32126
rect 27244 32060 27356 32116
rect 26964 29596 27076 29652
rect 26908 29586 26964 29596
rect 27020 29538 27076 29596
rect 27132 29986 27188 29998
rect 27132 29934 27134 29986
rect 27186 29934 27188 29986
rect 27132 29652 27188 29934
rect 27132 29558 27188 29596
rect 27020 29486 27022 29538
rect 27074 29486 27076 29538
rect 27020 29474 27076 29486
rect 26908 28196 26964 28206
rect 26908 26962 26964 28140
rect 27020 27970 27076 27982
rect 27020 27918 27022 27970
rect 27074 27918 27076 27970
rect 27020 27300 27076 27918
rect 27020 27234 27076 27244
rect 27244 27298 27300 32060
rect 27356 32050 27412 32060
rect 27692 31892 27748 33070
rect 27692 31826 27748 31836
rect 27468 31778 27524 31790
rect 27468 31726 27470 31778
rect 27522 31726 27524 31778
rect 27468 30436 27524 31726
rect 27468 30370 27524 30380
rect 27916 31778 27972 31790
rect 27916 31726 27918 31778
rect 27970 31726 27972 31778
rect 27916 29540 27972 31726
rect 27916 29474 27972 29484
rect 27356 29316 27412 29326
rect 27356 28756 27412 29260
rect 28028 29204 28084 38612
rect 28140 37490 28196 39116
rect 28252 38612 28308 38622
rect 28252 38162 28308 38556
rect 28364 38500 28420 44044
rect 28588 43652 28644 44156
rect 28700 44100 28756 44110
rect 29036 44100 29092 44268
rect 29148 44322 29316 44324
rect 29148 44270 29150 44322
rect 29202 44270 29316 44322
rect 29148 44268 29316 44270
rect 29484 44324 29540 47404
rect 29148 44258 29204 44268
rect 29484 44258 29540 44268
rect 29596 45778 29652 45790
rect 29596 45726 29598 45778
rect 29650 45726 29652 45778
rect 29260 44100 29316 44110
rect 29036 44098 29316 44100
rect 29036 44046 29262 44098
rect 29314 44046 29316 44098
rect 29036 44044 29316 44046
rect 28700 44006 28756 44044
rect 29260 43764 29316 44044
rect 29484 44100 29540 44110
rect 29484 44006 29540 44044
rect 29148 43708 29316 43764
rect 28812 43652 28868 43662
rect 28588 43650 28868 43652
rect 28588 43598 28814 43650
rect 28866 43598 28868 43650
rect 28588 43596 28868 43598
rect 28812 43586 28868 43596
rect 28812 42196 28868 42234
rect 28812 42130 28868 42140
rect 28924 40964 28980 40974
rect 28476 40628 28532 40638
rect 28476 40514 28532 40572
rect 28924 40626 28980 40908
rect 28924 40574 28926 40626
rect 28978 40574 28980 40626
rect 28924 40562 28980 40574
rect 28476 40462 28478 40514
rect 28530 40462 28532 40514
rect 28476 40450 28532 40462
rect 28924 40068 28980 40078
rect 28588 39732 28644 39742
rect 28588 39396 28644 39676
rect 28588 38668 28644 39340
rect 28364 38434 28420 38444
rect 28476 38612 28644 38668
rect 28700 38722 28756 38734
rect 28700 38670 28702 38722
rect 28754 38670 28756 38722
rect 28252 38110 28254 38162
rect 28306 38110 28308 38162
rect 28252 37940 28308 38110
rect 28252 37874 28308 37884
rect 28140 37438 28142 37490
rect 28194 37438 28196 37490
rect 28140 37426 28196 37438
rect 28476 37492 28532 38612
rect 28364 37268 28420 37278
rect 28476 37268 28532 37436
rect 28364 37266 28532 37268
rect 28364 37214 28366 37266
rect 28418 37214 28532 37266
rect 28364 37212 28532 37214
rect 28588 37380 28644 37390
rect 28588 37266 28644 37324
rect 28588 37214 28590 37266
rect 28642 37214 28644 37266
rect 28364 37202 28420 37212
rect 28588 37202 28644 37214
rect 28252 37154 28308 37166
rect 28252 37102 28254 37154
rect 28306 37102 28308 37154
rect 28252 36484 28308 37102
rect 28252 36418 28308 36428
rect 28588 36708 28644 36718
rect 28364 36260 28420 36270
rect 28140 36036 28196 36046
rect 28140 35922 28196 35980
rect 28140 35870 28142 35922
rect 28194 35870 28196 35922
rect 28140 35858 28196 35870
rect 28252 33346 28308 33358
rect 28252 33294 28254 33346
rect 28306 33294 28308 33346
rect 28252 32900 28308 33294
rect 28252 32834 28308 32844
rect 28252 32676 28308 32686
rect 28140 32450 28196 32462
rect 28140 32398 28142 32450
rect 28194 32398 28196 32450
rect 28140 31780 28196 32398
rect 28252 32002 28308 32620
rect 28252 31950 28254 32002
rect 28306 31950 28308 32002
rect 28252 31938 28308 31950
rect 28140 30996 28196 31724
rect 28140 30930 28196 30940
rect 27692 29148 28308 29204
rect 27356 28754 27524 28756
rect 27356 28702 27358 28754
rect 27410 28702 27524 28754
rect 27356 28700 27524 28702
rect 27356 28690 27412 28700
rect 27468 27858 27524 28700
rect 27692 28754 27748 29148
rect 27692 28702 27694 28754
rect 27746 28702 27748 28754
rect 27692 28690 27748 28702
rect 28252 28754 28308 29148
rect 28252 28702 28254 28754
rect 28306 28702 28308 28754
rect 28252 28690 28308 28702
rect 27804 28418 27860 28430
rect 27804 28366 27806 28418
rect 27858 28366 27860 28418
rect 27468 27806 27470 27858
rect 27522 27806 27524 27858
rect 27468 27794 27524 27806
rect 27692 27860 27748 27870
rect 27692 27766 27748 27804
rect 27244 27246 27246 27298
rect 27298 27246 27300 27298
rect 27244 27188 27300 27246
rect 27244 27122 27300 27132
rect 27692 27636 27748 27646
rect 26908 26910 26910 26962
rect 26962 26910 26964 26962
rect 26908 26628 26964 26910
rect 26908 26562 26964 26572
rect 27132 26908 27188 26918
rect 26572 25340 26852 25396
rect 26572 20132 26628 25340
rect 27020 24052 27076 24062
rect 27020 23958 27076 23996
rect 26796 23828 26852 23838
rect 26684 23044 26740 23054
rect 26684 21812 26740 22988
rect 26796 22482 26852 23772
rect 27020 23156 27076 23166
rect 27020 23062 27076 23100
rect 27020 22708 27076 22718
rect 26796 22430 26798 22482
rect 26850 22430 26852 22482
rect 26796 22418 26852 22430
rect 26908 22596 26964 22606
rect 26908 22260 26964 22540
rect 26908 22194 26964 22204
rect 26684 21746 26740 21756
rect 27020 20914 27076 22652
rect 27020 20862 27022 20914
rect 27074 20862 27076 20914
rect 27020 20850 27076 20862
rect 26572 20066 26628 20076
rect 26908 20018 26964 20030
rect 26908 19966 26910 20018
rect 26962 19966 26964 20018
rect 26460 17726 26462 17778
rect 26514 17726 26516 17778
rect 26460 17714 26516 17726
rect 26572 19908 26628 19918
rect 26908 19908 26964 19966
rect 26572 19906 26964 19908
rect 26572 19854 26574 19906
rect 26626 19854 26964 19906
rect 26572 19852 26964 19854
rect 25788 16146 25844 16156
rect 25900 17442 25956 17454
rect 25900 17390 25902 17442
rect 25954 17390 25956 17442
rect 24892 14644 24948 14654
rect 24892 14550 24948 14588
rect 24668 13972 24724 13982
rect 24724 13916 24836 13972
rect 24668 13878 24724 13916
rect 24668 13076 24724 13086
rect 24556 13074 24724 13076
rect 24556 13022 24670 13074
rect 24722 13022 24724 13074
rect 24556 13020 24724 13022
rect 24668 13010 24724 13020
rect 23996 12350 23998 12402
rect 24050 12350 24052 12402
rect 23996 12338 24052 12350
rect 24332 12460 24500 12516
rect 23660 11566 23662 11618
rect 23714 11566 23716 11618
rect 23660 11554 23716 11566
rect 24108 11396 24164 11406
rect 24108 11302 24164 11340
rect 23100 11116 23716 11172
rect 23324 10948 23380 10958
rect 23380 10892 23492 10948
rect 23324 10882 23380 10892
rect 23436 9940 23492 10892
rect 23548 9940 23604 9950
rect 23436 9884 23548 9940
rect 23548 9846 23604 9884
rect 22652 8372 23044 8428
rect 22652 8370 22708 8372
rect 22652 8318 22654 8370
rect 22706 8318 22708 8370
rect 22652 8306 22708 8318
rect 22988 8370 23044 8372
rect 22988 8318 22990 8370
rect 23042 8318 23044 8370
rect 22988 8306 23044 8318
rect 22652 7364 22708 7374
rect 22540 7362 22708 7364
rect 22540 7310 22654 7362
rect 22706 7310 22708 7362
rect 22540 7308 22708 7310
rect 22652 7298 22708 7308
rect 22204 6692 22260 6702
rect 22092 6690 22260 6692
rect 22092 6638 22206 6690
rect 22258 6638 22260 6690
rect 22092 6636 22260 6638
rect 19836 6234 20100 6244
rect 20188 6188 20468 6244
rect 20748 6580 20804 6590
rect 19628 6020 19684 6030
rect 19516 6018 19684 6020
rect 19516 5966 19630 6018
rect 19682 5966 19684 6018
rect 19516 5964 19684 5966
rect 19628 5124 19684 5964
rect 20188 6018 20244 6188
rect 20188 5966 20190 6018
rect 20242 5966 20244 6018
rect 20188 5954 20244 5966
rect 19964 5908 20020 5918
rect 20748 5908 20804 6524
rect 19628 5010 19684 5068
rect 19852 5124 19908 5134
rect 19964 5124 20020 5852
rect 20412 5906 20804 5908
rect 20412 5854 20750 5906
rect 20802 5854 20804 5906
rect 20412 5852 20804 5854
rect 20412 5236 20468 5852
rect 20748 5842 20804 5852
rect 21420 5348 21476 6636
rect 22204 6626 22260 6636
rect 21980 6468 22036 6478
rect 21532 6466 22036 6468
rect 21532 6414 21982 6466
rect 22034 6414 22036 6466
rect 21532 6412 22036 6414
rect 21532 6018 21588 6412
rect 21980 6402 22036 6412
rect 21532 5966 21534 6018
rect 21586 5966 21588 6018
rect 21532 5954 21588 5966
rect 23100 6020 23156 6030
rect 21532 5348 21588 5358
rect 21420 5292 21532 5348
rect 20412 5142 20468 5180
rect 21532 5234 21588 5292
rect 21532 5182 21534 5234
rect 21586 5182 21588 5234
rect 21532 5170 21588 5182
rect 22652 5236 22708 5246
rect 19852 5122 20020 5124
rect 19852 5070 19854 5122
rect 19906 5070 20020 5122
rect 19852 5068 20020 5070
rect 21868 5124 21924 5134
rect 19852 5058 19908 5068
rect 21868 5030 21924 5068
rect 19628 4958 19630 5010
rect 19682 4958 19684 5010
rect 19628 4946 19684 4958
rect 22428 5010 22484 5022
rect 22428 4958 22430 5010
rect 22482 4958 22484 5010
rect 19292 4900 19348 4910
rect 19180 4898 19348 4900
rect 19180 4846 19294 4898
rect 19346 4846 19348 4898
rect 19180 4844 19348 4846
rect 19292 4834 19348 4844
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19068 4162 19124 4172
rect 20300 4228 20356 4238
rect 20300 4134 20356 4172
rect 18956 3574 19012 3612
rect 19516 3668 19572 3678
rect 19516 3666 19908 3668
rect 19516 3614 19518 3666
rect 19570 3614 19908 3666
rect 19516 3612 19908 3614
rect 19516 3602 19572 3612
rect 19180 3554 19236 3566
rect 19180 3502 19182 3554
rect 19234 3502 19236 3554
rect 19180 3444 19236 3502
rect 19852 3554 19908 3612
rect 19852 3502 19854 3554
rect 19906 3502 19908 3554
rect 19852 3490 19908 3502
rect 18732 3388 19236 3444
rect 20188 3332 20244 3342
rect 20188 3330 20356 3332
rect 20188 3278 20190 3330
rect 20242 3278 20356 3330
rect 20188 3276 20356 3278
rect 20188 3266 20244 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 18284 2902 18340 2940
rect 19180 2996 19236 3006
rect 19180 2902 19236 2940
rect 19628 2996 19684 3006
rect 19628 2770 19684 2940
rect 20300 2882 20356 3276
rect 20300 2830 20302 2882
rect 20354 2830 20356 2882
rect 20300 2818 20356 2830
rect 19628 2718 19630 2770
rect 19682 2718 19684 2770
rect 19628 2706 19684 2718
rect 22428 2772 22484 4958
rect 22652 3668 22708 5180
rect 23100 5124 23156 5964
rect 23660 5794 23716 11116
rect 24220 9940 24276 9950
rect 24220 9846 24276 9884
rect 23884 9604 23940 9614
rect 24332 9604 24388 12460
rect 24444 12290 24500 12302
rect 24444 12238 24446 12290
rect 24498 12238 24500 12290
rect 24444 11508 24500 12238
rect 24556 12180 24612 12190
rect 24780 12180 24836 13916
rect 25116 13636 25172 13646
rect 25116 13074 25172 13580
rect 25116 13022 25118 13074
rect 25170 13022 25172 13074
rect 25116 13010 25172 13022
rect 25788 12964 25844 12974
rect 25900 12964 25956 17390
rect 26572 16884 26628 19852
rect 27132 19796 27188 26852
rect 27244 26516 27300 26526
rect 27244 22484 27300 26460
rect 27580 26404 27636 26414
rect 27580 26310 27636 26348
rect 27580 24052 27636 24062
rect 27580 23938 27636 23996
rect 27692 24050 27748 27580
rect 27804 27074 27860 28366
rect 27916 27860 27972 27870
rect 27916 27858 28308 27860
rect 27916 27806 27918 27858
rect 27970 27806 28308 27858
rect 27916 27804 28308 27806
rect 27916 27794 27972 27804
rect 28252 27186 28308 27804
rect 28252 27134 28254 27186
rect 28306 27134 28308 27186
rect 28252 27122 28308 27134
rect 27804 27022 27806 27074
rect 27858 27022 27860 27074
rect 27804 26514 27860 27022
rect 27804 26462 27806 26514
rect 27858 26462 27860 26514
rect 27804 26450 27860 26462
rect 28252 26852 28308 26862
rect 28252 26404 28308 26796
rect 27916 26068 27972 26078
rect 27916 26066 28084 26068
rect 27916 26014 27918 26066
rect 27970 26014 28084 26066
rect 27916 26012 28084 26014
rect 27916 26002 27972 26012
rect 27692 23998 27694 24050
rect 27746 23998 27748 24050
rect 27692 23986 27748 23998
rect 27804 24052 27860 24062
rect 27580 23886 27582 23938
rect 27634 23886 27636 23938
rect 27580 23874 27636 23886
rect 27804 23938 27860 23996
rect 27804 23886 27806 23938
rect 27858 23886 27860 23938
rect 27804 23874 27860 23886
rect 27916 23940 27972 23950
rect 27916 23846 27972 23884
rect 27356 23826 27412 23838
rect 27356 23774 27358 23826
rect 27410 23774 27412 23826
rect 27356 22708 27412 23774
rect 28028 23492 28084 26012
rect 28252 25618 28308 26348
rect 28252 25566 28254 25618
rect 28306 25566 28308 25618
rect 28252 25554 28308 25566
rect 27804 23436 28084 23492
rect 28252 24052 28308 24062
rect 27804 23266 27860 23436
rect 27804 23214 27806 23266
rect 27858 23214 27860 23266
rect 27804 23202 27860 23214
rect 27356 22642 27412 22652
rect 27244 22428 27412 22484
rect 27244 22260 27300 22270
rect 27244 22166 27300 22204
rect 26908 19740 27188 19796
rect 26908 18788 26964 19740
rect 27020 19460 27076 19470
rect 27356 19460 27412 22428
rect 28252 22482 28308 23996
rect 28252 22430 28254 22482
rect 28306 22430 28308 22482
rect 28252 22418 28308 22430
rect 28028 22370 28084 22382
rect 28028 22318 28030 22370
rect 28082 22318 28084 22370
rect 27692 22148 27748 22158
rect 28028 22148 28084 22318
rect 27692 22146 27972 22148
rect 27692 22094 27694 22146
rect 27746 22094 27972 22146
rect 27692 22092 27972 22094
rect 27692 22082 27748 22092
rect 27916 20802 27972 22092
rect 28028 22082 28084 22092
rect 28140 21476 28196 21486
rect 28140 21382 28196 21420
rect 27916 20750 27918 20802
rect 27970 20750 27972 20802
rect 27916 20738 27972 20750
rect 27692 20578 27748 20590
rect 27692 20526 27694 20578
rect 27746 20526 27748 20578
rect 27692 20130 27748 20526
rect 27692 20078 27694 20130
rect 27746 20078 27748 20130
rect 27692 20066 27748 20078
rect 27020 19458 27412 19460
rect 27020 19406 27022 19458
rect 27074 19406 27412 19458
rect 27020 19404 27412 19406
rect 27020 19394 27076 19404
rect 27132 19124 27188 19134
rect 27132 19122 28196 19124
rect 27132 19070 27134 19122
rect 27186 19070 28196 19122
rect 27132 19068 28196 19070
rect 27132 19058 27188 19068
rect 26908 18732 27076 18788
rect 26908 17444 26964 17454
rect 26908 17350 26964 17388
rect 26684 16884 26740 16894
rect 26572 16828 26684 16884
rect 26684 13636 26740 16828
rect 27020 15148 27076 18732
rect 28140 18338 28196 19068
rect 28140 18286 28142 18338
rect 28194 18286 28196 18338
rect 28140 18274 28196 18286
rect 27356 17444 27412 17454
rect 27356 17350 27412 17388
rect 28028 16884 28084 16894
rect 28028 16790 28084 16828
rect 27356 16772 27412 16782
rect 27356 16678 27412 16716
rect 28252 15426 28308 15438
rect 28252 15374 28254 15426
rect 28306 15374 28308 15426
rect 28252 15148 28308 15374
rect 27020 15092 27300 15148
rect 27132 14084 27188 14094
rect 26684 13542 26740 13580
rect 27020 14028 27132 14084
rect 25788 12962 25956 12964
rect 25788 12910 25790 12962
rect 25842 12910 25956 12962
rect 25788 12908 25956 12910
rect 25788 12898 25844 12908
rect 26012 12740 26068 12750
rect 26012 12646 26068 12684
rect 24556 12178 24836 12180
rect 24556 12126 24558 12178
rect 24610 12126 24836 12178
rect 24556 12124 24836 12126
rect 25228 12180 25284 12190
rect 24556 12114 24612 12124
rect 24444 9938 24500 11452
rect 24668 11506 24724 12124
rect 25228 12066 25284 12124
rect 25228 12014 25230 12066
rect 25282 12014 25284 12066
rect 25228 12002 25284 12014
rect 24668 11454 24670 11506
rect 24722 11454 24724 11506
rect 24668 11442 24724 11454
rect 25116 11732 25172 11742
rect 25116 11506 25172 11676
rect 25116 11454 25118 11506
rect 25170 11454 25172 11506
rect 25116 11442 25172 11454
rect 25452 11508 25508 11518
rect 25452 11414 25508 11452
rect 24444 9886 24446 9938
rect 24498 9886 24500 9938
rect 24444 9874 24500 9886
rect 25900 11396 25956 11406
rect 23884 9602 24052 9604
rect 23884 9550 23886 9602
rect 23938 9550 24052 9602
rect 23884 9548 24052 9550
rect 23884 9538 23940 9548
rect 23996 9154 24052 9548
rect 23996 9102 23998 9154
rect 24050 9102 24052 9154
rect 23996 9090 24052 9102
rect 24220 9548 24388 9604
rect 23660 5742 23662 5794
rect 23714 5742 23716 5794
rect 23660 5730 23716 5742
rect 23884 5908 23940 5918
rect 23100 5010 23156 5068
rect 23324 5348 23380 5358
rect 23324 5236 23380 5292
rect 23884 5236 23940 5852
rect 23324 5234 23940 5236
rect 23324 5182 23886 5234
rect 23938 5182 23940 5234
rect 23324 5180 23940 5182
rect 23324 5122 23380 5180
rect 23884 5170 23940 5180
rect 23324 5070 23326 5122
rect 23378 5070 23380 5122
rect 23324 5058 23380 5070
rect 23100 4958 23102 5010
rect 23154 4958 23156 5010
rect 23100 4946 23156 4958
rect 23436 5012 23492 5022
rect 23436 4918 23492 4956
rect 24220 5012 24276 9548
rect 24332 9154 24388 9166
rect 24332 9102 24334 9154
rect 24386 9102 24388 9154
rect 24332 8428 24388 9102
rect 24332 8372 25172 8428
rect 25116 8370 25172 8372
rect 25116 8318 25118 8370
rect 25170 8318 25172 8370
rect 25116 8306 25172 8318
rect 25900 8258 25956 11340
rect 26572 9716 26628 9726
rect 26572 9266 26628 9660
rect 26572 9214 26574 9266
rect 26626 9214 26628 9266
rect 26572 8428 26628 9214
rect 26908 9044 26964 9054
rect 26908 8950 26964 8988
rect 27020 8930 27076 14028
rect 27132 14018 27188 14028
rect 27132 13746 27188 13758
rect 27132 13694 27134 13746
rect 27186 13694 27188 13746
rect 27132 13636 27188 13694
rect 27132 13570 27188 13580
rect 27020 8878 27022 8930
rect 27074 8878 27076 8930
rect 27020 8866 27076 8878
rect 27132 9042 27188 9054
rect 27132 8990 27134 9042
rect 27186 8990 27188 9042
rect 27132 8932 27188 8990
rect 27132 8866 27188 8876
rect 27244 8708 27300 15092
rect 27804 15092 28308 15148
rect 27804 13858 27860 15092
rect 28364 14084 28420 36204
rect 28588 32900 28644 36652
rect 28588 32834 28644 32844
rect 28588 32676 28644 32686
rect 28588 32582 28644 32620
rect 28476 32562 28532 32574
rect 28476 32510 28478 32562
rect 28530 32510 28532 32562
rect 28476 32452 28532 32510
rect 28476 32396 28644 32452
rect 28588 32002 28644 32396
rect 28588 31950 28590 32002
rect 28642 31950 28644 32002
rect 28588 31938 28644 31950
rect 28476 31666 28532 31678
rect 28476 31614 28478 31666
rect 28530 31614 28532 31666
rect 28476 27636 28532 31614
rect 28700 31332 28756 38670
rect 28924 38276 28980 40012
rect 28924 38210 28980 38220
rect 28924 38052 28980 38062
rect 28812 37156 28868 37166
rect 28812 34018 28868 37100
rect 28924 35140 28980 37996
rect 29148 37380 29204 43708
rect 29372 43652 29428 43662
rect 29260 43428 29316 43438
rect 29260 42866 29316 43372
rect 29260 42814 29262 42866
rect 29314 42814 29316 42866
rect 29260 42420 29316 42814
rect 29260 42354 29316 42364
rect 29260 42082 29316 42094
rect 29260 42030 29262 42082
rect 29314 42030 29316 42082
rect 29260 41188 29316 42030
rect 29372 41970 29428 43596
rect 29372 41918 29374 41970
rect 29426 41918 29428 41970
rect 29372 41906 29428 41918
rect 29596 41300 29652 45726
rect 29596 41234 29652 41244
rect 29260 41122 29316 41132
rect 29708 41186 29764 48300
rect 29820 47572 29876 47582
rect 29820 47478 29876 47516
rect 29932 47236 29988 56252
rect 30044 54740 30100 54750
rect 30044 47460 30100 54684
rect 30156 54514 30212 54526
rect 30156 54462 30158 54514
rect 30210 54462 30212 54514
rect 30156 53956 30212 54462
rect 30156 53890 30212 53900
rect 30156 53730 30212 53742
rect 30156 53678 30158 53730
rect 30210 53678 30212 53730
rect 30156 52948 30212 53678
rect 30156 52882 30212 52892
rect 30268 51268 30324 57148
rect 30268 51174 30324 51212
rect 30380 51044 30436 58044
rect 30716 57540 30772 57550
rect 30716 57446 30772 57484
rect 30716 56980 30772 56990
rect 30772 56924 31108 56980
rect 30716 56886 30772 56924
rect 31052 56866 31108 56924
rect 31052 56814 31054 56866
rect 31106 56814 31108 56866
rect 31052 56802 31108 56814
rect 31164 56308 31220 60508
rect 31612 60452 31668 67564
rect 32060 65492 32116 65502
rect 32060 65398 32116 65436
rect 32396 65380 32452 69132
rect 32508 67284 32564 69470
rect 32956 69188 33012 69198
rect 32956 69094 33012 69132
rect 33068 68740 33124 68750
rect 32620 68738 33124 68740
rect 32620 68686 33070 68738
rect 33122 68686 33124 68738
rect 32620 68684 33124 68686
rect 32620 67954 32676 68684
rect 33068 68674 33124 68684
rect 32620 67902 32622 67954
rect 32674 67902 32676 67954
rect 32620 67890 32676 67902
rect 32508 67228 32788 67284
rect 32620 66946 32676 66958
rect 32620 66894 32622 66946
rect 32674 66894 32676 66946
rect 32620 66836 32676 66894
rect 32732 66948 32788 67228
rect 33292 67172 33348 70814
rect 33628 70196 33684 70206
rect 33628 70082 33684 70140
rect 33628 70030 33630 70082
rect 33682 70030 33684 70082
rect 33628 69188 33684 70030
rect 33852 70084 33908 71038
rect 33964 71428 34020 71438
rect 33964 70420 34020 71372
rect 34076 70420 34132 70430
rect 33964 70418 34468 70420
rect 33964 70366 34078 70418
rect 34130 70366 34468 70418
rect 33964 70364 34468 70366
rect 34076 70354 34132 70364
rect 34412 70306 34468 70364
rect 34412 70254 34414 70306
rect 34466 70254 34468 70306
rect 34412 70242 34468 70254
rect 33852 70028 34020 70084
rect 33628 69122 33684 69132
rect 33852 69412 33908 69422
rect 33404 68628 33460 68638
rect 33404 68626 33572 68628
rect 33404 68574 33406 68626
rect 33458 68574 33572 68626
rect 33404 68572 33572 68574
rect 33404 68562 33460 68572
rect 33516 67172 33572 68572
rect 33628 67172 33684 67182
rect 33292 67116 33460 67172
rect 33516 67170 33684 67172
rect 33516 67118 33630 67170
rect 33682 67118 33684 67170
rect 33516 67116 33684 67118
rect 33068 66948 33124 66958
rect 32732 66946 33124 66948
rect 32732 66894 33070 66946
rect 33122 66894 33124 66946
rect 32732 66892 33124 66894
rect 32620 65492 32676 66780
rect 32956 65492 33012 66892
rect 33068 66882 33124 66892
rect 33292 66836 33348 66846
rect 33292 66742 33348 66780
rect 33068 65492 33124 65502
rect 32956 65436 33068 65492
rect 33404 65492 33460 67116
rect 33628 67106 33684 67116
rect 33740 67060 33796 67070
rect 33628 66498 33684 66510
rect 33628 66446 33630 66498
rect 33682 66446 33684 66498
rect 33628 66386 33684 66446
rect 33628 66334 33630 66386
rect 33682 66334 33684 66386
rect 33628 66322 33684 66334
rect 33404 65436 33684 65492
rect 32620 65426 32676 65436
rect 33068 65426 33124 65436
rect 32508 65380 32564 65390
rect 32396 65378 32564 65380
rect 32396 65326 32510 65378
rect 32562 65326 32564 65378
rect 32396 65324 32564 65326
rect 32284 64820 32340 64830
rect 32284 64818 32452 64820
rect 32284 64766 32286 64818
rect 32338 64766 32452 64818
rect 32284 64764 32452 64766
rect 32284 64754 32340 64764
rect 31948 64036 32004 64046
rect 31948 63250 32004 63980
rect 31948 63198 31950 63250
rect 32002 63198 32004 63250
rect 31724 62356 31780 62366
rect 31724 62262 31780 62300
rect 31948 62188 32004 63198
rect 32396 63252 32452 64764
rect 32396 63138 32452 63196
rect 32396 63086 32398 63138
rect 32450 63086 32452 63138
rect 32396 63074 32452 63086
rect 32508 63924 32564 65324
rect 33180 65268 33236 65278
rect 33516 65268 33572 65278
rect 33180 65266 33460 65268
rect 33180 65214 33182 65266
rect 33234 65214 33460 65266
rect 33180 65212 33460 65214
rect 33180 65202 33236 65212
rect 32844 64706 32900 64718
rect 32844 64654 32846 64706
rect 32898 64654 32900 64706
rect 32844 64148 32900 64654
rect 32844 63924 32900 64092
rect 32508 63922 32900 63924
rect 32508 63870 32510 63922
rect 32562 63870 32900 63922
rect 32508 63868 32900 63870
rect 32956 64036 33012 64046
rect 33404 64036 33460 65212
rect 33516 65174 33572 65212
rect 33628 65044 33684 65436
rect 33740 65490 33796 67004
rect 33740 65438 33742 65490
rect 33794 65438 33796 65490
rect 33740 65426 33796 65438
rect 33852 65268 33908 69356
rect 33964 69188 34020 70028
rect 34524 69412 34580 73892
rect 34972 73108 35028 73118
rect 34860 72770 34916 72782
rect 34860 72718 34862 72770
rect 34914 72718 34916 72770
rect 34748 72322 34804 72334
rect 34748 72270 34750 72322
rect 34802 72270 34804 72322
rect 34748 71764 34804 72270
rect 34748 71698 34804 71708
rect 34860 71762 34916 72718
rect 34860 71710 34862 71762
rect 34914 71710 34916 71762
rect 34860 71090 34916 71710
rect 34860 71038 34862 71090
rect 34914 71038 34916 71090
rect 34636 70308 34692 70318
rect 34636 70214 34692 70252
rect 34748 70084 34804 70094
rect 34860 70084 34916 71038
rect 34972 70978 35028 73052
rect 35084 71762 35140 74956
rect 35196 74946 35252 74956
rect 35756 74786 35812 74798
rect 35756 74734 35758 74786
rect 35810 74734 35812 74786
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 35756 74226 35812 74734
rect 35756 74174 35758 74226
rect 35810 74174 35812 74226
rect 35756 74162 35812 74174
rect 35644 74114 35700 74126
rect 35644 74062 35646 74114
rect 35698 74062 35700 74114
rect 35308 74004 35364 74014
rect 35308 73910 35364 73948
rect 35644 73892 35700 74062
rect 35980 74004 36036 74014
rect 35980 73910 36036 73948
rect 35644 73108 35700 73836
rect 36316 73892 36372 75406
rect 36988 75012 37044 75022
rect 36988 74338 37044 74956
rect 37884 74788 37940 74798
rect 36988 74286 36990 74338
rect 37042 74286 37044 74338
rect 36988 74274 37044 74286
rect 37100 74786 37940 74788
rect 37100 74734 37886 74786
rect 37938 74734 37940 74786
rect 37100 74732 37940 74734
rect 37100 74226 37156 74732
rect 37884 74722 37940 74732
rect 37100 74174 37102 74226
rect 37154 74174 37156 74226
rect 37100 74162 37156 74174
rect 36316 73826 36372 73836
rect 37436 74004 37492 74014
rect 35644 73042 35700 73052
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 35196 72770 35252 72782
rect 35196 72718 35198 72770
rect 35250 72718 35252 72770
rect 35196 72658 35252 72718
rect 35196 72606 35198 72658
rect 35250 72606 35252 72658
rect 35196 72594 35252 72606
rect 37100 72322 37156 72334
rect 37100 72270 37102 72322
rect 37154 72270 37156 72322
rect 37100 71876 37156 72270
rect 37100 71810 37156 71820
rect 37436 72324 37492 73948
rect 37548 72324 37604 72334
rect 37436 72322 37604 72324
rect 37436 72270 37550 72322
rect 37602 72270 37604 72322
rect 37436 72268 37604 72270
rect 35084 71710 35086 71762
rect 35138 71710 35140 71762
rect 35084 71698 35140 71710
rect 35980 71764 36036 71774
rect 36092 71764 36148 71774
rect 36036 71762 36148 71764
rect 36036 71710 36094 71762
rect 36146 71710 36148 71762
rect 36036 71708 36148 71710
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 34972 70926 34974 70978
rect 35026 70926 35028 70978
rect 34972 70914 35028 70926
rect 35980 70978 36036 71708
rect 36092 71698 36148 71708
rect 36428 71764 36484 71774
rect 36204 71538 36260 71550
rect 36204 71486 36206 71538
rect 36258 71486 36260 71538
rect 35980 70926 35982 70978
rect 36034 70926 36036 70978
rect 35084 70644 35140 70654
rect 35084 70196 35140 70588
rect 35084 70102 35140 70140
rect 35644 70308 35700 70318
rect 34860 70028 35028 70084
rect 34748 69990 34804 70028
rect 34972 69522 35028 70028
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 34972 69470 34974 69522
rect 35026 69470 35028 69522
rect 34860 69412 34916 69422
rect 34524 69410 34916 69412
rect 34524 69358 34862 69410
rect 34914 69358 34916 69410
rect 34524 69356 34916 69358
rect 34860 69346 34916 69356
rect 34188 69188 34244 69198
rect 34972 69188 35028 69470
rect 35644 69412 35700 70252
rect 35868 70084 35924 70094
rect 35868 69990 35924 70028
rect 35980 69860 36036 70926
rect 33964 69186 35028 69188
rect 33964 69134 34190 69186
rect 34242 69134 35028 69186
rect 33964 69132 35028 69134
rect 35532 69410 35700 69412
rect 35532 69358 35646 69410
rect 35698 69358 35700 69410
rect 35532 69356 35700 69358
rect 33964 66948 34020 66958
rect 33964 66052 34020 66892
rect 34076 66276 34132 69132
rect 34188 69122 34244 69132
rect 35532 68850 35588 69356
rect 35644 69346 35700 69356
rect 35868 69804 36036 69860
rect 36092 71202 36148 71214
rect 36092 71150 36094 71202
rect 36146 71150 36148 71202
rect 35868 69412 35924 69804
rect 35868 69318 35924 69356
rect 35980 69634 36036 69646
rect 35980 69582 35982 69634
rect 36034 69582 36036 69634
rect 35532 68798 35534 68850
rect 35586 68798 35588 68850
rect 35532 68786 35588 68798
rect 35644 68516 35700 68526
rect 35644 68514 35924 68516
rect 35644 68462 35646 68514
rect 35698 68462 35924 68514
rect 35644 68460 35924 68462
rect 35644 68450 35700 68460
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 34748 67954 34804 67966
rect 34748 67902 34750 67954
rect 34802 67902 34804 67954
rect 34748 67060 34804 67902
rect 34748 66994 34804 67004
rect 35084 67170 35140 67182
rect 35084 67118 35086 67170
rect 35138 67118 35140 67170
rect 34188 66948 34244 66958
rect 34188 66854 34244 66892
rect 34524 66946 34580 66958
rect 34524 66894 34526 66946
rect 34578 66894 34580 66946
rect 34524 66836 34580 66894
rect 35084 66836 35140 67118
rect 35308 67060 35364 67070
rect 35308 66966 35364 67004
rect 34300 66780 35140 66836
rect 34188 66500 34244 66510
rect 34300 66500 34356 66780
rect 34188 66498 34356 66500
rect 34188 66446 34190 66498
rect 34242 66446 34356 66498
rect 34188 66444 34356 66446
rect 34188 66434 34244 66444
rect 34076 66220 34356 66276
rect 34076 66052 34132 66062
rect 33964 66050 34132 66052
rect 33964 65998 34078 66050
rect 34130 65998 34132 66050
rect 33964 65996 34132 65998
rect 34076 65986 34132 65996
rect 34188 65492 34244 65502
rect 34188 65398 34244 65436
rect 33852 65212 34244 65268
rect 33516 64988 33684 65044
rect 33516 64260 33572 64988
rect 33628 64596 33684 64606
rect 33628 64594 33908 64596
rect 33628 64542 33630 64594
rect 33682 64542 33908 64594
rect 33628 64540 33908 64542
rect 33628 64530 33684 64540
rect 33516 64204 33684 64260
rect 33516 64036 33572 64046
rect 33404 64034 33572 64036
rect 33404 63982 33518 64034
rect 33570 63982 33572 64034
rect 33404 63980 33572 63982
rect 32508 62356 32564 63868
rect 32956 63026 33012 63980
rect 33516 63970 33572 63980
rect 33180 63922 33236 63934
rect 33180 63870 33182 63922
rect 33234 63870 33236 63922
rect 33180 63252 33236 63870
rect 33180 63186 33236 63196
rect 33628 63140 33684 64204
rect 33852 64146 33908 64540
rect 33852 64094 33854 64146
rect 33906 64094 33908 64146
rect 33852 64082 33908 64094
rect 34076 63252 34132 63262
rect 33964 63140 34020 63150
rect 33628 63138 34020 63140
rect 33628 63086 33966 63138
rect 34018 63086 34020 63138
rect 33628 63084 34020 63086
rect 33964 63074 34020 63084
rect 32956 62974 32958 63026
rect 33010 62974 33012 63026
rect 32956 62962 33012 62974
rect 33180 63028 33236 63038
rect 32564 62300 32900 62356
rect 32508 62290 32564 62300
rect 31948 62132 32340 62188
rect 32172 60900 32228 60910
rect 31276 60396 31668 60452
rect 31948 60898 32228 60900
rect 31948 60846 32174 60898
rect 32226 60846 32228 60898
rect 31948 60844 32228 60846
rect 31276 60116 31332 60396
rect 31276 60002 31332 60060
rect 31276 59950 31278 60002
rect 31330 59950 31332 60002
rect 31276 59938 31332 59950
rect 31836 59890 31892 59902
rect 31836 59838 31838 59890
rect 31890 59838 31892 59890
rect 31836 59780 31892 59838
rect 31836 59714 31892 59724
rect 31948 59556 32004 60844
rect 32172 60834 32228 60844
rect 32284 60676 32340 62132
rect 32620 61348 32676 61358
rect 32508 61346 32676 61348
rect 32508 61294 32622 61346
rect 32674 61294 32676 61346
rect 32508 61292 32676 61294
rect 32508 60898 32564 61292
rect 32620 61282 32676 61292
rect 32508 60846 32510 60898
rect 32562 60846 32564 60898
rect 32508 60834 32564 60846
rect 32844 60788 32900 62300
rect 32956 62132 33012 62142
rect 32956 61794 33012 62076
rect 32956 61742 32958 61794
rect 33010 61742 33012 61794
rect 32956 61730 33012 61742
rect 33180 61682 33236 62972
rect 33180 61630 33182 61682
rect 33234 61630 33236 61682
rect 33180 61618 33236 61630
rect 33628 62132 33684 62142
rect 33628 61682 33684 62076
rect 33628 61630 33630 61682
rect 33682 61630 33684 61682
rect 33628 61618 33684 61630
rect 33180 60788 33236 60798
rect 32844 60786 33236 60788
rect 32844 60734 33182 60786
rect 33234 60734 33236 60786
rect 32844 60732 33236 60734
rect 31612 59500 32004 59556
rect 32060 60620 32340 60676
rect 31612 58546 31668 59500
rect 31612 58494 31614 58546
rect 31666 58494 31668 58546
rect 31612 58482 31668 58494
rect 31612 58324 31668 58334
rect 31668 58268 31892 58324
rect 31612 58258 31668 58268
rect 31836 57762 31892 58268
rect 31836 57710 31838 57762
rect 31890 57710 31892 57762
rect 31836 57698 31892 57710
rect 31500 57650 31556 57662
rect 32060 57652 32116 60620
rect 32732 59780 32788 59790
rect 32732 59686 32788 59724
rect 33180 59780 33236 60732
rect 33852 60676 33908 60686
rect 33180 59714 33236 59724
rect 33404 60674 33908 60676
rect 33404 60622 33854 60674
rect 33906 60622 33908 60674
rect 33404 60620 33908 60622
rect 33404 59442 33460 60620
rect 33852 60610 33908 60620
rect 33404 59390 33406 59442
rect 33458 59390 33460 59442
rect 33404 59378 33460 59390
rect 33068 59220 33124 59230
rect 32508 59218 33124 59220
rect 32508 59166 33070 59218
rect 33122 59166 33124 59218
rect 32508 59164 33124 59166
rect 32284 58548 32340 58558
rect 32284 57874 32340 58492
rect 32284 57822 32286 57874
rect 32338 57822 32340 57874
rect 32284 57810 32340 57822
rect 32396 57876 32452 57886
rect 32396 57782 32452 57820
rect 31500 57598 31502 57650
rect 31554 57598 31556 57650
rect 31500 57204 31556 57598
rect 31500 57138 31556 57148
rect 31948 57596 32060 57652
rect 31164 56252 31332 56308
rect 30492 54628 30548 54638
rect 30492 54626 30996 54628
rect 30492 54574 30494 54626
rect 30546 54574 30996 54626
rect 30492 54572 30996 54574
rect 30492 54562 30548 54572
rect 30940 53842 30996 54572
rect 30940 53790 30942 53842
rect 30994 53790 30996 53842
rect 30940 53778 30996 53790
rect 30716 52276 30772 52286
rect 30716 52182 30772 52220
rect 31164 51938 31220 51950
rect 31164 51886 31166 51938
rect 31218 51886 31220 51938
rect 30716 51604 30772 51614
rect 30716 51510 30772 51548
rect 31052 51268 31108 51278
rect 30268 50988 30436 51044
rect 30604 51154 30660 51166
rect 30604 51102 30606 51154
rect 30658 51102 30660 51154
rect 30156 50708 30212 50718
rect 30156 49698 30212 50652
rect 30156 49646 30158 49698
rect 30210 49646 30212 49698
rect 30156 49634 30212 49646
rect 30268 49140 30324 50988
rect 30492 50594 30548 50606
rect 30492 50542 30494 50594
rect 30546 50542 30548 50594
rect 30380 50370 30436 50382
rect 30380 50318 30382 50370
rect 30434 50318 30436 50370
rect 30380 49812 30436 50318
rect 30492 49924 30548 50542
rect 30492 49858 30548 49868
rect 30380 49252 30436 49756
rect 30380 49186 30436 49196
rect 30492 49700 30548 49710
rect 30156 49084 30324 49140
rect 30156 48692 30212 49084
rect 30268 48916 30324 48926
rect 30268 48822 30324 48860
rect 30380 48914 30436 48926
rect 30380 48862 30382 48914
rect 30434 48862 30436 48914
rect 30156 48636 30324 48692
rect 30044 47394 30100 47404
rect 29932 47180 30100 47236
rect 29932 47012 29988 47022
rect 29820 46564 29876 46574
rect 29820 46450 29876 46508
rect 29820 46398 29822 46450
rect 29874 46398 29876 46450
rect 29820 46386 29876 46398
rect 29932 45890 29988 46956
rect 29932 45838 29934 45890
rect 29986 45838 29988 45890
rect 29932 45826 29988 45838
rect 29932 45108 29988 45118
rect 29820 45106 29988 45108
rect 29820 45054 29934 45106
rect 29986 45054 29988 45106
rect 29820 45052 29988 45054
rect 29820 43764 29876 45052
rect 29932 45042 29988 45052
rect 29820 43698 29876 43708
rect 29932 44660 29988 44670
rect 29820 42980 29876 42990
rect 29820 42866 29876 42924
rect 29820 42814 29822 42866
rect 29874 42814 29876 42866
rect 29820 42802 29876 42814
rect 29932 42532 29988 44604
rect 30044 43652 30100 47180
rect 30156 47234 30212 47246
rect 30156 47182 30158 47234
rect 30210 47182 30212 47234
rect 30156 45892 30212 47182
rect 30156 45826 30212 45836
rect 30156 45666 30212 45678
rect 30156 45614 30158 45666
rect 30210 45614 30212 45666
rect 30156 43764 30212 45614
rect 30156 43698 30212 43708
rect 30044 43586 30100 43596
rect 30044 43428 30100 43438
rect 30044 43426 30212 43428
rect 30044 43374 30046 43426
rect 30098 43374 30212 43426
rect 30044 43372 30212 43374
rect 30044 43362 30100 43372
rect 30044 42532 30100 42542
rect 29932 42476 30044 42532
rect 30044 42466 30100 42476
rect 30044 41972 30100 41982
rect 30044 41878 30100 41916
rect 29932 41300 29988 41310
rect 29932 41206 29988 41244
rect 29708 41134 29710 41186
rect 29762 41134 29764 41186
rect 29260 40962 29316 40974
rect 29260 40910 29262 40962
rect 29314 40910 29316 40962
rect 29260 40852 29316 40910
rect 29708 40852 29764 41134
rect 30044 41188 30100 41198
rect 30156 41188 30212 43372
rect 30268 43204 30324 48636
rect 30380 48132 30436 48862
rect 30380 48066 30436 48076
rect 30492 48914 30548 49644
rect 30492 48862 30494 48914
rect 30546 48862 30548 48914
rect 30492 46676 30548 48862
rect 30604 48132 30660 51102
rect 30604 48066 30660 48076
rect 30716 50596 30772 50606
rect 30492 46610 30548 46620
rect 30380 46562 30436 46574
rect 30380 46510 30382 46562
rect 30434 46510 30436 46562
rect 30380 45890 30436 46510
rect 30604 46450 30660 46462
rect 30604 46398 30606 46450
rect 30658 46398 30660 46450
rect 30604 46228 30660 46398
rect 30716 46452 30772 50540
rect 30828 50036 30884 50046
rect 30828 49810 30884 49980
rect 31052 50034 31108 51212
rect 31164 50708 31220 51886
rect 31164 50642 31220 50652
rect 31052 49982 31054 50034
rect 31106 49982 31108 50034
rect 31052 49970 31108 49982
rect 31164 50260 31220 50270
rect 31164 50034 31220 50204
rect 31276 50148 31332 56252
rect 31388 52836 31444 52846
rect 31836 52836 31892 52846
rect 31388 52834 31892 52836
rect 31388 52782 31390 52834
rect 31442 52782 31838 52834
rect 31890 52782 31892 52834
rect 31388 52780 31892 52782
rect 31388 52770 31444 52780
rect 31388 51604 31444 51614
rect 31444 51548 31556 51604
rect 31388 51538 31444 51548
rect 31388 51266 31444 51278
rect 31388 51214 31390 51266
rect 31442 51214 31444 51266
rect 31388 51154 31444 51214
rect 31388 51102 31390 51154
rect 31442 51102 31444 51154
rect 31388 51090 31444 51102
rect 31500 50932 31556 51548
rect 31276 50082 31332 50092
rect 31388 50876 31556 50932
rect 31164 49982 31166 50034
rect 31218 49982 31220 50034
rect 31164 49970 31220 49982
rect 31276 49924 31332 49934
rect 31276 49830 31332 49868
rect 30828 49758 30830 49810
rect 30882 49758 30884 49810
rect 30828 49746 30884 49758
rect 31388 49810 31444 50876
rect 31500 50708 31556 50718
rect 31500 50482 31556 50652
rect 31500 50430 31502 50482
rect 31554 50430 31556 50482
rect 31500 50418 31556 50430
rect 31388 49758 31390 49810
rect 31442 49758 31444 49810
rect 31388 49746 31444 49758
rect 31052 49588 31108 49598
rect 31276 49588 31332 49598
rect 31052 49138 31108 49532
rect 31052 49086 31054 49138
rect 31106 49086 31108 49138
rect 31052 47348 31108 49086
rect 31052 47282 31108 47292
rect 31164 49532 31276 49588
rect 30716 46386 30772 46396
rect 30604 46172 30772 46228
rect 30380 45838 30382 45890
rect 30434 45838 30436 45890
rect 30380 45444 30436 45838
rect 30716 45780 30772 46172
rect 30716 45686 30772 45724
rect 30380 45378 30436 45388
rect 30604 45666 30660 45678
rect 30604 45614 30606 45666
rect 30658 45614 30660 45666
rect 30604 45444 30660 45614
rect 30604 45388 30996 45444
rect 30492 45220 30548 45230
rect 30492 45126 30548 45164
rect 30380 44436 30436 44446
rect 30380 44210 30436 44380
rect 30604 44322 30660 45388
rect 30940 45106 30996 45388
rect 31164 45332 31220 49532
rect 31276 49522 31332 49532
rect 31500 48802 31556 48814
rect 31500 48750 31502 48802
rect 31554 48750 31556 48802
rect 31500 48244 31556 48750
rect 31388 48132 31444 48142
rect 31388 47572 31444 48076
rect 31388 47346 31444 47516
rect 31500 47458 31556 48188
rect 31500 47406 31502 47458
rect 31554 47406 31556 47458
rect 31500 47394 31556 47406
rect 31388 47294 31390 47346
rect 31442 47294 31444 47346
rect 31388 47282 31444 47294
rect 31276 45892 31332 45902
rect 31276 45798 31332 45836
rect 31164 45238 31220 45276
rect 31500 45780 31556 45790
rect 30940 45054 30942 45106
rect 30994 45054 30996 45106
rect 30940 45042 30996 45054
rect 31388 45106 31444 45118
rect 31388 45054 31390 45106
rect 31442 45054 31444 45106
rect 30604 44270 30606 44322
rect 30658 44270 30660 44322
rect 30604 44258 30660 44270
rect 31276 44994 31332 45006
rect 31276 44942 31278 44994
rect 31330 44942 31332 44994
rect 30380 44158 30382 44210
rect 30434 44158 30436 44210
rect 30380 44146 30436 44158
rect 31164 44098 31220 44110
rect 31164 44046 31166 44098
rect 31218 44046 31220 44098
rect 30828 43764 30884 43774
rect 30380 43540 30436 43550
rect 30380 43446 30436 43484
rect 30716 43540 30772 43550
rect 30268 43148 30436 43204
rect 30268 42532 30324 42542
rect 30268 42438 30324 42476
rect 30268 42196 30324 42206
rect 30268 42082 30324 42140
rect 30268 42030 30270 42082
rect 30322 42030 30324 42082
rect 30268 42018 30324 42030
rect 30044 41186 30212 41188
rect 30044 41134 30046 41186
rect 30098 41134 30212 41186
rect 30044 41132 30212 41134
rect 30268 41858 30324 41870
rect 30268 41806 30270 41858
rect 30322 41806 30324 41858
rect 29820 40964 29876 40974
rect 29820 40870 29876 40908
rect 29260 38836 29316 40796
rect 29372 40796 29764 40852
rect 29372 39730 29428 40796
rect 29820 40740 29876 40750
rect 30044 40740 30100 41132
rect 30156 40964 30212 40974
rect 30156 40870 30212 40908
rect 29820 40514 29876 40684
rect 29820 40462 29822 40514
rect 29874 40462 29876 40514
rect 29820 40450 29876 40462
rect 29932 40684 30100 40740
rect 29372 39678 29374 39730
rect 29426 39678 29428 39730
rect 29372 39666 29428 39678
rect 29484 40402 29540 40414
rect 29484 40350 29486 40402
rect 29538 40350 29540 40402
rect 29484 39732 29540 40350
rect 29484 39666 29540 39676
rect 29596 40068 29652 40078
rect 29596 38946 29652 40012
rect 29932 39620 29988 40684
rect 30156 40404 30212 40414
rect 30156 40310 30212 40348
rect 30156 39844 30212 39854
rect 30156 39750 30212 39788
rect 29596 38894 29598 38946
rect 29650 38894 29652 38946
rect 29596 38882 29652 38894
rect 29820 39564 29988 39620
rect 30156 39620 30212 39630
rect 29260 38770 29316 38780
rect 29820 38668 29876 39564
rect 29932 39394 29988 39406
rect 29932 39342 29934 39394
rect 29986 39342 29988 39394
rect 29932 39172 29988 39342
rect 30044 39396 30100 39406
rect 30044 39302 30100 39340
rect 29932 39106 29988 39116
rect 29932 38836 29988 38846
rect 29988 38780 30100 38836
rect 29932 38770 29988 38780
rect 29372 38612 29876 38668
rect 29260 38276 29316 38286
rect 29260 38162 29316 38220
rect 29260 38110 29262 38162
rect 29314 38110 29316 38162
rect 29260 38098 29316 38110
rect 29260 37380 29316 37390
rect 29148 37378 29316 37380
rect 29148 37326 29262 37378
rect 29314 37326 29316 37378
rect 29148 37324 29316 37326
rect 29260 37314 29316 37324
rect 28924 35074 28980 35084
rect 29260 36258 29316 36270
rect 29260 36206 29262 36258
rect 29314 36206 29316 36258
rect 29260 34916 29316 36206
rect 29372 35588 29428 38612
rect 29932 38274 29988 38286
rect 29932 38222 29934 38274
rect 29986 38222 29988 38274
rect 29708 38164 29764 38174
rect 29708 38070 29764 38108
rect 29484 37492 29540 37502
rect 29484 37378 29540 37436
rect 29484 37326 29486 37378
rect 29538 37326 29540 37378
rect 29484 37314 29540 37326
rect 29596 37490 29652 37502
rect 29596 37438 29598 37490
rect 29650 37438 29652 37490
rect 29596 36482 29652 37438
rect 29820 37268 29876 37278
rect 29820 37174 29876 37212
rect 29596 36430 29598 36482
rect 29650 36430 29652 36482
rect 29596 36418 29652 36430
rect 29708 37042 29764 37054
rect 29708 36990 29710 37042
rect 29762 36990 29764 37042
rect 29596 35812 29652 35822
rect 29596 35718 29652 35756
rect 29372 35532 29652 35588
rect 28812 33966 28814 34018
rect 28866 33966 28868 34018
rect 28812 32116 28868 33966
rect 28812 32050 28868 32060
rect 28924 34860 29316 34916
rect 29484 35140 29540 35150
rect 28700 31266 28756 31276
rect 28812 30882 28868 30894
rect 28812 30830 28814 30882
rect 28866 30830 28868 30882
rect 28812 30772 28868 30830
rect 28588 29988 28644 29998
rect 28588 29894 28644 29932
rect 28812 29764 28868 30716
rect 28812 29698 28868 29708
rect 28476 27570 28532 27580
rect 28588 29652 28644 29662
rect 28476 27074 28532 27086
rect 28476 27022 28478 27074
rect 28530 27022 28532 27074
rect 28476 26964 28532 27022
rect 28476 26898 28532 26908
rect 28476 26628 28532 26638
rect 28476 26514 28532 26572
rect 28476 26462 28478 26514
rect 28530 26462 28532 26514
rect 28476 26404 28532 26462
rect 28476 26338 28532 26348
rect 28588 23548 28644 29596
rect 28812 29426 28868 29438
rect 28812 29374 28814 29426
rect 28866 29374 28868 29426
rect 28812 29204 28868 29374
rect 28812 29138 28868 29148
rect 28924 28084 28980 34860
rect 29148 34692 29204 34702
rect 29036 34468 29092 34478
rect 29036 34132 29092 34412
rect 29036 30772 29092 34076
rect 29148 34244 29204 34636
rect 29372 34692 29428 34702
rect 29148 31668 29204 34188
rect 29260 34356 29316 34366
rect 29372 34356 29428 34636
rect 29316 34300 29428 34356
rect 29260 34242 29316 34300
rect 29260 34190 29262 34242
rect 29314 34190 29316 34242
rect 29260 34178 29316 34190
rect 29372 34130 29428 34142
rect 29372 34078 29374 34130
rect 29426 34078 29428 34130
rect 29372 33796 29428 34078
rect 29372 33730 29428 33740
rect 29260 31892 29316 31902
rect 29260 31798 29316 31836
rect 29484 31778 29540 35084
rect 29484 31726 29486 31778
rect 29538 31726 29540 31778
rect 29484 31714 29540 31726
rect 29148 31612 29316 31668
rect 29148 30996 29204 31006
rect 29148 30902 29204 30940
rect 29036 30716 29204 30772
rect 29148 29428 29204 30716
rect 29148 29334 29204 29372
rect 29260 28756 29316 31612
rect 29372 31556 29428 31566
rect 29428 31500 29540 31556
rect 29372 31490 29428 31500
rect 29372 30772 29428 30782
rect 29372 30678 29428 30716
rect 29484 30434 29540 31500
rect 29484 30382 29486 30434
rect 29538 30382 29540 30434
rect 29484 30370 29540 30382
rect 29260 28690 29316 28700
rect 29372 29540 29428 29550
rect 28924 28018 28980 28028
rect 29036 27970 29092 27982
rect 29036 27918 29038 27970
rect 29090 27918 29092 27970
rect 28812 27188 28868 27198
rect 28812 26404 28868 27132
rect 29036 26628 29092 27918
rect 29260 27188 29316 27198
rect 29260 27074 29316 27132
rect 29372 27186 29428 29484
rect 29596 27524 29652 35532
rect 29708 34356 29764 36990
rect 29932 36820 29988 38222
rect 29932 36754 29988 36764
rect 29820 36484 29876 36494
rect 29820 36390 29876 36428
rect 30044 36148 30100 38780
rect 30156 37826 30212 39564
rect 30156 37774 30158 37826
rect 30210 37774 30212 37826
rect 30156 36708 30212 37774
rect 30156 36642 30212 36652
rect 30268 36596 30324 41806
rect 30380 36708 30436 43148
rect 30716 42866 30772 43484
rect 30716 42814 30718 42866
rect 30770 42814 30772 42866
rect 30716 42802 30772 42814
rect 30716 41972 30772 41982
rect 30604 41916 30716 41972
rect 30604 40180 30660 41916
rect 30716 41906 30772 41916
rect 30716 41186 30772 41198
rect 30716 41134 30718 41186
rect 30770 41134 30772 41186
rect 30716 40404 30772 41134
rect 30716 40338 30772 40348
rect 30716 40180 30772 40190
rect 30604 40178 30772 40180
rect 30604 40126 30718 40178
rect 30770 40126 30772 40178
rect 30604 40124 30772 40126
rect 30716 40114 30772 40124
rect 30604 39844 30660 39854
rect 30492 38946 30548 38958
rect 30492 38894 30494 38946
rect 30546 38894 30548 38946
rect 30492 38276 30548 38894
rect 30492 38210 30548 38220
rect 30604 38164 30660 39788
rect 30716 39394 30772 39406
rect 30716 39342 30718 39394
rect 30770 39342 30772 39394
rect 30716 38612 30772 39342
rect 30828 38834 30884 43708
rect 30940 43652 30996 43662
rect 30940 43558 30996 43596
rect 31164 43428 31220 44046
rect 31164 43362 31220 43372
rect 31164 43204 31220 43214
rect 31164 42866 31220 43148
rect 31164 42814 31166 42866
rect 31218 42814 31220 42866
rect 31164 41972 31220 42814
rect 31276 42868 31332 44942
rect 31388 43876 31444 45054
rect 31500 44996 31556 45724
rect 31612 45218 31668 52780
rect 31836 52770 31892 52780
rect 31836 51940 31892 51950
rect 31836 51846 31892 51884
rect 31836 51268 31892 51278
rect 31724 51266 31892 51268
rect 31724 51214 31838 51266
rect 31890 51214 31892 51266
rect 31724 51212 31892 51214
rect 31724 49028 31780 51212
rect 31836 51202 31892 51212
rect 31948 50428 32004 57596
rect 32060 57558 32116 57596
rect 32172 57538 32228 57550
rect 32172 57486 32174 57538
rect 32226 57486 32228 57538
rect 32060 57428 32116 57438
rect 32060 57090 32116 57372
rect 32060 57038 32062 57090
rect 32114 57038 32116 57090
rect 32060 52948 32116 57038
rect 32172 53060 32228 57486
rect 32508 55972 32564 59164
rect 33068 59154 33124 59164
rect 33740 58548 33796 58558
rect 33740 58454 33796 58492
rect 34076 57876 34132 63196
rect 33068 57652 33124 57662
rect 33124 57596 33236 57652
rect 33068 57586 33124 57596
rect 33180 57538 33236 57596
rect 33180 57486 33182 57538
rect 33234 57486 33236 57538
rect 33180 57474 33236 57486
rect 33740 57538 33796 57550
rect 33740 57486 33742 57538
rect 33794 57486 33796 57538
rect 33740 57204 33796 57486
rect 33740 57138 33796 57148
rect 33964 56644 34020 56654
rect 33740 56642 34020 56644
rect 33740 56590 33966 56642
rect 34018 56590 34020 56642
rect 33740 56588 34020 56590
rect 32284 55916 32564 55972
rect 33404 56194 33460 56206
rect 33404 56142 33406 56194
rect 33458 56142 33460 56194
rect 32284 53172 32340 55916
rect 33404 55412 33460 56142
rect 33740 56194 33796 56588
rect 33964 56578 34020 56588
rect 34076 56420 34132 57820
rect 33740 56142 33742 56194
rect 33794 56142 33796 56194
rect 33740 56130 33796 56142
rect 33964 56364 34132 56420
rect 33516 55412 33572 55422
rect 33404 55410 33572 55412
rect 33404 55358 33518 55410
rect 33570 55358 33572 55410
rect 33404 55356 33572 55358
rect 33516 55346 33572 55356
rect 32844 55298 32900 55310
rect 32844 55246 32846 55298
rect 32898 55246 32900 55298
rect 32396 55076 32452 55086
rect 32844 55076 32900 55246
rect 32396 55074 32900 55076
rect 32396 55022 32398 55074
rect 32450 55022 32900 55074
rect 32396 55020 32900 55022
rect 32396 55010 32452 55020
rect 32396 53172 32452 53182
rect 32284 53170 32452 53172
rect 32284 53118 32398 53170
rect 32450 53118 32452 53170
rect 32284 53116 32452 53118
rect 32396 53106 32452 53116
rect 32172 53004 32340 53060
rect 32284 52948 32340 53004
rect 32060 52892 32228 52948
rect 32284 52892 32676 52948
rect 32060 52724 32116 52734
rect 32060 52630 32116 52668
rect 31724 48962 31780 48972
rect 31836 50372 32004 50428
rect 31836 47124 31892 50372
rect 31948 49700 32004 49710
rect 32172 49700 32228 52892
rect 32284 51940 32340 51950
rect 32284 51846 32340 51884
rect 32004 49644 32228 49700
rect 32284 51266 32340 51278
rect 32284 51214 32286 51266
rect 32338 51214 32340 51266
rect 31948 49606 32004 49644
rect 32284 49028 32340 51214
rect 32396 50596 32452 50606
rect 32396 50502 32452 50540
rect 32508 49812 32564 49822
rect 32396 49700 32452 49710
rect 32396 49606 32452 49644
rect 32396 49028 32452 49038
rect 32284 49026 32452 49028
rect 32284 48974 32398 49026
rect 32450 48974 32452 49026
rect 32284 48972 32452 48974
rect 32172 47684 32228 47694
rect 32172 47458 32228 47628
rect 32172 47406 32174 47458
rect 32226 47406 32228 47458
rect 32172 47394 32228 47406
rect 32060 47348 32116 47358
rect 32060 47254 32116 47292
rect 31612 45166 31614 45218
rect 31666 45166 31668 45218
rect 31612 45154 31668 45166
rect 31724 47068 31892 47124
rect 31500 44940 31668 44996
rect 31388 43810 31444 43820
rect 31500 43428 31556 43438
rect 31276 42802 31332 42812
rect 31388 43426 31556 43428
rect 31388 43374 31502 43426
rect 31554 43374 31556 43426
rect 31388 43372 31556 43374
rect 31388 42644 31444 43372
rect 31500 43362 31556 43372
rect 31164 41906 31220 41916
rect 31276 42588 31444 42644
rect 31500 43092 31556 43102
rect 31276 40964 31332 42588
rect 31500 42532 31556 43036
rect 31276 40898 31332 40908
rect 31388 42196 31444 42206
rect 30828 38782 30830 38834
rect 30882 38782 30884 38834
rect 30828 38770 30884 38782
rect 30940 40068 30996 40078
rect 30716 38546 30772 38556
rect 30716 38164 30772 38174
rect 30604 38162 30772 38164
rect 30604 38110 30718 38162
rect 30770 38110 30772 38162
rect 30604 38108 30772 38110
rect 30716 38098 30772 38108
rect 30716 37828 30772 37838
rect 30772 37772 30884 37828
rect 30716 37762 30772 37772
rect 30604 37492 30660 37502
rect 30604 37398 30660 37436
rect 30828 36820 30884 37772
rect 30940 37490 30996 40012
rect 31276 39732 31332 39742
rect 31388 39732 31444 42140
rect 31276 39730 31444 39732
rect 31276 39678 31278 39730
rect 31330 39678 31444 39730
rect 31276 39676 31444 39678
rect 31500 41970 31556 42476
rect 31500 41918 31502 41970
rect 31554 41918 31556 41970
rect 31500 41860 31556 41918
rect 31276 39620 31332 39676
rect 31276 39554 31332 39564
rect 31500 39396 31556 41804
rect 31276 39340 31556 39396
rect 31276 38668 31332 39340
rect 31612 38668 31668 44940
rect 31724 43204 31780 47068
rect 31836 46900 31892 46910
rect 31892 46844 32004 46900
rect 31836 46806 31892 46844
rect 31948 44210 32004 46844
rect 32396 46788 32452 48972
rect 32508 48242 32564 49756
rect 32508 48190 32510 48242
rect 32562 48190 32564 48242
rect 32508 46900 32564 48190
rect 32620 47012 32676 52892
rect 32732 52052 32788 52062
rect 32732 50706 32788 51996
rect 32844 51940 32900 55020
rect 33292 54402 33348 54414
rect 33292 54350 33294 54402
rect 33346 54350 33348 54402
rect 33068 53844 33124 53854
rect 33292 53844 33348 54350
rect 33740 54402 33796 54414
rect 33740 54350 33742 54402
rect 33794 54350 33796 54402
rect 33740 53844 33796 54350
rect 33852 53844 33908 53854
rect 32844 51874 32900 51884
rect 32956 53842 33572 53844
rect 32956 53790 33070 53842
rect 33122 53790 33572 53842
rect 32956 53788 33572 53790
rect 33740 53842 33908 53844
rect 33740 53790 33854 53842
rect 33906 53790 33908 53842
rect 33740 53788 33908 53790
rect 32732 50654 32734 50706
rect 32786 50654 32788 50706
rect 32732 50596 32788 50654
rect 32732 50530 32788 50540
rect 32956 50428 33012 53788
rect 33068 53778 33124 53788
rect 33516 53732 33572 53788
rect 33628 53732 33684 53742
rect 33516 53730 33684 53732
rect 33516 53678 33630 53730
rect 33682 53678 33684 53730
rect 33516 53676 33684 53678
rect 33628 53666 33684 53676
rect 33628 52948 33684 52958
rect 33628 52854 33684 52892
rect 33180 52836 33236 52846
rect 33180 52834 33348 52836
rect 33180 52782 33182 52834
rect 33234 52782 33348 52834
rect 33180 52780 33348 52782
rect 33180 52770 33236 52780
rect 33292 52724 33348 52780
rect 33180 52276 33236 52286
rect 33068 51940 33124 51950
rect 33068 51378 33124 51884
rect 33068 51326 33070 51378
rect 33122 51326 33124 51378
rect 33068 50820 33124 51326
rect 33068 50754 33124 50764
rect 32620 46946 32676 46956
rect 32844 50372 33012 50428
rect 32508 46834 32564 46844
rect 32396 46694 32452 46732
rect 32284 46674 32340 46686
rect 32284 46622 32286 46674
rect 32338 46622 32340 46674
rect 32284 46564 32340 46622
rect 32284 46498 32340 46508
rect 32508 45332 32564 45342
rect 32508 45238 32564 45276
rect 32060 44996 32116 45006
rect 32060 44994 32228 44996
rect 32060 44942 32062 44994
rect 32114 44942 32228 44994
rect 32060 44940 32228 44942
rect 32060 44930 32116 44940
rect 31948 44158 31950 44210
rect 32002 44158 32004 44210
rect 31948 44146 32004 44158
rect 32060 44548 32116 44558
rect 31836 43428 31892 43438
rect 31892 43372 32004 43428
rect 31836 43334 31892 43372
rect 31724 43138 31780 43148
rect 31836 42756 31892 42766
rect 31836 41860 31892 42700
rect 31948 42196 32004 43372
rect 31948 42130 32004 42140
rect 32060 42980 32116 44492
rect 32172 44322 32228 44940
rect 32844 44548 32900 50372
rect 33068 49812 33124 49822
rect 33068 49718 33124 49756
rect 32956 49700 33012 49710
rect 32956 48916 33012 49644
rect 32956 48822 33012 48860
rect 33068 48244 33124 48254
rect 33068 48150 33124 48188
rect 33180 47570 33236 52220
rect 33292 52164 33348 52668
rect 33852 52500 33908 53788
rect 33516 52444 33908 52500
rect 33516 52164 33572 52444
rect 33964 52164 34020 56364
rect 34188 56308 34244 65212
rect 34300 58828 34356 66220
rect 34748 65604 34804 66780
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 35756 66052 35812 66062
rect 34524 65602 34804 65604
rect 34524 65550 34750 65602
rect 34802 65550 34804 65602
rect 34524 65548 34804 65550
rect 34524 64146 34580 65548
rect 34748 65538 34804 65548
rect 35644 65996 35756 66052
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 34524 64094 34526 64146
rect 34578 64094 34580 64146
rect 34524 64036 34580 64094
rect 35644 64148 35700 65996
rect 35756 65958 35812 65996
rect 35644 64082 35700 64092
rect 35756 64818 35812 64830
rect 35756 64766 35758 64818
rect 35810 64766 35812 64818
rect 34524 63970 34580 63980
rect 35196 64036 35252 64046
rect 35196 63942 35252 63980
rect 35308 63924 35364 63934
rect 35308 63830 35364 63868
rect 35756 63924 35812 64766
rect 35756 63858 35812 63868
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 35644 63028 35700 63038
rect 35644 62934 35700 62972
rect 34860 62916 34916 62926
rect 34860 62822 34916 62860
rect 35868 62188 35924 68460
rect 35980 65490 36036 69582
rect 36092 69076 36148 71150
rect 36092 69010 36148 69020
rect 36204 68964 36260 71486
rect 36428 70978 36484 71708
rect 36540 71762 36596 71774
rect 36540 71710 36542 71762
rect 36594 71710 36596 71762
rect 36540 71652 36596 71710
rect 36540 71586 36596 71596
rect 37212 71540 37268 71550
rect 37436 71540 37492 72268
rect 37548 72258 37604 72268
rect 37548 71764 37604 71802
rect 37548 71698 37604 71708
rect 38332 71764 38388 71774
rect 37996 71650 38052 71662
rect 37996 71598 37998 71650
rect 38050 71598 38052 71650
rect 37268 71484 37492 71540
rect 37548 71540 37604 71550
rect 37548 71538 37828 71540
rect 37548 71486 37550 71538
rect 37602 71486 37828 71538
rect 37548 71484 37828 71486
rect 37212 71446 37268 71484
rect 37548 71474 37604 71484
rect 37772 71090 37828 71484
rect 37772 71038 37774 71090
rect 37826 71038 37828 71090
rect 37772 71026 37828 71038
rect 36428 70926 36430 70978
rect 36482 70926 36484 70978
rect 36428 70914 36484 70926
rect 36988 70978 37044 70990
rect 36988 70926 36990 70978
rect 37042 70926 37044 70978
rect 36988 70644 37044 70926
rect 36988 70578 37044 70588
rect 37996 70644 38052 71598
rect 37996 70578 38052 70588
rect 38332 70418 38388 71708
rect 38332 70366 38334 70418
rect 38386 70366 38388 70418
rect 38332 70354 38388 70366
rect 38780 71652 38836 71662
rect 38780 70418 38836 71596
rect 39900 71092 39956 71102
rect 38780 70366 38782 70418
rect 38834 70366 38836 70418
rect 38780 70354 38836 70366
rect 38892 71090 39956 71092
rect 38892 71038 39902 71090
rect 39954 71038 39956 71090
rect 38892 71036 39956 71038
rect 38892 70306 38948 71036
rect 39900 71026 39956 71036
rect 38892 70254 38894 70306
rect 38946 70254 38948 70306
rect 38892 70242 38948 70254
rect 38444 70196 38500 70206
rect 37996 70194 38500 70196
rect 37996 70142 38446 70194
rect 38498 70142 38500 70194
rect 37996 70140 38500 70142
rect 37996 70082 38052 70140
rect 38444 70130 38500 70140
rect 37996 70030 37998 70082
rect 38050 70030 38052 70082
rect 37996 70018 38052 70030
rect 37100 69412 37156 69422
rect 37100 69318 37156 69356
rect 36204 68898 36260 68908
rect 36988 69076 37044 69086
rect 36988 67058 37044 69020
rect 36988 67006 36990 67058
rect 37042 67006 37044 67058
rect 36988 66994 37044 67006
rect 37100 68964 37156 68974
rect 35980 65438 35982 65490
rect 36034 65438 36036 65490
rect 35980 65426 36036 65438
rect 36204 66274 36260 66286
rect 36204 66222 36206 66274
rect 36258 66222 36260 66274
rect 36204 64932 36260 66222
rect 36988 66274 37044 66286
rect 36988 66222 36990 66274
rect 37042 66222 37044 66274
rect 36428 66164 36484 66174
rect 36428 66070 36484 66108
rect 36988 66052 37044 66222
rect 36988 65986 37044 65996
rect 36204 64866 36260 64876
rect 36988 64932 37044 64942
rect 36988 64838 37044 64876
rect 36428 64482 36484 64494
rect 36428 64430 36430 64482
rect 36482 64430 36484 64482
rect 35980 64148 36036 64158
rect 36428 64148 36484 64430
rect 36036 64092 36484 64148
rect 35980 62578 36036 64092
rect 37100 63922 37156 68908
rect 37100 63870 37102 63922
rect 37154 63870 37156 63922
rect 37100 63858 37156 63870
rect 37212 67170 37268 67182
rect 37212 67118 37214 67170
rect 37266 67118 37268 67170
rect 36428 63252 36484 63262
rect 36428 63138 36484 63196
rect 36428 63086 36430 63138
rect 36482 63086 36484 63138
rect 36428 63074 36484 63086
rect 35980 62526 35982 62578
rect 36034 62526 36036 62578
rect 35980 62514 36036 62526
rect 36316 63028 36372 63038
rect 36092 62244 36148 62254
rect 35868 62132 36036 62188
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 35980 60674 36036 62132
rect 35980 60622 35982 60674
rect 36034 60622 36036 60674
rect 35980 60610 36036 60622
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 34636 59780 34692 59790
rect 34636 59220 34692 59724
rect 35084 59220 35140 59230
rect 34636 59218 35140 59220
rect 34636 59166 34638 59218
rect 34690 59166 35086 59218
rect 35138 59166 35140 59218
rect 34636 59164 35140 59166
rect 34636 59154 34692 59164
rect 34300 58772 34468 58828
rect 34300 58436 34356 58446
rect 34300 58342 34356 58380
rect 34300 56980 34356 56990
rect 34300 56886 34356 56924
rect 33292 52108 33516 52164
rect 33516 52070 33572 52108
rect 33628 52108 34020 52164
rect 34076 56252 34244 56308
rect 33628 50932 33684 52108
rect 33964 51940 34020 51950
rect 33292 50876 33628 50932
rect 33292 50706 33348 50876
rect 33628 50866 33684 50876
rect 33852 51266 33908 51278
rect 33852 51214 33854 51266
rect 33906 51214 33908 51266
rect 33852 50818 33908 51214
rect 33852 50766 33854 50818
rect 33906 50766 33908 50818
rect 33852 50754 33908 50766
rect 33292 50654 33294 50706
rect 33346 50654 33348 50706
rect 33292 50642 33348 50654
rect 33628 50708 33684 50718
rect 33180 47518 33182 47570
rect 33234 47518 33236 47570
rect 33180 47506 33236 47518
rect 33292 46788 33348 46798
rect 33348 46732 33460 46788
rect 33292 46722 33348 46732
rect 33292 46564 33348 46574
rect 33292 45892 33348 46508
rect 32172 44270 32174 44322
rect 32226 44270 32228 44322
rect 32172 43540 32228 44270
rect 32732 44492 32900 44548
rect 33068 45836 33292 45892
rect 33068 45218 33124 45836
rect 33292 45826 33348 45836
rect 33068 45166 33070 45218
rect 33122 45166 33124 45218
rect 33068 44548 33124 45166
rect 33292 45108 33348 45118
rect 33404 45108 33460 46732
rect 33292 45106 33460 45108
rect 33292 45054 33294 45106
rect 33346 45054 33460 45106
rect 33292 45052 33460 45054
rect 33516 46002 33572 46014
rect 33516 45950 33518 46002
rect 33570 45950 33572 46002
rect 33292 45042 33348 45052
rect 33516 44548 33572 45950
rect 33628 45332 33684 50652
rect 33740 50596 33796 50606
rect 33740 49812 33796 50540
rect 33964 50482 34020 51884
rect 33964 50430 33966 50482
rect 34018 50430 34020 50482
rect 33964 50428 34020 50430
rect 33740 49364 33796 49756
rect 33852 50372 34020 50428
rect 33852 49476 33908 50372
rect 33964 49922 34020 49934
rect 33964 49870 33966 49922
rect 34018 49870 34020 49922
rect 33964 49700 34020 49870
rect 33964 49634 34020 49644
rect 34076 49698 34132 56252
rect 34188 54516 34244 54526
rect 34188 53954 34244 54460
rect 34188 53902 34190 53954
rect 34242 53902 34244 53954
rect 34188 53890 34244 53902
rect 34188 52164 34244 52174
rect 34188 51156 34244 52108
rect 34188 50818 34244 51100
rect 34188 50766 34190 50818
rect 34242 50766 34244 50818
rect 34188 50754 34244 50766
rect 34076 49646 34078 49698
rect 34130 49646 34132 49698
rect 34076 49634 34132 49646
rect 33852 49420 34244 49476
rect 33740 49308 33908 49364
rect 33628 45266 33684 45276
rect 33740 49028 33796 49038
rect 33628 45108 33684 45118
rect 33628 45014 33684 45052
rect 33628 44548 33684 44558
rect 33516 44492 33628 44548
rect 32284 43540 32340 43550
rect 32228 43538 32340 43540
rect 32228 43486 32286 43538
rect 32338 43486 32340 43538
rect 32228 43484 32340 43486
rect 32172 43474 32228 43484
rect 31276 38612 31444 38668
rect 31276 37940 31332 37950
rect 31276 37846 31332 37884
rect 31388 37604 31444 38612
rect 30940 37438 30942 37490
rect 30994 37438 30996 37490
rect 30940 37156 30996 37438
rect 30940 37090 30996 37100
rect 31276 37548 31444 37604
rect 31500 38612 31668 38668
rect 31724 41858 31892 41860
rect 31724 41806 31838 41858
rect 31890 41806 31892 41858
rect 31724 41804 31892 41806
rect 31276 36820 31332 37548
rect 31388 37268 31444 37278
rect 31388 37174 31444 37212
rect 30828 36764 31220 36820
rect 31276 36764 31444 36820
rect 30380 36652 30660 36708
rect 30268 36540 30548 36596
rect 30156 36484 30212 36494
rect 30156 36390 30212 36428
rect 30268 36370 30324 36382
rect 30268 36318 30270 36370
rect 30322 36318 30324 36370
rect 30044 36092 30212 36148
rect 30044 35924 30100 35934
rect 30044 35586 30100 35868
rect 30044 35534 30046 35586
rect 30098 35534 30100 35586
rect 30044 34916 30100 35534
rect 30156 35364 30212 36092
rect 30156 35298 30212 35308
rect 30268 35140 30324 36318
rect 29820 34860 30100 34916
rect 30156 35084 30324 35140
rect 29820 34580 29876 34860
rect 29932 34692 29988 34702
rect 29932 34598 29988 34636
rect 29820 34514 29876 34524
rect 30156 34468 30212 35084
rect 29932 34412 30212 34468
rect 30380 34914 30436 34926
rect 30380 34862 30382 34914
rect 30434 34862 30436 34914
rect 29708 34300 29876 34356
rect 29708 34132 29764 34142
rect 29708 34038 29764 34076
rect 29708 32564 29764 32574
rect 29708 31218 29764 32508
rect 29708 31166 29710 31218
rect 29762 31166 29764 31218
rect 29708 31154 29764 31166
rect 29708 29538 29764 29550
rect 29708 29486 29710 29538
rect 29762 29486 29764 29538
rect 29708 28756 29764 29486
rect 29820 29204 29876 34300
rect 29932 32786 29988 34412
rect 30156 34244 30212 34254
rect 30156 34150 30212 34188
rect 30380 33796 30436 34862
rect 30380 33730 30436 33740
rect 30268 33460 30324 33470
rect 30268 33366 30324 33404
rect 29932 32734 29934 32786
rect 29986 32734 29988 32786
rect 29932 32722 29988 32734
rect 30044 32674 30100 32686
rect 30044 32622 30046 32674
rect 30098 32622 30100 32674
rect 30044 31890 30100 32622
rect 30492 32676 30548 36540
rect 30604 33572 30660 36652
rect 30828 36594 30884 36764
rect 31164 36708 31220 36764
rect 31164 36652 31332 36708
rect 30828 36542 30830 36594
rect 30882 36542 30884 36594
rect 30828 36530 30884 36542
rect 30940 36482 30996 36494
rect 30940 36430 30942 36482
rect 30994 36430 30996 36482
rect 30828 36372 30884 36382
rect 30716 35812 30772 35850
rect 30716 35746 30772 35756
rect 30604 33506 30660 33516
rect 30716 35586 30772 35598
rect 30716 35534 30718 35586
rect 30770 35534 30772 35586
rect 30604 33348 30660 33358
rect 30604 33254 30660 33292
rect 30604 32676 30660 32686
rect 30492 32674 30660 32676
rect 30492 32622 30606 32674
rect 30658 32622 30660 32674
rect 30492 32620 30660 32622
rect 30604 32610 30660 32620
rect 30156 32562 30212 32574
rect 30156 32510 30158 32562
rect 30210 32510 30212 32562
rect 30156 32340 30212 32510
rect 30716 32562 30772 35534
rect 30716 32510 30718 32562
rect 30770 32510 30772 32562
rect 30716 32498 30772 32510
rect 30492 32340 30548 32350
rect 30156 32338 30548 32340
rect 30156 32286 30494 32338
rect 30546 32286 30548 32338
rect 30156 32284 30548 32286
rect 30492 32274 30548 32284
rect 30044 31838 30046 31890
rect 30098 31838 30100 31890
rect 30044 31826 30100 31838
rect 30156 31892 30212 31902
rect 30156 31778 30212 31836
rect 30828 31780 30884 36316
rect 30940 35924 30996 36430
rect 30940 35858 30996 35868
rect 31052 36372 31108 36382
rect 30940 35700 30996 35738
rect 30940 35634 30996 35644
rect 30940 35476 30996 35486
rect 30940 31892 30996 35420
rect 31052 34244 31108 36316
rect 31164 35698 31220 35710
rect 31164 35646 31166 35698
rect 31218 35646 31220 35698
rect 31164 35476 31220 35646
rect 31164 35410 31220 35420
rect 31276 34802 31332 36652
rect 31388 35924 31444 36764
rect 31388 35858 31444 35868
rect 31276 34750 31278 34802
rect 31330 34750 31332 34802
rect 31276 34738 31332 34750
rect 31052 34178 31108 34188
rect 31388 33236 31444 33246
rect 31276 33234 31444 33236
rect 31276 33182 31390 33234
rect 31442 33182 31444 33234
rect 31276 33180 31444 33182
rect 30940 31836 31108 31892
rect 30156 31726 30158 31778
rect 30210 31726 30212 31778
rect 30156 31714 30212 31726
rect 30716 31724 30884 31780
rect 31052 31778 31108 31836
rect 31052 31726 31054 31778
rect 31106 31726 31108 31778
rect 29932 31554 29988 31566
rect 29932 31502 29934 31554
rect 29986 31502 29988 31554
rect 29932 29764 29988 31502
rect 30492 31220 30548 31230
rect 30492 31126 30548 31164
rect 29932 29698 29988 29708
rect 30044 30210 30100 30222
rect 30044 30158 30046 30210
rect 30098 30158 30100 30210
rect 30044 29876 30100 30158
rect 30044 29428 30100 29820
rect 30044 29362 30100 29372
rect 29820 29148 30212 29204
rect 30156 28866 30212 29148
rect 30156 28814 30158 28866
rect 30210 28814 30212 28866
rect 30156 28802 30212 28814
rect 30604 28980 30660 28990
rect 29708 28690 29764 28700
rect 29932 28756 29988 28766
rect 29932 28662 29988 28700
rect 30380 28644 30436 28654
rect 30156 28084 30212 28094
rect 30156 27990 30212 28028
rect 30380 27972 30436 28588
rect 30604 28642 30660 28924
rect 30604 28590 30606 28642
rect 30658 28590 30660 28642
rect 30604 28578 30660 28590
rect 30492 27972 30548 27982
rect 30380 27970 30548 27972
rect 30380 27918 30494 27970
rect 30546 27918 30548 27970
rect 30380 27916 30548 27918
rect 30492 27906 30548 27916
rect 29932 27860 29988 27870
rect 29932 27766 29988 27804
rect 29596 27468 30212 27524
rect 29372 27134 29374 27186
rect 29426 27134 29428 27186
rect 29372 27122 29428 27134
rect 29260 27022 29262 27074
rect 29314 27022 29316 27074
rect 29260 27010 29316 27022
rect 29484 27076 29540 27086
rect 29484 26982 29540 27020
rect 29820 27076 29876 27086
rect 29708 26852 29764 26862
rect 29036 26562 29092 26572
rect 29372 26850 29764 26852
rect 29372 26798 29710 26850
rect 29762 26798 29764 26850
rect 29372 26796 29764 26798
rect 29036 26404 29092 26414
rect 28812 26402 28980 26404
rect 28812 26350 28814 26402
rect 28866 26350 28980 26402
rect 28812 26348 28980 26350
rect 28812 26338 28868 26348
rect 28924 25844 28980 26348
rect 29036 25956 29092 26348
rect 29148 26180 29204 26190
rect 29372 26180 29428 26796
rect 29708 26786 29764 26796
rect 29148 26178 29428 26180
rect 29148 26126 29150 26178
rect 29202 26126 29428 26178
rect 29148 26124 29428 26126
rect 29484 26180 29540 26190
rect 29820 26180 29876 27020
rect 29484 26178 29876 26180
rect 29484 26126 29486 26178
rect 29538 26126 29876 26178
rect 29484 26124 29876 26126
rect 29932 26962 29988 26974
rect 29932 26910 29934 26962
rect 29986 26910 29988 26962
rect 29148 26114 29204 26124
rect 29484 26114 29540 26124
rect 29036 25900 29764 25956
rect 28924 25788 29316 25844
rect 29260 25620 29316 25788
rect 29708 25620 29764 25900
rect 29260 25618 29652 25620
rect 29260 25566 29262 25618
rect 29314 25566 29652 25618
rect 29260 25564 29652 25566
rect 29260 25554 29316 25564
rect 29596 24946 29652 25564
rect 29708 25526 29764 25564
rect 29596 24894 29598 24946
rect 29650 24894 29652 24946
rect 29596 24882 29652 24894
rect 29708 25284 29764 25294
rect 28588 23492 28756 23548
rect 28700 22148 28756 23492
rect 29708 22932 29764 25228
rect 29932 23156 29988 26910
rect 30156 25508 30212 27468
rect 30604 27412 30660 27422
rect 30268 27300 30324 27310
rect 30604 27300 30660 27356
rect 30268 27206 30324 27244
rect 30492 27298 30660 27300
rect 30492 27246 30606 27298
rect 30658 27246 30660 27298
rect 30492 27244 30660 27246
rect 30492 25730 30548 27244
rect 30604 27234 30660 27244
rect 30716 27300 30772 31724
rect 30940 31668 30996 31678
rect 30940 31574 30996 31612
rect 31052 31220 31108 31726
rect 30828 30098 30884 30110
rect 30828 30046 30830 30098
rect 30882 30046 30884 30098
rect 30828 29876 30884 30046
rect 30828 29810 30884 29820
rect 31052 28756 31108 31164
rect 31276 31218 31332 33180
rect 31388 33170 31444 33180
rect 31500 32788 31556 38612
rect 31612 37156 31668 37166
rect 31612 36372 31668 37100
rect 31612 36278 31668 36316
rect 31724 36596 31780 41804
rect 31836 41794 31892 41804
rect 32060 41076 32116 42924
rect 32284 42082 32340 43484
rect 32284 42030 32286 42082
rect 32338 42030 32340 42082
rect 32172 41076 32228 41086
rect 32060 41074 32228 41076
rect 32060 41022 32174 41074
rect 32226 41022 32228 41074
rect 32060 41020 32228 41022
rect 32060 40740 32116 41020
rect 32172 41010 32228 41020
rect 32284 41076 32340 42030
rect 32620 42084 32676 42094
rect 32620 41748 32676 42028
rect 32508 41692 32676 41748
rect 32284 41010 32340 41020
rect 32396 41298 32452 41310
rect 32396 41246 32398 41298
rect 32450 41246 32452 41298
rect 31948 40516 32004 40526
rect 31948 40422 32004 40460
rect 31948 39172 32004 39182
rect 31836 39116 31948 39172
rect 31836 39058 31892 39116
rect 31948 39106 32004 39116
rect 31836 39006 31838 39058
rect 31890 39006 31892 39058
rect 31836 38994 31892 39006
rect 31948 38948 32004 38958
rect 32060 38948 32116 40684
rect 32284 40404 32340 40414
rect 32172 40180 32228 40190
rect 32172 39396 32228 40124
rect 32172 39330 32228 39340
rect 31948 38946 32116 38948
rect 31948 38894 31950 38946
rect 32002 38894 32116 38946
rect 31948 38892 32116 38894
rect 31948 37940 32004 38892
rect 32284 38836 32340 40348
rect 32060 38834 32340 38836
rect 32060 38782 32286 38834
rect 32338 38782 32340 38834
rect 32060 38780 32340 38782
rect 32060 38052 32116 38780
rect 32284 38770 32340 38780
rect 32396 38668 32452 41246
rect 32508 40626 32564 41692
rect 32508 40574 32510 40626
rect 32562 40574 32564 40626
rect 32508 40562 32564 40574
rect 32060 37986 32116 37996
rect 32172 38612 32452 38668
rect 32508 39508 32564 39518
rect 32508 38724 32564 39452
rect 32508 38658 32564 38668
rect 31836 37380 31892 37390
rect 31836 37286 31892 37324
rect 31948 37268 32004 37884
rect 31948 37156 32004 37212
rect 31612 35924 31668 35934
rect 31724 35924 31780 36540
rect 31612 35922 31780 35924
rect 31612 35870 31614 35922
rect 31666 35870 31780 35922
rect 31612 35868 31780 35870
rect 31836 37100 32004 37156
rect 31612 35858 31668 35868
rect 31388 32732 31556 32788
rect 31724 35476 31780 35486
rect 31724 34690 31780 35420
rect 31724 34638 31726 34690
rect 31778 34638 31780 34690
rect 31388 31444 31444 32732
rect 31500 32562 31556 32574
rect 31500 32510 31502 32562
rect 31554 32510 31556 32562
rect 31500 32002 31556 32510
rect 31500 31950 31502 32002
rect 31554 31950 31556 32002
rect 31500 31938 31556 31950
rect 31612 31780 31668 31790
rect 31612 31686 31668 31724
rect 31724 31556 31780 34638
rect 31836 34692 31892 37100
rect 32060 37044 32116 37054
rect 32060 35924 32116 36988
rect 31836 34626 31892 34636
rect 31948 35922 32116 35924
rect 31948 35870 32062 35922
rect 32114 35870 32116 35922
rect 31948 35868 32116 35870
rect 31836 33460 31892 33470
rect 31836 32562 31892 33404
rect 31836 32510 31838 32562
rect 31890 32510 31892 32562
rect 31836 32498 31892 32510
rect 31388 31378 31444 31388
rect 31612 31500 31780 31556
rect 31276 31166 31278 31218
rect 31330 31166 31332 31218
rect 31276 31154 31332 31166
rect 31500 30994 31556 31006
rect 31500 30942 31502 30994
rect 31554 30942 31556 30994
rect 31164 30770 31220 30782
rect 31164 30718 31166 30770
rect 31218 30718 31220 30770
rect 31164 30436 31220 30718
rect 31500 30548 31556 30942
rect 31220 30380 31444 30436
rect 31164 30370 31220 30380
rect 31388 28866 31444 30380
rect 31500 30100 31556 30492
rect 31500 30034 31556 30044
rect 31500 29876 31556 29886
rect 31500 29426 31556 29820
rect 31612 29764 31668 31500
rect 31836 31108 31892 31118
rect 31836 31014 31892 31052
rect 31948 30548 32004 35868
rect 32060 35858 32116 35868
rect 32060 34914 32116 34926
rect 32060 34862 32062 34914
rect 32114 34862 32116 34914
rect 32060 34692 32116 34862
rect 32060 34626 32116 34636
rect 32060 31778 32116 31790
rect 32060 31726 32062 31778
rect 32114 31726 32116 31778
rect 32060 31556 32116 31726
rect 32060 31490 32116 31500
rect 32060 30994 32116 31006
rect 32060 30942 32062 30994
rect 32114 30942 32116 30994
rect 32060 30660 32116 30942
rect 32060 30594 32116 30604
rect 31724 30492 32004 30548
rect 31724 30210 31780 30492
rect 32172 30436 32228 38612
rect 32284 38500 32340 38510
rect 32284 37938 32340 38444
rect 32284 37886 32286 37938
rect 32338 37886 32340 37938
rect 32284 37874 32340 37886
rect 32508 38388 32564 38398
rect 32508 37490 32564 38332
rect 32508 37438 32510 37490
rect 32562 37438 32564 37490
rect 32508 37268 32564 37438
rect 32732 37492 32788 44492
rect 33068 44482 33124 44492
rect 33404 44434 33460 44446
rect 33404 44382 33406 44434
rect 33458 44382 33460 44434
rect 33068 44322 33124 44334
rect 33068 44270 33070 44322
rect 33122 44270 33124 44322
rect 32956 44210 33012 44222
rect 32956 44158 32958 44210
rect 33010 44158 33012 44210
rect 32956 43764 33012 44158
rect 33068 44212 33124 44270
rect 33068 44156 33348 44212
rect 32956 43698 33012 43708
rect 33180 43426 33236 43438
rect 33180 43374 33182 43426
rect 33234 43374 33236 43426
rect 32956 43314 33012 43326
rect 32956 43262 32958 43314
rect 33010 43262 33012 43314
rect 32956 42866 33012 43262
rect 33180 43092 33236 43374
rect 33180 43026 33236 43036
rect 32956 42814 32958 42866
rect 33010 42814 33012 42866
rect 32956 38668 33012 42814
rect 33292 42754 33348 44156
rect 33292 42702 33294 42754
rect 33346 42702 33348 42754
rect 33068 42644 33124 42654
rect 33068 42082 33124 42588
rect 33180 42642 33236 42654
rect 33180 42590 33182 42642
rect 33234 42590 33236 42642
rect 33180 42196 33236 42590
rect 33180 42130 33236 42140
rect 33068 42030 33070 42082
rect 33122 42030 33124 42082
rect 33068 41076 33124 42030
rect 33292 41636 33348 42702
rect 33292 41186 33348 41580
rect 33292 41134 33294 41186
rect 33346 41134 33348 41186
rect 33292 41122 33348 41134
rect 33068 40982 33124 41020
rect 33404 39844 33460 44382
rect 33516 44324 33572 44334
rect 33516 43314 33572 44268
rect 33516 43262 33518 43314
rect 33570 43262 33572 43314
rect 33516 43250 33572 43262
rect 33516 42754 33572 42766
rect 33516 42702 33518 42754
rect 33570 42702 33572 42754
rect 33516 42644 33572 42702
rect 33516 42578 33572 42588
rect 33516 41636 33572 41646
rect 33516 40402 33572 41580
rect 33628 40516 33684 44492
rect 33740 41188 33796 48972
rect 33852 48914 33908 49308
rect 33852 48862 33854 48914
rect 33906 48862 33908 48914
rect 33852 48850 33908 48862
rect 33852 48132 33908 48142
rect 33852 48130 34020 48132
rect 33852 48078 33854 48130
rect 33906 48078 34020 48130
rect 33852 48076 34020 48078
rect 33852 48066 33908 48076
rect 33852 46900 33908 46910
rect 33964 46900 34020 48076
rect 33852 46898 34020 46900
rect 33852 46846 33854 46898
rect 33906 46846 34020 46898
rect 33852 46844 34020 46846
rect 34076 47234 34132 47246
rect 34076 47182 34078 47234
rect 34130 47182 34132 47234
rect 33852 46834 33908 46844
rect 34076 46674 34132 47182
rect 34076 46622 34078 46674
rect 34130 46622 34132 46674
rect 34076 46610 34132 46622
rect 33852 45108 33908 45118
rect 33852 42644 33908 45052
rect 33964 43316 34020 43326
rect 33964 43222 34020 43260
rect 33964 42644 34020 42654
rect 33852 42588 33964 42644
rect 33964 42550 34020 42588
rect 33852 41970 33908 41982
rect 33852 41918 33854 41970
rect 33906 41918 33908 41970
rect 33852 41860 33908 41918
rect 33852 41794 33908 41804
rect 33964 41858 34020 41870
rect 33964 41806 33966 41858
rect 34018 41806 34020 41858
rect 33740 41122 33796 41132
rect 33628 40422 33684 40460
rect 33964 40628 34020 41806
rect 33516 40350 33518 40402
rect 33570 40350 33572 40402
rect 33516 40068 33572 40350
rect 33516 40002 33572 40012
rect 33852 40404 33908 40414
rect 33404 39788 33572 39844
rect 33068 39620 33124 39630
rect 33404 39620 33460 39630
rect 33068 39618 33460 39620
rect 33068 39566 33070 39618
rect 33122 39566 33406 39618
rect 33458 39566 33460 39618
rect 33068 39564 33460 39566
rect 33068 39172 33124 39564
rect 33404 39554 33460 39564
rect 33068 39106 33124 39116
rect 33180 39396 33236 39406
rect 33516 39396 33572 39788
rect 33180 39058 33236 39340
rect 33180 39006 33182 39058
rect 33234 39006 33236 39058
rect 33180 38994 33236 39006
rect 33404 39340 33572 39396
rect 33740 39396 33796 39406
rect 32956 38612 33236 38668
rect 32732 37426 32788 37436
rect 33068 37268 33124 37278
rect 32508 37266 33124 37268
rect 32508 37214 33070 37266
rect 33122 37214 33124 37266
rect 32508 37212 33124 37214
rect 33068 37202 33124 37212
rect 32956 37044 33012 37054
rect 32620 36820 32676 36830
rect 32284 36596 32340 36606
rect 32284 32788 32340 36540
rect 32620 36482 32676 36764
rect 32620 36430 32622 36482
rect 32674 36430 32676 36482
rect 32620 35812 32676 36430
rect 32956 36258 33012 36988
rect 32956 36206 32958 36258
rect 33010 36206 33012 36258
rect 32956 36194 33012 36206
rect 33180 35924 33236 38612
rect 32956 35868 33236 35924
rect 33292 38052 33348 38062
rect 32732 35812 32788 35822
rect 32620 35756 32732 35812
rect 32732 35746 32788 35756
rect 32508 35588 32564 35626
rect 32508 35522 32564 35532
rect 32844 35476 32900 35486
rect 32508 35364 32564 35374
rect 32508 34244 32564 35308
rect 32620 34692 32676 34702
rect 32676 34636 32788 34692
rect 32620 34626 32676 34636
rect 32508 34188 32676 34244
rect 32508 34018 32564 34030
rect 32508 33966 32510 34018
rect 32562 33966 32564 34018
rect 32508 33572 32564 33966
rect 32508 33506 32564 33516
rect 32620 33012 32676 34188
rect 32620 32946 32676 32956
rect 32508 32788 32564 32798
rect 32284 32786 32564 32788
rect 32284 32734 32510 32786
rect 32562 32734 32564 32786
rect 32284 32732 32564 32734
rect 32284 31668 32340 32732
rect 32508 32722 32564 32732
rect 32620 32788 32676 32798
rect 32284 31602 32340 31612
rect 32284 31220 32340 31230
rect 32284 31126 32340 31164
rect 32508 31108 32564 31118
rect 32620 31108 32676 32732
rect 32732 31890 32788 34636
rect 32732 31838 32734 31890
rect 32786 31838 32788 31890
rect 32732 31220 32788 31838
rect 32732 31154 32788 31164
rect 32508 31106 32676 31108
rect 32508 31054 32510 31106
rect 32562 31054 32676 31106
rect 32508 31052 32676 31054
rect 32396 30772 32452 30782
rect 32396 30678 32452 30716
rect 31724 30158 31726 30210
rect 31778 30158 31780 30210
rect 31724 29988 31780 30158
rect 31724 29922 31780 29932
rect 31948 30380 32228 30436
rect 31948 29876 32004 30380
rect 31948 29810 32004 29820
rect 32060 30100 32116 30110
rect 31612 29708 31892 29764
rect 31500 29374 31502 29426
rect 31554 29374 31556 29426
rect 31500 29362 31556 29374
rect 31724 29204 31780 29214
rect 31388 28814 31390 28866
rect 31442 28814 31444 28866
rect 31388 28802 31444 28814
rect 31612 29202 31780 29204
rect 31612 29150 31726 29202
rect 31778 29150 31780 29202
rect 31612 29148 31780 29150
rect 31164 28756 31220 28766
rect 31108 28754 31220 28756
rect 31108 28702 31166 28754
rect 31218 28702 31220 28754
rect 31108 28700 31220 28702
rect 31052 28690 31108 28700
rect 31164 28690 31220 28700
rect 30828 28530 30884 28542
rect 30828 28478 30830 28530
rect 30882 28478 30884 28530
rect 30828 27636 30884 28478
rect 30828 27570 30884 27580
rect 31052 28530 31108 28542
rect 31052 28478 31054 28530
rect 31106 28478 31108 28530
rect 30492 25678 30494 25730
rect 30546 25678 30548 25730
rect 30492 25666 30548 25678
rect 30380 25620 30436 25630
rect 30268 25508 30324 25518
rect 30156 25506 30324 25508
rect 30156 25454 30270 25506
rect 30322 25454 30324 25506
rect 30156 25452 30324 25454
rect 29932 23042 29988 23100
rect 29932 22990 29934 23042
rect 29986 22990 29988 23042
rect 29932 22978 29988 22990
rect 30044 24612 30100 24622
rect 30268 24612 30324 25452
rect 30044 24610 30324 24612
rect 30044 24558 30046 24610
rect 30098 24558 30324 24610
rect 30044 24556 30324 24558
rect 29596 22876 29764 22932
rect 28700 22082 28756 22092
rect 29260 22148 29316 22158
rect 29148 17556 29204 17566
rect 28588 17444 28644 17454
rect 29148 17444 29204 17500
rect 28588 17442 29204 17444
rect 28588 17390 28590 17442
rect 28642 17390 29204 17442
rect 28588 17388 29204 17390
rect 28588 17378 28644 17388
rect 28588 15316 28644 15354
rect 28588 15250 28644 15260
rect 28700 15148 28756 17388
rect 28812 16996 28868 17006
rect 28812 16902 28868 16940
rect 29148 16660 29204 16670
rect 28924 16658 29204 16660
rect 28924 16606 29150 16658
rect 29202 16606 29204 16658
rect 28924 16604 29204 16606
rect 28924 15876 28980 16604
rect 29148 16594 29204 16604
rect 29260 16436 29316 22092
rect 28364 14018 28420 14028
rect 28588 15092 28756 15148
rect 28812 15820 28980 15876
rect 29036 16380 29316 16436
rect 29372 20802 29428 20814
rect 29372 20750 29374 20802
rect 29426 20750 29428 20802
rect 27804 13806 27806 13858
rect 27858 13806 27860 13858
rect 27804 13794 27860 13806
rect 28028 13636 28084 13646
rect 27356 12740 27412 12750
rect 27356 12290 27412 12684
rect 27356 12238 27358 12290
rect 27410 12238 27412 12290
rect 27356 12226 27412 12238
rect 28028 12178 28084 13580
rect 28588 12964 28644 15092
rect 28700 14644 28756 14654
rect 28700 14550 28756 14588
rect 28588 12908 28756 12964
rect 28588 12738 28644 12750
rect 28588 12686 28590 12738
rect 28642 12686 28644 12738
rect 28588 12404 28644 12686
rect 28588 12338 28644 12348
rect 28476 12292 28532 12302
rect 28028 12126 28030 12178
rect 28082 12126 28084 12178
rect 28028 12114 28084 12126
rect 28140 12290 28532 12292
rect 28140 12238 28478 12290
rect 28530 12238 28532 12290
rect 28140 12236 28532 12238
rect 28140 11732 28196 12236
rect 28476 12226 28532 12236
rect 27580 11676 28196 11732
rect 27580 11506 27636 11676
rect 27580 11454 27582 11506
rect 27634 11454 27636 11506
rect 27580 11442 27636 11454
rect 28252 11396 28308 11406
rect 28252 11302 28308 11340
rect 27916 9940 27972 9950
rect 27356 9604 27412 9614
rect 27356 9266 27412 9548
rect 27356 9214 27358 9266
rect 27410 9214 27412 9266
rect 27356 9202 27412 9214
rect 27804 9044 27860 9054
rect 27692 8988 27804 9044
rect 27020 8652 27300 8708
rect 27468 8932 27524 8942
rect 26572 8372 26740 8428
rect 25900 8206 25902 8258
rect 25954 8206 25956 8258
rect 25900 7364 25956 8206
rect 26348 7474 26404 7486
rect 26348 7422 26350 7474
rect 26402 7422 26404 7474
rect 26012 7364 26068 7374
rect 26348 7364 26404 7422
rect 25900 7362 26404 7364
rect 25900 7310 26014 7362
rect 26066 7310 26404 7362
rect 25900 7308 26404 7310
rect 25788 6020 25844 6030
rect 25788 5926 25844 5964
rect 25228 5796 25284 5806
rect 24220 4946 24276 4956
rect 24444 5124 24500 5134
rect 23548 4452 23604 4462
rect 23548 4450 23828 4452
rect 23548 4398 23550 4450
rect 23602 4398 23828 4450
rect 23548 4396 23828 4398
rect 23548 4386 23604 4396
rect 22652 3666 23044 3668
rect 22652 3614 22654 3666
rect 22706 3614 23044 3666
rect 22652 3612 23044 3614
rect 22652 3602 22708 3612
rect 22988 3554 23044 3612
rect 23772 3666 23828 4396
rect 23772 3614 23774 3666
rect 23826 3614 23828 3666
rect 23772 3602 23828 3614
rect 23884 4338 23940 4350
rect 23884 4286 23886 4338
rect 23938 4286 23940 4338
rect 22988 3502 22990 3554
rect 23042 3502 23044 3554
rect 22988 3490 23044 3502
rect 23772 2996 23828 3006
rect 23884 2996 23940 4286
rect 24444 4338 24500 5068
rect 24892 5124 24948 5134
rect 25228 5124 25284 5740
rect 26012 5796 26068 7308
rect 26012 5730 26068 5740
rect 26348 6018 26404 6030
rect 26348 5966 26350 6018
rect 26402 5966 26404 6018
rect 24892 5122 25284 5124
rect 24892 5070 24894 5122
rect 24946 5070 25284 5122
rect 24892 5068 25284 5070
rect 24892 5058 24948 5068
rect 24668 4452 24724 4462
rect 24668 4358 24724 4396
rect 24444 4286 24446 4338
rect 24498 4286 24500 4338
rect 24444 4274 24500 4286
rect 25228 4340 25284 5068
rect 25452 5124 25508 5134
rect 25452 5030 25508 5068
rect 25788 5124 25844 5134
rect 26012 5124 26068 5134
rect 26348 5124 26404 5966
rect 26684 6020 26740 8372
rect 26908 6916 26964 6926
rect 26908 6822 26964 6860
rect 27020 6130 27076 8652
rect 27468 8372 27524 8876
rect 27356 8316 27524 8372
rect 27132 8034 27188 8046
rect 27132 7982 27134 8034
rect 27186 7982 27188 8034
rect 27132 7586 27188 7982
rect 27132 7534 27134 7586
rect 27186 7534 27188 7586
rect 27132 7522 27188 7534
rect 27356 6804 27412 8316
rect 27468 8148 27524 8158
rect 27468 8146 27636 8148
rect 27468 8094 27470 8146
rect 27522 8094 27636 8146
rect 27468 8092 27636 8094
rect 27468 8082 27524 8092
rect 27580 6916 27636 8092
rect 27580 6850 27636 6860
rect 27468 6804 27524 6814
rect 27356 6802 27524 6804
rect 27356 6750 27470 6802
rect 27522 6750 27524 6802
rect 27356 6748 27524 6750
rect 27244 6692 27300 6702
rect 27020 6078 27022 6130
rect 27074 6078 27076 6130
rect 27020 6066 27076 6078
rect 27132 6636 27244 6692
rect 26684 5926 26740 5964
rect 25340 4340 25396 4350
rect 25228 4338 25396 4340
rect 25228 4286 25342 4338
rect 25394 4286 25396 4338
rect 25228 4284 25396 4286
rect 23772 2994 23940 2996
rect 23772 2942 23774 2994
rect 23826 2942 23940 2994
rect 23772 2940 23940 2942
rect 23772 2930 23828 2940
rect 23212 2772 23268 2782
rect 22428 2770 23268 2772
rect 22428 2718 23214 2770
rect 23266 2718 23268 2770
rect 22428 2716 23268 2718
rect 22428 2658 22484 2716
rect 23212 2706 23268 2716
rect 23436 2772 23492 2782
rect 23436 2678 23492 2716
rect 24220 2772 24276 2782
rect 24220 2678 24276 2716
rect 25340 2772 25396 4284
rect 25788 2884 25844 5068
rect 25900 5122 26404 5124
rect 25900 5070 26014 5122
rect 26066 5070 26404 5122
rect 25900 5068 26404 5070
rect 26460 5124 26516 5134
rect 25900 3666 25956 5068
rect 26012 5058 26068 5068
rect 26460 5030 26516 5068
rect 27132 5124 27188 6636
rect 27244 6598 27300 6636
rect 27244 6132 27300 6142
rect 27244 5906 27300 6076
rect 27244 5854 27246 5906
rect 27298 5854 27300 5906
rect 27244 5842 27300 5854
rect 27132 5058 27188 5068
rect 26012 4452 26068 4462
rect 26012 4358 26068 4396
rect 27468 4228 27524 6748
rect 27692 6132 27748 8988
rect 27804 8950 27860 8988
rect 27916 6802 27972 9884
rect 28588 9604 28644 9614
rect 28588 9266 28644 9548
rect 28588 9214 28590 9266
rect 28642 9214 28644 9266
rect 28588 9202 28644 9214
rect 27916 6750 27918 6802
rect 27970 6750 27972 6802
rect 27916 6692 27972 6750
rect 28700 6692 28756 12908
rect 28812 12290 28868 15820
rect 29036 15148 29092 16380
rect 29148 15874 29204 15886
rect 29148 15822 29150 15874
rect 29202 15822 29204 15874
rect 29148 15316 29204 15822
rect 29148 15250 29204 15260
rect 29372 15148 29428 20750
rect 29484 20692 29540 20702
rect 29484 20598 29540 20636
rect 29596 18564 29652 22876
rect 30044 22820 30100 24556
rect 30380 23380 30436 25564
rect 29484 18508 29652 18564
rect 29708 22764 30100 22820
rect 30268 23324 30436 23380
rect 30604 23380 30660 23390
rect 29484 16884 29540 18508
rect 29596 18340 29652 18350
rect 29708 18340 29764 22764
rect 30268 21588 30324 23324
rect 30380 23156 30436 23166
rect 30380 23062 30436 23100
rect 30604 23154 30660 23324
rect 30604 23102 30606 23154
rect 30658 23102 30660 23154
rect 30604 23090 30660 23102
rect 30716 21924 30772 27244
rect 31052 27188 31108 28478
rect 31612 28084 31668 29148
rect 31724 29138 31780 29148
rect 31052 27122 31108 27132
rect 31388 28028 31668 28084
rect 31724 28866 31780 28878
rect 31724 28814 31726 28866
rect 31778 28814 31780 28866
rect 31724 28754 31780 28814
rect 31836 28868 31892 29708
rect 31948 29428 32004 29438
rect 31948 29334 32004 29372
rect 31836 28812 32004 28868
rect 31724 28702 31726 28754
rect 31778 28702 31780 28754
rect 30828 27076 30884 27086
rect 30828 26982 30884 27020
rect 31276 26964 31332 27002
rect 31276 26898 31332 26908
rect 31388 26516 31444 28028
rect 31724 27972 31780 28702
rect 31500 27916 31780 27972
rect 31500 26852 31556 27916
rect 31948 27860 32004 28812
rect 32060 28420 32116 30044
rect 32172 29652 32228 29662
rect 32172 29558 32228 29596
rect 32396 29540 32452 29550
rect 32396 29446 32452 29484
rect 32508 29428 32564 31052
rect 32172 29314 32228 29326
rect 32172 29262 32174 29314
rect 32226 29262 32228 29314
rect 32172 28868 32228 29262
rect 32172 28802 32228 28812
rect 32284 28980 32340 28990
rect 32172 28420 32228 28430
rect 32060 28418 32228 28420
rect 32060 28366 32174 28418
rect 32226 28366 32228 28418
rect 32060 28364 32228 28366
rect 31836 27804 32004 27860
rect 32172 27860 32228 28364
rect 32284 28082 32340 28924
rect 32508 28756 32564 29372
rect 32620 30660 32676 30670
rect 32620 29986 32676 30604
rect 32620 29934 32622 29986
rect 32674 29934 32676 29986
rect 32620 29204 32676 29934
rect 32620 29138 32676 29148
rect 32620 28756 32676 28766
rect 32508 28754 32676 28756
rect 32508 28702 32622 28754
rect 32674 28702 32676 28754
rect 32508 28700 32676 28702
rect 32620 28308 32676 28700
rect 32620 28242 32676 28252
rect 32284 28030 32286 28082
rect 32338 28030 32340 28082
rect 32284 28018 32340 28030
rect 32172 27804 32340 27860
rect 31836 27748 31892 27804
rect 31500 26786 31556 26796
rect 31724 27692 31892 27748
rect 31388 26450 31444 26460
rect 31612 26180 31668 26190
rect 31500 26178 31668 26180
rect 31500 26126 31614 26178
rect 31666 26126 31668 26178
rect 31500 26124 31668 26126
rect 30828 25396 30884 25406
rect 31164 25396 31220 25406
rect 30828 25394 31220 25396
rect 30828 25342 30830 25394
rect 30882 25342 31166 25394
rect 31218 25342 31220 25394
rect 30828 25340 31220 25342
rect 30828 25330 30884 25340
rect 31164 25330 31220 25340
rect 31500 25394 31556 26124
rect 31612 26114 31668 26124
rect 31500 25342 31502 25394
rect 31554 25342 31556 25394
rect 31500 25330 31556 25342
rect 31612 25844 31668 25854
rect 31164 25060 31220 25070
rect 30940 25004 31164 25060
rect 30940 24052 30996 25004
rect 31164 24994 31220 25004
rect 30828 24050 31332 24052
rect 30828 23998 30942 24050
rect 30994 23998 31332 24050
rect 30828 23996 31332 23998
rect 30828 22036 30884 23996
rect 30940 23986 30996 23996
rect 31164 23716 31220 23726
rect 31164 23044 31220 23660
rect 31276 23266 31332 23996
rect 31612 23716 31668 25788
rect 31612 23622 31668 23660
rect 31276 23214 31278 23266
rect 31330 23214 31332 23266
rect 31276 23202 31332 23214
rect 31612 23156 31668 23166
rect 31164 22988 31332 23044
rect 30940 22932 30996 22942
rect 30940 22930 31108 22932
rect 30940 22878 30942 22930
rect 30994 22878 31108 22930
rect 30940 22876 31108 22878
rect 30940 22866 30996 22876
rect 31052 22370 31108 22876
rect 31052 22318 31054 22370
rect 31106 22318 31108 22370
rect 31052 22306 31108 22318
rect 30828 21980 31108 22036
rect 30716 21868 30996 21924
rect 30380 21812 30436 21822
rect 30716 21812 30772 21868
rect 30380 21810 30772 21812
rect 30380 21758 30382 21810
rect 30434 21758 30772 21810
rect 30380 21756 30772 21758
rect 30380 21746 30436 21756
rect 30828 21700 30884 21710
rect 30492 21588 30548 21598
rect 30268 21532 30492 21588
rect 30548 21532 30660 21588
rect 30492 21494 30548 21532
rect 30492 20916 30548 20926
rect 30268 20914 30548 20916
rect 30268 20862 30494 20914
rect 30546 20862 30548 20914
rect 30268 20860 30548 20862
rect 30268 20242 30324 20860
rect 30492 20850 30548 20860
rect 30604 20804 30660 21532
rect 30828 21586 30884 21644
rect 30828 21534 30830 21586
rect 30882 21534 30884 21586
rect 30716 21028 30772 21038
rect 30828 21028 30884 21534
rect 30716 21026 30884 21028
rect 30716 20974 30718 21026
rect 30770 20974 30884 21026
rect 30716 20972 30884 20974
rect 30716 20962 30772 20972
rect 30604 20748 30884 20804
rect 30268 20190 30270 20242
rect 30322 20190 30324 20242
rect 30268 20178 30324 20190
rect 30380 20580 30436 20590
rect 29596 18338 29764 18340
rect 29596 18286 29598 18338
rect 29650 18286 29764 18338
rect 29596 18284 29764 18286
rect 29820 19908 29876 19918
rect 30156 19908 30212 19918
rect 29820 19906 30212 19908
rect 29820 19854 29822 19906
rect 29874 19854 30158 19906
rect 30210 19854 30212 19906
rect 29820 19852 30212 19854
rect 29596 18274 29652 18284
rect 29708 16996 29764 17006
rect 29708 16902 29764 16940
rect 29484 16828 29652 16884
rect 29484 16660 29540 16670
rect 29484 16566 29540 16604
rect 29484 16098 29540 16110
rect 29484 16046 29486 16098
rect 29538 16046 29540 16098
rect 29484 15652 29540 16046
rect 29596 15988 29652 16828
rect 29708 16212 29764 16222
rect 29820 16212 29876 19852
rect 30156 19842 30212 19852
rect 29932 17554 29988 17566
rect 29932 17502 29934 17554
rect 29986 17502 29988 17554
rect 29932 17444 29988 17502
rect 29932 16660 29988 17388
rect 30268 17108 30324 17118
rect 30268 17014 30324 17052
rect 29932 16594 29988 16604
rect 30268 16660 30324 16670
rect 29708 16210 29876 16212
rect 29708 16158 29710 16210
rect 29762 16158 29876 16210
rect 29708 16156 29876 16158
rect 30268 16210 30324 16604
rect 30268 16158 30270 16210
rect 30322 16158 30324 16210
rect 29708 16146 29764 16156
rect 30268 16146 30324 16158
rect 29596 15932 30100 15988
rect 29484 15596 29988 15652
rect 29932 15538 29988 15596
rect 29932 15486 29934 15538
rect 29986 15486 29988 15538
rect 29932 15148 29988 15486
rect 28812 12238 28814 12290
rect 28866 12238 28868 12290
rect 28812 12226 28868 12238
rect 28924 15092 29092 15148
rect 29148 15092 29428 15148
rect 29820 15092 29988 15148
rect 28924 9940 28980 15092
rect 29148 10164 29204 15092
rect 29820 14756 29876 15092
rect 29820 14690 29876 14700
rect 29260 14644 29316 14654
rect 29260 14530 29316 14588
rect 29260 14478 29262 14530
rect 29314 14478 29316 14530
rect 29260 14466 29316 14478
rect 29372 14532 29428 14542
rect 29372 14418 29428 14476
rect 29372 14366 29374 14418
rect 29426 14366 29428 14418
rect 29372 14354 29428 14366
rect 29932 14532 29988 14542
rect 29596 14308 29652 14318
rect 29820 14308 29876 14318
rect 29596 14214 29652 14252
rect 29708 14306 29876 14308
rect 29708 14254 29822 14306
rect 29874 14254 29876 14306
rect 29708 14252 29876 14254
rect 29708 13524 29764 14252
rect 29820 14242 29876 14252
rect 29932 13634 29988 14476
rect 29932 13582 29934 13634
rect 29986 13582 29988 13634
rect 29932 13570 29988 13582
rect 29372 13468 29764 13524
rect 29372 12962 29428 13468
rect 29372 12910 29374 12962
rect 29426 12910 29428 12962
rect 29372 12898 29428 12910
rect 29932 13188 29988 13198
rect 29932 12850 29988 13132
rect 29932 12798 29934 12850
rect 29986 12798 29988 12850
rect 29596 12740 29652 12750
rect 29596 12646 29652 12684
rect 29932 12404 29988 12798
rect 29932 12338 29988 12348
rect 29708 12292 29764 12302
rect 29708 12178 29764 12236
rect 29708 12126 29710 12178
rect 29762 12126 29764 12178
rect 29708 12114 29764 12126
rect 28924 9874 28980 9884
rect 29036 10108 29204 10164
rect 29932 11620 29988 11630
rect 28924 9604 28980 9614
rect 28924 9266 28980 9548
rect 28924 9214 28926 9266
rect 28978 9214 28980 9266
rect 28924 9202 28980 9214
rect 29036 8930 29092 10108
rect 29932 10050 29988 11564
rect 29932 9998 29934 10050
rect 29986 9998 29988 10050
rect 29932 9986 29988 9998
rect 30044 10836 30100 15932
rect 30380 15148 30436 20524
rect 30604 20468 30660 20748
rect 30828 20690 30884 20748
rect 30828 20638 30830 20690
rect 30882 20638 30884 20690
rect 30828 20626 30884 20638
rect 30604 20402 30660 20412
rect 30492 17108 30548 17118
rect 30492 17106 30884 17108
rect 30492 17054 30494 17106
rect 30546 17054 30884 17106
rect 30492 17052 30884 17054
rect 30492 17042 30548 17052
rect 30604 16884 30660 16894
rect 30604 16882 30772 16884
rect 30604 16830 30606 16882
rect 30658 16830 30772 16882
rect 30604 16828 30772 16830
rect 30604 16818 30660 16828
rect 30380 15092 30660 15148
rect 30156 14756 30212 14766
rect 30156 14530 30212 14700
rect 30156 14478 30158 14530
rect 30210 14478 30212 14530
rect 30156 14420 30212 14478
rect 30380 14532 30436 14542
rect 30380 14438 30436 14476
rect 30156 14354 30212 14364
rect 30492 14308 30548 14318
rect 30492 13858 30548 14252
rect 30604 13970 30660 15092
rect 30604 13918 30606 13970
rect 30658 13918 30660 13970
rect 30604 13906 30660 13918
rect 30492 13806 30494 13858
rect 30546 13806 30548 13858
rect 30492 13794 30548 13806
rect 30268 13746 30324 13758
rect 30268 13694 30270 13746
rect 30322 13694 30324 13746
rect 30268 11620 30324 13694
rect 30380 12740 30436 12750
rect 30380 12290 30436 12684
rect 30380 12238 30382 12290
rect 30434 12238 30436 12290
rect 30380 12226 30436 12238
rect 30268 11554 30324 11564
rect 30156 10836 30212 10846
rect 30044 10834 30212 10836
rect 30044 10782 30158 10834
rect 30210 10782 30212 10834
rect 30044 10780 30212 10782
rect 29372 9828 29428 9838
rect 29372 9154 29428 9772
rect 29820 9716 29876 9726
rect 30044 9716 30100 10780
rect 30156 10770 30212 10780
rect 30492 9828 30548 9838
rect 30716 9828 30772 16828
rect 30828 16322 30884 17052
rect 30828 16270 30830 16322
rect 30882 16270 30884 16322
rect 30828 16258 30884 16270
rect 30940 16324 30996 21868
rect 31052 17780 31108 21980
rect 31164 21588 31220 21598
rect 31164 20242 31220 21532
rect 31164 20190 31166 20242
rect 31218 20190 31220 20242
rect 31164 20178 31220 20190
rect 31052 17714 31108 17724
rect 31052 17554 31108 17566
rect 31052 17502 31054 17554
rect 31106 17502 31108 17554
rect 31052 17106 31108 17502
rect 31052 17054 31054 17106
rect 31106 17054 31108 17106
rect 31052 17042 31108 17054
rect 31164 16324 31220 16334
rect 30940 16322 31220 16324
rect 30940 16270 31166 16322
rect 31218 16270 31220 16322
rect 30940 16268 31220 16270
rect 30940 16098 30996 16268
rect 31164 16258 31220 16268
rect 30940 16046 30942 16098
rect 30994 16046 30996 16098
rect 30828 15876 30884 15886
rect 30828 15782 30884 15820
rect 30940 15428 30996 16046
rect 31276 15988 31332 22988
rect 31612 22372 31668 23100
rect 31724 22596 31780 27692
rect 31948 27636 32004 27646
rect 31836 27580 31948 27636
rect 31836 27186 31892 27580
rect 31948 27570 32004 27580
rect 31836 27134 31838 27186
rect 31890 27134 31892 27186
rect 31836 27122 31892 27134
rect 31948 27412 32004 27422
rect 31948 25618 32004 27356
rect 32172 27300 32228 27310
rect 31948 25566 31950 25618
rect 32002 25566 32004 25618
rect 31948 24836 32004 25566
rect 31948 24770 32004 24780
rect 32060 27188 32116 27198
rect 31948 24052 32004 24062
rect 32060 24052 32116 27132
rect 32172 27186 32228 27244
rect 32172 27134 32174 27186
rect 32226 27134 32228 27186
rect 32172 27122 32228 27134
rect 32284 26964 32340 27804
rect 32844 27748 32900 35420
rect 32956 29652 33012 35868
rect 33068 35700 33124 35710
rect 33068 34244 33124 35644
rect 33180 34468 33236 34478
rect 33292 34468 33348 37996
rect 33404 36036 33460 39340
rect 33628 39060 33684 39070
rect 33628 37380 33684 39004
rect 33740 38276 33796 39340
rect 33852 38836 33908 40348
rect 33964 39508 34020 40572
rect 34076 41748 34132 41758
rect 34076 39732 34132 41692
rect 34188 40292 34244 49420
rect 34412 49250 34468 58772
rect 34524 58548 34580 58558
rect 34524 56978 34580 58492
rect 35084 58436 35140 59164
rect 35756 59106 35812 59118
rect 35756 59054 35758 59106
rect 35810 59054 35812 59106
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 35084 58370 35140 58380
rect 35644 58434 35700 58446
rect 35644 58382 35646 58434
rect 35698 58382 35700 58434
rect 35644 57874 35700 58382
rect 35756 58324 35812 59054
rect 35868 58324 35924 58334
rect 35756 58322 35924 58324
rect 35756 58270 35870 58322
rect 35922 58270 35924 58322
rect 35756 58268 35924 58270
rect 35868 58258 35924 58268
rect 36092 57876 36148 62188
rect 36316 62242 36372 62972
rect 36316 62190 36318 62242
rect 36370 62190 36372 62242
rect 36316 62178 36372 62190
rect 36988 62914 37044 62926
rect 36988 62862 36990 62914
rect 37042 62862 37044 62914
rect 36988 62188 37044 62862
rect 36988 62132 37156 62188
rect 37100 61570 37156 62132
rect 37100 61518 37102 61570
rect 37154 61518 37156 61570
rect 37100 61506 37156 61518
rect 35644 57822 35646 57874
rect 35698 57822 35700 57874
rect 35644 57810 35700 57822
rect 35756 57874 36148 57876
rect 35756 57822 36094 57874
rect 36146 57822 36148 57874
rect 35756 57820 36148 57822
rect 35308 57652 35364 57662
rect 35756 57652 35812 57820
rect 36092 57810 36148 57820
rect 35308 57650 35812 57652
rect 35308 57598 35310 57650
rect 35362 57598 35812 57650
rect 35308 57596 35812 57598
rect 35308 57586 35364 57596
rect 35084 57538 35140 57550
rect 35084 57486 35086 57538
rect 35138 57486 35140 57538
rect 34524 56926 34526 56978
rect 34578 56926 34580 56978
rect 34524 56914 34580 56926
rect 34972 56980 35028 56990
rect 34972 56886 35028 56924
rect 34860 54516 34916 54526
rect 34860 54422 34916 54460
rect 34636 53506 34692 53518
rect 34636 53454 34638 53506
rect 34690 53454 34692 53506
rect 34636 52948 34692 53454
rect 34636 52882 34692 52892
rect 35084 52388 35140 57486
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 35420 57092 35476 57102
rect 35420 56308 35476 57036
rect 35420 56082 35476 56252
rect 35420 56030 35422 56082
rect 35474 56030 35476 56082
rect 35420 56018 35476 56030
rect 35532 56980 35588 57596
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35196 55524 35252 55534
rect 35196 54738 35252 55468
rect 35532 55188 35588 56924
rect 36092 55970 36148 55982
rect 36092 55918 36094 55970
rect 36146 55918 36148 55970
rect 36092 55524 36148 55918
rect 36092 55458 36148 55468
rect 35644 55412 35700 55422
rect 35644 55410 35924 55412
rect 35644 55358 35646 55410
rect 35698 55358 35924 55410
rect 35644 55356 35924 55358
rect 35644 55346 35700 55356
rect 35532 55132 35700 55188
rect 35196 54686 35198 54738
rect 35250 54686 35252 54738
rect 35196 54674 35252 54686
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35532 53172 35588 53182
rect 35532 52948 35588 53116
rect 35532 52854 35588 52892
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35644 52500 35700 55132
rect 34972 52332 35140 52388
rect 35644 52386 35700 52444
rect 35644 52334 35646 52386
rect 35698 52334 35700 52386
rect 34524 51940 34580 51950
rect 34524 51846 34580 51884
rect 34972 51268 35028 52332
rect 35644 52322 35700 52334
rect 34860 50932 34916 50942
rect 34748 50594 34804 50606
rect 34748 50542 34750 50594
rect 34802 50542 34804 50594
rect 34748 50484 34804 50542
rect 34860 50596 34916 50876
rect 34972 50596 35028 51212
rect 35084 52164 35140 52174
rect 35420 52164 35476 52174
rect 35084 52162 35476 52164
rect 35084 52110 35086 52162
rect 35138 52110 35422 52162
rect 35474 52110 35476 52162
rect 35084 52108 35476 52110
rect 35084 50820 35140 52108
rect 35420 52098 35476 52108
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35084 50764 35252 50820
rect 35084 50596 35140 50606
rect 34972 50594 35140 50596
rect 34972 50542 35086 50594
rect 35138 50542 35140 50594
rect 34972 50540 35140 50542
rect 34860 50502 34916 50540
rect 35084 50530 35140 50540
rect 35196 50428 35252 50764
rect 35756 50708 35812 50718
rect 35756 50614 35812 50652
rect 34748 50418 34804 50428
rect 34972 50370 35028 50382
rect 34972 50318 34974 50370
rect 35026 50318 35028 50370
rect 34748 49812 34804 49822
rect 34748 49718 34804 49756
rect 34412 49198 34414 49250
rect 34466 49198 34468 49250
rect 34412 49186 34468 49198
rect 34972 48804 35028 50318
rect 34972 48738 35028 48748
rect 35084 50372 35252 50428
rect 35308 50594 35364 50606
rect 35308 50542 35310 50594
rect 35362 50542 35364 50594
rect 35308 50428 35364 50542
rect 35868 50484 35924 55356
rect 35980 53618 36036 53630
rect 35980 53566 35982 53618
rect 36034 53566 36036 53618
rect 35980 52386 36036 53566
rect 36316 53506 36372 53518
rect 36316 53454 36318 53506
rect 36370 53454 36372 53506
rect 36316 53058 36372 53454
rect 36316 53006 36318 53058
rect 36370 53006 36372 53058
rect 36316 52994 36372 53006
rect 36204 52500 36260 52510
rect 36260 52444 36484 52500
rect 36204 52434 36260 52444
rect 35980 52334 35982 52386
rect 36034 52334 36036 52386
rect 35980 52322 36036 52334
rect 35980 51268 36036 51278
rect 35980 51174 36036 51212
rect 36204 50596 36260 50606
rect 36204 50502 36260 50540
rect 35308 50372 35700 50428
rect 35868 50418 35924 50428
rect 35084 47796 35140 50372
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35644 49252 35700 50372
rect 36204 49698 36260 49710
rect 36204 49646 36206 49698
rect 36258 49646 36260 49698
rect 35756 49252 35812 49262
rect 35644 49250 35812 49252
rect 35644 49198 35758 49250
rect 35810 49198 35812 49250
rect 35644 49196 35812 49198
rect 35756 49186 35812 49196
rect 35868 48916 35924 48926
rect 36204 48916 36260 49646
rect 35756 48914 36260 48916
rect 35756 48862 35870 48914
rect 35922 48862 36260 48914
rect 35756 48860 36260 48862
rect 35644 48804 35700 48814
rect 34972 47740 35140 47796
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 34412 47460 34468 47470
rect 34412 47366 34468 47404
rect 34636 47458 34692 47470
rect 34636 47406 34638 47458
rect 34690 47406 34692 47458
rect 34636 47124 34692 47406
rect 34636 47058 34692 47068
rect 34636 46788 34692 46798
rect 34636 45778 34692 46732
rect 34636 45726 34638 45778
rect 34690 45726 34692 45778
rect 34300 45666 34356 45678
rect 34300 45614 34302 45666
rect 34354 45614 34356 45666
rect 34300 45332 34356 45614
rect 34636 45332 34692 45726
rect 34300 45238 34356 45276
rect 34524 45276 34636 45332
rect 34524 41636 34580 45276
rect 34636 45266 34692 45276
rect 34636 44994 34692 45006
rect 34636 44942 34638 44994
rect 34690 44942 34692 44994
rect 34636 44772 34692 44942
rect 34636 43538 34692 44716
rect 34972 44996 35028 47740
rect 35084 47572 35140 47582
rect 35084 47234 35140 47516
rect 35084 47182 35086 47234
rect 35138 47182 35140 47234
rect 35084 45668 35140 47182
rect 35532 47236 35588 47246
rect 35532 46674 35588 47180
rect 35532 46622 35534 46674
rect 35586 46622 35588 46674
rect 35532 46610 35588 46622
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35196 45892 35252 45902
rect 35196 45798 35252 45836
rect 35532 45892 35588 45902
rect 35084 45602 35140 45612
rect 35084 45332 35140 45342
rect 35084 45238 35140 45276
rect 35532 45330 35588 45836
rect 35532 45278 35534 45330
rect 35586 45278 35588 45330
rect 35532 45266 35588 45278
rect 34972 44322 35028 44940
rect 35532 44882 35588 44894
rect 35532 44830 35534 44882
rect 35586 44830 35588 44882
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34972 44270 34974 44322
rect 35026 44270 35028 44322
rect 34972 44258 35028 44270
rect 35420 44324 35476 44334
rect 35532 44324 35588 44830
rect 35420 44322 35588 44324
rect 35420 44270 35422 44322
rect 35474 44270 35588 44322
rect 35420 44268 35588 44270
rect 35420 44258 35476 44268
rect 35196 44100 35252 44110
rect 35084 44044 35196 44100
rect 34636 43486 34638 43538
rect 34690 43486 34692 43538
rect 34636 43474 34692 43486
rect 34748 43650 34804 43662
rect 34748 43598 34750 43650
rect 34802 43598 34804 43650
rect 34748 42532 34804 43598
rect 34748 42466 34804 42476
rect 34972 42420 35028 42430
rect 34524 41570 34580 41580
rect 34860 42196 34916 42206
rect 34412 41186 34468 41198
rect 34412 41134 34414 41186
rect 34466 41134 34468 41186
rect 34188 40236 34356 40292
rect 34300 40068 34356 40236
rect 34300 40002 34356 40012
rect 34076 39666 34132 39676
rect 34188 39956 34244 39966
rect 33964 39414 34020 39452
rect 34076 39060 34132 39070
rect 34188 39060 34244 39900
rect 34076 39058 34244 39060
rect 34076 39006 34078 39058
rect 34130 39006 34244 39058
rect 34076 39004 34244 39006
rect 34076 38994 34132 39004
rect 33852 38780 34132 38836
rect 33740 38220 33908 38276
rect 33740 38050 33796 38062
rect 33740 37998 33742 38050
rect 33794 37998 33796 38050
rect 33740 37940 33796 37998
rect 33740 37874 33796 37884
rect 33628 36482 33684 37324
rect 33628 36430 33630 36482
rect 33682 36430 33684 36482
rect 33628 36418 33684 36430
rect 33740 37268 33796 37278
rect 33404 35476 33460 35980
rect 33404 35410 33460 35420
rect 33236 34412 33348 34468
rect 33180 34402 33236 34412
rect 33628 34356 33684 34366
rect 33628 34262 33684 34300
rect 33068 34242 33236 34244
rect 33068 34190 33070 34242
rect 33122 34190 33236 34242
rect 33068 34188 33236 34190
rect 33068 34178 33124 34188
rect 33180 34132 33236 34188
rect 33180 34076 33572 34132
rect 33292 33906 33348 33918
rect 33292 33854 33294 33906
rect 33346 33854 33348 33906
rect 33068 33796 33124 33806
rect 33068 30994 33124 33740
rect 33292 33572 33348 33854
rect 33180 33012 33236 33022
rect 33180 32450 33236 32956
rect 33180 32398 33182 32450
rect 33234 32398 33236 32450
rect 33180 31556 33236 32398
rect 33180 31490 33236 31500
rect 33068 30942 33070 30994
rect 33122 30942 33124 30994
rect 33068 30660 33124 30942
rect 33068 30594 33124 30604
rect 33292 30212 33348 33516
rect 33516 33458 33572 34076
rect 33516 33406 33518 33458
rect 33570 33406 33572 33458
rect 33516 33394 33572 33406
rect 33740 32676 33796 37212
rect 33628 32620 33796 32676
rect 33404 32452 33460 32462
rect 33404 31778 33460 32396
rect 33628 32004 33684 32620
rect 33628 31938 33684 31948
rect 33740 32450 33796 32462
rect 33740 32398 33742 32450
rect 33794 32398 33796 32450
rect 33404 31726 33406 31778
rect 33458 31726 33460 31778
rect 33404 31714 33460 31726
rect 33740 31780 33796 32398
rect 33628 31668 33684 31678
rect 33628 31108 33684 31612
rect 33516 31106 33684 31108
rect 33516 31054 33630 31106
rect 33682 31054 33684 31106
rect 33516 31052 33684 31054
rect 32956 29586 33012 29596
rect 33068 30156 33348 30212
rect 33404 30772 33460 30782
rect 33404 30212 33460 30716
rect 33516 30324 33572 31052
rect 33628 31042 33684 31052
rect 33740 30660 33796 31724
rect 33740 30594 33796 30604
rect 33740 30324 33796 30334
rect 33516 30268 33684 30324
rect 33404 30156 33572 30212
rect 32956 27748 33012 27758
rect 32844 27692 32956 27748
rect 32956 27682 33012 27692
rect 32620 27300 32676 27310
rect 32620 27186 32676 27244
rect 32620 27134 32622 27186
rect 32674 27134 32676 27186
rect 32620 27122 32676 27134
rect 32172 26908 32340 26964
rect 32172 25060 32228 26908
rect 32620 26628 32676 26638
rect 32284 26290 32340 26302
rect 32284 26238 32286 26290
rect 32338 26238 32340 26290
rect 32284 25284 32340 26238
rect 32396 26292 32452 26302
rect 32396 25620 32452 26236
rect 32396 25618 32564 25620
rect 32396 25566 32398 25618
rect 32450 25566 32564 25618
rect 32396 25564 32564 25566
rect 32396 25554 32452 25564
rect 32284 25218 32340 25228
rect 32172 25004 32340 25060
rect 31948 24050 32116 24052
rect 31948 23998 31950 24050
rect 32002 23998 32116 24050
rect 31948 23996 32116 23998
rect 31948 23986 32004 23996
rect 32172 23940 32228 23950
rect 32060 23938 32228 23940
rect 32060 23886 32174 23938
rect 32226 23886 32228 23938
rect 32060 23884 32228 23886
rect 32060 23716 32116 23884
rect 32172 23874 32228 23884
rect 31724 22540 31892 22596
rect 31724 22372 31780 22382
rect 31612 22370 31780 22372
rect 31612 22318 31726 22370
rect 31778 22318 31780 22370
rect 31612 22316 31780 22318
rect 31724 22306 31780 22316
rect 31388 22146 31444 22158
rect 31388 22094 31390 22146
rect 31442 22094 31444 22146
rect 31388 20916 31444 22094
rect 31500 21588 31556 21598
rect 31500 21494 31556 21532
rect 31388 20850 31444 20860
rect 31612 20802 31668 20814
rect 31612 20750 31614 20802
rect 31666 20750 31668 20802
rect 31612 19906 31668 20750
rect 31612 19854 31614 19906
rect 31666 19854 31668 19906
rect 31612 18564 31668 19854
rect 31612 18498 31668 18508
rect 31724 18340 31780 18350
rect 31388 18338 31780 18340
rect 31388 18286 31726 18338
rect 31778 18286 31780 18338
rect 31388 18284 31780 18286
rect 31388 17554 31444 18284
rect 31724 18274 31780 18284
rect 31836 18116 31892 22540
rect 32060 22148 32116 23660
rect 32172 23156 32228 23166
rect 32172 23042 32228 23100
rect 32172 22990 32174 23042
rect 32226 22990 32228 23042
rect 32172 22978 32228 22990
rect 32284 22260 32340 25004
rect 32396 24610 32452 24622
rect 32396 24558 32398 24610
rect 32450 24558 32452 24610
rect 32396 24500 32452 24558
rect 32508 24500 32564 25564
rect 32620 25506 32676 26572
rect 33068 26292 33124 30156
rect 33516 30098 33572 30156
rect 33516 30046 33518 30098
rect 33570 30046 33572 30098
rect 33516 30034 33572 30046
rect 33292 29988 33348 29998
rect 33292 29894 33348 29932
rect 33404 29986 33460 29998
rect 33404 29934 33406 29986
rect 33458 29934 33460 29986
rect 33180 29876 33236 29886
rect 33180 29650 33236 29820
rect 33180 29598 33182 29650
rect 33234 29598 33236 29650
rect 33180 28084 33236 29598
rect 33292 28756 33348 28766
rect 33404 28756 33460 29934
rect 33628 29650 33684 30268
rect 33740 30230 33796 30268
rect 33852 30212 33908 38220
rect 33964 37492 34020 37502
rect 33964 37378 34020 37436
rect 33964 37326 33966 37378
rect 34018 37326 34020 37378
rect 33964 37314 34020 37326
rect 33964 34020 34020 34030
rect 33964 33458 34020 33964
rect 33964 33406 33966 33458
rect 34018 33406 34020 33458
rect 33964 33348 34020 33406
rect 33964 33282 34020 33292
rect 34076 32676 34132 38780
rect 34188 37044 34244 39004
rect 34300 39172 34356 39182
rect 34300 38164 34356 39116
rect 34412 38612 34468 41134
rect 34636 41188 34692 41198
rect 34692 41132 34804 41188
rect 34636 41122 34692 41132
rect 34524 40964 34580 40974
rect 34524 40870 34580 40908
rect 34636 40962 34692 40974
rect 34636 40910 34638 40962
rect 34690 40910 34692 40962
rect 34636 40740 34692 40910
rect 34412 38546 34468 38556
rect 34524 40684 34692 40740
rect 34300 38108 34468 38164
rect 34300 37940 34356 37950
rect 34300 37846 34356 37884
rect 34412 37716 34468 38108
rect 34188 36978 34244 36988
rect 34300 37660 34468 37716
rect 34188 35812 34244 35822
rect 34188 33570 34244 35756
rect 34300 35028 34356 37660
rect 34524 37268 34580 40684
rect 34748 40404 34804 41132
rect 34860 40740 34916 42140
rect 34972 42194 35028 42364
rect 34972 42142 34974 42194
rect 35026 42142 35028 42194
rect 34972 42130 35028 42142
rect 35084 41524 35140 44044
rect 35196 44006 35252 44044
rect 35308 44098 35364 44110
rect 35532 44100 35588 44110
rect 35308 44046 35310 44098
rect 35362 44046 35364 44098
rect 35308 43316 35364 44046
rect 35420 44098 35588 44100
rect 35420 44046 35534 44098
rect 35586 44046 35588 44098
rect 35420 44044 35588 44046
rect 35420 43652 35476 44044
rect 35532 44034 35588 44044
rect 35420 43586 35476 43596
rect 35532 43650 35588 43662
rect 35532 43598 35534 43650
rect 35586 43598 35588 43650
rect 35532 43540 35588 43598
rect 35532 43474 35588 43484
rect 35308 43260 35588 43316
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35196 42868 35252 42878
rect 35196 42774 35252 42812
rect 35532 42754 35588 43260
rect 35532 42702 35534 42754
rect 35586 42702 35588 42754
rect 35532 42690 35588 42702
rect 35420 42642 35476 42654
rect 35420 42590 35422 42642
rect 35474 42590 35476 42642
rect 35420 42532 35476 42590
rect 35644 42532 35700 48748
rect 35756 45444 35812 48860
rect 35868 48850 35924 48860
rect 36316 48802 36372 52444
rect 36428 52274 36484 52444
rect 36428 52222 36430 52274
rect 36482 52222 36484 52274
rect 36428 52210 36484 52222
rect 36540 51266 36596 51278
rect 36540 51214 36542 51266
rect 36594 51214 36596 51266
rect 36540 50428 36596 51214
rect 37100 50818 37156 50830
rect 37100 50766 37102 50818
rect 37154 50766 37156 50818
rect 37100 50706 37156 50766
rect 37100 50654 37102 50706
rect 37154 50654 37156 50706
rect 37100 50428 37156 50654
rect 36316 48750 36318 48802
rect 36370 48750 36372 48802
rect 35980 48132 36036 48142
rect 35756 45378 35812 45388
rect 35868 48130 36036 48132
rect 35868 48078 35982 48130
rect 36034 48078 36036 48130
rect 35868 48076 36036 48078
rect 35868 47458 35924 48076
rect 35980 48066 36036 48076
rect 35868 47406 35870 47458
rect 35922 47406 35924 47458
rect 35868 44882 35924 47406
rect 36092 47460 36148 47470
rect 36316 47460 36372 48750
rect 36428 50372 36596 50428
rect 36988 50372 37156 50428
rect 37212 50428 37268 67118
rect 39228 67170 39284 67182
rect 39228 67118 39230 67170
rect 39282 67118 39284 67170
rect 38556 67060 38612 67070
rect 38332 67058 38612 67060
rect 38332 67006 38558 67058
rect 38610 67006 38612 67058
rect 38332 67004 38612 67006
rect 38332 66948 38388 67004
rect 38556 66994 38612 67004
rect 37772 66164 37828 66174
rect 37772 66070 37828 66108
rect 38108 65714 38164 65726
rect 38108 65662 38110 65714
rect 38162 65662 38164 65714
rect 37436 65602 37492 65614
rect 37436 65550 37438 65602
rect 37490 65550 37492 65602
rect 37324 64706 37380 64718
rect 37324 64654 37326 64706
rect 37378 64654 37380 64706
rect 37324 63140 37380 64654
rect 37324 62244 37380 63084
rect 37324 62178 37380 62188
rect 37436 64708 37492 65550
rect 37996 64820 38052 64830
rect 37772 64818 38052 64820
rect 37772 64766 37998 64818
rect 38050 64766 38052 64818
rect 37772 64764 38052 64766
rect 37548 64708 37604 64718
rect 37436 64706 37604 64708
rect 37436 64654 37550 64706
rect 37602 64654 37604 64706
rect 37436 64652 37604 64654
rect 37436 62188 37492 64652
rect 37548 64642 37604 64652
rect 37772 64036 37828 64764
rect 37996 64754 38052 64764
rect 37548 63980 37828 64036
rect 37548 63250 37604 63980
rect 37772 63922 37828 63980
rect 37772 63870 37774 63922
rect 37826 63870 37828 63922
rect 37772 63858 37828 63870
rect 37548 63198 37550 63250
rect 37602 63198 37604 63250
rect 37548 63186 37604 63198
rect 37660 63810 37716 63822
rect 37660 63758 37662 63810
rect 37714 63758 37716 63810
rect 37660 63140 37716 63758
rect 37996 63252 38052 63262
rect 37996 63158 38052 63196
rect 37660 63084 37828 63140
rect 37772 62916 37828 63084
rect 37772 62860 37940 62916
rect 37884 62188 37940 62860
rect 37436 62132 37716 62188
rect 37884 62132 38052 62188
rect 37548 61460 37604 61470
rect 37436 61404 37548 61460
rect 37436 61346 37492 61404
rect 37548 61394 37604 61404
rect 37436 61294 37438 61346
rect 37490 61294 37492 61346
rect 37436 61282 37492 61294
rect 37660 59108 37716 62132
rect 37884 59108 37940 59118
rect 37660 59106 37940 59108
rect 37660 59054 37886 59106
rect 37938 59054 37940 59106
rect 37660 59052 37940 59054
rect 37884 59042 37940 59052
rect 37548 58436 37604 58446
rect 37884 58436 37940 58446
rect 37604 58434 37940 58436
rect 37604 58382 37886 58434
rect 37938 58382 37940 58434
rect 37604 58380 37940 58382
rect 37548 58342 37604 58380
rect 37884 58212 37940 58380
rect 37884 58146 37940 58156
rect 37660 57988 37716 57998
rect 37996 57988 38052 62132
rect 37548 57932 37660 57988
rect 37324 54628 37380 54638
rect 37324 52386 37380 54572
rect 37324 52334 37326 52386
rect 37378 52334 37380 52386
rect 37324 50818 37380 52334
rect 37436 51940 37492 51950
rect 37436 51846 37492 51884
rect 37324 50766 37326 50818
rect 37378 50766 37380 50818
rect 37324 50754 37380 50766
rect 37212 50372 37380 50428
rect 36428 48468 36484 50372
rect 36540 49700 36596 49710
rect 36540 48804 36596 49644
rect 36540 48738 36596 48748
rect 36428 48412 36596 48468
rect 36428 48242 36484 48254
rect 36428 48190 36430 48242
rect 36482 48190 36484 48242
rect 36428 47682 36484 48190
rect 36428 47630 36430 47682
rect 36482 47630 36484 47682
rect 36428 47618 36484 47630
rect 36148 47404 36372 47460
rect 36092 47366 36148 47404
rect 36540 47124 36596 48412
rect 36764 48356 36820 48366
rect 36764 48262 36820 48300
rect 36988 48018 37044 50372
rect 37100 48804 37156 48814
rect 37100 48710 37156 48748
rect 36988 47966 36990 48018
rect 37042 47966 37044 48018
rect 36988 47954 37044 47966
rect 37100 48468 37156 48478
rect 37100 47458 37156 48412
rect 37100 47406 37102 47458
rect 37154 47406 37156 47458
rect 37100 47394 37156 47406
rect 37212 48130 37268 48142
rect 37212 48078 37214 48130
rect 37266 48078 37268 48130
rect 37212 47460 37268 48078
rect 37324 47572 37380 50372
rect 37324 47506 37380 47516
rect 36204 46900 36260 46910
rect 36204 46786 36260 46844
rect 36204 46734 36206 46786
rect 36258 46734 36260 46786
rect 36204 46722 36260 46734
rect 35868 44830 35870 44882
rect 35922 44830 35924 44882
rect 35868 44818 35924 44830
rect 35980 46116 36036 46126
rect 35980 44994 36036 46060
rect 36092 45892 36148 45902
rect 36092 45798 36148 45836
rect 35980 44942 35982 44994
rect 36034 44942 36036 44994
rect 35980 44436 36036 44942
rect 35980 44370 36036 44380
rect 35980 44210 36036 44222
rect 35980 44158 35982 44210
rect 36034 44158 36036 44210
rect 35868 43652 35924 43662
rect 35420 42476 35700 42532
rect 35756 42754 35812 42766
rect 35756 42702 35758 42754
rect 35810 42702 35812 42754
rect 35644 42196 35700 42206
rect 35532 41970 35588 41982
rect 35532 41918 35534 41970
rect 35586 41918 35588 41970
rect 34860 40514 34916 40684
rect 34860 40462 34862 40514
rect 34914 40462 34916 40514
rect 34860 40450 34916 40462
rect 34972 41468 35140 41524
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 34636 40402 34804 40404
rect 34636 40350 34750 40402
rect 34802 40350 34804 40402
rect 34636 40348 34804 40350
rect 34636 39060 34692 40348
rect 34748 40338 34804 40348
rect 34636 38994 34692 39004
rect 34748 40068 34804 40078
rect 34524 37202 34580 37212
rect 34636 38722 34692 38734
rect 34636 38670 34638 38722
rect 34690 38670 34692 38722
rect 34412 37044 34468 37054
rect 34412 37042 34580 37044
rect 34412 36990 34414 37042
rect 34466 36990 34580 37042
rect 34412 36988 34580 36990
rect 34412 36978 34468 36988
rect 34300 34962 34356 34972
rect 34412 34802 34468 34814
rect 34412 34750 34414 34802
rect 34466 34750 34468 34802
rect 34412 34356 34468 34750
rect 34412 34290 34468 34300
rect 34300 34020 34356 34030
rect 34300 33926 34356 33964
rect 34188 33518 34190 33570
rect 34242 33518 34244 33570
rect 34188 33506 34244 33518
rect 34524 33348 34580 36988
rect 34636 36708 34692 38670
rect 34748 37604 34804 40012
rect 34972 39396 35028 41468
rect 35532 41412 35588 41918
rect 35532 41346 35588 41356
rect 35644 41186 35700 42140
rect 35644 41134 35646 41186
rect 35698 41134 35700 41186
rect 35644 41122 35700 41134
rect 35532 41076 35588 41086
rect 35532 40982 35588 41020
rect 34972 39302 35028 39340
rect 35084 40964 35140 40974
rect 34972 37828 35028 37838
rect 35084 37828 35140 40908
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35196 39732 35252 39742
rect 35196 39638 35252 39676
rect 35756 38668 35812 42702
rect 35868 42196 35924 43596
rect 35868 42130 35924 42140
rect 35980 42084 36036 44158
rect 36316 44098 36372 44110
rect 36316 44046 36318 44098
rect 36370 44046 36372 44098
rect 36204 43764 36260 43774
rect 35980 42018 36036 42028
rect 36092 43708 36204 43764
rect 36092 42082 36148 43708
rect 36204 43698 36260 43708
rect 36316 43652 36372 44046
rect 36316 43586 36372 43596
rect 36092 42030 36094 42082
rect 36146 42030 36148 42082
rect 36092 42018 36148 42030
rect 36204 42530 36260 42542
rect 36204 42478 36206 42530
rect 36258 42478 36260 42530
rect 35980 41858 36036 41870
rect 35980 41806 35982 41858
rect 36034 41806 36036 41858
rect 35868 40516 35924 40526
rect 35868 40290 35924 40460
rect 35868 40238 35870 40290
rect 35922 40238 35924 40290
rect 35868 40226 35924 40238
rect 35532 38612 35812 38668
rect 35868 38612 35924 38622
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34972 37826 35140 37828
rect 34972 37774 34974 37826
rect 35026 37774 35140 37826
rect 34972 37772 35140 37774
rect 34748 37548 34916 37604
rect 34748 37378 34804 37390
rect 34748 37326 34750 37378
rect 34802 37326 34804 37378
rect 34748 37156 34804 37326
rect 34748 37090 34804 37100
rect 34636 36642 34692 36652
rect 34860 37044 34916 37548
rect 34636 36260 34692 36270
rect 34748 36260 34804 36270
rect 34636 36258 34748 36260
rect 34636 36206 34638 36258
rect 34690 36206 34748 36258
rect 34636 36204 34748 36206
rect 34636 36194 34692 36204
rect 34748 35586 34804 36204
rect 34748 35534 34750 35586
rect 34802 35534 34804 35586
rect 34748 35474 34804 35534
rect 34748 35422 34750 35474
rect 34802 35422 34804 35474
rect 34748 35410 34804 35422
rect 34748 34690 34804 34702
rect 34748 34638 34750 34690
rect 34802 34638 34804 34690
rect 34748 34244 34804 34638
rect 34748 34178 34804 34188
rect 34636 34130 34692 34142
rect 34636 34078 34638 34130
rect 34690 34078 34692 34130
rect 34636 34020 34692 34078
rect 34748 34020 34804 34030
rect 34636 33964 34748 34020
rect 34748 33954 34804 33964
rect 33964 32620 34132 32676
rect 34188 33292 34580 33348
rect 34636 33684 34692 33694
rect 33964 31108 34020 32620
rect 34076 32452 34132 32462
rect 34076 32358 34132 32396
rect 34188 32004 34244 33292
rect 34300 33124 34356 33134
rect 34300 32452 34356 33068
rect 34412 33122 34468 33134
rect 34412 33070 34414 33122
rect 34466 33070 34468 33122
rect 34412 32788 34468 33070
rect 34524 33124 34580 33134
rect 34636 33124 34692 33628
rect 34524 33122 34692 33124
rect 34524 33070 34526 33122
rect 34578 33070 34692 33122
rect 34524 33068 34692 33070
rect 34524 33058 34580 33068
rect 34636 32900 34692 32910
rect 34524 32788 34580 32798
rect 34468 32786 34580 32788
rect 34468 32734 34526 32786
rect 34578 32734 34580 32786
rect 34468 32732 34580 32734
rect 34412 32694 34468 32732
rect 34524 32722 34580 32732
rect 34300 32386 34356 32396
rect 33964 31042 34020 31052
rect 34076 31948 34244 32004
rect 33964 30548 34020 30558
rect 33964 30434 34020 30492
rect 33964 30382 33966 30434
rect 34018 30382 34020 30434
rect 33964 30370 34020 30382
rect 34076 30212 34132 31948
rect 34188 31668 34244 31678
rect 34188 31666 34580 31668
rect 34188 31614 34190 31666
rect 34242 31614 34580 31666
rect 34188 31612 34580 31614
rect 34188 31602 34244 31612
rect 34188 31444 34244 31454
rect 34188 30434 34244 31388
rect 34300 31108 34356 31118
rect 34356 31052 34468 31108
rect 34300 31042 34356 31052
rect 34188 30382 34190 30434
rect 34242 30382 34244 30434
rect 34188 30324 34244 30382
rect 34300 30324 34356 30334
rect 34188 30268 34300 30324
rect 34300 30258 34356 30268
rect 33852 30156 34020 30212
rect 34076 30156 34244 30212
rect 33628 29598 33630 29650
rect 33682 29598 33684 29650
rect 33628 29586 33684 29598
rect 33740 29876 33796 29886
rect 33740 29428 33796 29820
rect 33964 29428 34020 30156
rect 34076 29876 34132 29886
rect 34076 29650 34132 29820
rect 34076 29598 34078 29650
rect 34130 29598 34132 29650
rect 34076 29586 34132 29598
rect 33628 29372 33796 29428
rect 33852 29372 34020 29428
rect 33516 28868 33572 28878
rect 33516 28774 33572 28812
rect 33292 28754 33460 28756
rect 33292 28702 33294 28754
rect 33346 28702 33460 28754
rect 33292 28700 33460 28702
rect 33292 28690 33348 28700
rect 33628 28532 33684 29372
rect 33740 28756 33796 28766
rect 33740 28662 33796 28700
rect 33628 28476 33796 28532
rect 33628 28308 33684 28318
rect 33180 28082 33572 28084
rect 33180 28030 33182 28082
rect 33234 28030 33572 28082
rect 33180 28028 33572 28030
rect 33180 28018 33236 28028
rect 33516 27300 33572 28028
rect 33628 28082 33684 28252
rect 33628 28030 33630 28082
rect 33682 28030 33684 28082
rect 33628 28018 33684 28030
rect 33516 27244 33684 27300
rect 33516 27076 33572 27086
rect 33068 26198 33124 26236
rect 33180 27074 33572 27076
rect 33180 27022 33518 27074
rect 33570 27022 33572 27074
rect 33180 27020 33572 27022
rect 33180 26850 33236 27020
rect 33516 27010 33572 27020
rect 33628 26908 33684 27244
rect 33180 26798 33182 26850
rect 33234 26798 33236 26850
rect 32620 25454 32622 25506
rect 32674 25454 32676 25506
rect 32620 25442 32676 25454
rect 33180 25508 33236 26798
rect 33516 26852 33684 26908
rect 33180 25452 33460 25508
rect 32956 25396 33012 25406
rect 32956 25394 33348 25396
rect 32956 25342 32958 25394
rect 33010 25342 33348 25394
rect 32956 25340 33348 25342
rect 32956 25330 33012 25340
rect 32844 25282 32900 25294
rect 32844 25230 32846 25282
rect 32898 25230 32900 25282
rect 32844 24500 32900 25230
rect 32508 24444 32676 24500
rect 32396 23828 32452 24444
rect 32508 24050 32564 24062
rect 32508 23998 32510 24050
rect 32562 23998 32564 24050
rect 32508 23940 32564 23998
rect 32508 23874 32564 23884
rect 32396 23762 32452 23772
rect 32508 23716 32564 23726
rect 32508 22482 32564 23660
rect 32620 23548 32676 24444
rect 32844 24434 32900 24444
rect 32956 24948 33012 24958
rect 32844 23716 32900 23726
rect 32844 23622 32900 23660
rect 32620 23492 32788 23548
rect 32508 22430 32510 22482
rect 32562 22430 32564 22482
rect 32508 22418 32564 22430
rect 32284 22204 32564 22260
rect 32060 22092 32452 22148
rect 31948 21812 32004 21822
rect 32004 21756 32228 21812
rect 31948 21718 32004 21756
rect 32172 20242 32228 21756
rect 32284 20916 32340 20926
rect 32284 20822 32340 20860
rect 32396 20692 32452 22092
rect 32172 20190 32174 20242
rect 32226 20190 32228 20242
rect 32172 20178 32228 20190
rect 32284 20636 32452 20692
rect 31388 17502 31390 17554
rect 31442 17502 31444 17554
rect 31388 17490 31444 17502
rect 31724 18060 31892 18116
rect 32060 20132 32116 20142
rect 31612 16770 31668 16782
rect 31612 16718 31614 16770
rect 31666 16718 31668 16770
rect 31388 16660 31444 16670
rect 31388 16566 31444 16604
rect 31388 16322 31444 16334
rect 31388 16270 31390 16322
rect 31442 16270 31444 16322
rect 31388 16210 31444 16270
rect 31388 16158 31390 16210
rect 31442 16158 31444 16210
rect 31388 16146 31444 16158
rect 31276 15932 31444 15988
rect 30828 15372 30996 15428
rect 30828 14644 30884 15372
rect 31164 15204 31220 15242
rect 30828 14578 30884 14588
rect 30940 15092 31220 15148
rect 30828 14420 30884 14430
rect 30828 14326 30884 14364
rect 30940 13186 30996 15092
rect 31276 13748 31332 13758
rect 30940 13134 30942 13186
rect 30994 13134 30996 13186
rect 30940 12292 30996 13134
rect 30940 12226 30996 12236
rect 31052 13746 31332 13748
rect 31052 13694 31278 13746
rect 31330 13694 31332 13746
rect 31052 13692 31332 13694
rect 31052 10050 31108 13692
rect 31276 13682 31332 13692
rect 31388 13634 31444 15932
rect 31612 15876 31668 16718
rect 31612 15148 31668 15820
rect 31500 15092 31668 15148
rect 31500 14642 31556 15092
rect 31724 14868 31780 18060
rect 31500 14590 31502 14642
rect 31554 14590 31556 14642
rect 31500 14578 31556 14590
rect 31612 14812 31780 14868
rect 32060 17106 32116 20076
rect 32060 17054 32062 17106
rect 32114 17054 32116 17106
rect 32060 16660 32116 17054
rect 31612 14084 31668 14812
rect 31388 13582 31390 13634
rect 31442 13582 31444 13634
rect 31388 13570 31444 13582
rect 31500 14028 31668 14084
rect 31724 14644 31780 14654
rect 31500 10948 31556 14028
rect 31612 13858 31668 13870
rect 31612 13806 31614 13858
rect 31666 13806 31668 13858
rect 31612 13186 31668 13806
rect 31612 13134 31614 13186
rect 31666 13134 31668 13186
rect 31612 13122 31668 13134
rect 31724 12964 31780 14588
rect 32060 14420 32116 16604
rect 32060 13748 32116 14364
rect 32060 13682 32116 13692
rect 32284 13076 32340 20636
rect 32396 18450 32452 18462
rect 32396 18398 32398 18450
rect 32450 18398 32452 18450
rect 32396 18340 32452 18398
rect 32396 18274 32452 18284
rect 32508 15148 32564 22204
rect 32620 17556 32676 17566
rect 32732 17556 32788 23492
rect 32956 20916 33012 24892
rect 33180 24836 33236 24846
rect 33068 23940 33124 23950
rect 33068 23846 33124 23884
rect 32956 20850 33012 20860
rect 33180 23380 33236 24780
rect 33180 20132 33236 23324
rect 33180 20066 33236 20076
rect 32676 17500 32788 17556
rect 33068 18340 33124 18350
rect 33180 18340 33236 18350
rect 33124 18338 33236 18340
rect 33124 18286 33182 18338
rect 33234 18286 33236 18338
rect 33124 18284 33236 18286
rect 32620 17490 32676 17500
rect 33068 15204 33124 18284
rect 33180 18274 33236 18284
rect 33180 17780 33236 17790
rect 33180 17686 33236 17724
rect 33292 17106 33348 25340
rect 33404 25284 33460 25452
rect 33404 23156 33460 25228
rect 33404 23090 33460 23100
rect 33516 21812 33572 26852
rect 33516 21746 33572 21756
rect 33740 19908 33796 28476
rect 33740 19842 33796 19852
rect 33516 17780 33572 17790
rect 33516 17666 33572 17724
rect 33516 17614 33518 17666
rect 33570 17614 33572 17666
rect 33516 17602 33572 17614
rect 33292 17054 33294 17106
rect 33346 17054 33348 17106
rect 33292 17042 33348 17054
rect 33628 17220 33684 17230
rect 33516 16996 33572 17006
rect 33516 16902 33572 16940
rect 33628 16994 33684 17164
rect 33852 17108 33908 29372
rect 33964 29204 34020 29214
rect 33964 28866 34020 29148
rect 34188 29092 34244 30156
rect 33964 28814 33966 28866
rect 34018 28814 34020 28866
rect 33964 28802 34020 28814
rect 34076 29036 34244 29092
rect 34412 30100 34468 31052
rect 34524 30434 34580 31612
rect 34636 31106 34692 32844
rect 34636 31054 34638 31106
rect 34690 31054 34692 31106
rect 34636 30772 34692 31054
rect 34748 31220 34804 31230
rect 34748 30994 34804 31164
rect 34748 30942 34750 30994
rect 34802 30942 34804 30994
rect 34748 30930 34804 30942
rect 34860 30772 34916 36988
rect 34972 36484 35028 37772
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35308 36708 35364 36718
rect 35084 36484 35140 36494
rect 34972 36482 35140 36484
rect 34972 36430 35086 36482
rect 35138 36430 35140 36482
rect 34972 36428 35140 36430
rect 35084 36418 35140 36428
rect 35308 36482 35364 36652
rect 35420 36596 35476 36606
rect 35532 36596 35588 38612
rect 35868 38164 35924 38556
rect 35868 38070 35924 38108
rect 35420 36594 35588 36596
rect 35420 36542 35422 36594
rect 35474 36542 35588 36594
rect 35420 36540 35588 36542
rect 35644 38052 35700 38062
rect 35420 36530 35476 36540
rect 35308 36430 35310 36482
rect 35362 36430 35364 36482
rect 35308 36418 35364 36430
rect 35532 36260 35588 36270
rect 35532 36166 35588 36204
rect 35196 35700 35252 35710
rect 35196 35606 35252 35644
rect 35644 35588 35700 37996
rect 35756 36370 35812 36382
rect 35756 36318 35758 36370
rect 35810 36318 35812 36370
rect 35756 35700 35812 36318
rect 35980 35812 36036 41806
rect 36092 41524 36148 41534
rect 36092 41410 36148 41468
rect 36092 41358 36094 41410
rect 36146 41358 36148 41410
rect 36092 41346 36148 41358
rect 36092 38052 36148 38062
rect 36092 37958 36148 37996
rect 36204 37492 36260 42478
rect 36316 41298 36372 41310
rect 36316 41246 36318 41298
rect 36370 41246 36372 41298
rect 36316 41188 36372 41246
rect 36316 41122 36372 41132
rect 36540 41076 36596 47068
rect 37212 47012 37268 47404
rect 36988 46956 37268 47012
rect 36540 41010 36596 41020
rect 36652 44996 36708 45006
rect 36316 40962 36372 40974
rect 36316 40910 36318 40962
rect 36370 40910 36372 40962
rect 36316 40852 36372 40910
rect 36316 40786 36372 40796
rect 36652 40628 36708 44940
rect 36764 44994 36820 45006
rect 36764 44942 36766 44994
rect 36818 44942 36820 44994
rect 36764 42756 36820 44942
rect 36988 43316 37044 46956
rect 37100 46788 37156 46798
rect 37100 46694 37156 46732
rect 37548 46564 37604 57932
rect 37660 57922 37716 57932
rect 37772 57932 38052 57988
rect 38108 57988 38164 65662
rect 38332 65492 38388 66892
rect 39228 66388 39284 67118
rect 38332 65490 38612 65492
rect 38332 65438 38334 65490
rect 38386 65438 38612 65490
rect 38332 65436 38612 65438
rect 38332 65426 38388 65436
rect 38556 63924 38612 65436
rect 39228 65490 39284 66332
rect 39900 66388 39956 66398
rect 39900 66294 39956 66332
rect 39228 65438 39230 65490
rect 39282 65438 39284 65490
rect 39228 65426 39284 65438
rect 39004 65380 39060 65390
rect 39004 65286 39060 65324
rect 39676 65380 39732 65390
rect 38444 63922 38612 63924
rect 38444 63870 38558 63922
rect 38610 63870 38612 63922
rect 38444 63868 38612 63870
rect 38444 63252 38500 63868
rect 38556 63858 38612 63868
rect 38668 65266 38724 65278
rect 38668 65214 38670 65266
rect 38722 65214 38724 65266
rect 38668 63700 38724 65214
rect 39676 64148 39732 65324
rect 40796 64706 40852 64718
rect 40796 64654 40798 64706
rect 40850 64654 40852 64706
rect 40124 64596 40180 64606
rect 38444 63186 38500 63196
rect 38556 63644 38724 63700
rect 39228 64146 39732 64148
rect 39228 64094 39678 64146
rect 39730 64094 39732 64146
rect 39228 64092 39732 64094
rect 38556 63138 38612 63644
rect 39228 63252 39284 64092
rect 39676 64082 39732 64092
rect 39788 64594 40180 64596
rect 39788 64542 40126 64594
rect 40178 64542 40180 64594
rect 39788 64540 40180 64542
rect 39228 63158 39284 63196
rect 39788 63140 39844 64540
rect 40124 64530 40180 64540
rect 38556 63086 38558 63138
rect 38610 63086 38612 63138
rect 38556 63074 38612 63086
rect 39340 63084 39844 63140
rect 38780 63028 38836 63038
rect 39340 63028 39396 63084
rect 38780 63026 39396 63028
rect 38780 62974 38782 63026
rect 38834 62974 39396 63026
rect 38780 62972 39396 62974
rect 38780 62962 38836 62972
rect 39116 62354 39172 62366
rect 39116 62302 39118 62354
rect 39170 62302 39172 62354
rect 38444 62242 38500 62254
rect 38444 62190 38446 62242
rect 38498 62190 38500 62242
rect 38444 61460 38500 62190
rect 38444 61394 38500 61404
rect 39116 61684 39172 62302
rect 39564 61684 39620 61694
rect 39116 61682 39956 61684
rect 39116 61630 39566 61682
rect 39618 61630 39956 61682
rect 39116 61628 39956 61630
rect 38556 58324 38612 58334
rect 38444 58322 38612 58324
rect 38444 58270 38558 58322
rect 38610 58270 38612 58322
rect 38444 58268 38612 58270
rect 37660 52164 37716 52174
rect 37660 52070 37716 52108
rect 37660 51604 37716 51614
rect 37660 50708 37716 51548
rect 37660 50614 37716 50652
rect 37772 50428 37828 57932
rect 38108 57922 38164 57932
rect 38220 58100 38276 58110
rect 38108 57540 38164 57550
rect 38220 57540 38276 58044
rect 38108 57538 38276 57540
rect 38108 57486 38110 57538
rect 38162 57486 38276 57538
rect 38108 57484 38276 57486
rect 38444 57538 38500 58268
rect 38556 58258 38612 58268
rect 39116 58212 39172 61628
rect 39564 61618 39620 61628
rect 39900 61572 39956 61628
rect 40124 61572 40180 61582
rect 39900 61570 40124 61572
rect 39900 61518 39902 61570
rect 39954 61518 40124 61570
rect 39900 61516 40124 61518
rect 39900 61506 39956 61516
rect 39116 58146 39172 58156
rect 39676 60674 39732 60686
rect 39676 60622 39678 60674
rect 39730 60622 39732 60674
rect 39676 60564 39732 60622
rect 40012 60564 40068 60574
rect 39676 60562 40068 60564
rect 39676 60510 40014 60562
rect 40066 60510 40068 60562
rect 39676 60508 40068 60510
rect 39676 59780 39732 60508
rect 40012 60498 40068 60508
rect 40124 60114 40180 61516
rect 40796 61572 40852 64654
rect 42812 61684 42868 61694
rect 40684 61460 40740 61470
rect 40348 61458 40740 61460
rect 40348 61406 40686 61458
rect 40738 61406 40740 61458
rect 40348 61404 40740 61406
rect 40236 60898 40292 60910
rect 40236 60846 40238 60898
rect 40290 60846 40292 60898
rect 40236 60452 40292 60846
rect 40348 60674 40404 61404
rect 40684 61394 40740 61404
rect 40796 60788 40852 61516
rect 42364 61682 42868 61684
rect 42364 61630 42814 61682
rect 42866 61630 42868 61682
rect 42364 61628 42868 61630
rect 40908 60788 40964 60798
rect 40796 60786 40964 60788
rect 40796 60734 40910 60786
rect 40962 60734 40964 60786
rect 40796 60732 40964 60734
rect 40908 60722 40964 60732
rect 41692 60676 41748 60686
rect 40348 60622 40350 60674
rect 40402 60622 40404 60674
rect 40348 60610 40404 60622
rect 41244 60674 41748 60676
rect 41244 60622 41694 60674
rect 41746 60622 41748 60674
rect 41244 60620 41748 60622
rect 40236 60396 40516 60452
rect 40124 60062 40126 60114
rect 40178 60062 40180 60114
rect 40124 60050 40180 60062
rect 38444 57486 38446 57538
rect 38498 57486 38500 57538
rect 38108 57474 38164 57484
rect 38444 57474 38500 57486
rect 38556 57762 38612 57774
rect 38556 57710 38558 57762
rect 38610 57710 38612 57762
rect 38444 56756 38500 56766
rect 38220 56754 38500 56756
rect 38220 56702 38446 56754
rect 38498 56702 38500 56754
rect 38220 56700 38500 56702
rect 38220 55970 38276 56700
rect 38444 56690 38500 56700
rect 38220 55918 38222 55970
rect 38274 55918 38276 55970
rect 38220 55906 38276 55918
rect 38556 56642 38612 57710
rect 38780 57764 38836 57774
rect 38780 57670 38836 57708
rect 39676 57764 39732 59724
rect 40460 58324 40516 60396
rect 41244 60226 41300 60620
rect 41692 60610 41748 60620
rect 41244 60174 41246 60226
rect 41298 60174 41300 60226
rect 41244 60162 41300 60174
rect 42364 60114 42420 61628
rect 42812 61618 42868 61628
rect 42364 60062 42366 60114
rect 42418 60062 42420 60114
rect 42364 60050 42420 60062
rect 42812 60676 42868 60686
rect 42812 60114 42868 60620
rect 43820 60676 43876 60686
rect 43820 60582 43876 60620
rect 42812 60062 42814 60114
rect 42866 60062 42868 60114
rect 42812 60050 42868 60062
rect 41244 60004 41300 60014
rect 41244 60002 41524 60004
rect 41244 59950 41246 60002
rect 41298 59950 41524 60002
rect 41244 59948 41524 59950
rect 41244 59938 41300 59948
rect 40908 59890 40964 59902
rect 40908 59838 40910 59890
rect 40962 59838 40964 59890
rect 40572 59780 40628 59790
rect 40908 59780 40964 59838
rect 40628 59724 40964 59780
rect 41468 59780 41524 59948
rect 40572 59686 40628 59724
rect 40684 58548 40740 58558
rect 41132 58548 41188 58558
rect 40684 58546 41188 58548
rect 40684 58494 40686 58546
rect 40738 58494 41134 58546
rect 41186 58494 41188 58546
rect 40684 58492 41188 58494
rect 40684 58482 40740 58492
rect 41132 58482 41188 58492
rect 41020 58324 41076 58334
rect 40460 58322 41188 58324
rect 40460 58270 41022 58322
rect 41074 58270 41188 58322
rect 40460 58268 41188 58270
rect 41020 58258 41076 58268
rect 39676 57698 39732 57708
rect 38556 56590 38558 56642
rect 38610 56590 38612 56642
rect 38556 55524 38612 56590
rect 41020 56642 41076 56654
rect 41020 56590 41022 56642
rect 41074 56590 41076 56642
rect 38220 55468 38612 55524
rect 38668 56308 38724 56318
rect 38220 52274 38276 55468
rect 38444 55300 38500 55310
rect 38668 55300 38724 56252
rect 41020 56308 41076 56590
rect 38444 55298 38724 55300
rect 38444 55246 38446 55298
rect 38498 55246 38724 55298
rect 38444 55244 38724 55246
rect 40684 56084 40740 56094
rect 38444 55234 38500 55244
rect 39116 55188 39172 55198
rect 39004 55186 39172 55188
rect 39004 55134 39118 55186
rect 39170 55134 39172 55186
rect 39004 55132 39172 55134
rect 38332 54628 38388 54638
rect 38332 54534 38388 54572
rect 38892 54626 38948 54638
rect 38892 54574 38894 54626
rect 38946 54574 38948 54626
rect 38668 54404 38724 54414
rect 38668 54310 38724 54348
rect 38556 53620 38612 53630
rect 38444 53618 38612 53620
rect 38444 53566 38558 53618
rect 38610 53566 38612 53618
rect 38444 53564 38612 53566
rect 38444 52834 38500 53564
rect 38556 53554 38612 53564
rect 38668 53506 38724 53518
rect 38668 53454 38670 53506
rect 38722 53454 38724 53506
rect 38668 53396 38724 53454
rect 38892 53396 38948 54574
rect 39004 54402 39060 55132
rect 39116 55122 39172 55132
rect 39004 54350 39006 54402
rect 39058 54350 39060 54402
rect 39004 54338 39060 54350
rect 40236 53508 40292 53518
rect 40236 53506 40404 53508
rect 40236 53454 40238 53506
rect 40290 53454 40404 53506
rect 40236 53452 40404 53454
rect 40236 53442 40292 53452
rect 38668 53340 39396 53396
rect 38892 53172 38948 53182
rect 38892 53078 38948 53116
rect 38444 52782 38446 52834
rect 38498 52782 38500 52834
rect 38444 52770 38500 52782
rect 38220 52222 38222 52274
rect 38274 52222 38276 52274
rect 38220 52210 38276 52222
rect 38332 52276 38388 52286
rect 38332 52162 38388 52220
rect 38332 52110 38334 52162
rect 38386 52110 38388 52162
rect 38332 52098 38388 52110
rect 39228 52162 39284 52174
rect 39228 52110 39230 52162
rect 39282 52110 39284 52162
rect 38668 51940 38724 51950
rect 38668 51490 38724 51884
rect 39228 51604 39284 52110
rect 39340 52164 39396 53340
rect 40236 52836 40292 52846
rect 39676 52388 39732 52398
rect 39676 52386 40068 52388
rect 39676 52334 39678 52386
rect 39730 52334 40068 52386
rect 39676 52332 40068 52334
rect 39676 52322 39732 52332
rect 39564 52164 39620 52174
rect 39340 52162 39620 52164
rect 39340 52110 39566 52162
rect 39618 52110 39620 52162
rect 39340 52108 39620 52110
rect 39564 52098 39620 52108
rect 39900 52052 39956 52062
rect 39900 51604 39956 51996
rect 39228 51538 39284 51548
rect 39452 51602 39956 51604
rect 39452 51550 39902 51602
rect 39954 51550 39956 51602
rect 39452 51548 39956 51550
rect 38668 51438 38670 51490
rect 38722 51438 38724 51490
rect 38668 51426 38724 51438
rect 38332 51380 38388 51390
rect 37772 50372 38052 50428
rect 37660 49028 37716 49038
rect 37660 48468 37716 48972
rect 37660 48374 37716 48412
rect 37772 48356 37828 48366
rect 37772 47570 37828 48300
rect 37772 47518 37774 47570
rect 37826 47518 37828 47570
rect 37772 47506 37828 47518
rect 37212 46508 37828 46564
rect 37100 44996 37156 45006
rect 37100 44902 37156 44940
rect 37212 44772 37268 46508
rect 37772 46002 37828 46508
rect 37772 45950 37774 46002
rect 37826 45950 37828 46002
rect 37772 45938 37828 45950
rect 37884 46562 37940 46574
rect 37884 46510 37886 46562
rect 37938 46510 37940 46562
rect 37100 44716 37268 44772
rect 37324 45666 37380 45678
rect 37324 45614 37326 45666
rect 37378 45614 37380 45666
rect 37100 43538 37156 44716
rect 37212 44100 37268 44110
rect 37212 44006 37268 44044
rect 37324 43652 37380 45614
rect 37772 45668 37828 45678
rect 37548 45444 37604 45454
rect 37548 45106 37604 45388
rect 37548 45054 37550 45106
rect 37602 45054 37604 45106
rect 37548 44324 37604 45054
rect 37548 44258 37604 44268
rect 37660 44322 37716 44334
rect 37660 44270 37662 44322
rect 37714 44270 37716 44322
rect 37100 43486 37102 43538
rect 37154 43486 37156 43538
rect 37100 43474 37156 43486
rect 37212 43596 37380 43652
rect 37660 44212 37716 44270
rect 37212 43540 37268 43596
rect 37436 43540 37492 43550
rect 37212 43474 37268 43484
rect 37324 43538 37492 43540
rect 37324 43486 37438 43538
rect 37490 43486 37492 43538
rect 37324 43484 37492 43486
rect 36988 43260 37268 43316
rect 36764 42690 36820 42700
rect 36988 42530 37044 42542
rect 36988 42478 36990 42530
rect 37042 42478 37044 42530
rect 36988 42196 37044 42478
rect 36988 42130 37044 42140
rect 37100 41412 37156 41422
rect 37100 41298 37156 41356
rect 37100 41246 37102 41298
rect 37154 41246 37156 41298
rect 37100 41234 37156 41246
rect 36540 40572 36708 40628
rect 36764 40740 36820 40750
rect 36428 40180 36484 40190
rect 36428 39730 36484 40124
rect 36428 39678 36430 39730
rect 36482 39678 36484 39730
rect 36428 39666 36484 39678
rect 36540 38668 36596 40572
rect 36652 40402 36708 40414
rect 36652 40350 36654 40402
rect 36706 40350 36708 40402
rect 36652 39172 36708 40350
rect 36764 40180 36820 40684
rect 37212 40404 37268 43260
rect 37324 42308 37380 43484
rect 37436 43474 37492 43484
rect 37548 42756 37604 42766
rect 37436 42644 37492 42654
rect 37436 42550 37492 42588
rect 37548 42420 37604 42700
rect 37660 42754 37716 44156
rect 37772 44210 37828 45612
rect 37772 44158 37774 44210
rect 37826 44158 37828 44210
rect 37772 44146 37828 44158
rect 37660 42702 37662 42754
rect 37714 42702 37716 42754
rect 37660 42690 37716 42702
rect 37548 42364 37716 42420
rect 37324 42252 37604 42308
rect 37324 42084 37380 42094
rect 37324 41990 37380 42028
rect 37548 41186 37604 42252
rect 37548 41134 37550 41186
rect 37602 41134 37604 41186
rect 37436 40404 37492 40414
rect 37212 40402 37492 40404
rect 37212 40350 37438 40402
rect 37490 40350 37492 40402
rect 37212 40348 37492 40350
rect 36764 40114 36820 40124
rect 37100 39732 37156 39742
rect 37100 39638 37156 39676
rect 37436 39620 37492 40348
rect 37548 39844 37604 41134
rect 37660 41076 37716 42364
rect 37660 41010 37716 41020
rect 37548 39778 37604 39788
rect 37772 40292 37828 40302
rect 37436 39564 37604 39620
rect 36652 39106 36708 39116
rect 37436 38834 37492 38846
rect 37436 38782 37438 38834
rect 37490 38782 37492 38834
rect 36092 37436 36260 37492
rect 36316 38612 36596 38668
rect 36764 38722 36820 38734
rect 36764 38670 36766 38722
rect 36818 38670 36820 38722
rect 36764 38668 36820 38670
rect 36764 38612 37044 38668
rect 36092 36484 36148 37436
rect 36204 37268 36260 37278
rect 36204 37174 36260 37212
rect 36092 36418 36148 36428
rect 36204 36258 36260 36270
rect 36204 36206 36206 36258
rect 36258 36206 36260 36258
rect 35980 35756 36148 35812
rect 35756 35644 36036 35700
rect 34972 35474 35028 35486
rect 34972 35422 34974 35474
rect 35026 35422 35028 35474
rect 34972 34916 35028 35422
rect 35084 35476 35140 35486
rect 35084 35140 35140 35420
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 35140 35252 35150
rect 35084 35084 35196 35140
rect 35196 35074 35252 35084
rect 34972 34860 35140 34916
rect 34972 34692 35028 34702
rect 34972 33684 35028 34636
rect 34972 33346 35028 33628
rect 34972 33294 34974 33346
rect 35026 33294 35028 33346
rect 34972 33282 35028 33294
rect 35084 33348 35140 34860
rect 35420 34244 35476 34254
rect 35420 34150 35476 34188
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35644 33460 35700 35532
rect 35980 35586 36036 35644
rect 35980 35534 35982 35586
rect 36034 35534 36036 35586
rect 35756 33460 35812 33470
rect 35644 33458 35812 33460
rect 35644 33406 35758 33458
rect 35810 33406 35812 33458
rect 35644 33404 35812 33406
rect 35084 33292 35308 33348
rect 35252 33236 35308 33292
rect 35252 33180 35364 33236
rect 35308 32900 35364 33180
rect 35084 32844 35364 32900
rect 34636 30716 34804 30772
rect 34524 30382 34526 30434
rect 34578 30382 34580 30434
rect 34524 30370 34580 30382
rect 34636 30548 34692 30558
rect 34636 30212 34692 30492
rect 34076 22260 34132 29036
rect 34412 28980 34468 30044
rect 34412 28914 34468 28924
rect 34524 30156 34692 30212
rect 34748 30212 34804 30716
rect 34860 30706 34916 30716
rect 34972 31444 35028 31454
rect 34972 30996 35028 31388
rect 34860 30436 34916 30446
rect 34860 30342 34916 30380
rect 34748 30156 34916 30212
rect 34524 29540 34580 30156
rect 34636 29988 34692 29998
rect 34692 29932 34804 29988
rect 34636 29894 34692 29932
rect 34524 28868 34580 29484
rect 34636 29428 34692 29438
rect 34636 29334 34692 29372
rect 34748 28868 34804 29932
rect 34860 29540 34916 30156
rect 34972 29650 35028 30940
rect 34972 29598 34974 29650
rect 35026 29598 35028 29650
rect 34972 29586 35028 29598
rect 34860 29474 34916 29484
rect 34860 28868 34916 28878
rect 34524 28812 34692 28868
rect 34748 28812 34860 28868
rect 34412 28644 34468 28654
rect 34636 28644 34692 28812
rect 34860 28802 34916 28812
rect 34860 28644 34916 28654
rect 34636 28642 34916 28644
rect 34636 28590 34862 28642
rect 34914 28590 34916 28642
rect 34636 28588 34916 28590
rect 34412 28550 34468 28588
rect 34860 28578 34916 28588
rect 35084 28084 35140 32844
rect 35532 32564 35588 32574
rect 35532 32470 35588 32508
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35532 31892 35588 31902
rect 35588 31836 35700 31892
rect 35532 31826 35588 31836
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35308 30100 35364 30110
rect 35308 30006 35364 30044
rect 35532 29652 35588 29662
rect 35532 29558 35588 29596
rect 35644 29428 35700 31836
rect 35756 30884 35812 33404
rect 35868 32674 35924 32686
rect 35868 32622 35870 32674
rect 35922 32622 35924 32674
rect 35868 31108 35924 32622
rect 35868 31042 35924 31052
rect 35756 30818 35812 30828
rect 35980 30548 36036 35534
rect 36092 33236 36148 35756
rect 36204 35476 36260 36206
rect 36204 35410 36260 35420
rect 36092 33170 36148 33180
rect 36316 31890 36372 38612
rect 36764 38052 36820 38062
rect 36428 37940 36484 37950
rect 36428 37846 36484 37884
rect 36764 37490 36820 37996
rect 36988 37938 37044 38612
rect 37436 38612 37492 38782
rect 36988 37886 36990 37938
rect 37042 37886 37044 37938
rect 36988 37874 37044 37886
rect 37212 38050 37268 38062
rect 37212 37998 37214 38050
rect 37266 37998 37268 38050
rect 37212 37940 37268 37998
rect 37212 37874 37268 37884
rect 36764 37438 36766 37490
rect 36818 37438 36820 37490
rect 36764 37426 36820 37438
rect 37212 37156 37268 37194
rect 37268 37100 37380 37156
rect 37212 37090 37268 37100
rect 37100 37042 37156 37054
rect 37100 36990 37102 37042
rect 37154 36990 37156 37042
rect 36988 36708 37044 36718
rect 36988 36594 37044 36652
rect 36988 36542 36990 36594
rect 37042 36542 37044 36594
rect 36988 36530 37044 36542
rect 36652 35588 36708 35598
rect 36652 35494 36708 35532
rect 36540 34916 36596 34926
rect 37100 34916 37156 36990
rect 37212 36932 37268 36942
rect 37212 36482 37268 36876
rect 37212 36430 37214 36482
rect 37266 36430 37268 36482
rect 37212 35588 37268 36430
rect 37212 35522 37268 35532
rect 37212 34916 37268 34926
rect 37100 34860 37212 34916
rect 36428 34692 36484 34702
rect 36540 34692 36596 34860
rect 37212 34822 37268 34860
rect 36428 34690 36596 34692
rect 36428 34638 36430 34690
rect 36482 34638 36596 34690
rect 36428 34636 36596 34638
rect 36428 34626 36484 34636
rect 36540 34020 36596 34636
rect 36316 31838 36318 31890
rect 36370 31838 36372 31890
rect 36316 31826 36372 31838
rect 36428 32452 36484 32462
rect 36428 31106 36484 32396
rect 36428 31054 36430 31106
rect 36482 31054 36484 31106
rect 36428 31042 36484 31054
rect 35868 30492 36036 30548
rect 36540 30996 36596 33964
rect 36652 30996 36708 31006
rect 36540 30994 36708 30996
rect 36540 30942 36654 30994
rect 36706 30942 36708 30994
rect 36540 30940 36708 30942
rect 35756 30324 35812 30334
rect 35868 30324 35924 30492
rect 35868 30268 36036 30324
rect 35756 30210 35812 30268
rect 35756 30158 35758 30210
rect 35810 30158 35812 30210
rect 35756 30146 35812 30158
rect 35532 29372 35700 29428
rect 35980 29428 36036 30268
rect 36204 30212 36260 30222
rect 36204 30118 36260 30156
rect 36428 30212 36484 30222
rect 36204 29764 36260 29774
rect 35980 29372 36148 29428
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35532 28868 35588 29372
rect 35868 29316 35924 29326
rect 34972 28028 35140 28084
rect 35308 28812 35588 28868
rect 35644 29314 35924 29316
rect 35644 29262 35870 29314
rect 35922 29262 35924 29314
rect 35644 29260 35924 29262
rect 35308 28530 35364 28812
rect 35420 28644 35476 28654
rect 35420 28550 35476 28588
rect 35308 28478 35310 28530
rect 35362 28478 35364 28530
rect 34412 27748 34468 27758
rect 34748 27748 34804 27758
rect 34076 22194 34132 22204
rect 34188 27746 34804 27748
rect 34188 27694 34414 27746
rect 34466 27694 34750 27746
rect 34802 27694 34804 27746
rect 34188 27692 34804 27694
rect 33964 21812 34020 21822
rect 34188 21812 34244 27692
rect 34412 27682 34468 27692
rect 34748 27682 34804 27692
rect 34860 27746 34916 27758
rect 34860 27694 34862 27746
rect 34914 27694 34916 27746
rect 34860 27300 34916 27694
rect 34300 27244 34916 27300
rect 34300 27186 34356 27244
rect 34300 27134 34302 27186
rect 34354 27134 34356 27186
rect 34300 27122 34356 27134
rect 34972 23548 35028 28028
rect 35084 27860 35140 27870
rect 35084 27766 35140 27804
rect 35308 27636 35364 28478
rect 35532 28530 35588 28542
rect 35532 28478 35534 28530
rect 35586 28478 35588 28530
rect 35532 28420 35588 28478
rect 35420 28364 35588 28420
rect 35420 27860 35476 28364
rect 35420 27794 35476 27804
rect 35532 27746 35588 27758
rect 35532 27694 35534 27746
rect 35586 27694 35588 27746
rect 35532 27636 35588 27694
rect 35308 27580 35588 27636
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 26852 35252 26862
rect 35196 26178 35252 26796
rect 35196 26126 35198 26178
rect 35250 26126 35252 26178
rect 35196 26114 35252 26126
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35532 24164 35588 27580
rect 35644 26852 35700 29260
rect 35868 29250 35924 29260
rect 35980 28644 36036 28654
rect 35980 28550 36036 28588
rect 35644 26786 35700 26796
rect 35532 24108 35924 24164
rect 34972 23492 35140 23548
rect 34300 23156 34356 23166
rect 34748 23156 34804 23166
rect 34356 23154 34804 23156
rect 34356 23102 34750 23154
rect 34802 23102 34804 23154
rect 34356 23100 34804 23102
rect 34300 23062 34356 23100
rect 33964 17220 34020 21756
rect 34076 21756 34244 21812
rect 34636 22482 34692 22494
rect 34636 22430 34638 22482
rect 34690 22430 34692 22482
rect 34076 20020 34132 21756
rect 34076 19954 34132 19964
rect 34188 21588 34244 21598
rect 34636 21588 34692 22430
rect 34748 22372 34804 23100
rect 35084 22596 35140 23492
rect 35420 23044 35476 23054
rect 35420 23042 35812 23044
rect 35420 22990 35422 23042
rect 35474 22990 35812 23042
rect 35420 22988 35812 22990
rect 35420 22978 35476 22988
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35084 22540 35252 22596
rect 35084 22372 35140 22382
rect 34748 22316 35084 22372
rect 35084 22278 35140 22316
rect 35196 21812 35252 22540
rect 35756 22258 35812 22988
rect 35756 22206 35758 22258
rect 35810 22206 35812 22258
rect 35756 22194 35812 22206
rect 35084 21700 35140 21710
rect 35196 21700 35252 21756
rect 35084 21698 35252 21700
rect 35084 21646 35086 21698
rect 35138 21646 35252 21698
rect 35084 21644 35252 21646
rect 35868 21700 35924 24108
rect 35084 21634 35140 21644
rect 35868 21634 35924 21644
rect 35980 22370 36036 22382
rect 35980 22318 35982 22370
rect 36034 22318 36036 22370
rect 34188 21586 34692 21588
rect 34188 21534 34190 21586
rect 34242 21534 34692 21586
rect 34188 21532 34692 21534
rect 33964 17108 34020 17164
rect 34076 17108 34132 17118
rect 33964 17106 34132 17108
rect 33964 17054 34078 17106
rect 34130 17054 34132 17106
rect 33964 17052 34132 17054
rect 33852 17042 33908 17052
rect 34076 17042 34132 17052
rect 33628 16942 33630 16994
rect 33682 16942 33684 16994
rect 33628 16930 33684 16942
rect 33740 16772 33796 16782
rect 33516 16212 33572 16222
rect 33516 16118 33572 16156
rect 33740 16098 33796 16716
rect 34076 16212 34132 16222
rect 33740 16046 33742 16098
rect 33794 16046 33796 16098
rect 33740 16034 33796 16046
rect 33964 16100 34020 16110
rect 33964 15986 34020 16044
rect 34076 16098 34132 16156
rect 34076 16046 34078 16098
rect 34130 16046 34132 16098
rect 34076 16034 34132 16046
rect 33964 15934 33966 15986
rect 34018 15934 34020 15986
rect 33964 15922 34020 15934
rect 34076 15540 34132 15550
rect 34076 15446 34132 15484
rect 33404 15426 33460 15438
rect 33404 15374 33406 15426
rect 33458 15374 33460 15426
rect 32508 15092 33012 15148
rect 33068 15138 33124 15148
rect 33180 15314 33236 15326
rect 33180 15262 33182 15314
rect 33234 15262 33236 15314
rect 33180 15148 33236 15262
rect 33404 15148 33460 15374
rect 33180 15092 33348 15148
rect 33404 15092 33684 15148
rect 32956 13860 33012 15092
rect 33292 14308 33348 15092
rect 33628 14642 33684 15092
rect 33628 14590 33630 14642
rect 33682 14590 33684 14642
rect 33628 14578 33684 14590
rect 33292 14252 33684 14308
rect 33628 13970 33684 14252
rect 33628 13918 33630 13970
rect 33682 13918 33684 13970
rect 33628 13906 33684 13918
rect 32956 13804 33236 13860
rect 33068 13636 33124 13646
rect 32284 13010 32340 13020
rect 32508 13634 33124 13636
rect 32508 13582 33070 13634
rect 33122 13582 33124 13634
rect 32508 13580 33124 13582
rect 32172 12964 32228 12974
rect 31724 12962 32228 12964
rect 31724 12910 31726 12962
rect 31778 12910 32174 12962
rect 32226 12910 32228 12962
rect 31724 12908 32228 12910
rect 31724 12898 31780 12908
rect 32172 12898 32228 12908
rect 31612 12852 31668 12862
rect 31612 12758 31668 12796
rect 32508 12852 32564 13580
rect 33068 13570 33124 13580
rect 32508 12066 32564 12796
rect 32508 12014 32510 12066
rect 32562 12014 32564 12066
rect 32508 12002 32564 12014
rect 33068 13076 33124 13086
rect 31164 10892 32004 10948
rect 31164 10834 31220 10892
rect 31164 10782 31166 10834
rect 31218 10782 31220 10834
rect 31164 10770 31220 10782
rect 31052 9998 31054 10050
rect 31106 9998 31108 10050
rect 31052 9986 31108 9998
rect 31164 10050 31220 10062
rect 31164 9998 31166 10050
rect 31218 9998 31220 10050
rect 31164 9828 31220 9998
rect 30548 9772 30660 9828
rect 30716 9772 31220 9828
rect 31388 9940 31444 9950
rect 30492 9734 30548 9772
rect 29820 9714 30100 9716
rect 29820 9662 29822 9714
rect 29874 9662 30100 9714
rect 29820 9660 30100 9662
rect 29820 9650 29876 9660
rect 29596 9604 29652 9614
rect 30044 9604 30100 9660
rect 29596 9602 29764 9604
rect 29596 9550 29598 9602
rect 29650 9550 29764 9602
rect 29596 9548 29764 9550
rect 29596 9538 29652 9548
rect 29372 9102 29374 9154
rect 29426 9102 29428 9154
rect 29372 9090 29428 9102
rect 29036 8878 29038 8930
rect 29090 8878 29092 8930
rect 29036 8866 29092 8878
rect 29148 9042 29204 9054
rect 29148 8990 29150 9042
rect 29202 8990 29204 9042
rect 29148 7364 29204 8990
rect 29596 8148 29652 8158
rect 29596 7474 29652 8092
rect 29596 7422 29598 7474
rect 29650 7422 29652 7474
rect 29596 7410 29652 7422
rect 29260 7364 29316 7374
rect 29148 7362 29316 7364
rect 29148 7310 29262 7362
rect 29314 7310 29316 7362
rect 29148 7308 29316 7310
rect 27916 6626 27972 6636
rect 28140 6636 28868 6692
rect 27692 6038 27748 6076
rect 28140 5460 28196 6636
rect 28140 5234 28196 5404
rect 28140 5182 28142 5234
rect 28194 5182 28196 5234
rect 28140 5170 28196 5182
rect 28812 6132 28868 6636
rect 28812 4338 28868 6076
rect 29036 4452 29092 4462
rect 29260 4452 29316 7308
rect 29036 4450 29316 4452
rect 29036 4398 29038 4450
rect 29090 4398 29316 4450
rect 29036 4396 29316 4398
rect 29596 6020 29652 6030
rect 29036 4386 29092 4396
rect 28812 4286 28814 4338
rect 28866 4286 28868 4338
rect 28812 4274 28868 4286
rect 27468 4162 27524 4172
rect 28140 4228 28196 4238
rect 28140 4134 28196 4172
rect 25900 3614 25902 3666
rect 25954 3614 25956 3666
rect 25900 3602 25956 3614
rect 28476 4114 28532 4126
rect 28476 4062 28478 4114
rect 28530 4062 28532 4114
rect 28476 3554 28532 4062
rect 29596 3668 29652 5964
rect 29708 4340 29764 9548
rect 30044 9538 30100 9548
rect 30156 9268 30212 9278
rect 30604 9268 30660 9772
rect 30156 9266 30660 9268
rect 30156 9214 30158 9266
rect 30210 9214 30606 9266
rect 30658 9214 30660 9266
rect 30156 9212 30660 9214
rect 30156 9202 30212 9212
rect 30604 9202 30660 9212
rect 30716 9602 30772 9614
rect 30716 9550 30718 9602
rect 30770 9550 30772 9602
rect 30380 7364 30436 7374
rect 30380 7362 30548 7364
rect 30380 7310 30382 7362
rect 30434 7310 30548 7362
rect 30380 7308 30548 7310
rect 30380 7298 30436 7308
rect 30492 6578 30548 7308
rect 30492 6526 30494 6578
rect 30546 6526 30548 6578
rect 30492 6514 30548 6526
rect 30380 6132 30436 6142
rect 30380 6038 30436 6076
rect 30716 6020 30772 9550
rect 30940 9604 30996 9614
rect 31276 9604 31332 9614
rect 30996 9602 31332 9604
rect 30996 9550 31278 9602
rect 31330 9550 31332 9602
rect 30996 9548 31332 9550
rect 30940 9266 30996 9548
rect 31276 9538 31332 9548
rect 30940 9214 30942 9266
rect 30994 9214 30996 9266
rect 30940 9202 30996 9214
rect 31388 9268 31444 9884
rect 31724 9828 31780 10892
rect 31948 10834 32004 10892
rect 31948 10782 31950 10834
rect 32002 10782 32004 10834
rect 31948 10770 32004 10782
rect 32508 9828 32564 9838
rect 31724 9734 31780 9772
rect 32396 9826 32564 9828
rect 32396 9774 32510 9826
rect 32562 9774 32564 9826
rect 32396 9772 32564 9774
rect 31500 9604 31556 9614
rect 31500 9602 31668 9604
rect 31500 9550 31502 9602
rect 31554 9550 31668 9602
rect 31500 9548 31668 9550
rect 31500 9538 31556 9548
rect 31500 9268 31556 9278
rect 31388 9266 31556 9268
rect 31388 9214 31502 9266
rect 31554 9214 31556 9266
rect 31388 9212 31556 9214
rect 31500 9044 31556 9212
rect 31500 8978 31556 8988
rect 31612 8932 31668 9548
rect 32284 9602 32340 9614
rect 32284 9550 32286 9602
rect 32338 9550 32340 9602
rect 32060 9044 32116 9054
rect 31836 8932 31892 8942
rect 31612 8930 31892 8932
rect 31612 8878 31838 8930
rect 31890 8878 31892 8930
rect 31612 8876 31892 8878
rect 31612 8258 31668 8270
rect 31612 8206 31614 8258
rect 31666 8206 31668 8258
rect 31164 8148 31220 8158
rect 31164 8054 31220 8092
rect 31612 8148 31668 8206
rect 31612 8082 31668 8092
rect 31836 7364 31892 8876
rect 32060 8260 32116 8988
rect 32284 8370 32340 9550
rect 32396 9266 32452 9772
rect 32508 9762 32564 9772
rect 32396 9214 32398 9266
rect 32450 9214 32452 9266
rect 32396 9202 32452 9214
rect 32284 8318 32286 8370
rect 32338 8318 32340 8370
rect 32284 8306 32340 8318
rect 32060 8194 32116 8204
rect 32732 8148 32788 8158
rect 32508 7364 32564 7374
rect 31836 7362 32564 7364
rect 31836 7310 32510 7362
rect 32562 7310 32564 7362
rect 31836 7308 32564 7310
rect 32508 7298 32564 7308
rect 30828 6580 30884 6590
rect 30828 6578 31332 6580
rect 30828 6526 30830 6578
rect 30882 6526 31332 6578
rect 30828 6524 31332 6526
rect 30828 6514 30884 6524
rect 30716 5926 30772 5964
rect 30940 6132 30996 6142
rect 30940 5906 30996 6076
rect 31276 6130 31332 6524
rect 31276 6078 31278 6130
rect 31330 6078 31332 6130
rect 31276 6066 31332 6078
rect 30940 5854 30942 5906
rect 30994 5854 30996 5906
rect 30940 5842 30996 5854
rect 32732 5236 32788 8092
rect 33068 5348 33124 13020
rect 33180 12404 33236 13804
rect 33292 13748 33348 13758
rect 33292 13654 33348 13692
rect 34076 13748 34132 13758
rect 34076 13654 34132 13692
rect 33404 13076 33460 13086
rect 33404 12982 33460 13020
rect 34076 13076 34132 13086
rect 34188 13076 34244 21532
rect 34412 21364 34468 21374
rect 34412 20914 34468 21308
rect 34412 20862 34414 20914
rect 34466 20862 34468 20914
rect 34412 20850 34468 20862
rect 35084 21364 35140 21374
rect 34860 20132 34916 20142
rect 34860 20018 34916 20076
rect 34860 19966 34862 20018
rect 34914 19966 34916 20018
rect 34860 19954 34916 19966
rect 35084 20018 35140 21308
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35868 21028 35924 21038
rect 35980 21028 36036 22318
rect 36092 21588 36148 29372
rect 36204 28866 36260 29708
rect 36428 29428 36484 30156
rect 36428 29362 36484 29372
rect 36540 29988 36596 30940
rect 36652 30930 36708 30940
rect 36764 30884 36820 30894
rect 36204 28814 36206 28866
rect 36258 28814 36260 28866
rect 36204 28802 36260 28814
rect 36316 28530 36372 28542
rect 36316 28478 36318 28530
rect 36370 28478 36372 28530
rect 36092 21522 36148 21532
rect 36204 27860 36260 27870
rect 36204 21476 36260 27804
rect 36316 27188 36372 28478
rect 36428 27746 36484 27758
rect 36428 27694 36430 27746
rect 36482 27694 36484 27746
rect 36428 27636 36484 27694
rect 36428 27570 36484 27580
rect 36428 27188 36484 27198
rect 36316 27186 36484 27188
rect 36316 27134 36430 27186
rect 36482 27134 36484 27186
rect 36316 27132 36484 27134
rect 36428 27122 36484 27132
rect 36540 26908 36596 29932
rect 36652 30100 36708 30110
rect 36652 29650 36708 30044
rect 36652 29598 36654 29650
rect 36706 29598 36708 29650
rect 36652 28980 36708 29598
rect 36652 28914 36708 28924
rect 36764 28084 36820 30828
rect 37212 30324 37268 30334
rect 37100 29988 37156 29998
rect 37100 29894 37156 29932
rect 37212 28980 37268 30268
rect 37100 28924 37268 28980
rect 37100 28868 37156 28924
rect 36988 28812 37156 28868
rect 36876 28644 36932 28654
rect 36876 28550 36932 28588
rect 36988 28642 37044 28812
rect 36988 28590 36990 28642
rect 37042 28590 37044 28642
rect 36988 28578 37044 28590
rect 37100 28644 37156 28654
rect 36876 28084 36932 28094
rect 36764 28028 36876 28084
rect 36876 27990 36932 28028
rect 36988 27188 37044 27198
rect 36988 27094 37044 27132
rect 37100 26908 37156 28588
rect 37212 28420 37268 28430
rect 37212 28326 37268 28364
rect 36540 26852 36820 26908
rect 36652 26180 36708 26190
rect 36764 26180 36820 26852
rect 36652 26178 36820 26180
rect 36652 26126 36654 26178
rect 36706 26126 36820 26178
rect 36652 26124 36820 26126
rect 36988 26852 37156 26908
rect 37212 27634 37268 27646
rect 37212 27582 37214 27634
rect 37266 27582 37268 27634
rect 37212 26908 37268 27582
rect 37324 27188 37380 37100
rect 37436 37042 37492 38556
rect 37436 36990 37438 37042
rect 37490 36990 37492 37042
rect 37436 36978 37492 36990
rect 37548 36484 37604 39564
rect 37772 39618 37828 40236
rect 37772 39566 37774 39618
rect 37826 39566 37828 39618
rect 37772 39554 37828 39566
rect 37884 37940 37940 46510
rect 37996 44436 38052 50372
rect 38332 49028 38388 51324
rect 39452 51380 39508 51548
rect 39900 51538 39956 51548
rect 39452 51286 39508 51324
rect 38332 48934 38388 48972
rect 38668 50484 38724 50494
rect 38220 48130 38276 48142
rect 38220 48078 38222 48130
rect 38274 48078 38276 48130
rect 38220 48020 38276 48078
rect 38556 48020 38612 48030
rect 38220 48018 38612 48020
rect 38220 47966 38222 48018
rect 38274 47966 38558 48018
rect 38610 47966 38612 48018
rect 38220 47964 38612 47966
rect 38108 46452 38164 46462
rect 38108 45106 38164 46396
rect 38220 46116 38276 47964
rect 38556 47954 38612 47964
rect 38556 47572 38612 47582
rect 38556 46674 38612 47516
rect 38556 46622 38558 46674
rect 38610 46622 38612 46674
rect 38556 46610 38612 46622
rect 38668 46116 38724 50428
rect 39004 48914 39060 48926
rect 39004 48862 39006 48914
rect 39058 48862 39060 48914
rect 38780 48354 38836 48366
rect 38780 48302 38782 48354
rect 38834 48302 38836 48354
rect 38780 46900 38836 48302
rect 38892 48132 38948 48142
rect 39004 48132 39060 48862
rect 38892 48130 39060 48132
rect 38892 48078 38894 48130
rect 38946 48078 39060 48130
rect 38892 48076 39060 48078
rect 39340 48130 39396 48142
rect 39340 48078 39342 48130
rect 39394 48078 39396 48130
rect 38892 48066 38948 48076
rect 39116 47236 39172 47246
rect 39004 47180 39116 47236
rect 38892 46900 38948 46910
rect 38780 46898 38948 46900
rect 38780 46846 38894 46898
rect 38946 46846 38948 46898
rect 38780 46844 38948 46846
rect 38780 46452 38836 46844
rect 38892 46834 38948 46844
rect 39004 46786 39060 47180
rect 39116 47170 39172 47180
rect 39004 46734 39006 46786
rect 39058 46734 39060 46786
rect 39004 46722 39060 46734
rect 39340 46788 39396 48078
rect 39900 47570 39956 47582
rect 39900 47518 39902 47570
rect 39954 47518 39956 47570
rect 39900 47236 39956 47518
rect 39900 47170 39956 47180
rect 40012 47012 40068 52332
rect 40236 52162 40292 52780
rect 40236 52110 40238 52162
rect 40290 52110 40292 52162
rect 40236 52098 40292 52110
rect 40348 51604 40404 53452
rect 40348 51510 40404 51548
rect 40124 49028 40180 49038
rect 40124 48466 40180 48972
rect 40124 48414 40126 48466
rect 40178 48414 40180 48466
rect 40124 47068 40180 48414
rect 40348 47572 40404 47582
rect 40348 47478 40404 47516
rect 40124 47012 40292 47068
rect 39788 46956 40068 47012
rect 39564 46788 39620 46798
rect 39340 46732 39564 46788
rect 38780 46386 38836 46396
rect 38668 46060 38948 46116
rect 38220 46050 38276 46060
rect 38332 46004 38388 46014
rect 38220 45668 38276 45678
rect 38332 45668 38388 45948
rect 38276 45612 38388 45668
rect 38668 45666 38724 45678
rect 38668 45614 38670 45666
rect 38722 45614 38724 45666
rect 38220 45574 38276 45612
rect 38668 45444 38724 45614
rect 38668 45378 38724 45388
rect 38108 45054 38110 45106
rect 38162 45054 38164 45106
rect 38108 45042 38164 45054
rect 38780 45106 38836 45118
rect 38780 45054 38782 45106
rect 38834 45054 38836 45106
rect 38556 44994 38612 45006
rect 38556 44942 38558 44994
rect 38610 44942 38612 44994
rect 37996 44370 38052 44380
rect 38444 44436 38500 44446
rect 38332 44322 38388 44334
rect 38332 44270 38334 44322
rect 38386 44270 38388 44322
rect 38332 43876 38388 44270
rect 38332 43810 38388 43820
rect 38220 43652 38276 43662
rect 38220 43558 38276 43596
rect 38220 42532 38276 42542
rect 38220 42438 38276 42476
rect 38444 41972 38500 44380
rect 38556 43708 38612 44942
rect 38780 44546 38836 45054
rect 38780 44494 38782 44546
rect 38834 44494 38836 44546
rect 38780 44482 38836 44494
rect 38556 43652 38724 43708
rect 38668 42642 38724 43652
rect 38668 42590 38670 42642
rect 38722 42590 38724 42642
rect 38668 42578 38724 42590
rect 38780 42084 38836 42094
rect 38668 41972 38724 41982
rect 38444 41970 38724 41972
rect 38444 41918 38670 41970
rect 38722 41918 38724 41970
rect 38444 41916 38724 41918
rect 38668 41906 38724 41916
rect 38780 41860 38836 42028
rect 38892 41972 38948 46060
rect 39452 45890 39508 45902
rect 39452 45838 39454 45890
rect 39506 45838 39508 45890
rect 39452 45780 39508 45838
rect 39452 45714 39508 45724
rect 39116 44994 39172 45006
rect 39116 44942 39118 44994
rect 39170 44942 39172 44994
rect 39004 44548 39060 44558
rect 39004 44322 39060 44492
rect 39004 44270 39006 44322
rect 39058 44270 39060 44322
rect 39004 44258 39060 44270
rect 39116 43876 39172 44942
rect 39340 44996 39396 45006
rect 39340 44902 39396 44940
rect 39452 44212 39508 44222
rect 39452 44118 39508 44156
rect 39116 43810 39172 43820
rect 39116 41972 39172 41982
rect 38892 41970 39172 41972
rect 38892 41918 39118 41970
rect 39170 41918 39172 41970
rect 38892 41916 39172 41918
rect 39116 41906 39172 41916
rect 38780 41804 39060 41860
rect 38332 41188 38388 41198
rect 38332 41094 38388 41132
rect 38556 40852 38612 40862
rect 38332 40516 38388 40526
rect 38332 40402 38388 40460
rect 38332 40350 38334 40402
rect 38386 40350 38388 40402
rect 38332 40338 38388 40350
rect 38556 40402 38612 40796
rect 38892 40628 38948 40638
rect 38556 40350 38558 40402
rect 38610 40350 38612 40402
rect 38332 39844 38388 39854
rect 38332 39750 38388 39788
rect 38444 39172 38500 39182
rect 38444 39058 38500 39116
rect 38444 39006 38446 39058
rect 38498 39006 38500 39058
rect 38444 38836 38500 39006
rect 38444 38770 38500 38780
rect 38108 38722 38164 38734
rect 38108 38670 38110 38722
rect 38162 38670 38164 38722
rect 38108 38612 38164 38670
rect 38108 38546 38164 38556
rect 37996 38164 38052 38174
rect 37996 38070 38052 38108
rect 37772 37884 37940 37940
rect 37660 37268 37716 37278
rect 37660 37174 37716 37212
rect 37436 36428 37604 36484
rect 37436 31332 37492 36428
rect 37548 36258 37604 36270
rect 37548 36206 37550 36258
rect 37602 36206 37604 36258
rect 37548 35810 37604 36206
rect 37772 36260 37828 37884
rect 38108 37156 38164 37166
rect 38108 37042 38164 37100
rect 38108 36990 38110 37042
rect 38162 36990 38164 37042
rect 38108 36978 38164 36990
rect 38556 36820 38612 40350
rect 38108 36764 38612 36820
rect 38780 40572 38892 40628
rect 38108 36706 38164 36764
rect 38108 36654 38110 36706
rect 38162 36654 38164 36706
rect 38108 36642 38164 36654
rect 37996 36596 38052 36634
rect 37996 36530 38052 36540
rect 38332 36484 38388 36494
rect 37996 36372 38052 36382
rect 37772 36194 37828 36204
rect 37884 36316 37996 36372
rect 37884 36036 37940 36316
rect 37996 36306 38052 36316
rect 38108 36260 38164 36270
rect 37884 35980 38052 36036
rect 37548 35758 37550 35810
rect 37602 35758 37604 35810
rect 37548 35746 37604 35758
rect 37884 35810 37940 35822
rect 37884 35758 37886 35810
rect 37938 35758 37940 35810
rect 37884 35026 37940 35758
rect 37884 34974 37886 35026
rect 37938 34974 37940 35026
rect 37884 34962 37940 34974
rect 37996 34804 38052 35980
rect 37548 34748 38052 34804
rect 37548 34018 37604 34748
rect 37548 33966 37550 34018
rect 37602 33966 37604 34018
rect 37548 33954 37604 33966
rect 38108 31780 38164 36204
rect 38108 31714 38164 31724
rect 37660 31668 37716 31678
rect 37660 31574 37716 31612
rect 38108 31554 38164 31566
rect 38108 31502 38110 31554
rect 38162 31502 38164 31554
rect 38108 31444 38164 31502
rect 38108 31378 38164 31388
rect 38220 31556 38276 31566
rect 37436 31276 37716 31332
rect 37436 31108 37492 31118
rect 37436 31014 37492 31052
rect 37548 28642 37604 28654
rect 37548 28590 37550 28642
rect 37602 28590 37604 28642
rect 37548 28532 37604 28590
rect 37548 28466 37604 28476
rect 37436 28418 37492 28430
rect 37436 28366 37438 28418
rect 37490 28366 37492 28418
rect 37436 27636 37492 28366
rect 37548 28084 37604 28094
rect 37548 27858 37604 28028
rect 37548 27806 37550 27858
rect 37602 27806 37604 27858
rect 37548 27794 37604 27806
rect 37436 27570 37492 27580
rect 37660 27412 37716 31276
rect 38220 30324 38276 31500
rect 38108 29988 38164 29998
rect 38108 29650 38164 29932
rect 38108 29598 38110 29650
rect 38162 29598 38164 29650
rect 38108 29586 38164 29598
rect 38108 28756 38164 28766
rect 38220 28756 38276 30268
rect 38108 28754 38276 28756
rect 38108 28702 38110 28754
rect 38162 28702 38276 28754
rect 38108 28700 38276 28702
rect 38108 28690 38164 28700
rect 37772 28420 37828 28430
rect 37772 27858 37828 28364
rect 37772 27806 37774 27858
rect 37826 27806 37828 27858
rect 37772 27794 37828 27806
rect 37660 27346 37716 27356
rect 37324 27132 38052 27188
rect 37212 26852 37380 26908
rect 36652 25284 36708 26124
rect 36652 25218 36708 25228
rect 36428 24948 36484 24958
rect 36428 24722 36484 24892
rect 36428 24670 36430 24722
rect 36482 24670 36484 24722
rect 36428 24658 36484 24670
rect 36652 24834 36708 24846
rect 36652 24782 36654 24834
rect 36706 24782 36708 24834
rect 36652 22484 36708 24782
rect 36988 24162 37044 26852
rect 37324 26402 37380 26852
rect 37772 26740 37828 26750
rect 37660 26516 37716 26526
rect 37660 26422 37716 26460
rect 37324 26350 37326 26402
rect 37378 26350 37380 26402
rect 37324 26338 37380 26350
rect 37212 24948 37268 24958
rect 37212 24854 37268 24892
rect 36988 24110 36990 24162
rect 37042 24110 37044 24162
rect 36988 24098 37044 24110
rect 37100 23828 37156 23838
rect 37100 23826 37604 23828
rect 37100 23774 37102 23826
rect 37154 23774 37604 23826
rect 37100 23772 37604 23774
rect 37100 23762 37156 23772
rect 37548 23042 37604 23772
rect 37548 22990 37550 23042
rect 37602 22990 37604 23042
rect 37548 22978 37604 22990
rect 37772 22708 37828 26684
rect 36652 22418 36708 22428
rect 37660 22652 37828 22708
rect 37100 22372 37156 22382
rect 36204 21410 36260 21420
rect 36540 21586 36596 21598
rect 36540 21534 36542 21586
rect 36594 21534 36596 21586
rect 35868 21026 36036 21028
rect 35868 20974 35870 21026
rect 35922 20974 36036 21026
rect 35868 20972 36036 20974
rect 36540 21028 36596 21534
rect 36876 21586 36932 21598
rect 36876 21534 36878 21586
rect 36930 21534 36932 21586
rect 36876 21364 36932 21534
rect 36876 21298 36932 21308
rect 35868 20962 35924 20972
rect 36540 20962 36596 20972
rect 37100 20916 37156 22316
rect 37212 20916 37268 20926
rect 37100 20914 37268 20916
rect 37100 20862 37214 20914
rect 37266 20862 37268 20914
rect 37100 20860 37268 20862
rect 37212 20850 37268 20860
rect 36204 20802 36260 20814
rect 36204 20750 36206 20802
rect 36258 20750 36260 20802
rect 35532 20132 35588 20142
rect 35532 20038 35588 20076
rect 36204 20132 36260 20750
rect 36204 20066 36260 20076
rect 36428 20802 36484 20814
rect 36428 20750 36430 20802
rect 36482 20750 36484 20802
rect 35084 19966 35086 20018
rect 35138 19966 35140 20018
rect 35084 19954 35140 19966
rect 35196 20020 35252 20030
rect 34524 19796 34580 19806
rect 35196 19796 35252 19964
rect 34524 19794 34804 19796
rect 34524 19742 34526 19794
rect 34578 19742 34804 19794
rect 34524 19740 34804 19742
rect 34524 19730 34580 19740
rect 34748 19460 34804 19740
rect 35084 19740 35252 19796
rect 34748 19404 35028 19460
rect 34972 19234 35028 19404
rect 34972 19182 34974 19234
rect 35026 19182 35028 19234
rect 34972 19170 35028 19182
rect 34748 19012 34804 19022
rect 34300 19010 34804 19012
rect 34300 18958 34750 19010
rect 34802 18958 34804 19010
rect 34300 18956 34804 18958
rect 34300 17778 34356 18956
rect 34748 18946 34804 18956
rect 34300 17726 34302 17778
rect 34354 17726 34356 17778
rect 34300 17714 34356 17726
rect 34412 16996 34468 17006
rect 34300 15204 34356 15214
rect 34300 14532 34356 15148
rect 34412 15148 34468 16940
rect 34972 16772 35028 16782
rect 34524 16324 34580 16334
rect 34524 15538 34580 16268
rect 34972 16100 35028 16716
rect 34524 15486 34526 15538
rect 34578 15486 34580 15538
rect 34524 15474 34580 15486
rect 34748 16098 35028 16100
rect 34748 16046 34974 16098
rect 35026 16046 35028 16098
rect 34748 16044 35028 16046
rect 34748 15540 34804 16044
rect 34972 16034 35028 16044
rect 35084 15876 35140 19740
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 36428 18564 36484 20750
rect 37548 20578 37604 20590
rect 37548 20526 37550 20578
rect 37602 20526 37604 20578
rect 37548 20132 37604 20526
rect 37660 20580 37716 22652
rect 37772 22484 37828 22494
rect 37772 22390 37828 22428
rect 37996 21028 38052 27132
rect 38332 26908 38388 36428
rect 38668 31778 38724 31790
rect 38668 31726 38670 31778
rect 38722 31726 38724 31778
rect 38668 31220 38724 31726
rect 38668 31154 38724 31164
rect 38444 28754 38500 28766
rect 38444 28702 38446 28754
rect 38498 28702 38500 28754
rect 38444 28420 38500 28702
rect 38444 28354 38500 28364
rect 38108 26852 38388 26908
rect 38108 21810 38164 26852
rect 38780 24948 38836 40572
rect 38892 40562 38948 40572
rect 38892 39732 38948 39742
rect 38892 39058 38948 39676
rect 38892 39006 38894 39058
rect 38946 39006 38948 39058
rect 38892 38836 38948 39006
rect 38892 38770 38948 38780
rect 39004 39508 39060 41804
rect 39340 41746 39396 41758
rect 39340 41694 39342 41746
rect 39394 41694 39396 41746
rect 39340 39732 39396 41694
rect 39452 40404 39508 40414
rect 39452 40290 39508 40348
rect 39452 40238 39454 40290
rect 39506 40238 39508 40290
rect 39452 40226 39508 40238
rect 39340 39666 39396 39676
rect 39116 39508 39172 39518
rect 39004 39506 39172 39508
rect 39004 39454 39118 39506
rect 39170 39454 39172 39506
rect 39004 39452 39172 39454
rect 38892 33124 38948 33134
rect 38892 33030 38948 33068
rect 38892 32562 38948 32574
rect 38892 32510 38894 32562
rect 38946 32510 38948 32562
rect 38892 32002 38948 32510
rect 38892 31950 38894 32002
rect 38946 31950 38948 32002
rect 38892 31938 38948 31950
rect 38892 31668 38948 31678
rect 38892 31574 38948 31612
rect 38892 29314 38948 29326
rect 38892 29262 38894 29314
rect 38946 29262 38948 29314
rect 38892 29204 38948 29262
rect 38892 29138 38948 29148
rect 38780 24882 38836 24892
rect 38556 24052 38612 24062
rect 38556 23958 38612 23996
rect 38220 23714 38276 23726
rect 38220 23662 38222 23714
rect 38274 23662 38276 23714
rect 38220 23492 38276 23662
rect 38220 22372 38276 23436
rect 38220 22306 38276 22316
rect 38108 21758 38110 21810
rect 38162 21758 38164 21810
rect 38108 21746 38164 21758
rect 38892 21700 38948 21710
rect 38332 21586 38388 21598
rect 38332 21534 38334 21586
rect 38386 21534 38388 21586
rect 38332 21476 38388 21534
rect 38332 21410 38388 21420
rect 38780 21476 38836 21486
rect 38780 21382 38836 21420
rect 37660 20514 37716 20524
rect 37772 20972 38052 21028
rect 37324 20076 37548 20132
rect 37324 18564 37380 20076
rect 37548 20066 37604 20076
rect 36428 18508 37044 18564
rect 36652 18340 36708 18350
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 36428 17778 36484 17790
rect 36428 17726 36430 17778
rect 36482 17726 36484 17778
rect 35644 17220 35700 17230
rect 35196 17108 35252 17118
rect 35196 17014 35252 17052
rect 35644 17106 35700 17164
rect 36204 17220 36260 17230
rect 35644 17054 35646 17106
rect 35698 17054 35700 17106
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35196 16100 35252 16110
rect 35196 16006 35252 16044
rect 34748 15474 34804 15484
rect 34860 15820 35140 15876
rect 34412 15092 34580 15148
rect 34412 14532 34468 14542
rect 34300 14476 34412 14532
rect 34412 14438 34468 14476
rect 34300 13076 34356 13086
rect 34188 13074 34356 13076
rect 34188 13022 34302 13074
rect 34354 13022 34356 13074
rect 34188 13020 34356 13022
rect 34076 12982 34132 13020
rect 34300 13010 34356 13020
rect 33740 12740 33796 12750
rect 33740 12738 34020 12740
rect 33740 12686 33742 12738
rect 33794 12686 34020 12738
rect 33740 12684 34020 12686
rect 33740 12674 33796 12684
rect 33180 12348 33348 12404
rect 33180 12180 33236 12190
rect 33180 12086 33236 12124
rect 33292 10050 33348 12348
rect 33404 12180 33460 12190
rect 33404 11508 33460 12124
rect 33740 12180 33796 12190
rect 33740 12086 33796 12124
rect 33404 11506 33572 11508
rect 33404 11454 33406 11506
rect 33458 11454 33572 11506
rect 33404 11452 33572 11454
rect 33404 11442 33460 11452
rect 33292 9998 33294 10050
rect 33346 9998 33348 10050
rect 33292 9986 33348 9998
rect 33516 10052 33572 11452
rect 33964 11394 34020 12684
rect 34524 12292 34580 15092
rect 33964 11342 33966 11394
rect 34018 11342 34020 11394
rect 33964 11330 34020 11342
rect 34076 12236 34580 12292
rect 33516 9996 33908 10052
rect 33404 9716 33460 9726
rect 33404 9714 33572 9716
rect 33404 9662 33406 9714
rect 33458 9662 33572 9714
rect 33404 9660 33572 9662
rect 33404 9650 33460 9660
rect 33404 9044 33460 9054
rect 33404 8148 33460 8988
rect 33516 8372 33572 9660
rect 33628 9044 33684 9996
rect 33852 9938 33908 9996
rect 33852 9886 33854 9938
rect 33906 9886 33908 9938
rect 33852 9874 33908 9886
rect 33628 8978 33684 8988
rect 33516 8306 33572 8316
rect 33180 8092 33404 8148
rect 33180 7698 33236 8092
rect 33404 8082 33460 8092
rect 33180 7646 33182 7698
rect 33234 7646 33236 7698
rect 33180 7634 33236 7646
rect 34076 7588 34132 12236
rect 34524 12066 34580 12078
rect 34524 12014 34526 12066
rect 34578 12014 34580 12066
rect 34524 11508 34580 12014
rect 34860 12068 34916 15820
rect 35644 15540 35700 17054
rect 35196 15484 35700 15540
rect 35196 15148 35252 15484
rect 35644 15426 35700 15484
rect 35644 15374 35646 15426
rect 35698 15374 35700 15426
rect 35644 15362 35700 15374
rect 35756 17108 35812 17118
rect 35308 15316 35364 15326
rect 35308 15222 35364 15260
rect 34972 15092 35252 15148
rect 34972 14644 35028 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35756 14868 35812 17052
rect 36204 16994 36260 17164
rect 36204 16942 36206 16994
rect 36258 16942 36260 16994
rect 36204 16930 36260 16942
rect 36204 16324 36260 16334
rect 36204 16210 36260 16268
rect 36204 16158 36206 16210
rect 36258 16158 36260 16210
rect 36204 16146 36260 16158
rect 35756 14802 35812 14812
rect 35868 16098 35924 16110
rect 35868 16046 35870 16098
rect 35922 16046 35924 16098
rect 34972 14550 35028 14588
rect 35420 14756 35476 14766
rect 35420 14642 35476 14700
rect 35420 14590 35422 14642
rect 35474 14590 35476 14642
rect 35420 14578 35476 14590
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35644 13188 35700 13198
rect 35644 13074 35700 13132
rect 35644 13022 35646 13074
rect 35698 13022 35700 13074
rect 35644 13010 35700 13022
rect 35868 13076 35924 16046
rect 35980 15988 36036 15998
rect 35980 15894 36036 15932
rect 36428 15876 36484 17726
rect 36652 17780 36708 18284
rect 36988 18338 37044 18508
rect 36988 18286 36990 18338
rect 37042 18286 37044 18338
rect 36988 18116 37044 18286
rect 36988 18060 37268 18116
rect 36652 17714 36708 17724
rect 36764 17220 36820 17230
rect 36820 17164 36932 17220
rect 36764 17154 36820 17164
rect 36540 16884 36596 16894
rect 36540 16790 36596 16828
rect 35980 15764 36036 15774
rect 35980 13186 36036 15708
rect 36428 15148 36484 15820
rect 36652 15988 36708 15998
rect 36876 15988 36932 17164
rect 37100 16098 37156 16110
rect 37100 16046 37102 16098
rect 37154 16046 37156 16098
rect 36988 15988 37044 15998
rect 36876 15986 37044 15988
rect 36876 15934 36990 15986
rect 37042 15934 37044 15986
rect 36876 15932 37044 15934
rect 36652 15314 36708 15932
rect 36988 15922 37044 15932
rect 36652 15262 36654 15314
rect 36706 15262 36708 15314
rect 36652 15250 36708 15262
rect 37100 15148 37156 16046
rect 37212 15316 37268 18060
rect 37324 17778 37380 18508
rect 37324 17726 37326 17778
rect 37378 17726 37380 17778
rect 37324 17714 37380 17726
rect 37660 17666 37716 17678
rect 37660 17614 37662 17666
rect 37714 17614 37716 17666
rect 37660 16996 37716 17614
rect 37660 16930 37716 16940
rect 37548 15540 37604 15550
rect 37772 15540 37828 20972
rect 38220 20916 38276 20926
rect 38220 20356 38276 20860
rect 38892 20804 38948 21644
rect 37996 20300 38220 20356
rect 37548 15538 37828 15540
rect 37548 15486 37550 15538
rect 37602 15486 37828 15538
rect 37548 15484 37828 15486
rect 37884 18564 37940 18574
rect 37884 17890 37940 18508
rect 37884 17838 37886 17890
rect 37938 17838 37940 17890
rect 37548 15474 37604 15484
rect 37660 15316 37716 15326
rect 37212 15314 37716 15316
rect 37212 15262 37662 15314
rect 37714 15262 37716 15314
rect 37212 15260 37716 15262
rect 37660 15250 37716 15260
rect 36428 15092 36932 15148
rect 36540 14644 36596 14654
rect 36540 14550 36596 14588
rect 36876 13746 36932 15092
rect 36876 13694 36878 13746
rect 36930 13694 36932 13746
rect 36876 13682 36932 13694
rect 36988 15092 37156 15148
rect 35980 13134 35982 13186
rect 36034 13134 36036 13186
rect 35980 13122 36036 13134
rect 36764 13188 36820 13198
rect 36988 13188 37044 15092
rect 37212 14868 37268 14878
rect 37212 14642 37268 14812
rect 37212 14590 37214 14642
rect 37266 14590 37268 14642
rect 37212 14578 37268 14590
rect 37884 13972 37940 17838
rect 37100 13970 37940 13972
rect 37100 13918 37886 13970
rect 37938 13918 37940 13970
rect 37100 13916 37940 13918
rect 37100 13746 37156 13916
rect 37884 13906 37940 13916
rect 37996 16772 38052 20300
rect 38220 20290 38276 20300
rect 38444 20802 38948 20804
rect 38444 20750 38894 20802
rect 38946 20750 38948 20802
rect 38444 20748 38948 20750
rect 38444 19906 38500 20748
rect 38892 20738 38948 20748
rect 39004 20188 39060 39452
rect 39116 39442 39172 39452
rect 39452 39396 39508 39406
rect 39452 39302 39508 39340
rect 39340 38948 39396 38958
rect 39340 38854 39396 38892
rect 39228 38836 39284 38846
rect 39116 34356 39172 34366
rect 39228 34356 39284 38780
rect 39452 34356 39508 34366
rect 39116 34354 39452 34356
rect 39116 34302 39118 34354
rect 39170 34302 39452 34354
rect 39116 34300 39452 34302
rect 39116 27860 39172 34300
rect 39452 34242 39508 34300
rect 39452 34190 39454 34242
rect 39506 34190 39508 34242
rect 39452 34178 39508 34190
rect 39228 33346 39284 33358
rect 39228 33294 39230 33346
rect 39282 33294 39284 33346
rect 39228 33124 39284 33294
rect 39228 33058 39284 33068
rect 39340 32452 39396 32462
rect 39340 32358 39396 32396
rect 39564 31948 39620 46732
rect 39676 46674 39732 46686
rect 39676 46622 39678 46674
rect 39730 46622 39732 46674
rect 39676 45330 39732 46622
rect 39676 45278 39678 45330
rect 39730 45278 39732 45330
rect 39676 45266 39732 45278
rect 39788 42754 39844 46956
rect 39900 46788 39956 46798
rect 39900 46786 40180 46788
rect 39900 46734 39902 46786
rect 39954 46734 40180 46786
rect 39900 46732 40180 46734
rect 39900 46722 39956 46732
rect 40124 46002 40180 46732
rect 40236 46564 40292 47012
rect 40348 46564 40404 46574
rect 40236 46562 40404 46564
rect 40236 46510 40350 46562
rect 40402 46510 40404 46562
rect 40236 46508 40404 46510
rect 40124 45950 40126 46002
rect 40178 45950 40180 46002
rect 40124 45938 40180 45950
rect 40348 45780 40404 46508
rect 40348 45714 40404 45724
rect 40012 44996 40068 45006
rect 40124 44996 40180 45006
rect 40068 44994 40180 44996
rect 40068 44942 40126 44994
rect 40178 44942 40180 44994
rect 40068 44940 40180 44942
rect 39900 44436 39956 44446
rect 39900 44342 39956 44380
rect 39788 42702 39790 42754
rect 39842 42702 39844 42754
rect 39788 42690 39844 42702
rect 40012 41860 40068 44940
rect 40124 44930 40180 44940
rect 40348 44548 40404 44558
rect 40684 44548 40740 56028
rect 41020 55524 41076 56252
rect 41020 54738 41076 55468
rect 41020 54686 41022 54738
rect 41074 54686 41076 54738
rect 41020 54516 41076 54686
rect 41020 54450 41076 54460
rect 40908 53954 40964 53966
rect 40908 53902 40910 53954
rect 40962 53902 40964 53954
rect 40908 52388 40964 53902
rect 41132 53842 41188 58268
rect 41356 56978 41412 56990
rect 41356 56926 41358 56978
rect 41410 56926 41412 56978
rect 41244 55970 41300 55982
rect 41244 55918 41246 55970
rect 41298 55918 41300 55970
rect 41244 55858 41300 55918
rect 41244 55806 41246 55858
rect 41298 55806 41300 55858
rect 41244 55794 41300 55806
rect 41244 55412 41300 55422
rect 41244 55318 41300 55356
rect 41356 54740 41412 56926
rect 41356 54674 41412 54684
rect 41356 54516 41412 54526
rect 41356 54422 41412 54460
rect 41468 53844 41524 59724
rect 42252 59780 42308 59790
rect 42252 59686 42308 59724
rect 42700 59778 42756 59790
rect 42700 59726 42702 59778
rect 42754 59726 42756 59778
rect 41916 57204 41972 57214
rect 41916 56308 41972 57148
rect 42700 57204 42756 59726
rect 42700 57138 42756 57148
rect 44156 56866 44212 56878
rect 44156 56814 44158 56866
rect 44210 56814 44212 56866
rect 43484 56756 43540 56766
rect 41692 56306 41972 56308
rect 41692 56254 41918 56306
rect 41970 56254 41972 56306
rect 41692 56252 41972 56254
rect 41580 55858 41636 55870
rect 41580 55806 41582 55858
rect 41634 55806 41636 55858
rect 41580 55186 41636 55806
rect 41580 55134 41582 55186
rect 41634 55134 41636 55186
rect 41580 54404 41636 55134
rect 41580 54338 41636 54348
rect 41692 53956 41748 56252
rect 41916 56242 41972 56252
rect 42140 56754 43540 56756
rect 42140 56702 43486 56754
rect 43538 56702 43540 56754
rect 42140 56700 43540 56702
rect 42140 56306 42196 56700
rect 43484 56690 43540 56700
rect 42140 56254 42142 56306
rect 42194 56254 42196 56306
rect 42140 56242 42196 56254
rect 41804 56084 41860 56094
rect 41804 55990 41860 56028
rect 42476 56084 42532 56094
rect 42476 55990 42532 56028
rect 41916 55412 41972 55422
rect 42364 55412 42420 55422
rect 41916 55410 42196 55412
rect 41916 55358 41918 55410
rect 41970 55358 42196 55410
rect 41916 55356 42196 55358
rect 41916 55346 41972 55356
rect 41804 55186 41860 55198
rect 41804 55134 41806 55186
rect 41858 55134 41860 55186
rect 41804 55076 41860 55134
rect 41916 55076 41972 55086
rect 41804 55020 41916 55076
rect 41916 55010 41972 55020
rect 42140 54626 42196 55356
rect 42364 55318 42420 55356
rect 42812 55412 42868 55422
rect 42812 55318 42868 55356
rect 44156 55412 44212 56814
rect 44156 55346 44212 55356
rect 42140 54574 42142 54626
rect 42194 54574 42196 54626
rect 42140 54562 42196 54574
rect 42252 55076 42308 55086
rect 41692 53900 41860 53956
rect 41132 53790 41134 53842
rect 41186 53790 41188 53842
rect 41132 53778 41188 53790
rect 41244 53788 41524 53844
rect 41020 53730 41076 53742
rect 41020 53678 41022 53730
rect 41074 53678 41076 53730
rect 41020 53060 41076 53678
rect 41020 53004 41188 53060
rect 41020 52836 41076 52846
rect 41020 52742 41076 52780
rect 40796 52332 40964 52388
rect 40796 46676 40852 52332
rect 41132 52276 41188 53004
rect 41132 52162 41188 52220
rect 41132 52110 41134 52162
rect 41186 52110 41188 52162
rect 41132 52098 41188 52110
rect 41132 51380 41188 51390
rect 41244 51380 41300 53788
rect 41692 53730 41748 53742
rect 41692 53678 41694 53730
rect 41746 53678 41748 53730
rect 41468 52836 41524 52846
rect 41692 52836 41748 53678
rect 41468 52834 41748 52836
rect 41468 52782 41470 52834
rect 41522 52782 41748 52834
rect 41468 52780 41748 52782
rect 41132 51378 41300 51380
rect 41132 51326 41134 51378
rect 41186 51326 41300 51378
rect 41132 51324 41300 51326
rect 41356 52276 41412 52286
rect 41356 51378 41412 52220
rect 41468 51940 41524 52780
rect 41804 52276 41860 53900
rect 41692 52220 41860 52276
rect 42140 53842 42196 53854
rect 42140 53790 42142 53842
rect 42194 53790 42196 53842
rect 42140 53508 42196 53790
rect 42252 53730 42308 55020
rect 42252 53678 42254 53730
rect 42306 53678 42308 53730
rect 42252 53666 42308 53678
rect 42364 54516 42420 54526
rect 42140 52836 42196 53452
rect 42364 53172 42420 54460
rect 42812 54404 42868 54414
rect 44268 54404 44324 54414
rect 42812 53844 42868 54348
rect 44044 54402 44324 54404
rect 44044 54350 44270 54402
rect 44322 54350 44324 54402
rect 44044 54348 44324 54350
rect 42420 53116 42644 53172
rect 42364 53078 42420 53116
rect 42140 52274 42196 52780
rect 42476 52388 42532 52398
rect 42476 52294 42532 52332
rect 42140 52222 42142 52274
rect 42194 52222 42196 52274
rect 41692 52162 41748 52220
rect 41692 52110 41694 52162
rect 41746 52110 41748 52162
rect 41692 52098 41748 52110
rect 42028 52162 42084 52174
rect 42028 52110 42030 52162
rect 42082 52110 42084 52162
rect 42028 51940 42084 52110
rect 41468 51884 42084 51940
rect 41468 51604 41524 51884
rect 41468 51538 41524 51548
rect 41356 51326 41358 51378
rect 41410 51326 41412 51378
rect 41132 51314 41188 51324
rect 41356 51314 41412 51326
rect 42028 51380 42084 51884
rect 42028 51314 42084 51324
rect 42140 51604 42196 52222
rect 42364 52164 42420 52174
rect 42364 52070 42420 52108
rect 42140 51378 42196 51548
rect 42140 51326 42142 51378
rect 42194 51326 42196 51378
rect 41356 51156 41412 51166
rect 42140 51156 42196 51326
rect 42252 51380 42308 51390
rect 42252 51286 42308 51324
rect 41356 50484 41412 51100
rect 41356 50390 41412 50428
rect 41804 51100 42196 51156
rect 41692 49810 41748 49822
rect 41692 49758 41694 49810
rect 41746 49758 41748 49810
rect 41132 49700 41188 49710
rect 41020 49698 41188 49700
rect 41020 49646 41134 49698
rect 41186 49646 41188 49698
rect 41020 49644 41188 49646
rect 41020 48916 41076 49644
rect 41132 49634 41188 49644
rect 41132 49140 41188 49150
rect 41580 49140 41636 49150
rect 41132 49138 41636 49140
rect 41132 49086 41134 49138
rect 41186 49086 41582 49138
rect 41634 49086 41636 49138
rect 41132 49084 41636 49086
rect 41132 49074 41188 49084
rect 41580 49074 41636 49084
rect 41020 48860 41412 48916
rect 41020 48692 41076 48702
rect 41020 48242 41076 48636
rect 41020 48190 41022 48242
rect 41074 48190 41076 48242
rect 41020 48178 41076 48190
rect 41244 48356 41300 48366
rect 40908 48018 40964 48030
rect 40908 47966 40910 48018
rect 40962 47966 40964 48018
rect 40908 47458 40964 47966
rect 40908 47406 40910 47458
rect 40962 47406 40964 47458
rect 40908 47394 40964 47406
rect 41132 47570 41188 47582
rect 41132 47518 41134 47570
rect 41186 47518 41188 47570
rect 41132 46786 41188 47518
rect 41244 47124 41300 48300
rect 41356 47572 41412 48860
rect 41692 48802 41748 49758
rect 41692 48750 41694 48802
rect 41746 48750 41748 48802
rect 41580 48244 41636 48254
rect 41580 48150 41636 48188
rect 41468 47572 41524 47582
rect 41356 47570 41524 47572
rect 41356 47518 41470 47570
rect 41522 47518 41524 47570
rect 41356 47516 41524 47518
rect 41356 47124 41412 47134
rect 41244 47068 41356 47124
rect 41356 47058 41412 47068
rect 41244 46900 41300 46910
rect 41244 46806 41300 46844
rect 41132 46734 41134 46786
rect 41186 46734 41188 46786
rect 41132 46722 41188 46734
rect 41020 46676 41076 46686
rect 40796 46674 41076 46676
rect 40796 46622 41022 46674
rect 41074 46622 41076 46674
rect 40796 46620 41076 46622
rect 41020 46610 41076 46620
rect 41132 45780 41188 45790
rect 41132 44772 41188 45724
rect 41244 45332 41300 45342
rect 41468 45332 41524 47516
rect 41692 47458 41748 48750
rect 41692 47406 41694 47458
rect 41746 47406 41748 47458
rect 41692 47394 41748 47406
rect 41804 46900 41860 51100
rect 42028 50820 42084 50830
rect 42028 50708 42084 50764
rect 42028 50706 42420 50708
rect 42028 50654 42030 50706
rect 42082 50654 42420 50706
rect 42028 50652 42420 50654
rect 42028 50642 42084 50652
rect 42028 50484 42084 50494
rect 42028 49922 42084 50428
rect 42028 49870 42030 49922
rect 42082 49870 42084 49922
rect 41916 49700 41972 49710
rect 41916 49606 41972 49644
rect 41300 45276 41524 45332
rect 41580 46844 41860 46900
rect 41244 44996 41300 45276
rect 41580 45220 41636 46844
rect 41916 46788 41972 46798
rect 41804 46732 41916 46788
rect 41244 44902 41300 44940
rect 41356 45164 41636 45220
rect 41692 45332 41748 45342
rect 41132 44716 41300 44772
rect 41244 44660 41300 44716
rect 41132 44548 41188 44558
rect 40684 44492 41076 44548
rect 40348 44434 40404 44492
rect 40348 44382 40350 44434
rect 40402 44382 40404 44434
rect 40348 44370 40404 44382
rect 40796 44212 40852 44222
rect 40796 44118 40852 44156
rect 40908 44100 40964 44110
rect 40348 43876 40404 43886
rect 40124 43652 40180 43662
rect 40124 42196 40180 43596
rect 40348 43426 40404 43820
rect 40348 43374 40350 43426
rect 40402 43374 40404 43426
rect 40348 43362 40404 43374
rect 40236 42756 40292 42766
rect 40236 42754 40628 42756
rect 40236 42702 40238 42754
rect 40290 42702 40628 42754
rect 40236 42700 40628 42702
rect 40236 42690 40292 42700
rect 40124 42082 40180 42140
rect 40124 42030 40126 42082
rect 40178 42030 40180 42082
rect 40124 42018 40180 42030
rect 40236 42082 40292 42094
rect 40236 42030 40238 42082
rect 40290 42030 40292 42082
rect 40236 41972 40292 42030
rect 40292 41916 40404 41972
rect 40236 41906 40292 41916
rect 40012 41804 40180 41860
rect 39676 41746 39732 41758
rect 39676 41694 39678 41746
rect 39730 41694 39732 41746
rect 39676 40628 39732 41694
rect 39676 40562 39732 40572
rect 39788 41524 39844 41534
rect 39676 40402 39732 40414
rect 39676 40350 39678 40402
rect 39730 40350 39732 40402
rect 39676 39060 39732 40350
rect 39676 38994 39732 39004
rect 39676 38836 39732 38846
rect 39788 38836 39844 41468
rect 39900 39842 39956 39854
rect 39900 39790 39902 39842
rect 39954 39790 39956 39842
rect 39900 39730 39956 39790
rect 39900 39678 39902 39730
rect 39954 39678 39956 39730
rect 39900 39666 39956 39678
rect 39676 38834 39788 38836
rect 39676 38782 39678 38834
rect 39730 38782 39788 38834
rect 39676 38780 39788 38782
rect 39676 38770 39732 38780
rect 39788 38742 39844 38780
rect 40012 39620 40068 39630
rect 40012 38834 40068 39564
rect 40124 39284 40180 41804
rect 40236 41748 40292 41758
rect 40236 41654 40292 41692
rect 40348 41412 40404 41916
rect 40236 41356 40404 41412
rect 40236 40626 40292 41356
rect 40236 40574 40238 40626
rect 40290 40574 40292 40626
rect 40236 40562 40292 40574
rect 40460 41298 40516 41310
rect 40460 41246 40462 41298
rect 40514 41246 40516 41298
rect 40348 40516 40404 40526
rect 40460 40516 40516 41246
rect 40348 40514 40516 40516
rect 40348 40462 40350 40514
rect 40402 40462 40516 40514
rect 40348 40460 40516 40462
rect 40348 40450 40404 40460
rect 40348 40292 40404 40302
rect 40348 40068 40404 40236
rect 40348 39730 40404 40012
rect 40348 39678 40350 39730
rect 40402 39678 40404 39730
rect 40348 39666 40404 39678
rect 40124 39218 40180 39228
rect 40012 38782 40014 38834
rect 40066 38782 40068 38834
rect 40012 38770 40068 38782
rect 40012 38612 40068 38622
rect 40012 38610 40180 38612
rect 40012 38558 40014 38610
rect 40066 38558 40180 38610
rect 40012 38556 40180 38558
rect 40012 38546 40068 38556
rect 40124 38162 40180 38556
rect 40124 38110 40126 38162
rect 40178 38110 40180 38162
rect 40124 38098 40180 38110
rect 40572 36484 40628 42700
rect 40684 42642 40740 42654
rect 40684 42590 40686 42642
rect 40738 42590 40740 42642
rect 40684 40404 40740 42590
rect 40908 41188 40964 44044
rect 41020 43652 41076 44492
rect 41020 43558 41076 43596
rect 40684 40338 40740 40348
rect 40796 41186 40964 41188
rect 40796 41134 40910 41186
rect 40962 41134 40964 41186
rect 40796 41132 40964 41134
rect 40796 40628 40852 41132
rect 40908 41122 40964 41132
rect 40796 39844 40852 40572
rect 40908 40964 40964 40974
rect 40908 40514 40964 40908
rect 40908 40462 40910 40514
rect 40962 40462 40964 40514
rect 40908 39956 40964 40462
rect 41020 40740 41076 40750
rect 41020 40402 41076 40684
rect 41020 40350 41022 40402
rect 41074 40350 41076 40402
rect 41020 40338 41076 40350
rect 40908 39900 41076 39956
rect 40852 39788 40964 39844
rect 40796 39778 40852 39788
rect 40908 39730 40964 39788
rect 40908 39678 40910 39730
rect 40962 39678 40964 39730
rect 40908 39666 40964 39678
rect 40348 36428 40628 36484
rect 40684 39284 40740 39294
rect 40684 36484 40740 39228
rect 41020 39058 41076 39900
rect 41132 39396 41188 44492
rect 41244 44100 41300 44604
rect 41244 44006 41300 44044
rect 41244 41970 41300 41982
rect 41244 41918 41246 41970
rect 41298 41918 41300 41970
rect 41244 41860 41300 41918
rect 41244 40516 41300 41804
rect 41244 40450 41300 40460
rect 41356 40290 41412 45164
rect 41692 45106 41748 45276
rect 41692 45054 41694 45106
rect 41746 45054 41748 45106
rect 41580 44882 41636 44894
rect 41580 44830 41582 44882
rect 41634 44830 41636 44882
rect 41580 44322 41636 44830
rect 41692 44548 41748 45054
rect 41692 44482 41748 44492
rect 41580 44270 41582 44322
rect 41634 44270 41636 44322
rect 41580 44258 41636 44270
rect 41804 44212 41860 46732
rect 41916 46722 41972 46732
rect 41916 45556 41972 45566
rect 41916 45218 41972 45500
rect 41916 45166 41918 45218
rect 41970 45166 41972 45218
rect 41916 45154 41972 45166
rect 42028 44436 42084 49870
rect 42364 49810 42420 50652
rect 42364 49758 42366 49810
rect 42418 49758 42420 49810
rect 42252 49250 42308 49262
rect 42252 49198 42254 49250
rect 42306 49198 42308 49250
rect 42140 48802 42196 48814
rect 42140 48750 42142 48802
rect 42194 48750 42196 48802
rect 42140 48356 42196 48750
rect 42140 48290 42196 48300
rect 42252 48242 42308 49198
rect 42252 48190 42254 48242
rect 42306 48190 42308 48242
rect 42252 47908 42308 48190
rect 42252 47842 42308 47852
rect 42364 47684 42420 49758
rect 42588 49138 42644 53116
rect 42812 53170 42868 53788
rect 43596 53844 43652 53854
rect 43148 53508 43204 53518
rect 43148 53414 43204 53452
rect 42812 53118 42814 53170
rect 42866 53118 42868 53170
rect 42812 53106 42868 53118
rect 43148 53172 43204 53182
rect 43148 52946 43204 53116
rect 43148 52894 43150 52946
rect 43202 52894 43204 52946
rect 43148 52882 43204 52894
rect 43372 52388 43428 52398
rect 43428 52332 43540 52388
rect 43372 52322 43428 52332
rect 42812 52164 42868 52174
rect 42812 51378 42868 52108
rect 42812 51326 42814 51378
rect 42866 51326 42868 51378
rect 42812 51314 42868 51326
rect 42700 51156 42756 51166
rect 42700 51154 42868 51156
rect 42700 51102 42702 51154
rect 42754 51102 42868 51154
rect 42700 51100 42868 51102
rect 42700 51090 42756 51100
rect 42588 49086 42590 49138
rect 42642 49086 42644 49138
rect 42588 49074 42644 49086
rect 42140 47628 42420 47684
rect 42476 48692 42532 48702
rect 42140 45780 42196 47628
rect 42252 47236 42308 47246
rect 42252 46002 42308 47180
rect 42252 45950 42254 46002
rect 42306 45950 42308 46002
rect 42252 45938 42308 45950
rect 42364 47124 42420 47134
rect 42140 45724 42308 45780
rect 42028 44370 42084 44380
rect 42252 44212 42308 45724
rect 42364 45556 42420 47068
rect 42364 45490 42420 45500
rect 42476 46114 42532 48636
rect 42700 48244 42756 48254
rect 42700 47570 42756 48188
rect 42700 47518 42702 47570
rect 42754 47518 42756 47570
rect 42700 47460 42756 47518
rect 42700 47394 42756 47404
rect 42476 46062 42478 46114
rect 42530 46062 42532 46114
rect 42476 45332 42532 46062
rect 42588 47348 42644 47358
rect 42812 47348 42868 51100
rect 43148 49700 43204 49710
rect 43148 49606 43204 49644
rect 43036 49250 43092 49262
rect 43036 49198 43038 49250
rect 43090 49198 43092 49250
rect 43036 49138 43092 49198
rect 43036 49086 43038 49138
rect 43090 49086 43092 49138
rect 43036 49074 43092 49086
rect 42924 48692 42980 48702
rect 42924 48466 42980 48636
rect 42924 48414 42926 48466
rect 42978 48414 42980 48466
rect 42924 48402 42980 48414
rect 43372 48130 43428 48142
rect 43372 48078 43374 48130
rect 43426 48078 43428 48130
rect 42924 47572 42980 47582
rect 43372 47572 43428 48078
rect 42924 47570 43428 47572
rect 42924 47518 42926 47570
rect 42978 47518 43428 47570
rect 42924 47516 43428 47518
rect 42924 47506 42980 47516
rect 43260 47348 43316 47358
rect 42812 47292 43204 47348
rect 42588 45668 42644 47292
rect 43148 47012 43204 47292
rect 43260 47234 43316 47292
rect 43260 47182 43262 47234
rect 43314 47182 43316 47234
rect 43260 47170 43316 47182
rect 43148 46956 43316 47012
rect 43148 46114 43204 46126
rect 43148 46062 43150 46114
rect 43202 46062 43204 46114
rect 43148 46002 43204 46062
rect 43148 45950 43150 46002
rect 43202 45950 43204 46002
rect 43148 45938 43204 45950
rect 42588 45602 42644 45612
rect 42700 45666 42756 45678
rect 42700 45614 42702 45666
rect 42754 45614 42756 45666
rect 42700 45556 42756 45614
rect 42700 45490 42756 45500
rect 42924 45668 42980 45678
rect 42476 45266 42532 45276
rect 42364 45220 42420 45230
rect 42364 45106 42420 45164
rect 42364 45054 42366 45106
rect 42418 45054 42420 45106
rect 42364 45042 42420 45054
rect 42924 45106 42980 45612
rect 43148 45556 43204 45566
rect 42924 45054 42926 45106
rect 42978 45054 42980 45106
rect 42700 44996 42756 45006
rect 42700 44434 42756 44940
rect 42700 44382 42702 44434
rect 42754 44382 42756 44434
rect 42588 44324 42644 44334
rect 42588 44230 42644 44268
rect 41804 44156 41972 44212
rect 41804 43764 41860 43774
rect 41804 43670 41860 43708
rect 41468 41972 41524 41982
rect 41468 41878 41524 41916
rect 41692 41748 41748 41758
rect 41692 41298 41748 41692
rect 41916 41746 41972 44156
rect 41916 41694 41918 41746
rect 41970 41694 41972 41746
rect 41916 41682 41972 41694
rect 42028 44156 42308 44212
rect 41692 41246 41694 41298
rect 41746 41246 41748 41298
rect 41692 41234 41748 41246
rect 41692 40740 41748 40750
rect 41356 40238 41358 40290
rect 41410 40238 41412 40290
rect 41356 39956 41412 40238
rect 41356 39890 41412 39900
rect 41468 40404 41524 40414
rect 41244 39844 41300 39854
rect 41244 39732 41300 39788
rect 41356 39732 41412 39742
rect 41244 39730 41412 39732
rect 41244 39678 41358 39730
rect 41410 39678 41412 39730
rect 41244 39676 41412 39678
rect 41356 39666 41412 39676
rect 41132 39330 41188 39340
rect 41468 39618 41524 40348
rect 41468 39566 41470 39618
rect 41522 39566 41524 39618
rect 41020 39006 41022 39058
rect 41074 39006 41076 39058
rect 41020 38994 41076 39006
rect 41468 39060 41524 39566
rect 41468 38994 41524 39004
rect 41468 38836 41524 38846
rect 41468 38742 41524 38780
rect 41132 38610 41188 38622
rect 41132 38558 41134 38610
rect 41186 38558 41188 38610
rect 40908 38050 40964 38062
rect 40908 37998 40910 38050
rect 40962 37998 40964 38050
rect 40908 37156 40964 37998
rect 41132 37490 41188 38558
rect 41356 38612 41412 38622
rect 41356 38162 41412 38556
rect 41356 38110 41358 38162
rect 41410 38110 41412 38162
rect 41356 38098 41412 38110
rect 41692 38610 41748 40684
rect 42028 40068 42084 44156
rect 42476 42530 42532 42542
rect 42476 42478 42478 42530
rect 42530 42478 42532 42530
rect 42252 41972 42308 41982
rect 42476 41972 42532 42478
rect 42308 41916 42532 41972
rect 42028 40002 42084 40012
rect 42140 40516 42196 40526
rect 42140 39730 42196 40460
rect 42252 40404 42308 41916
rect 42252 40338 42308 40348
rect 42140 39678 42142 39730
rect 42194 39678 42196 39730
rect 42140 39666 42196 39678
rect 42588 39620 42644 39630
rect 42588 39526 42644 39564
rect 42364 39396 42420 39406
rect 41916 39060 41972 39070
rect 42364 39060 42420 39340
rect 41916 38966 41972 39004
rect 42028 39058 42420 39060
rect 42028 39006 42366 39058
rect 42418 39006 42420 39058
rect 42028 39004 42420 39006
rect 41692 38558 41694 38610
rect 41746 38558 41748 38610
rect 41132 37438 41134 37490
rect 41186 37438 41188 37490
rect 41132 37426 41188 37438
rect 41580 37492 41636 37502
rect 41580 37398 41636 37436
rect 40908 37090 40964 37100
rect 41356 36596 41412 36606
rect 41356 36502 41412 36540
rect 41132 36484 41188 36494
rect 41692 36484 41748 38558
rect 42028 38500 42084 39004
rect 42364 38994 42420 39004
rect 42700 38724 42756 44382
rect 42812 44210 42868 44222
rect 42812 44158 42814 44210
rect 42866 44158 42868 44210
rect 42812 43650 42868 44158
rect 42924 44212 42980 45054
rect 42924 44146 42980 44156
rect 43036 45332 43092 45342
rect 42812 43598 42814 43650
rect 42866 43598 42868 43650
rect 42812 43586 42868 43598
rect 42924 42530 42980 42542
rect 42924 42478 42926 42530
rect 42978 42478 42980 42530
rect 42812 41972 42868 41982
rect 42924 41972 42980 42478
rect 42868 41916 42980 41972
rect 42812 41878 42868 41916
rect 42812 40740 42868 40750
rect 42812 40626 42868 40684
rect 42812 40574 42814 40626
rect 42866 40574 42868 40626
rect 42812 40562 42868 40574
rect 42924 39506 42980 39518
rect 42924 39454 42926 39506
rect 42978 39454 42980 39506
rect 42812 38724 42868 38734
rect 42700 38722 42868 38724
rect 42700 38670 42814 38722
rect 42866 38670 42868 38722
rect 42700 38668 42868 38670
rect 41916 38444 42084 38500
rect 42140 38612 42196 38622
rect 41916 38050 41972 38444
rect 41916 37998 41918 38050
rect 41970 37998 41972 38050
rect 41916 37986 41972 37998
rect 42140 38050 42196 38556
rect 42140 37998 42142 38050
rect 42194 37998 42196 38050
rect 42140 37986 42196 37998
rect 42476 38610 42532 38622
rect 42476 38558 42478 38610
rect 42530 38558 42532 38610
rect 42476 37940 42532 38558
rect 42812 38052 42868 38668
rect 42924 38388 42980 39454
rect 43036 38388 43092 45276
rect 43148 38612 43204 45500
rect 43260 43538 43316 46956
rect 43372 45108 43428 47516
rect 43484 45332 43540 52332
rect 43596 52386 43652 53788
rect 44044 53842 44100 54348
rect 44268 54338 44324 54348
rect 44044 53790 44046 53842
rect 44098 53790 44100 53842
rect 44044 53778 44100 53790
rect 43932 53508 43988 53518
rect 43932 53506 44100 53508
rect 43932 53454 43934 53506
rect 43986 53454 44100 53506
rect 43932 53452 44100 53454
rect 43932 53442 43988 53452
rect 43596 52334 43598 52386
rect 43650 52334 43652 52386
rect 43596 52322 43652 52334
rect 43932 52834 43988 52846
rect 43932 52782 43934 52834
rect 43986 52782 43988 52834
rect 43932 52386 43988 52782
rect 43932 52334 43934 52386
rect 43986 52334 43988 52386
rect 43932 52322 43988 52334
rect 43932 52164 43988 52174
rect 44044 52164 44100 53452
rect 45164 52836 45220 52846
rect 45052 52276 45108 52286
rect 45052 52182 45108 52220
rect 45164 52274 45220 52780
rect 46060 52836 46116 52846
rect 46060 52742 46116 52780
rect 45164 52222 45166 52274
rect 45218 52222 45220 52274
rect 45164 52210 45220 52222
rect 43988 52108 44100 52164
rect 43932 52070 43988 52108
rect 43708 51604 43764 51614
rect 43708 51510 43764 51548
rect 44156 51604 44212 51614
rect 44156 51510 44212 51548
rect 45276 49700 45332 49710
rect 44940 49698 45332 49700
rect 44940 49646 45278 49698
rect 45330 49646 45332 49698
rect 44940 49644 45332 49646
rect 44940 49138 44996 49644
rect 45276 49634 45332 49644
rect 44940 49086 44942 49138
rect 44994 49086 44996 49138
rect 44940 49074 44996 49086
rect 44828 48802 44884 48814
rect 44828 48750 44830 48802
rect 44882 48750 44884 48802
rect 43820 47348 43876 47358
rect 43820 47254 43876 47292
rect 44156 47234 44212 47246
rect 44156 47182 44158 47234
rect 44210 47182 44212 47234
rect 43596 46788 43652 46798
rect 43596 46694 43652 46732
rect 44156 46788 44212 47182
rect 44156 46722 44212 46732
rect 44716 46676 44772 46686
rect 44380 46674 44772 46676
rect 44380 46622 44718 46674
rect 44770 46622 44772 46674
rect 44380 46620 44772 46622
rect 43484 45266 43540 45276
rect 43596 45666 43652 45678
rect 43596 45614 43598 45666
rect 43650 45614 43652 45666
rect 43596 45556 43652 45614
rect 44044 45668 44100 45678
rect 44044 45574 44100 45612
rect 43372 45042 43428 45052
rect 43484 45108 43540 45118
rect 43596 45108 43652 45500
rect 43484 45106 43652 45108
rect 43484 45054 43486 45106
rect 43538 45054 43652 45106
rect 43484 45052 43652 45054
rect 43484 44660 43540 45052
rect 44268 44996 44324 45006
rect 43484 44594 43540 44604
rect 44044 44994 44324 44996
rect 44044 44942 44270 44994
rect 44322 44942 44324 44994
rect 44044 44940 44324 44942
rect 44044 44546 44100 44940
rect 44268 44930 44324 44940
rect 44044 44494 44046 44546
rect 44098 44494 44100 44546
rect 44044 44482 44100 44494
rect 43372 44436 43428 44446
rect 43708 44436 43764 44446
rect 43428 44434 43764 44436
rect 43428 44382 43710 44434
rect 43762 44382 43764 44434
rect 43428 44380 43764 44382
rect 43372 44342 43428 44380
rect 43260 43486 43262 43538
rect 43314 43486 43316 43538
rect 43260 43474 43316 43486
rect 43372 44212 43428 44222
rect 43372 43316 43428 44156
rect 43260 43260 43428 43316
rect 43260 40516 43316 43260
rect 43372 41860 43428 41870
rect 43372 41766 43428 41804
rect 43260 40460 43428 40516
rect 43260 40292 43316 40302
rect 43260 40198 43316 40236
rect 43148 38546 43204 38556
rect 43036 38332 43316 38388
rect 42924 38322 42980 38332
rect 42924 38052 42980 38062
rect 42812 38050 42980 38052
rect 42812 37998 42926 38050
rect 42978 37998 42980 38050
rect 42812 37996 42980 37998
rect 42924 37986 42980 37996
rect 42588 37940 42644 37950
rect 42476 37938 42644 37940
rect 42476 37886 42590 37938
rect 42642 37886 42644 37938
rect 42476 37884 42644 37886
rect 42588 37874 42644 37884
rect 42364 37826 42420 37838
rect 42364 37774 42366 37826
rect 42418 37774 42420 37826
rect 42364 36596 42420 37774
rect 42700 37828 42756 37838
rect 42700 37734 42756 37772
rect 43036 37826 43092 37838
rect 43036 37774 43038 37826
rect 43090 37774 43092 37826
rect 42588 37380 42644 37390
rect 43036 37380 43092 37774
rect 43148 37826 43204 37838
rect 43148 37774 43150 37826
rect 43202 37774 43204 37826
rect 43148 37716 43204 37774
rect 43148 37650 43204 37660
rect 42588 37378 43092 37380
rect 42588 37326 42590 37378
rect 42642 37326 43092 37378
rect 42588 37324 43092 37326
rect 42588 37314 42644 37324
rect 43148 37268 43204 37278
rect 43260 37268 43316 38332
rect 43372 38052 43428 40460
rect 43484 39058 43540 44380
rect 43708 44370 43764 44380
rect 44044 44324 44100 44334
rect 44044 44230 44100 44268
rect 43596 43652 43652 43662
rect 43596 41746 43652 43596
rect 44268 43652 44324 43662
rect 44268 43558 44324 43596
rect 43596 41694 43598 41746
rect 43650 41694 43652 41746
rect 43596 41682 43652 41694
rect 43708 43538 43764 43550
rect 43708 43486 43710 43538
rect 43762 43486 43764 43538
rect 43596 40628 43652 40638
rect 43596 40404 43652 40572
rect 43596 40310 43652 40348
rect 43484 39006 43486 39058
rect 43538 39006 43540 39058
rect 43484 38276 43540 39006
rect 43484 38210 43540 38220
rect 43372 37996 43540 38052
rect 43372 37828 43428 37838
rect 43372 37734 43428 37772
rect 43148 37266 43316 37268
rect 43148 37214 43150 37266
rect 43202 37214 43316 37266
rect 43148 37212 43316 37214
rect 43148 37202 43204 37212
rect 42364 36530 42420 36540
rect 43484 36594 43540 37996
rect 43484 36542 43486 36594
rect 43538 36542 43540 36594
rect 40684 36482 41188 36484
rect 40684 36430 41134 36482
rect 41186 36430 41188 36482
rect 40684 36428 41188 36430
rect 40012 35028 40068 35038
rect 40012 35026 40292 35028
rect 40012 34974 40014 35026
rect 40066 34974 40292 35026
rect 40012 34972 40292 34974
rect 40012 34962 40068 34972
rect 39676 34242 39732 34254
rect 39676 34190 39678 34242
rect 39730 34190 39732 34242
rect 39676 34132 39732 34190
rect 40236 34242 40292 34972
rect 40236 34190 40238 34242
rect 40290 34190 40292 34242
rect 40236 34178 40292 34190
rect 40124 34132 40180 34142
rect 39676 34130 40180 34132
rect 39676 34078 40126 34130
rect 40178 34078 40180 34130
rect 39676 34076 40180 34078
rect 39676 32562 39732 34076
rect 40124 34066 40180 34076
rect 39788 33908 39844 33918
rect 39788 33906 40068 33908
rect 39788 33854 39790 33906
rect 39842 33854 40068 33906
rect 39788 33852 40068 33854
rect 39788 33842 39844 33852
rect 40012 33458 40068 33852
rect 40348 33572 40404 36428
rect 40460 36260 40516 36270
rect 40684 36260 40740 36428
rect 40460 36258 40740 36260
rect 40460 36206 40462 36258
rect 40514 36206 40740 36258
rect 40460 36204 40740 36206
rect 40796 36258 40852 36270
rect 40796 36206 40798 36258
rect 40850 36206 40852 36258
rect 40460 36194 40516 36204
rect 40796 34914 40852 36206
rect 40796 34862 40798 34914
rect 40850 34862 40852 34914
rect 40796 34850 40852 34862
rect 40012 33406 40014 33458
rect 40066 33406 40068 33458
rect 40012 33394 40068 33406
rect 40124 33516 40404 33572
rect 40572 34690 40628 34702
rect 40572 34638 40574 34690
rect 40626 34638 40628 34690
rect 40124 32674 40180 33516
rect 40124 32622 40126 32674
rect 40178 32622 40180 32674
rect 40124 32610 40180 32622
rect 39676 32510 39678 32562
rect 39730 32510 39732 32562
rect 39676 32498 39732 32510
rect 40572 31948 40628 34638
rect 40908 32452 40964 32462
rect 39564 31892 39732 31948
rect 40572 31892 40740 31948
rect 39340 31778 39396 31790
rect 39340 31726 39342 31778
rect 39394 31726 39396 31778
rect 39340 30884 39396 31726
rect 39564 30884 39620 30894
rect 39340 30882 39620 30884
rect 39340 30830 39566 30882
rect 39618 30830 39620 30882
rect 39340 30828 39620 30830
rect 39228 29540 39284 29550
rect 39564 29540 39620 30828
rect 39228 29538 39620 29540
rect 39228 29486 39230 29538
rect 39282 29486 39620 29538
rect 39228 29484 39620 29486
rect 39228 29474 39284 29484
rect 39452 29204 39508 29214
rect 39452 29110 39508 29148
rect 39676 27972 39732 31892
rect 40124 31778 40180 31790
rect 40124 31726 40126 31778
rect 40178 31726 40180 31778
rect 40124 31556 40180 31726
rect 40124 31490 40180 31500
rect 40572 31556 40628 31566
rect 40572 31462 40628 31500
rect 40348 30212 40404 30222
rect 40348 30118 40404 30156
rect 39788 29204 39844 29214
rect 39788 29202 40068 29204
rect 39788 29150 39790 29202
rect 39842 29150 40068 29202
rect 39788 29148 40068 29150
rect 39788 29138 39844 29148
rect 39340 27916 39732 27972
rect 40012 27970 40068 29148
rect 40572 28756 40628 28766
rect 40684 28756 40740 31892
rect 40796 31220 40852 31230
rect 40796 30322 40852 31164
rect 40796 30270 40798 30322
rect 40850 30270 40852 30322
rect 40796 30258 40852 30270
rect 40908 30884 40964 32396
rect 40908 29650 40964 30828
rect 40908 29598 40910 29650
rect 40962 29598 40964 29650
rect 40908 29586 40964 29598
rect 41132 29652 41188 36428
rect 41468 36482 41748 36484
rect 41468 36430 41694 36482
rect 41746 36430 41748 36482
rect 41468 36428 41748 36430
rect 41356 35924 41412 35934
rect 41468 35924 41524 36428
rect 41692 36418 41748 36428
rect 41356 35922 41524 35924
rect 41356 35870 41358 35922
rect 41410 35870 41524 35922
rect 41356 35868 41524 35870
rect 41356 35858 41412 35868
rect 42028 35700 42084 35710
rect 42028 33348 42084 35644
rect 43260 35698 43316 35710
rect 43260 35646 43262 35698
rect 43314 35646 43316 35698
rect 42924 35588 42980 35598
rect 43260 35588 43316 35646
rect 43484 35700 43540 36542
rect 43484 35634 43540 35644
rect 42924 35586 43316 35588
rect 42924 35534 42926 35586
rect 42978 35534 43316 35586
rect 42924 35532 43316 35534
rect 42700 34356 42756 34366
rect 42700 34262 42756 34300
rect 42140 33460 42196 33470
rect 42140 33458 42420 33460
rect 42140 33406 42142 33458
rect 42194 33406 42420 33458
rect 42140 33404 42420 33406
rect 42140 33394 42196 33404
rect 41916 33292 42084 33348
rect 41916 31778 41972 33292
rect 42028 33124 42084 33134
rect 42028 32786 42084 33068
rect 42028 32734 42030 32786
rect 42082 32734 42084 32786
rect 42028 32722 42084 32734
rect 42364 32674 42420 33404
rect 42588 33346 42644 33358
rect 42588 33294 42590 33346
rect 42642 33294 42644 33346
rect 42476 32788 42532 32798
rect 42476 32694 42532 32732
rect 42364 32622 42366 32674
rect 42418 32622 42420 32674
rect 42364 32610 42420 32622
rect 42588 32002 42644 33294
rect 42924 33124 42980 35532
rect 43036 34356 43092 34366
rect 43036 34242 43092 34300
rect 43036 34190 43038 34242
rect 43090 34190 43092 34242
rect 43036 34178 43092 34190
rect 43260 34242 43316 34254
rect 43260 34190 43262 34242
rect 43314 34190 43316 34242
rect 43260 33346 43316 34190
rect 43372 33908 43428 33918
rect 43372 33906 43652 33908
rect 43372 33854 43374 33906
rect 43426 33854 43652 33906
rect 43372 33852 43652 33854
rect 43372 33842 43428 33852
rect 43372 33460 43428 33470
rect 43372 33458 43540 33460
rect 43372 33406 43374 33458
rect 43426 33406 43540 33458
rect 43372 33404 43540 33406
rect 43372 33394 43428 33404
rect 43260 33294 43262 33346
rect 43314 33294 43316 33346
rect 43036 33124 43092 33134
rect 42924 33068 43036 33124
rect 43036 32564 43092 33068
rect 43148 32788 43204 32798
rect 43260 32788 43316 33294
rect 43204 32732 43316 32788
rect 43148 32722 43204 32732
rect 43036 32470 43092 32508
rect 42588 31950 42590 32002
rect 42642 31950 42644 32002
rect 42588 31938 42644 31950
rect 43484 31948 43540 33404
rect 43596 32788 43652 33852
rect 43708 33012 43764 43486
rect 43820 41972 43876 41982
rect 43820 41970 44324 41972
rect 43820 41918 43822 41970
rect 43874 41918 44324 41970
rect 43820 41916 44324 41918
rect 43820 41906 43876 41916
rect 44268 41410 44324 41916
rect 44268 41358 44270 41410
rect 44322 41358 44324 41410
rect 43820 41300 43876 41310
rect 44156 41300 44212 41310
rect 43820 41298 44212 41300
rect 43820 41246 43822 41298
rect 43874 41246 44158 41298
rect 44210 41246 44212 41298
rect 43820 41244 44212 41246
rect 43820 41234 43876 41244
rect 44156 41234 44212 41244
rect 44268 40964 44324 41358
rect 44268 40898 44324 40908
rect 44380 40740 44436 46620
rect 44716 46610 44772 46620
rect 44828 44324 44884 48750
rect 45948 46788 46004 46798
rect 45948 46694 46004 46732
rect 45164 46674 45220 46686
rect 45164 46622 45166 46674
rect 45218 46622 45220 46674
rect 44940 45668 44996 45678
rect 45164 45668 45220 46622
rect 44940 45666 45220 45668
rect 44940 45614 44942 45666
rect 44994 45614 45220 45666
rect 44940 45612 45220 45614
rect 48076 46562 48132 46574
rect 48076 46510 48078 46562
rect 48130 46510 48132 46562
rect 44940 45556 44996 45612
rect 44940 45490 44996 45500
rect 45164 45220 45220 45230
rect 48076 45220 48132 46510
rect 45220 45164 45332 45220
rect 45164 45154 45220 45164
rect 44828 44258 44884 44268
rect 44604 41858 44660 41870
rect 44604 41806 44606 41858
rect 44658 41806 44660 41858
rect 44604 41524 44660 41806
rect 44604 41458 44660 41468
rect 45164 41524 45220 41534
rect 45164 41410 45220 41468
rect 45164 41358 45166 41410
rect 45218 41358 45220 41410
rect 45164 41346 45220 41358
rect 43932 40684 44436 40740
rect 44828 41298 44884 41310
rect 44828 41246 44830 41298
rect 44882 41246 44884 41298
rect 43820 38276 43876 38286
rect 43820 38182 43876 38220
rect 43932 38052 43988 40684
rect 44828 40628 44884 41246
rect 44940 40964 44996 40974
rect 44940 40870 44996 40908
rect 44380 40572 44884 40628
rect 44380 40514 44436 40572
rect 44380 40462 44382 40514
rect 44434 40462 44436 40514
rect 44380 40450 44436 40462
rect 45052 39844 45108 39854
rect 44268 39842 45108 39844
rect 44268 39790 45054 39842
rect 45106 39790 45108 39842
rect 44268 39788 45108 39790
rect 44268 39730 44324 39788
rect 45052 39778 45108 39788
rect 45276 39732 45332 45164
rect 48076 45154 48132 45164
rect 46396 44996 46452 45006
rect 45948 44994 46452 44996
rect 45948 44942 46398 44994
rect 46450 44942 46452 44994
rect 45948 44940 46452 44942
rect 45948 43650 46004 44940
rect 46396 44930 46452 44940
rect 45948 43598 45950 43650
rect 46002 43598 46004 43650
rect 45948 43586 46004 43598
rect 44268 39678 44270 39730
rect 44322 39678 44324 39730
rect 44156 38612 44212 38622
rect 43820 37996 43988 38052
rect 44044 38556 44156 38612
rect 43820 33234 43876 37996
rect 44044 37940 44100 38556
rect 44156 38546 44212 38556
rect 44044 37846 44100 37884
rect 44156 38388 44212 38398
rect 43932 37826 43988 37838
rect 43932 37774 43934 37826
rect 43986 37774 43988 37826
rect 43932 35812 43988 37774
rect 44044 37380 44100 37390
rect 44156 37380 44212 38332
rect 44044 37378 44212 37380
rect 44044 37326 44046 37378
rect 44098 37326 44212 37378
rect 44044 37324 44212 37326
rect 44044 37314 44100 37324
rect 44268 36932 44324 39678
rect 45164 39676 45332 39732
rect 45836 43314 45892 43326
rect 45836 43262 45838 43314
rect 45890 43262 45892 43314
rect 44828 39620 44884 39630
rect 45164 39620 45220 39676
rect 44828 39618 45220 39620
rect 44828 39566 44830 39618
rect 44882 39566 45220 39618
rect 44828 39564 45220 39566
rect 44828 39554 44884 39564
rect 45388 39508 45444 39518
rect 45724 39508 45780 39518
rect 45388 39506 45780 39508
rect 45388 39454 45390 39506
rect 45442 39454 45726 39506
rect 45778 39454 45780 39506
rect 45388 39452 45780 39454
rect 45388 39442 45444 39452
rect 45724 39442 45780 39452
rect 45836 38612 45892 43262
rect 46508 40290 46564 40302
rect 46508 40238 46510 40290
rect 46562 40238 46564 40290
rect 46508 39730 46564 40238
rect 46508 39678 46510 39730
rect 46562 39678 46564 39730
rect 46508 39666 46564 39678
rect 46396 39620 46452 39630
rect 46396 39526 46452 39564
rect 45836 38546 45892 38556
rect 46060 39394 46116 39406
rect 46060 39342 46062 39394
rect 46114 39342 46116 39394
rect 45164 37268 45220 37278
rect 44268 36866 44324 36876
rect 44716 37266 45220 37268
rect 44716 37214 45166 37266
rect 45218 37214 45220 37266
rect 44716 37212 45220 37214
rect 44044 35812 44100 35822
rect 43932 35810 44100 35812
rect 43932 35758 44046 35810
rect 44098 35758 44100 35810
rect 43932 35756 44100 35758
rect 44044 35746 44100 35756
rect 44268 34356 44324 34366
rect 44268 33684 44324 34300
rect 44268 33458 44324 33628
rect 44268 33406 44270 33458
rect 44322 33406 44324 33458
rect 44268 33394 44324 33406
rect 43820 33182 43822 33234
rect 43874 33182 43876 33234
rect 43820 33170 43876 33182
rect 43708 32956 43988 33012
rect 43596 32732 43876 32788
rect 43820 32674 43876 32732
rect 43820 32622 43822 32674
rect 43874 32622 43876 32674
rect 43820 32610 43876 32622
rect 43372 31892 43540 31948
rect 43596 32116 43652 32126
rect 41916 31726 41918 31778
rect 41970 31726 41972 31778
rect 41356 31668 41412 31678
rect 41244 31554 41300 31566
rect 41244 31502 41246 31554
rect 41298 31502 41300 31554
rect 41244 31220 41300 31502
rect 41244 31154 41300 31164
rect 41356 30884 41412 31612
rect 41804 31668 41860 31678
rect 41804 31574 41860 31612
rect 41916 31556 41972 31726
rect 41468 30884 41524 30894
rect 41356 30882 41524 30884
rect 41356 30830 41470 30882
rect 41522 30830 41524 30882
rect 41356 30828 41524 30830
rect 41356 30436 41412 30828
rect 41468 30818 41524 30828
rect 41356 30380 41748 30436
rect 41244 30324 41300 30334
rect 41356 30324 41412 30380
rect 41244 30322 41412 30324
rect 41244 30270 41246 30322
rect 41298 30270 41412 30322
rect 41244 30268 41412 30270
rect 41692 30324 41748 30380
rect 41244 30258 41300 30268
rect 41580 30212 41636 30222
rect 41580 30118 41636 30156
rect 41692 30098 41748 30268
rect 41692 30046 41694 30098
rect 41746 30046 41748 30098
rect 41692 30034 41748 30046
rect 41916 29876 41972 31500
rect 42700 31778 42756 31790
rect 42700 31726 42702 31778
rect 42754 31726 42756 31778
rect 41804 29820 41972 29876
rect 42028 31220 42084 31230
rect 41132 29596 41300 29652
rect 41132 29426 41188 29438
rect 41132 29374 41134 29426
rect 41186 29374 41188 29426
rect 41020 29316 41076 29326
rect 41020 29222 41076 29260
rect 40572 28754 40740 28756
rect 40572 28702 40574 28754
rect 40626 28702 40740 28754
rect 40572 28700 40740 28702
rect 40572 28690 40628 28700
rect 41020 28644 41076 28654
rect 40012 27918 40014 27970
rect 40066 27918 40068 27970
rect 39116 27804 39284 27860
rect 39116 26962 39172 26974
rect 39116 26910 39118 26962
rect 39170 26910 39172 26962
rect 39116 26516 39172 26910
rect 39228 26852 39284 27804
rect 39228 26786 39284 26796
rect 39116 26450 39172 26460
rect 39228 21812 39284 21822
rect 39228 21718 39284 21756
rect 39228 21028 39284 21038
rect 39228 20934 39284 20972
rect 38444 19854 38446 19906
rect 38498 19854 38500 19906
rect 38332 19012 38388 19022
rect 38332 18340 38388 18956
rect 38332 18274 38388 18284
rect 38444 17780 38500 19854
rect 38780 20132 39060 20188
rect 38668 19234 38724 19246
rect 38668 19182 38670 19234
rect 38722 19182 38724 19234
rect 38668 19012 38724 19182
rect 38668 18946 38724 18956
rect 38444 17724 38724 17780
rect 38220 17556 38276 17566
rect 38556 17556 38612 17566
rect 38220 17554 38612 17556
rect 38220 17502 38222 17554
rect 38274 17502 38558 17554
rect 38610 17502 38612 17554
rect 38220 17500 38612 17502
rect 38220 17490 38276 17500
rect 38556 17490 38612 17500
rect 38668 17332 38724 17724
rect 38668 17266 38724 17276
rect 38332 17220 38388 17230
rect 37996 14306 38052 16716
rect 37996 14254 37998 14306
rect 38050 14254 38052 14306
rect 37100 13694 37102 13746
rect 37154 13694 37156 13746
rect 37100 13682 37156 13694
rect 37996 13748 38052 14254
rect 37996 13682 38052 13692
rect 38108 16884 38164 16894
rect 37436 13524 37492 13534
rect 37324 13522 37492 13524
rect 37324 13470 37438 13522
rect 37490 13470 37492 13522
rect 37324 13468 37492 13470
rect 36820 13132 36932 13188
rect 36988 13132 37156 13188
rect 36764 13122 36820 13132
rect 35868 13010 35924 13020
rect 36092 12964 36148 12974
rect 36876 12964 36932 13132
rect 36988 12964 37044 12974
rect 36092 12962 36708 12964
rect 36092 12910 36094 12962
rect 36146 12910 36708 12962
rect 36092 12908 36708 12910
rect 36876 12962 37044 12964
rect 36876 12910 36990 12962
rect 37042 12910 37044 12962
rect 36876 12908 37044 12910
rect 36092 12898 36148 12908
rect 35756 12628 35812 12638
rect 34860 12012 35028 12068
rect 34972 11788 35028 12012
rect 34524 11442 34580 11452
rect 34748 11732 35028 11788
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 34748 11284 34804 11732
rect 35196 11722 35460 11732
rect 35084 11508 35140 11518
rect 35084 11414 35140 11452
rect 35308 11396 35364 11406
rect 35308 11302 35364 11340
rect 35756 11396 35812 12572
rect 36092 12628 36148 12638
rect 35756 11330 35812 11340
rect 35868 12516 35924 12526
rect 34972 11284 35028 11294
rect 34748 11282 35028 11284
rect 34748 11230 34974 11282
rect 35026 11230 35028 11282
rect 34748 11228 35028 11230
rect 34300 11170 34356 11182
rect 34300 11118 34302 11170
rect 34354 11118 34356 11170
rect 34188 9156 34244 9166
rect 34300 9156 34356 11118
rect 34636 10724 34692 10734
rect 34636 10630 34692 10668
rect 34972 10724 35028 11228
rect 34972 10658 35028 10668
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 34188 9154 34356 9156
rect 34188 9102 34190 9154
rect 34242 9102 34356 9154
rect 34188 9100 34356 9102
rect 34188 9090 34244 9100
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 34412 8372 34468 8382
rect 34412 8278 34468 8316
rect 35756 8260 35812 8270
rect 35756 8166 35812 8204
rect 35644 8148 35700 8158
rect 35644 7698 35700 8092
rect 35644 7646 35646 7698
rect 35698 7646 35700 7698
rect 35644 7634 35700 7646
rect 33964 7532 34132 7588
rect 33068 5282 33124 5292
rect 33516 5348 33572 5358
rect 32732 5234 33012 5236
rect 32732 5182 32734 5234
rect 32786 5182 33012 5234
rect 32732 5180 33012 5182
rect 32732 5170 32788 5180
rect 30156 5012 30212 5022
rect 29932 4340 29988 4350
rect 29708 4338 29988 4340
rect 29708 4286 29934 4338
rect 29986 4286 29988 4338
rect 29708 4284 29988 4286
rect 29708 3668 29764 3678
rect 29596 3666 29764 3668
rect 29596 3614 29710 3666
rect 29762 3614 29764 3666
rect 29596 3612 29764 3614
rect 29708 3602 29764 3612
rect 28476 3502 28478 3554
rect 28530 3502 28532 3554
rect 28476 3490 28532 3502
rect 28140 3332 28196 3342
rect 25788 2818 25844 2828
rect 27916 3330 28196 3332
rect 27916 3278 28142 3330
rect 28194 3278 28196 3330
rect 27916 3276 28196 3278
rect 27916 2882 27972 3276
rect 28140 3266 28196 3276
rect 27916 2830 27918 2882
rect 27970 2830 27972 2882
rect 27916 2818 27972 2830
rect 25340 2706 25396 2716
rect 26796 2772 26852 2782
rect 27132 2772 27188 2782
rect 26852 2770 27188 2772
rect 26852 2718 27134 2770
rect 27186 2718 27188 2770
rect 26852 2716 27188 2718
rect 26796 2678 26852 2716
rect 27132 2706 27188 2716
rect 22428 2606 22430 2658
rect 22482 2606 22484 2658
rect 22428 2594 22484 2606
rect 29932 2660 29988 4284
rect 30156 4338 30212 4956
rect 30940 5012 30996 5022
rect 30940 4562 30996 4956
rect 30940 4510 30942 4562
rect 30994 4510 30996 4562
rect 30940 4498 30996 4510
rect 32508 4452 32564 4462
rect 32508 4358 32564 4396
rect 30156 4286 30158 4338
rect 30210 4286 30212 4338
rect 30156 4274 30212 4286
rect 32284 4338 32340 4350
rect 32284 4286 32286 4338
rect 32338 4286 32340 4338
rect 30492 4114 30548 4126
rect 30492 4062 30494 4114
rect 30546 4062 30548 4114
rect 30492 2770 30548 4062
rect 31836 3442 31892 3454
rect 31836 3390 31838 3442
rect 31890 3390 31892 3442
rect 31836 3388 31892 3390
rect 30716 3332 31892 3388
rect 32284 3388 32340 4286
rect 32956 4340 33012 5180
rect 33516 5234 33572 5292
rect 33516 5182 33518 5234
rect 33570 5182 33572 5234
rect 33516 5170 33572 5182
rect 33628 5012 33684 5022
rect 33068 4340 33124 4350
rect 32956 4338 33124 4340
rect 32956 4286 33070 4338
rect 33122 4286 33124 4338
rect 32956 4284 33124 4286
rect 33068 3668 33124 4284
rect 33628 3780 33684 4956
rect 33740 4898 33796 4910
rect 33740 4846 33742 4898
rect 33794 4846 33796 4898
rect 33740 4564 33796 4846
rect 33740 4498 33796 4508
rect 33852 4452 33908 4462
rect 33852 4358 33908 4396
rect 33964 4116 34020 7532
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 34972 5794 35028 5806
rect 34972 5742 34974 5794
rect 35026 5742 35028 5794
rect 34076 5348 34132 5358
rect 34076 5254 34132 5292
rect 34972 5348 35028 5742
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34972 5282 35028 5292
rect 35644 5348 35700 5358
rect 35644 5254 35700 5292
rect 34300 5236 34356 5246
rect 34300 5142 34356 5180
rect 34748 5236 34804 5246
rect 34748 5142 34804 5180
rect 35868 5234 35924 12460
rect 36092 11788 36148 12572
rect 36652 12066 36708 12908
rect 36988 12898 37044 12908
rect 36652 12014 36654 12066
rect 36706 12014 36708 12066
rect 36652 12002 36708 12014
rect 35980 11732 36148 11788
rect 35980 8708 36036 11732
rect 36316 8932 36372 8942
rect 36316 8838 36372 8876
rect 37100 8932 37156 13132
rect 37324 12178 37380 13468
rect 37436 13458 37492 13468
rect 37772 12852 37828 12862
rect 37548 12850 37828 12852
rect 37548 12798 37774 12850
rect 37826 12798 37828 12850
rect 37548 12796 37828 12798
rect 37548 12402 37604 12796
rect 37772 12786 37828 12796
rect 37548 12350 37550 12402
rect 37602 12350 37604 12402
rect 37548 12338 37604 12350
rect 37324 12126 37326 12178
rect 37378 12126 37380 12178
rect 37324 12114 37380 12126
rect 37660 9826 37716 9838
rect 37660 9774 37662 9826
rect 37714 9774 37716 9826
rect 37100 8866 37156 8876
rect 37324 9604 37380 9614
rect 37660 9604 37716 9774
rect 37324 9602 37716 9604
rect 37324 9550 37326 9602
rect 37378 9550 37716 9602
rect 37324 9548 37716 9550
rect 37324 9156 37380 9548
rect 35980 8652 36148 8708
rect 35868 5182 35870 5234
rect 35922 5182 35924 5234
rect 35868 5012 35924 5182
rect 35868 4946 35924 4956
rect 35980 8484 36036 8494
rect 35980 8148 36036 8428
rect 35980 7474 36036 8092
rect 35980 7422 35982 7474
rect 36034 7422 36036 7474
rect 35308 4900 35364 4910
rect 35308 4898 35588 4900
rect 35308 4846 35310 4898
rect 35362 4846 35588 4898
rect 35308 4844 35588 4846
rect 35308 4834 35364 4844
rect 33740 3780 33796 3790
rect 33628 3724 33740 3780
rect 33740 3686 33796 3724
rect 32620 3666 33124 3668
rect 32620 3614 33070 3666
rect 33122 3614 33124 3666
rect 32620 3612 33124 3614
rect 32620 3554 32676 3612
rect 33068 3602 33124 3612
rect 33964 3666 34020 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 33964 3614 33966 3666
rect 34018 3614 34020 3666
rect 33964 3602 34020 3614
rect 34412 3780 34468 3790
rect 34412 3666 34468 3724
rect 34412 3614 34414 3666
rect 34466 3614 34468 3666
rect 34412 3602 34468 3614
rect 32620 3502 32622 3554
rect 32674 3502 32676 3554
rect 32620 3490 32676 3502
rect 35532 3554 35588 4844
rect 35980 4452 36036 7422
rect 35980 4386 36036 4396
rect 36092 5236 36148 8652
rect 37324 8484 37380 9100
rect 37324 8418 37380 8428
rect 37548 8932 37604 8942
rect 37548 8370 37604 8876
rect 37548 8318 37550 8370
rect 37602 8318 37604 8370
rect 37548 8306 37604 8318
rect 36204 8258 36260 8270
rect 36204 8206 36206 8258
rect 36258 8206 36260 8258
rect 36204 8148 36260 8206
rect 36204 8082 36260 8092
rect 36316 8260 36372 8270
rect 36316 5236 36372 8204
rect 37324 8260 37380 8270
rect 37380 8204 37492 8260
rect 37324 8166 37380 8204
rect 36988 8148 37044 8158
rect 36988 8054 37044 8092
rect 36428 8036 36484 8046
rect 36428 8034 36820 8036
rect 36428 7982 36430 8034
rect 36482 7982 36820 8034
rect 36428 7980 36820 7982
rect 36428 7970 36484 7980
rect 36764 7586 36820 7980
rect 36764 7534 36766 7586
rect 36818 7534 36820 7586
rect 36764 7522 36820 7534
rect 37212 7028 37268 7038
rect 36428 5236 36484 5246
rect 36316 5234 36484 5236
rect 36316 5182 36430 5234
rect 36482 5182 36484 5234
rect 36316 5180 36484 5182
rect 35532 3502 35534 3554
rect 35586 3502 35588 3554
rect 35532 3490 35588 3502
rect 35756 4228 35812 4238
rect 33404 3442 33460 3454
rect 33404 3390 33406 3442
rect 33458 3390 33460 3442
rect 33404 3388 33460 3390
rect 32284 3332 33460 3388
rect 35756 3442 35812 4172
rect 35980 4228 36036 4238
rect 36092 4228 36148 5180
rect 36428 5170 36484 5180
rect 37212 5234 37268 6972
rect 37436 5346 37492 8204
rect 38108 7028 38164 16828
rect 38332 16324 38388 17164
rect 38332 14644 38388 16268
rect 38444 17108 38500 17118
rect 38444 15314 38500 17052
rect 38780 17106 38836 20132
rect 38892 20020 38948 20030
rect 39228 20020 39284 20030
rect 38948 20018 39284 20020
rect 38948 19966 39230 20018
rect 39282 19966 39284 20018
rect 38948 19964 39284 19966
rect 38892 19926 38948 19964
rect 39228 19954 39284 19964
rect 39116 18340 39172 18350
rect 38892 18338 39172 18340
rect 38892 18286 39118 18338
rect 39170 18286 39172 18338
rect 38892 18284 39172 18286
rect 38892 17554 38948 18284
rect 39116 18274 39172 18284
rect 39340 18004 39396 27916
rect 40012 27906 40068 27918
rect 40348 27970 40404 27982
rect 40348 27918 40350 27970
rect 40402 27918 40404 27970
rect 39900 27860 39956 27870
rect 39676 27804 39900 27860
rect 39676 27746 39732 27804
rect 39676 27694 39678 27746
rect 39730 27694 39732 27746
rect 39676 27682 39732 27694
rect 39900 27074 39956 27804
rect 40348 27636 40404 27918
rect 40348 27570 40404 27580
rect 41020 27860 41076 28588
rect 39900 27022 39902 27074
rect 39954 27022 39956 27074
rect 39900 27010 39956 27022
rect 40572 27186 40628 27198
rect 40572 27134 40574 27186
rect 40626 27134 40628 27186
rect 40236 26962 40292 26974
rect 40236 26910 40238 26962
rect 40290 26910 40292 26962
rect 39900 26852 39956 26862
rect 40236 26852 40292 26910
rect 40460 26964 40516 26974
rect 40460 26870 40516 26908
rect 39956 26796 40292 26852
rect 39900 26514 39956 26796
rect 39900 26462 39902 26514
rect 39954 26462 39956 26514
rect 39900 26450 39956 26462
rect 40572 24052 40628 27134
rect 41020 24948 41076 27804
rect 41132 26964 41188 29374
rect 41244 29204 41300 29596
rect 41580 29428 41636 29438
rect 41580 29426 41748 29428
rect 41580 29374 41582 29426
rect 41634 29374 41748 29426
rect 41580 29372 41748 29374
rect 41580 29362 41636 29372
rect 41244 29138 41300 29148
rect 41580 29204 41636 29214
rect 41356 28644 41412 28654
rect 41356 28550 41412 28588
rect 41580 28308 41636 29148
rect 41692 28754 41748 29372
rect 41692 28702 41694 28754
rect 41746 28702 41748 28754
rect 41692 28690 41748 28702
rect 41804 28644 41860 29820
rect 41916 29652 41972 29662
rect 42028 29652 42084 31164
rect 41916 29650 42028 29652
rect 41916 29598 41918 29650
rect 41970 29598 42028 29650
rect 41916 29596 42028 29598
rect 41916 29586 41972 29596
rect 42028 29558 42084 29596
rect 42252 30324 42308 30334
rect 42252 28756 42308 30268
rect 42476 30212 42532 30222
rect 42476 30210 42644 30212
rect 42476 30158 42478 30210
rect 42530 30158 42644 30210
rect 42476 30156 42644 30158
rect 42476 30146 42532 30156
rect 41804 28642 41972 28644
rect 41804 28590 41806 28642
rect 41858 28590 41972 28642
rect 41804 28588 41972 28590
rect 41804 28578 41860 28588
rect 41916 28308 41972 28588
rect 42252 28642 42308 28700
rect 42252 28590 42254 28642
rect 42306 28590 42308 28642
rect 42252 28578 42308 28590
rect 42364 29652 42420 29662
rect 42364 28642 42420 29596
rect 42364 28590 42366 28642
rect 42418 28590 42420 28642
rect 42364 28578 42420 28590
rect 41580 28252 41860 28308
rect 41692 27746 41748 27758
rect 41692 27694 41694 27746
rect 41746 27694 41748 27746
rect 41692 27636 41748 27694
rect 41692 27570 41748 27580
rect 41132 26898 41188 26908
rect 41020 24882 41076 24892
rect 41468 24948 41524 24958
rect 40684 24052 40740 24062
rect 40572 24050 40740 24052
rect 40572 23998 40686 24050
rect 40738 23998 40740 24050
rect 40572 23996 40740 23998
rect 40684 23986 40740 23996
rect 41468 23938 41524 24892
rect 41468 23886 41470 23938
rect 41522 23886 41524 23938
rect 41468 23874 41524 23886
rect 40348 23604 40404 23614
rect 40348 23378 40404 23548
rect 40348 23326 40350 23378
rect 40402 23326 40404 23378
rect 40348 23314 40404 23326
rect 40908 23044 40964 23054
rect 40908 22950 40964 22988
rect 39900 22484 39956 22494
rect 40348 22484 40404 22494
rect 39900 22482 40404 22484
rect 39900 22430 39902 22482
rect 39954 22430 40350 22482
rect 40402 22430 40404 22482
rect 39900 22428 40404 22430
rect 39900 22418 39956 22428
rect 40348 22418 40404 22428
rect 40236 22148 40292 22158
rect 39452 22146 40292 22148
rect 39452 22094 40238 22146
rect 40290 22094 40292 22146
rect 39452 22092 40292 22094
rect 39452 20802 39508 22092
rect 40236 22082 40292 22092
rect 41804 21588 41860 28252
rect 41916 28242 41972 28252
rect 42028 28418 42084 28430
rect 42028 28366 42030 28418
rect 42082 28366 42084 28418
rect 42028 24948 42084 28366
rect 41916 24892 42084 24948
rect 41916 24500 41972 24892
rect 42252 24836 42308 24846
rect 42252 24834 42532 24836
rect 42252 24782 42254 24834
rect 42306 24782 42532 24834
rect 42252 24780 42532 24782
rect 42252 24770 42308 24780
rect 42028 24724 42084 24734
rect 42028 24722 42196 24724
rect 42028 24670 42030 24722
rect 42082 24670 42196 24722
rect 42028 24668 42196 24670
rect 42028 24658 42084 24668
rect 41916 24444 42084 24500
rect 41916 24164 41972 24174
rect 41916 24050 41972 24108
rect 41916 23998 41918 24050
rect 41970 23998 41972 24050
rect 41916 23986 41972 23998
rect 42028 23044 42084 24444
rect 42140 24164 42196 24668
rect 42252 24164 42308 24174
rect 42140 24162 42308 24164
rect 42140 24110 42254 24162
rect 42306 24110 42308 24162
rect 42140 24108 42308 24110
rect 42252 24098 42308 24108
rect 42476 23828 42532 24780
rect 42588 24388 42644 30156
rect 42700 27188 42756 31726
rect 43148 31778 43204 31790
rect 43148 31726 43150 31778
rect 43202 31726 43204 31778
rect 43148 31220 43204 31726
rect 43148 31154 43204 31164
rect 43036 30994 43092 31006
rect 43036 30942 43038 30994
rect 43090 30942 43092 30994
rect 42812 30210 42868 30222
rect 42812 30158 42814 30210
rect 42866 30158 42868 30210
rect 42812 29652 42868 30158
rect 42868 29596 42980 29652
rect 42812 29586 42868 29596
rect 42924 29426 42980 29596
rect 43036 29650 43092 30942
rect 43372 30884 43428 31892
rect 43596 30994 43652 32060
rect 43596 30942 43598 30994
rect 43650 30942 43652 30994
rect 43596 30930 43652 30942
rect 43708 31554 43764 31566
rect 43708 31502 43710 31554
rect 43762 31502 43764 31554
rect 43372 30790 43428 30828
rect 43148 30436 43204 30446
rect 43148 30342 43204 30380
rect 43036 29598 43038 29650
rect 43090 29598 43092 29650
rect 43036 29586 43092 29598
rect 42924 29374 42926 29426
rect 42978 29374 42980 29426
rect 42924 29362 42980 29374
rect 43148 29538 43204 29550
rect 43148 29486 43150 29538
rect 43202 29486 43204 29538
rect 42924 28756 42980 28766
rect 43148 28756 43204 29486
rect 43596 29426 43652 29438
rect 43596 29374 43598 29426
rect 43650 29374 43652 29426
rect 43372 28756 43428 28766
rect 42980 28754 43428 28756
rect 42980 28702 43374 28754
rect 43426 28702 43428 28754
rect 42980 28700 43428 28702
rect 42924 28662 42980 28700
rect 43372 28690 43428 28700
rect 42700 27122 42756 27132
rect 43036 27748 43092 27758
rect 43036 27186 43092 27692
rect 43036 27134 43038 27186
rect 43090 27134 43092 27186
rect 43036 27076 43092 27134
rect 43372 27748 43428 27758
rect 43372 27188 43428 27692
rect 43596 27300 43652 29374
rect 43708 29428 43764 31502
rect 43932 31106 43988 32956
rect 44268 32564 44324 32574
rect 44268 32004 44324 32508
rect 44268 31890 44324 31948
rect 44268 31838 44270 31890
rect 44322 31838 44324 31890
rect 44268 31826 44324 31838
rect 43932 31054 43934 31106
rect 43986 31054 43988 31106
rect 43932 31042 43988 31054
rect 44380 30994 44436 31006
rect 44380 30942 44382 30994
rect 44434 30942 44436 30994
rect 44380 30436 44436 30942
rect 44716 30882 44772 37212
rect 45164 37202 45220 37212
rect 45724 37268 45780 37278
rect 45724 37266 45892 37268
rect 45724 37214 45726 37266
rect 45778 37214 45892 37266
rect 45724 37212 45892 37214
rect 45724 37202 45780 37212
rect 45276 37156 45332 37166
rect 45276 36484 45332 37100
rect 45612 37044 45668 37054
rect 45612 36950 45668 36988
rect 44940 36482 45332 36484
rect 44940 36430 45278 36482
rect 45330 36430 45332 36482
rect 44940 36428 45332 36430
rect 44940 35026 44996 36428
rect 45276 36418 45332 36428
rect 45836 35588 45892 37212
rect 45948 36596 46004 36606
rect 46060 36596 46116 39342
rect 45948 36594 46116 36596
rect 45948 36542 45950 36594
rect 46002 36542 46116 36594
rect 45948 36540 46116 36542
rect 48076 36596 48132 36606
rect 45948 36530 46004 36540
rect 48076 36502 48132 36540
rect 46172 35588 46228 35598
rect 45836 35586 46228 35588
rect 45836 35534 46174 35586
rect 46226 35534 46228 35586
rect 45836 35532 46228 35534
rect 46172 35522 46228 35532
rect 44940 34974 44942 35026
rect 44994 34974 44996 35026
rect 44940 34962 44996 34974
rect 44828 33684 44884 33694
rect 44828 33572 44884 33628
rect 44828 33570 44996 33572
rect 44828 33518 44830 33570
rect 44882 33518 44996 33570
rect 44828 33516 44996 33518
rect 44828 33506 44884 33516
rect 44828 32004 44884 32014
rect 44828 31778 44884 31948
rect 44828 31726 44830 31778
rect 44882 31726 44884 31778
rect 44828 31714 44884 31726
rect 44716 30830 44718 30882
rect 44770 30830 44772 30882
rect 44716 30818 44772 30830
rect 44380 30370 44436 30380
rect 44940 30212 44996 33516
rect 45164 33460 45220 33470
rect 45164 33458 45332 33460
rect 45164 33406 45166 33458
rect 45218 33406 45332 33458
rect 45164 33404 45332 33406
rect 45164 33394 45220 33404
rect 45052 33122 45108 33134
rect 45052 33070 45054 33122
rect 45106 33070 45108 33122
rect 45052 32116 45108 33070
rect 45052 32050 45108 32060
rect 45276 31948 45332 33404
rect 46396 32564 46452 32574
rect 45948 32562 46452 32564
rect 45948 32510 46398 32562
rect 46450 32510 46452 32562
rect 45948 32508 46452 32510
rect 45948 32450 46004 32508
rect 46396 32498 46452 32508
rect 45948 32398 45950 32450
rect 46002 32398 46004 32450
rect 45948 32386 46004 32398
rect 46284 32338 46340 32350
rect 46284 32286 46286 32338
rect 46338 32286 46340 32338
rect 46284 32116 46340 32286
rect 46284 32050 46340 32060
rect 45276 31892 45668 31948
rect 45612 31890 45668 31892
rect 45612 31838 45614 31890
rect 45666 31838 45668 31890
rect 45612 31826 45668 31838
rect 46396 31892 46452 31902
rect 46396 31106 46452 31836
rect 47740 31892 47796 31902
rect 47740 31798 47796 31836
rect 46396 31054 46398 31106
rect 46450 31054 46452 31106
rect 46396 31042 46452 31054
rect 45500 30996 45556 31006
rect 45052 30884 45108 30894
rect 45052 30790 45108 30828
rect 44940 30210 45220 30212
rect 44940 30158 44942 30210
rect 44994 30158 45220 30210
rect 44940 30156 45220 30158
rect 44940 30146 44996 30156
rect 45164 29538 45220 30156
rect 45164 29486 45166 29538
rect 45218 29486 45220 29538
rect 45164 29474 45220 29486
rect 44156 29428 44212 29438
rect 44828 29428 44884 29438
rect 43708 29426 44884 29428
rect 43708 29374 44158 29426
rect 44210 29374 44830 29426
rect 44882 29374 44884 29426
rect 43708 29372 44884 29374
rect 43820 28754 43876 29372
rect 44156 29362 44212 29372
rect 44828 29362 44884 29372
rect 45500 29426 45556 30940
rect 46284 30996 46340 31006
rect 46284 30902 46340 30940
rect 45500 29374 45502 29426
rect 45554 29374 45556 29426
rect 45500 29362 45556 29374
rect 45500 29204 45556 29214
rect 45500 29202 45780 29204
rect 45500 29150 45502 29202
rect 45554 29150 45780 29202
rect 45500 29148 45780 29150
rect 45500 29138 45556 29148
rect 43820 28702 43822 28754
rect 43874 28702 43876 28754
rect 43820 28308 43876 28702
rect 45724 28754 45780 29148
rect 47852 28756 47908 28766
rect 45724 28702 45726 28754
rect 45778 28702 45780 28754
rect 45724 28690 45780 28702
rect 47292 28754 47908 28756
rect 47292 28702 47854 28754
rect 47906 28702 47908 28754
rect 47292 28700 47908 28702
rect 44268 28644 44324 28654
rect 44268 28550 44324 28588
rect 44940 28644 44996 28654
rect 44940 28550 44996 28588
rect 43820 28242 43876 28252
rect 47292 27970 47348 28700
rect 47852 28690 47908 28700
rect 47292 27918 47294 27970
rect 47346 27918 47348 27970
rect 47292 27906 47348 27918
rect 43820 27748 43876 27758
rect 43820 27654 43876 27692
rect 47180 27634 47236 27646
rect 47180 27582 47182 27634
rect 47234 27582 47236 27634
rect 43596 27234 43652 27244
rect 45388 27300 45444 27310
rect 43372 27094 43428 27132
rect 43036 27010 43092 27020
rect 43596 27076 43652 27086
rect 43596 26982 43652 27020
rect 44268 27076 44324 27086
rect 43932 26852 43988 26862
rect 43932 26850 44100 26852
rect 43932 26798 43934 26850
rect 43986 26798 44100 26850
rect 43932 26796 44100 26798
rect 43932 26786 43988 26796
rect 43820 26402 43876 26414
rect 43820 26350 43822 26402
rect 43874 26350 43876 26402
rect 42812 24948 42868 24958
rect 42812 24854 42868 24892
rect 43260 24948 43316 24958
rect 43260 24724 43316 24892
rect 43820 24836 43876 26350
rect 44044 26290 44100 26796
rect 44044 26238 44046 26290
rect 44098 26238 44100 26290
rect 44044 26226 44100 26238
rect 44268 25282 44324 27020
rect 45388 25620 45444 27244
rect 47180 26964 47236 27582
rect 47180 26898 47236 26908
rect 45388 25618 46116 25620
rect 45388 25566 45390 25618
rect 45442 25566 46116 25618
rect 45388 25564 46116 25566
rect 45388 25554 45444 25564
rect 45164 25506 45220 25518
rect 45164 25454 45166 25506
rect 45218 25454 45220 25506
rect 44268 25230 44270 25282
rect 44322 25230 44324 25282
rect 44268 25172 44324 25230
rect 44828 25284 44884 25294
rect 44828 25282 44996 25284
rect 44828 25230 44830 25282
rect 44882 25230 44996 25282
rect 44828 25228 44996 25230
rect 44828 25218 44884 25228
rect 43932 24836 43988 24846
rect 43820 24834 43988 24836
rect 43820 24782 43934 24834
rect 43986 24782 43988 24834
rect 43820 24780 43988 24782
rect 43932 24770 43988 24780
rect 43260 24722 43540 24724
rect 43260 24670 43262 24722
rect 43314 24670 43540 24722
rect 43260 24668 43540 24670
rect 43260 24658 43316 24668
rect 42588 24332 42868 24388
rect 42588 24164 42644 24174
rect 42588 24070 42644 24108
rect 42812 24052 42868 24332
rect 42812 23958 42868 23996
rect 42476 23772 43092 23828
rect 43036 23266 43092 23772
rect 43484 23548 43540 24668
rect 43932 24164 43988 24174
rect 44268 24164 44324 25116
rect 43988 24108 44324 24164
rect 43708 23940 43764 23950
rect 43708 23548 43764 23884
rect 43484 23492 43764 23548
rect 43036 23214 43038 23266
rect 43090 23214 43092 23266
rect 43036 23202 43092 23214
rect 43708 23156 43764 23492
rect 43708 23062 43764 23100
rect 42084 22988 42308 23044
rect 42028 22978 42084 22988
rect 42252 21698 42308 22988
rect 42252 21646 42254 21698
rect 42306 21646 42308 21698
rect 42252 21634 42308 21646
rect 41916 21588 41972 21598
rect 41804 21532 41916 21588
rect 41916 21494 41972 21532
rect 42476 21588 42532 21598
rect 42476 21494 42532 21532
rect 39452 20750 39454 20802
rect 39506 20750 39508 20802
rect 39452 20242 39508 20750
rect 39452 20190 39454 20242
rect 39506 20190 39508 20242
rect 39452 20178 39508 20190
rect 40012 21476 40068 21486
rect 39452 19906 39508 19918
rect 39452 19854 39454 19906
rect 39506 19854 39508 19906
rect 39452 19346 39508 19854
rect 39452 19294 39454 19346
rect 39506 19294 39508 19346
rect 39452 19282 39508 19294
rect 39788 18450 39844 18462
rect 39788 18398 39790 18450
rect 39842 18398 39844 18450
rect 39788 18340 39844 18398
rect 39788 18274 39844 18284
rect 40012 18004 40068 21420
rect 42812 21362 42868 21374
rect 42812 21310 42814 21362
rect 42866 21310 42868 21362
rect 40236 20914 40292 20926
rect 40236 20862 40238 20914
rect 40290 20862 40292 20914
rect 40124 20802 40180 20814
rect 40124 20750 40126 20802
rect 40178 20750 40180 20802
rect 40124 20356 40180 20750
rect 40124 20290 40180 20300
rect 38892 17502 38894 17554
rect 38946 17502 38948 17554
rect 38892 17490 38948 17502
rect 39228 17948 39396 18004
rect 39788 17948 40068 18004
rect 38780 17054 38782 17106
rect 38834 17054 38836 17106
rect 38780 17042 38836 17054
rect 38444 15262 38446 15314
rect 38498 15262 38500 15314
rect 38444 14868 38500 15262
rect 38556 16882 38612 16894
rect 38556 16830 38558 16882
rect 38610 16830 38612 16882
rect 38556 15204 38612 16830
rect 38892 16884 38948 16894
rect 38892 16790 38948 16828
rect 39228 15986 39284 17948
rect 39340 17666 39396 17678
rect 39340 17614 39342 17666
rect 39394 17614 39396 17666
rect 39340 17332 39396 17614
rect 39340 17266 39396 17276
rect 39676 17554 39732 17566
rect 39676 17502 39678 17554
rect 39730 17502 39732 17554
rect 39676 17108 39732 17502
rect 39340 17052 39732 17108
rect 39788 17108 39844 17948
rect 39340 16098 39396 17052
rect 39340 16046 39342 16098
rect 39394 16046 39396 16098
rect 39340 16034 39396 16046
rect 39564 16884 39620 16894
rect 39228 15934 39230 15986
rect 39282 15934 39284 15986
rect 39228 15922 39284 15934
rect 38556 15148 38724 15204
rect 38444 14802 38500 14812
rect 38444 14644 38500 14654
rect 38332 14642 38500 14644
rect 38332 14590 38446 14642
rect 38498 14590 38500 14642
rect 38332 14588 38500 14590
rect 38444 13748 38500 14588
rect 38668 14084 38724 15148
rect 39004 14532 39060 14542
rect 39004 14438 39060 14476
rect 39452 14532 39508 14542
rect 39452 14438 39508 14476
rect 38668 14028 39060 14084
rect 39004 13858 39060 14028
rect 39004 13806 39006 13858
rect 39058 13806 39060 13858
rect 39004 13794 39060 13806
rect 38668 13748 38724 13758
rect 38444 13746 38724 13748
rect 38444 13694 38670 13746
rect 38722 13694 38724 13746
rect 38444 13692 38724 13694
rect 38668 13682 38724 13692
rect 39116 13746 39172 13758
rect 39116 13694 39118 13746
rect 39170 13694 39172 13746
rect 38556 10836 38612 10846
rect 39116 10836 39172 13694
rect 39564 13076 39620 16828
rect 39788 16884 39844 17052
rect 39788 16790 39844 16828
rect 39900 17668 39956 17678
rect 39788 16212 39844 16222
rect 39676 16098 39732 16110
rect 39676 16046 39678 16098
rect 39730 16046 39732 16098
rect 39676 15988 39732 16046
rect 39676 15922 39732 15932
rect 39788 15538 39844 16156
rect 39788 15486 39790 15538
rect 39842 15486 39844 15538
rect 39788 15428 39844 15486
rect 39788 15362 39844 15372
rect 39900 14420 39956 17612
rect 40236 17108 40292 20862
rect 42812 20802 42868 21310
rect 42812 20750 42814 20802
rect 42866 20750 42868 20802
rect 42812 20738 42868 20750
rect 42476 20578 42532 20590
rect 42476 20526 42478 20578
rect 42530 20526 42532 20578
rect 40348 20356 40404 20366
rect 40348 18452 40404 20300
rect 42476 20130 42532 20526
rect 42476 20078 42478 20130
rect 42530 20078 42532 20130
rect 42476 20066 42532 20078
rect 41804 20018 41860 20030
rect 41804 19966 41806 20018
rect 41858 19966 41860 20018
rect 41356 19908 41412 19918
rect 41804 19908 41860 19966
rect 41356 19906 41860 19908
rect 41356 19854 41358 19906
rect 41410 19854 41860 19906
rect 41356 19852 41860 19854
rect 41356 19842 41412 19852
rect 41580 19348 41636 19358
rect 41020 19346 41636 19348
rect 41020 19294 41582 19346
rect 41634 19294 41636 19346
rect 41020 19292 41636 19294
rect 41020 18562 41076 19292
rect 41580 19282 41636 19292
rect 41020 18510 41022 18562
rect 41074 18510 41076 18562
rect 41020 18498 41076 18510
rect 40348 18450 40628 18452
rect 40348 18398 40350 18450
rect 40402 18398 40628 18450
rect 40348 18396 40628 18398
rect 40348 18386 40404 18396
rect 40572 17666 40628 18396
rect 40572 17614 40574 17666
rect 40626 17614 40628 17666
rect 40572 17602 40628 17614
rect 40908 18226 40964 18238
rect 40908 18174 40910 18226
rect 40962 18174 40964 18226
rect 40908 17668 40964 18174
rect 41804 18116 41860 19852
rect 43820 19348 43876 19358
rect 43932 19348 43988 24108
rect 44268 23940 44324 23950
rect 44828 23940 44884 23950
rect 44324 23938 44884 23940
rect 44324 23886 44830 23938
rect 44882 23886 44884 23938
rect 44324 23884 44884 23886
rect 44268 23846 44324 23884
rect 44828 23874 44884 23884
rect 44940 23154 44996 25228
rect 45164 25172 45220 25454
rect 45164 25106 45220 25116
rect 46060 24610 46116 25564
rect 46060 24558 46062 24610
rect 46114 24558 46116 24610
rect 46060 24546 46116 24558
rect 47740 24052 47796 24062
rect 47740 23958 47796 23996
rect 45612 23828 45668 23838
rect 45164 23826 45668 23828
rect 45164 23774 45614 23826
rect 45666 23774 45668 23826
rect 45164 23772 45668 23774
rect 45164 23378 45220 23772
rect 45612 23762 45668 23772
rect 45164 23326 45166 23378
rect 45218 23326 45220 23378
rect 45164 23314 45220 23326
rect 44940 23102 44942 23154
rect 44994 23102 44996 23154
rect 44940 23090 44996 23102
rect 44604 19908 44660 19918
rect 43820 19346 43932 19348
rect 43820 19294 43822 19346
rect 43874 19294 43932 19346
rect 43820 19292 43932 19294
rect 43820 19282 43876 19292
rect 43932 19254 43988 19292
rect 44380 19852 44604 19908
rect 44660 19852 44884 19908
rect 44380 19346 44436 19852
rect 44604 19814 44660 19852
rect 44380 19294 44382 19346
rect 44434 19294 44436 19346
rect 44380 19282 44436 19294
rect 44828 19346 44884 19852
rect 45052 19458 45108 19470
rect 45052 19406 45054 19458
rect 45106 19406 45108 19458
rect 44828 19294 44830 19346
rect 44882 19294 44884 19346
rect 44828 19282 44884 19294
rect 44940 19348 44996 19358
rect 45052 19348 45108 19406
rect 44996 19292 45108 19348
rect 44940 19282 44996 19292
rect 44492 19012 44548 19022
rect 44156 18562 44212 18574
rect 44156 18510 44158 18562
rect 44210 18510 44212 18562
rect 41804 18060 42084 18116
rect 41916 17892 41972 17902
rect 40908 17602 40964 17612
rect 41020 17668 41076 17678
rect 41020 17666 41188 17668
rect 41020 17614 41022 17666
rect 41074 17614 41188 17666
rect 41020 17612 41188 17614
rect 41020 17602 41076 17612
rect 40236 17042 40292 17052
rect 40460 16884 40516 16894
rect 40460 16098 40516 16828
rect 40460 16046 40462 16098
rect 40514 16046 40516 16098
rect 40460 16034 40516 16046
rect 41020 16770 41076 16782
rect 41020 16718 41022 16770
rect 41074 16718 41076 16770
rect 41020 16658 41076 16718
rect 41020 16606 41022 16658
rect 41074 16606 41076 16658
rect 40012 15428 40068 15438
rect 40012 15334 40068 15372
rect 40124 15428 40180 15438
rect 41020 15428 41076 16606
rect 41132 16324 41188 17612
rect 41468 17442 41524 17454
rect 41468 17390 41470 17442
rect 41522 17390 41524 17442
rect 41468 17332 41524 17390
rect 41468 17266 41524 17276
rect 41916 17108 41972 17836
rect 41916 17014 41972 17052
rect 41804 16882 41860 16894
rect 41804 16830 41806 16882
rect 41858 16830 41860 16882
rect 41468 16772 41524 16782
rect 41804 16772 41860 16830
rect 41468 16770 41860 16772
rect 41468 16718 41470 16770
rect 41522 16718 41860 16770
rect 41468 16716 41860 16718
rect 42028 16772 42084 18060
rect 44156 16994 44212 18510
rect 44492 18450 44548 18956
rect 45388 19012 45444 19022
rect 45388 18918 45444 18956
rect 44492 18398 44494 18450
rect 44546 18398 44548 18450
rect 44492 18386 44548 18398
rect 45276 17892 45332 17902
rect 45276 17798 45332 17836
rect 45388 17556 45444 17566
rect 45388 17554 46340 17556
rect 45388 17502 45390 17554
rect 45442 17502 46340 17554
rect 45388 17500 46340 17502
rect 45388 17490 45444 17500
rect 44156 16942 44158 16994
rect 44210 16942 44212 16994
rect 44156 16930 44212 16942
rect 42140 16884 42196 16894
rect 42140 16882 42420 16884
rect 42140 16830 42142 16882
rect 42194 16830 42420 16882
rect 42140 16828 42420 16830
rect 42140 16818 42196 16828
rect 41468 16658 41524 16716
rect 41468 16606 41470 16658
rect 41522 16606 41524 16658
rect 41468 16594 41524 16606
rect 41132 15538 41188 16268
rect 41468 16100 41524 16110
rect 41468 16006 41524 16044
rect 41580 15988 41636 15998
rect 41580 15986 41972 15988
rect 41580 15934 41582 15986
rect 41634 15934 41972 15986
rect 41580 15932 41972 15934
rect 41580 15922 41636 15932
rect 41132 15486 41134 15538
rect 41186 15486 41188 15538
rect 41132 15474 41188 15486
rect 40124 15426 40292 15428
rect 40124 15374 40126 15426
rect 40178 15374 40292 15426
rect 40124 15372 40292 15374
rect 40124 15362 40180 15372
rect 40124 15090 40180 15102
rect 40124 15038 40126 15090
rect 40178 15038 40180 15090
rect 40124 14642 40180 15038
rect 40124 14590 40126 14642
rect 40178 14590 40180 14642
rect 40124 14578 40180 14590
rect 39900 14364 40180 14420
rect 39900 13748 39956 13758
rect 39900 13654 39956 13692
rect 39900 13076 39956 13086
rect 39564 13074 39956 13076
rect 39564 13022 39902 13074
rect 39954 13022 39956 13074
rect 39564 13020 39956 13022
rect 39900 13010 39956 13020
rect 39452 11396 39508 11406
rect 39452 11302 39508 11340
rect 38556 10834 38948 10836
rect 38556 10782 38558 10834
rect 38610 10782 38948 10834
rect 38556 10780 38948 10782
rect 38556 10724 38612 10780
rect 38556 10658 38612 10668
rect 38892 10724 38948 10780
rect 39116 10742 39172 10780
rect 39564 11282 39620 11294
rect 39564 11230 39566 11282
rect 39618 11230 39620 11282
rect 38892 10630 38948 10668
rect 39004 10498 39060 10510
rect 39004 10446 39006 10498
rect 39058 10446 39060 10498
rect 39004 10164 39060 10446
rect 38444 10108 39060 10164
rect 38444 9938 38500 10108
rect 39564 10052 39620 11230
rect 40012 11170 40068 11182
rect 40012 11118 40014 11170
rect 40066 11118 40068 11170
rect 39788 10724 39844 10734
rect 40012 10724 40068 11118
rect 39844 10668 40068 10724
rect 39788 10630 39844 10668
rect 40124 10610 40180 14364
rect 40236 14308 40292 15372
rect 41020 15334 41076 15372
rect 41356 15316 41412 15326
rect 41580 15316 41636 15326
rect 41356 15314 41524 15316
rect 41356 15262 41358 15314
rect 41410 15262 41524 15314
rect 41356 15260 41524 15262
rect 41356 15250 41412 15260
rect 40236 13634 40292 14252
rect 40908 14532 40964 14542
rect 40908 13748 40964 14476
rect 41468 14308 41524 15260
rect 41580 14532 41636 15260
rect 41916 15092 41972 15932
rect 42028 15874 42084 16716
rect 42028 15822 42030 15874
rect 42082 15822 42084 15874
rect 42028 15316 42084 15822
rect 42364 15426 42420 16828
rect 43484 16882 43540 16894
rect 43484 16830 43486 16882
rect 43538 16830 43540 16882
rect 43036 16772 43092 16782
rect 43036 16678 43092 16716
rect 43484 16772 43540 16830
rect 43484 16706 43540 16716
rect 46284 16770 46340 17500
rect 46284 16718 46286 16770
rect 46338 16718 46340 16770
rect 46284 16706 46340 16718
rect 43708 16324 43764 16334
rect 43708 16230 43764 16268
rect 43820 15988 43876 15998
rect 43820 15986 44548 15988
rect 43820 15934 43822 15986
rect 43874 15934 44548 15986
rect 43820 15932 44548 15934
rect 43820 15922 43876 15932
rect 42364 15374 42366 15426
rect 42418 15374 42420 15426
rect 42364 15362 42420 15374
rect 42028 15250 42084 15260
rect 44492 15202 44548 15932
rect 44492 15150 44494 15202
rect 44546 15150 44548 15202
rect 44492 15138 44548 15150
rect 41916 15036 42308 15092
rect 42252 14642 42308 15036
rect 42252 14590 42254 14642
rect 42306 14590 42308 14642
rect 42252 14578 42308 14590
rect 41580 14466 41636 14476
rect 42924 14420 42980 14430
rect 42924 14326 42980 14364
rect 43820 14420 43876 14430
rect 42812 14308 42868 14318
rect 41468 14252 41748 14308
rect 41692 13858 41748 14252
rect 42812 14214 42868 14252
rect 41692 13806 41694 13858
rect 41746 13806 41748 13858
rect 41692 13794 41748 13806
rect 40236 13582 40238 13634
rect 40290 13582 40292 13634
rect 40236 13570 40292 13582
rect 40572 13746 40964 13748
rect 40572 13694 40910 13746
rect 40962 13694 40964 13746
rect 40572 13692 40964 13694
rect 40572 13074 40628 13692
rect 40908 13682 40964 13692
rect 43820 13634 43876 14364
rect 43820 13582 43822 13634
rect 43874 13582 43876 13634
rect 43820 13570 43876 13582
rect 40572 13022 40574 13074
rect 40626 13022 40628 13074
rect 40572 13010 40628 13022
rect 40908 10836 40964 10846
rect 40908 10742 40964 10780
rect 40124 10558 40126 10610
rect 40178 10558 40180 10610
rect 40124 10546 40180 10558
rect 41020 10498 41076 10510
rect 41020 10446 41022 10498
rect 41074 10446 41076 10498
rect 39564 9986 39620 9996
rect 40124 10386 40180 10398
rect 40124 10334 40126 10386
rect 40178 10334 40180 10386
rect 38444 9886 38446 9938
rect 38498 9886 38500 9938
rect 38444 9874 38500 9886
rect 40124 9940 40180 10334
rect 40124 9874 40180 9884
rect 40572 10052 40628 10062
rect 40572 9938 40628 9996
rect 40572 9886 40574 9938
rect 40626 9886 40628 9938
rect 40572 9874 40628 9886
rect 40908 9940 40964 9950
rect 41020 9940 41076 10446
rect 40908 9938 41076 9940
rect 40908 9886 40910 9938
rect 40962 9886 41076 9938
rect 40908 9884 41076 9886
rect 43036 9940 43092 9950
rect 40908 9874 40964 9884
rect 43036 9846 43092 9884
rect 43708 9826 43764 9838
rect 43708 9774 43710 9826
rect 43762 9774 43764 9826
rect 43708 9268 43764 9774
rect 43708 9202 43764 9212
rect 41020 9156 41076 9166
rect 41020 9062 41076 9100
rect 38108 6962 38164 6972
rect 38892 7362 38948 7374
rect 38892 7310 38894 7362
rect 38946 7310 38948 7362
rect 38892 7028 38948 7310
rect 38892 6962 38948 6972
rect 37436 5294 37438 5346
rect 37490 5294 37492 5346
rect 37436 5282 37492 5294
rect 37212 5182 37214 5234
rect 37266 5182 37268 5234
rect 37212 5170 37268 5182
rect 37772 5124 37828 5134
rect 38108 5124 38164 5134
rect 37772 5122 38164 5124
rect 37772 5070 37774 5122
rect 37826 5070 38110 5122
rect 38162 5070 38164 5122
rect 37772 5068 38164 5070
rect 37772 5058 37828 5068
rect 38108 5058 38164 5068
rect 36988 5012 37044 5022
rect 35980 4226 36148 4228
rect 35980 4174 35982 4226
rect 36034 4174 36148 4226
rect 35980 4172 36148 4174
rect 36204 4452 36260 4462
rect 35980 4162 36036 4172
rect 36204 3666 36260 4396
rect 36764 4452 36820 4462
rect 36316 4226 36372 4238
rect 36316 4174 36318 4226
rect 36370 4174 36372 4226
rect 36316 4116 36372 4174
rect 36316 4050 36372 4060
rect 36204 3614 36206 3666
rect 36258 3614 36260 3666
rect 36204 3602 36260 3614
rect 35756 3390 35758 3442
rect 35810 3390 35812 3442
rect 35756 3378 35812 3390
rect 30716 2994 30772 3332
rect 30716 2942 30718 2994
rect 30770 2942 30772 2994
rect 30716 2930 30772 2942
rect 36764 2994 36820 4396
rect 36988 3666 37044 4956
rect 38444 4900 38500 4910
rect 38444 4898 39060 4900
rect 38444 4846 38446 4898
rect 38498 4846 39060 4898
rect 38444 4844 39060 4846
rect 38444 4834 38500 4844
rect 38444 4228 38500 4238
rect 38444 4134 38500 4172
rect 36988 3614 36990 3666
rect 37042 3614 37044 3666
rect 36988 3602 37044 3614
rect 39004 3668 39060 4844
rect 39116 4340 39172 4350
rect 39116 4246 39172 4284
rect 39788 4340 39844 4350
rect 39116 3668 39172 3678
rect 39004 3666 39172 3668
rect 39004 3614 39118 3666
rect 39170 3614 39172 3666
rect 39004 3612 39172 3614
rect 39116 3602 39172 3612
rect 39788 3554 39844 4284
rect 39788 3502 39790 3554
rect 39842 3502 39844 3554
rect 39788 3490 39844 3502
rect 36764 2942 36766 2994
rect 36818 2942 36820 2994
rect 36764 2930 36820 2942
rect 30492 2718 30494 2770
rect 30546 2718 30548 2770
rect 30492 2706 30548 2718
rect 30044 2660 30100 2670
rect 29932 2658 30100 2660
rect 29932 2606 30046 2658
rect 30098 2606 30100 2658
rect 29932 2604 30100 2606
rect 30044 2594 30100 2604
rect 10332 2492 10724 2548
rect 10108 2454 10164 2492
rect 35196 2380 35460 2390
rect 35252 2324 35300 2380
rect 35356 2324 35404 2380
rect 35196 2314 35460 2324
rect 6860 2100 6916 2110
rect 6748 2098 6916 2100
rect 6748 2046 6862 2098
rect 6914 2046 6916 2098
rect 6748 2044 6916 2046
rect 6860 2034 6916 2044
rect 19836 1596 20100 1606
rect 19892 1540 19940 1596
rect 19996 1540 20044 1596
rect 19836 1530 20100 1540
<< via2 >>
rect 19836 78426 19892 78428
rect 19836 78374 19838 78426
rect 19838 78374 19890 78426
rect 19890 78374 19892 78426
rect 19836 78372 19892 78374
rect 19940 78426 19996 78428
rect 19940 78374 19942 78426
rect 19942 78374 19994 78426
rect 19994 78374 19996 78426
rect 19940 78372 19996 78374
rect 20044 78426 20100 78428
rect 20044 78374 20046 78426
rect 20046 78374 20098 78426
rect 20098 78374 20100 78426
rect 20044 78372 20100 78374
rect 4476 77642 4532 77644
rect 4476 77590 4478 77642
rect 4478 77590 4530 77642
rect 4530 77590 4532 77642
rect 4476 77588 4532 77590
rect 4580 77642 4636 77644
rect 4580 77590 4582 77642
rect 4582 77590 4634 77642
rect 4634 77590 4636 77642
rect 4580 77588 4636 77590
rect 4684 77642 4740 77644
rect 4684 77590 4686 77642
rect 4686 77590 4738 77642
rect 4738 77590 4740 77642
rect 4684 77588 4740 77590
rect 35196 77642 35252 77644
rect 35196 77590 35198 77642
rect 35198 77590 35250 77642
rect 35250 77590 35252 77642
rect 35196 77588 35252 77590
rect 35300 77642 35356 77644
rect 35300 77590 35302 77642
rect 35302 77590 35354 77642
rect 35354 77590 35356 77642
rect 35300 77588 35356 77590
rect 35404 77642 35460 77644
rect 35404 77590 35406 77642
rect 35406 77590 35458 77642
rect 35458 77590 35460 77642
rect 35404 77588 35460 77590
rect 3052 76690 3108 76692
rect 3052 76638 3054 76690
rect 3054 76638 3106 76690
rect 3106 76638 3108 76690
rect 3052 76636 3108 76638
rect 7532 77026 7588 77028
rect 7532 76974 7534 77026
rect 7534 76974 7586 77026
rect 7586 76974 7588 77026
rect 7532 76972 7588 76974
rect 3276 75628 3332 75684
rect 3388 76860 3444 76916
rect 3164 72380 3220 72436
rect 2940 72156 2996 72212
rect 1820 70924 1876 70980
rect 2380 70978 2436 70980
rect 2380 70926 2382 70978
rect 2382 70926 2434 70978
rect 2434 70926 2436 70978
rect 2380 70924 2436 70926
rect 2716 70924 2772 70980
rect 3612 76690 3668 76692
rect 3612 76638 3614 76690
rect 3614 76638 3666 76690
rect 3666 76638 3668 76690
rect 3612 76636 3668 76638
rect 4284 76636 4340 76692
rect 4956 76636 5012 76692
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 4284 75122 4340 75124
rect 4284 75070 4286 75122
rect 4286 75070 4338 75122
rect 4338 75070 4340 75122
rect 4284 75068 4340 75070
rect 4396 75628 4452 75684
rect 4956 75068 5012 75124
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 4060 72380 4116 72436
rect 3500 72156 3556 72212
rect 3724 71932 3780 71988
rect 3612 70866 3668 70868
rect 3612 70814 3614 70866
rect 3614 70814 3666 70866
rect 3666 70814 3668 70866
rect 3612 70812 3668 70814
rect 3948 71932 4004 71988
rect 5740 75122 5796 75124
rect 5740 75070 5742 75122
rect 5742 75070 5794 75122
rect 5794 75070 5796 75122
rect 5740 75068 5796 75070
rect 8204 76972 8260 77028
rect 8876 76972 8932 77028
rect 30492 77250 30548 77252
rect 30492 77198 30494 77250
rect 30494 77198 30546 77250
rect 30546 77198 30548 77250
rect 30492 77196 30548 77198
rect 31276 77196 31332 77252
rect 10108 76972 10164 77028
rect 11228 76972 11284 77028
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 10444 76466 10500 76468
rect 10444 76414 10446 76466
rect 10446 76414 10498 76466
rect 10498 76414 10500 76466
rect 10444 76412 10500 76414
rect 5068 71986 5124 71988
rect 5068 71934 5070 71986
rect 5070 71934 5122 71986
rect 5122 71934 5124 71986
rect 5068 71932 5124 71934
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 4172 70978 4228 70980
rect 4172 70926 4174 70978
rect 4174 70926 4226 70978
rect 4226 70926 4228 70978
rect 4172 70924 4228 70926
rect 4060 70812 4116 70868
rect 5628 70866 5684 70868
rect 5628 70814 5630 70866
rect 5630 70814 5682 70866
rect 5682 70814 5684 70866
rect 5628 70812 5684 70814
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 3836 69468 3892 69524
rect 4284 69468 4340 69524
rect 2604 67452 2660 67508
rect 2492 67004 2548 67060
rect 2940 67842 2996 67844
rect 2940 67790 2942 67842
rect 2942 67790 2994 67842
rect 2994 67790 2996 67842
rect 2940 67788 2996 67790
rect 2940 67452 2996 67508
rect 3164 67116 3220 67172
rect 3052 67058 3108 67060
rect 3052 67006 3054 67058
rect 3054 67006 3106 67058
rect 3106 67006 3108 67058
rect 3052 67004 3108 67006
rect 2940 66946 2996 66948
rect 2940 66894 2942 66946
rect 2942 66894 2994 66946
rect 2994 66894 2996 66946
rect 2940 66892 2996 66894
rect 3052 63196 3108 63252
rect 2716 63026 2772 63028
rect 2716 62974 2718 63026
rect 2718 62974 2770 63026
rect 2770 62974 2772 63026
rect 2716 62972 2772 62974
rect 3276 60620 3332 60676
rect 2716 58434 2772 58436
rect 2716 58382 2718 58434
rect 2718 58382 2770 58434
rect 2770 58382 2772 58434
rect 2716 58380 2772 58382
rect 1932 57650 1988 57652
rect 1932 57598 1934 57650
rect 1934 57598 1986 57650
rect 1986 57598 1988 57650
rect 1932 57596 1988 57598
rect 3052 57538 3108 57540
rect 3052 57486 3054 57538
rect 3054 57486 3106 57538
rect 3106 57486 3108 57538
rect 3052 57484 3108 57486
rect 3276 57650 3332 57652
rect 3276 57598 3278 57650
rect 3278 57598 3330 57650
rect 3330 57598 3332 57650
rect 3276 57596 3332 57598
rect 2940 56866 2996 56868
rect 2940 56814 2942 56866
rect 2942 56814 2994 56866
rect 2994 56814 2996 56866
rect 2940 56812 2996 56814
rect 1932 55298 1988 55300
rect 1932 55246 1934 55298
rect 1934 55246 1986 55298
rect 1986 55246 1988 55298
rect 1932 55244 1988 55246
rect 1932 54348 1988 54404
rect 2604 54684 2660 54740
rect 2492 54402 2548 54404
rect 2492 54350 2494 54402
rect 2494 54350 2546 54402
rect 2546 54350 2548 54402
rect 2492 54348 2548 54350
rect 2268 52834 2324 52836
rect 2268 52782 2270 52834
rect 2270 52782 2322 52834
rect 2322 52782 2324 52834
rect 2268 52780 2324 52782
rect 2044 50988 2100 51044
rect 2268 52556 2324 52612
rect 1596 42028 1652 42084
rect 3276 54460 3332 54516
rect 2604 52668 2660 52724
rect 2716 51938 2772 51940
rect 2716 51886 2718 51938
rect 2718 51886 2770 51938
rect 2770 51886 2772 51938
rect 2716 51884 2772 51886
rect 2716 50428 2772 50484
rect 1820 49810 1876 49812
rect 1820 49758 1822 49810
rect 1822 49758 1874 49810
rect 1874 49758 1876 49810
rect 1820 49756 1876 49758
rect 1932 48914 1988 48916
rect 1932 48862 1934 48914
rect 1934 48862 1986 48914
rect 1986 48862 1988 48914
rect 1932 48860 1988 48862
rect 2156 48972 2212 49028
rect 1932 47740 1988 47796
rect 3164 53730 3220 53732
rect 3164 53678 3166 53730
rect 3166 53678 3218 53730
rect 3218 53678 3220 53730
rect 3164 53676 3220 53678
rect 3276 52834 3332 52836
rect 3276 52782 3278 52834
rect 3278 52782 3330 52834
rect 3330 52782 3332 52834
rect 3276 52780 3332 52782
rect 3500 67842 3556 67844
rect 3500 67790 3502 67842
rect 3502 67790 3554 67842
rect 3554 67790 3556 67842
rect 3500 67788 3556 67790
rect 3612 67170 3668 67172
rect 3612 67118 3614 67170
rect 3614 67118 3666 67170
rect 3666 67118 3668 67170
rect 3612 67116 3668 67118
rect 3500 65772 3556 65828
rect 3724 66050 3780 66052
rect 3724 65998 3726 66050
rect 3726 65998 3778 66050
rect 3778 65998 3780 66050
rect 3724 65996 3780 65998
rect 4620 69522 4676 69524
rect 4620 69470 4622 69522
rect 4622 69470 4674 69522
rect 4674 69470 4676 69522
rect 4620 69468 4676 69470
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 5740 69522 5796 69524
rect 5740 69470 5742 69522
rect 5742 69470 5794 69522
rect 5794 69470 5796 69522
rect 5740 69468 5796 69470
rect 4956 68012 5012 68068
rect 5740 68066 5796 68068
rect 5740 68014 5742 68066
rect 5742 68014 5794 68066
rect 5794 68014 5796 68066
rect 5740 68012 5796 68014
rect 13020 76466 13076 76468
rect 13020 76414 13022 76466
rect 13022 76414 13074 76466
rect 13074 76414 13076 76466
rect 13020 76412 13076 76414
rect 12572 76242 12628 76244
rect 12572 76190 12574 76242
rect 12574 76190 12626 76242
rect 12626 76190 12628 76242
rect 12572 76188 12628 76190
rect 18508 76466 18564 76468
rect 18508 76414 18510 76466
rect 18510 76414 18562 76466
rect 18562 76414 18564 76466
rect 18508 76412 18564 76414
rect 21756 76466 21812 76468
rect 21756 76414 21758 76466
rect 21758 76414 21810 76466
rect 21810 76414 21812 76466
rect 21756 76412 21812 76414
rect 13804 76188 13860 76244
rect 15148 76242 15204 76244
rect 15148 76190 15150 76242
rect 15150 76190 15202 76242
rect 15202 76190 15204 76242
rect 15148 76188 15204 76190
rect 9660 73948 9716 74004
rect 10668 73948 10724 74004
rect 12236 73836 12292 73892
rect 21420 76354 21476 76356
rect 21420 76302 21422 76354
rect 21422 76302 21474 76354
rect 21474 76302 21476 76354
rect 21420 76300 21476 76302
rect 19292 75852 19348 75908
rect 21308 75906 21364 75908
rect 21308 75854 21310 75906
rect 21310 75854 21362 75906
rect 21362 75854 21364 75906
rect 21308 75852 21364 75854
rect 23548 76300 23604 76356
rect 24556 75740 24612 75796
rect 20748 75682 20804 75684
rect 20748 75630 20750 75682
rect 20750 75630 20802 75682
rect 20802 75630 20804 75682
rect 20748 75628 20804 75630
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 6636 70140 6692 70196
rect 6188 69522 6244 69524
rect 6188 69470 6190 69522
rect 6190 69470 6242 69522
rect 6242 69470 6244 69522
rect 6188 69468 6244 69470
rect 6076 67842 6132 67844
rect 6076 67790 6078 67842
rect 6078 67790 6130 67842
rect 6130 67790 6132 67842
rect 6076 67788 6132 67790
rect 4844 66946 4900 66948
rect 4844 66894 4846 66946
rect 4846 66894 4898 66946
rect 4898 66894 4900 66946
rect 4844 66892 4900 66894
rect 5516 66892 5572 66948
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 4172 66050 4228 66052
rect 4172 65998 4174 66050
rect 4174 65998 4226 66050
rect 4226 65998 4228 66050
rect 4172 65996 4228 65998
rect 3612 65324 3668 65380
rect 3724 62972 3780 63028
rect 3948 65324 4004 65380
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 4508 63250 4564 63252
rect 4508 63198 4510 63250
rect 4510 63198 4562 63250
rect 4562 63198 4564 63250
rect 4508 63196 4564 63198
rect 5292 63196 5348 63252
rect 3948 61740 4004 61796
rect 4060 61852 4116 61908
rect 3500 58828 3556 58884
rect 3500 57372 3556 57428
rect 3724 60674 3780 60676
rect 3724 60622 3726 60674
rect 3726 60622 3778 60674
rect 3778 60622 3780 60674
rect 3724 60620 3780 60622
rect 4732 62130 4788 62132
rect 4732 62078 4734 62130
rect 4734 62078 4786 62130
rect 4786 62078 4788 62130
rect 4732 62076 4788 62078
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 4284 61404 4340 61460
rect 4620 61740 4676 61796
rect 3724 55356 3780 55412
rect 4172 60620 4228 60676
rect 4620 60620 4676 60676
rect 5852 62076 5908 62132
rect 5628 61458 5684 61460
rect 5628 61406 5630 61458
rect 5630 61406 5682 61458
rect 5682 61406 5684 61458
rect 5628 61404 5684 61406
rect 6412 67228 6468 67284
rect 7532 70194 7588 70196
rect 7532 70142 7534 70194
rect 7534 70142 7586 70194
rect 7586 70142 7588 70194
rect 7532 70140 7588 70142
rect 13020 73052 13076 73108
rect 9884 70194 9940 70196
rect 9884 70142 9886 70194
rect 9886 70142 9938 70194
rect 9938 70142 9940 70194
rect 9884 70140 9940 70142
rect 10668 70140 10724 70196
rect 8316 67954 8372 67956
rect 8316 67902 8318 67954
rect 8318 67902 8370 67954
rect 8370 67902 8372 67954
rect 8316 67900 8372 67902
rect 10332 69186 10388 69188
rect 10332 69134 10334 69186
rect 10334 69134 10386 69186
rect 10386 69134 10388 69186
rect 10332 69132 10388 69134
rect 10332 68012 10388 68068
rect 9436 67900 9492 67956
rect 7644 67842 7700 67844
rect 7644 67790 7646 67842
rect 7646 67790 7698 67842
rect 7698 67790 7700 67842
rect 7644 67788 7700 67790
rect 7196 67228 7252 67284
rect 6076 66946 6132 66948
rect 6076 66894 6078 66946
rect 6078 66894 6130 66946
rect 6130 66894 6132 66946
rect 6076 66892 6132 66894
rect 6748 66892 6804 66948
rect 6972 66834 7028 66836
rect 6972 66782 6974 66834
rect 6974 66782 7026 66834
rect 7026 66782 7028 66834
rect 6972 66780 7028 66782
rect 8764 67004 8820 67060
rect 7532 66780 7588 66836
rect 10780 69132 10836 69188
rect 11452 69132 11508 69188
rect 14252 73106 14308 73108
rect 14252 73054 14254 73106
rect 14254 73054 14306 73106
rect 14306 73054 14308 73106
rect 14252 73052 14308 73054
rect 12348 70194 12404 70196
rect 12348 70142 12350 70194
rect 12350 70142 12402 70194
rect 12402 70142 12404 70194
rect 12348 70140 12404 70142
rect 16828 70588 16884 70644
rect 13356 70194 13412 70196
rect 13356 70142 13358 70194
rect 13358 70142 13410 70194
rect 13410 70142 13412 70194
rect 13356 70140 13412 70142
rect 14700 70194 14756 70196
rect 14700 70142 14702 70194
rect 14702 70142 14754 70194
rect 14754 70142 14756 70194
rect 14700 70140 14756 70142
rect 11900 69132 11956 69188
rect 10668 67004 10724 67060
rect 10780 68066 10836 68068
rect 10780 68014 10782 68066
rect 10782 68014 10834 68066
rect 10834 68014 10836 68066
rect 10780 68012 10836 68014
rect 6860 66220 6916 66276
rect 7308 66220 7364 66276
rect 7644 66274 7700 66276
rect 7644 66222 7646 66274
rect 7646 66222 7698 66274
rect 7698 66222 7700 66274
rect 7644 66220 7700 66222
rect 6748 65436 6804 65492
rect 7756 65490 7812 65492
rect 7756 65438 7758 65490
rect 7758 65438 7810 65490
rect 7810 65438 7812 65490
rect 7756 65436 7812 65438
rect 9660 65996 9716 66052
rect 10220 66050 10276 66052
rect 10220 65998 10222 66050
rect 10222 65998 10274 66050
rect 10274 65998 10276 66050
rect 10220 65996 10276 65998
rect 11676 67058 11732 67060
rect 11676 67006 11678 67058
rect 11678 67006 11730 67058
rect 11730 67006 11732 67058
rect 11676 67004 11732 67006
rect 10780 65996 10836 66052
rect 9436 65436 9492 65492
rect 6636 65324 6692 65380
rect 8204 65378 8260 65380
rect 8204 65326 8206 65378
rect 8206 65326 8258 65378
rect 8258 65326 8260 65378
rect 8204 65324 8260 65326
rect 6076 63196 6132 63252
rect 6412 63196 6468 63252
rect 7420 63196 7476 63252
rect 7420 62578 7476 62580
rect 7420 62526 7422 62578
rect 7422 62526 7474 62578
rect 7474 62526 7476 62578
rect 7420 62524 7476 62526
rect 8988 65378 9044 65380
rect 8988 65326 8990 65378
rect 8990 65326 9042 65378
rect 9042 65326 9044 65378
rect 8988 65324 9044 65326
rect 10780 65490 10836 65492
rect 10780 65438 10782 65490
rect 10782 65438 10834 65490
rect 10834 65438 10836 65490
rect 10780 65436 10836 65438
rect 9548 65324 9604 65380
rect 10108 64652 10164 64708
rect 10780 64706 10836 64708
rect 10780 64654 10782 64706
rect 10782 64654 10834 64706
rect 10834 64654 10836 64706
rect 10780 64652 10836 64654
rect 10668 64482 10724 64484
rect 10668 64430 10670 64482
rect 10670 64430 10722 64482
rect 10722 64430 10724 64482
rect 10668 64428 10724 64430
rect 11116 65324 11172 65380
rect 11116 64652 11172 64708
rect 11340 66050 11396 66052
rect 11340 65998 11342 66050
rect 11342 65998 11394 66050
rect 11394 65998 11396 66050
rect 11340 65996 11396 65998
rect 11452 64428 11508 64484
rect 7644 61570 7700 61572
rect 7644 61518 7646 61570
rect 7646 61518 7698 61570
rect 7698 61518 7700 61570
rect 7644 61516 7700 61518
rect 5068 60674 5124 60676
rect 5068 60622 5070 60674
rect 5070 60622 5122 60674
rect 5122 60622 5124 60674
rect 5068 60620 5124 60622
rect 4956 60508 5012 60564
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 3724 55186 3780 55188
rect 3724 55134 3726 55186
rect 3726 55134 3778 55186
rect 3778 55134 3780 55186
rect 3724 55132 3780 55134
rect 3612 54684 3668 54740
rect 3612 54514 3668 54516
rect 3612 54462 3614 54514
rect 3614 54462 3666 54514
rect 3666 54462 3668 54514
rect 3612 54460 3668 54462
rect 3612 53788 3668 53844
rect 3948 58828 4004 58884
rect 3724 53452 3780 53508
rect 3500 52668 3556 52724
rect 3276 51884 3332 51940
rect 3164 51212 3220 51268
rect 2268 48914 2324 48916
rect 2268 48862 2270 48914
rect 2270 48862 2322 48914
rect 2322 48862 2324 48914
rect 2268 48860 2324 48862
rect 2380 48130 2436 48132
rect 2380 48078 2382 48130
rect 2382 48078 2434 48130
rect 2434 48078 2436 48130
rect 2380 48076 2436 48078
rect 2492 47964 2548 48020
rect 2268 47404 2324 47460
rect 2380 47346 2436 47348
rect 2380 47294 2382 47346
rect 2382 47294 2434 47346
rect 2434 47294 2436 47346
rect 2380 47292 2436 47294
rect 2940 49196 2996 49252
rect 2716 47740 2772 47796
rect 2828 48466 2884 48468
rect 2828 48414 2830 48466
rect 2830 48414 2882 48466
rect 2882 48414 2884 48466
rect 2828 48412 2884 48414
rect 3276 50316 3332 50372
rect 3388 50988 3444 51044
rect 3052 48972 3108 49028
rect 3276 49026 3332 49028
rect 3276 48974 3278 49026
rect 3278 48974 3330 49026
rect 3330 48974 3332 49026
rect 3276 48972 3332 48974
rect 2940 46956 2996 47012
rect 2604 46562 2660 46564
rect 2604 46510 2606 46562
rect 2606 46510 2658 46562
rect 2658 46510 2660 46562
rect 2604 46508 2660 46510
rect 2156 46284 2212 46340
rect 2380 46060 2436 46116
rect 3164 47964 3220 48020
rect 3276 48076 3332 48132
rect 3164 47458 3220 47460
rect 3164 47406 3166 47458
rect 3166 47406 3218 47458
rect 3218 47406 3220 47458
rect 3164 47404 3220 47406
rect 3276 46620 3332 46676
rect 3052 46508 3108 46564
rect 2940 46284 2996 46340
rect 2940 46114 2996 46116
rect 2940 46062 2942 46114
rect 2942 46062 2994 46114
rect 2994 46062 2996 46114
rect 2940 46060 2996 46062
rect 3276 45890 3332 45892
rect 3276 45838 3278 45890
rect 3278 45838 3330 45890
rect 3330 45838 3332 45890
rect 3276 45836 3332 45838
rect 3052 45500 3108 45556
rect 2380 44994 2436 44996
rect 2380 44942 2382 44994
rect 2382 44942 2434 44994
rect 2434 44942 2436 44994
rect 2380 44940 2436 44942
rect 2044 44492 2100 44548
rect 2492 44322 2548 44324
rect 2492 44270 2494 44322
rect 2494 44270 2546 44322
rect 2546 44270 2548 44322
rect 2492 44268 2548 44270
rect 2940 44940 2996 44996
rect 2940 44322 2996 44324
rect 2940 44270 2942 44322
rect 2942 44270 2994 44322
rect 2994 44270 2996 44322
rect 2940 44268 2996 44270
rect 2828 44210 2884 44212
rect 2828 44158 2830 44210
rect 2830 44158 2882 44210
rect 2882 44158 2884 44210
rect 2828 44156 2884 44158
rect 2940 43932 2996 43988
rect 2044 41580 2100 41636
rect 1820 41186 1876 41188
rect 1820 41134 1822 41186
rect 1822 41134 1874 41186
rect 1874 41134 1876 41186
rect 1820 41132 1876 41134
rect 2380 42588 2436 42644
rect 2940 42642 2996 42644
rect 2940 42590 2942 42642
rect 2942 42590 2994 42642
rect 2994 42590 2996 42642
rect 2940 42588 2996 42590
rect 3500 50540 3556 50596
rect 3500 50316 3556 50372
rect 3500 48076 3556 48132
rect 3500 47458 3556 47460
rect 3500 47406 3502 47458
rect 3502 47406 3554 47458
rect 3554 47406 3556 47458
rect 3500 47404 3556 47406
rect 3724 52332 3780 52388
rect 3724 52162 3780 52164
rect 3724 52110 3726 52162
rect 3726 52110 3778 52162
rect 3778 52110 3780 52162
rect 3724 52108 3780 52110
rect 3724 51266 3780 51268
rect 3724 51214 3726 51266
rect 3726 51214 3778 51266
rect 3778 51214 3780 51266
rect 3724 51212 3780 51214
rect 3724 50428 3780 50484
rect 4060 58434 4116 58436
rect 4060 58382 4062 58434
rect 4062 58382 4114 58434
rect 4114 58382 4116 58434
rect 4060 58380 4116 58382
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 5852 60508 5908 60564
rect 6300 59836 6356 59892
rect 4284 58380 4340 58436
rect 4060 57484 4116 57540
rect 4508 57372 4564 57428
rect 5740 58940 5796 58996
rect 5292 58380 5348 58436
rect 5292 57874 5348 57876
rect 5292 57822 5294 57874
rect 5294 57822 5346 57874
rect 5346 57822 5348 57874
rect 5292 57820 5348 57822
rect 5180 57596 5236 57652
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4172 55356 4228 55412
rect 4060 55132 4116 55188
rect 4172 55074 4228 55076
rect 4172 55022 4174 55074
rect 4174 55022 4226 55074
rect 4226 55022 4228 55074
rect 4172 55020 4228 55022
rect 4172 53900 4228 53956
rect 4620 55298 4676 55300
rect 4620 55246 4622 55298
rect 4622 55246 4674 55298
rect 4674 55246 4676 55298
rect 4620 55244 4676 55246
rect 4732 55020 4788 55076
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4060 53116 4116 53172
rect 4172 53676 4228 53732
rect 4284 53564 4340 53620
rect 4284 53058 4340 53060
rect 4284 53006 4286 53058
rect 4286 53006 4338 53058
rect 4338 53006 4340 53058
rect 4284 53004 4340 53006
rect 4060 52556 4116 52612
rect 4172 52780 4228 52836
rect 4060 52386 4116 52388
rect 4060 52334 4062 52386
rect 4062 52334 4114 52386
rect 4114 52334 4116 52386
rect 4060 52332 4116 52334
rect 4508 53900 4564 53956
rect 7644 60732 7700 60788
rect 7532 59890 7588 59892
rect 7532 59838 7534 59890
rect 7534 59838 7586 59890
rect 7586 59838 7588 59890
rect 7532 59836 7588 59838
rect 6300 58940 6356 58996
rect 6524 58434 6580 58436
rect 6524 58382 6526 58434
rect 6526 58382 6578 58434
rect 6578 58382 6580 58434
rect 6524 58380 6580 58382
rect 6412 57874 6468 57876
rect 6412 57822 6414 57874
rect 6414 57822 6466 57874
rect 6466 57822 6468 57874
rect 6412 57820 6468 57822
rect 7196 58380 7252 58436
rect 6748 57820 6804 57876
rect 7308 57484 7364 57540
rect 6748 56924 6804 56980
rect 5852 56866 5908 56868
rect 5852 56814 5854 56866
rect 5854 56814 5906 56866
rect 5906 56814 5908 56866
rect 5852 56812 5908 56814
rect 5740 55074 5796 55076
rect 5740 55022 5742 55074
rect 5742 55022 5794 55074
rect 5794 55022 5796 55074
rect 5740 55020 5796 55022
rect 5180 54908 5236 54964
rect 6188 55186 6244 55188
rect 6188 55134 6190 55186
rect 6190 55134 6242 55186
rect 6242 55134 6244 55186
rect 6188 55132 6244 55134
rect 6076 55074 6132 55076
rect 6076 55022 6078 55074
rect 6078 55022 6130 55074
rect 6130 55022 6132 55074
rect 6076 55020 6132 55022
rect 5964 54908 6020 54964
rect 4508 52892 4564 52948
rect 4172 51266 4228 51268
rect 4172 51214 4174 51266
rect 4174 51214 4226 51266
rect 4226 51214 4228 51266
rect 4172 51212 4228 51214
rect 5516 53564 5572 53620
rect 4844 53340 4900 53396
rect 5292 53116 5348 53172
rect 3948 50594 4004 50596
rect 3948 50542 3950 50594
rect 3950 50542 4002 50594
rect 4002 50542 4004 50594
rect 3948 50540 4004 50542
rect 3948 49868 4004 49924
rect 3948 49644 4004 49700
rect 3612 46956 3668 47012
rect 4060 48412 4116 48468
rect 3612 46620 3668 46676
rect 3500 46060 3556 46116
rect 3724 46060 3780 46116
rect 3612 45890 3668 45892
rect 3612 45838 3614 45890
rect 3614 45838 3666 45890
rect 3666 45838 3668 45890
rect 3612 45836 3668 45838
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4844 52444 4900 52500
rect 4396 51884 4452 51940
rect 4508 51212 4564 51268
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4844 50594 4900 50596
rect 4844 50542 4846 50594
rect 4846 50542 4898 50594
rect 4898 50542 4900 50594
rect 4844 50540 4900 50542
rect 4732 50428 4788 50484
rect 4844 49868 4900 49924
rect 4396 49644 4452 49700
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4284 49196 4340 49252
rect 4508 49138 4564 49140
rect 4508 49086 4510 49138
rect 4510 49086 4562 49138
rect 4562 49086 4564 49138
rect 4508 49084 4564 49086
rect 4284 48972 4340 49028
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4620 47628 4676 47684
rect 4060 47458 4116 47460
rect 4060 47406 4062 47458
rect 4062 47406 4114 47458
rect 4114 47406 4116 47458
rect 4060 47404 4116 47406
rect 3836 44940 3892 44996
rect 3052 42140 3108 42196
rect 3388 44268 3444 44324
rect 3500 44044 3556 44100
rect 3836 44098 3892 44100
rect 3836 44046 3838 44098
rect 3838 44046 3890 44098
rect 3890 44046 3892 44098
rect 3836 44044 3892 44046
rect 4060 46956 4116 47012
rect 5292 52220 5348 52276
rect 5292 49810 5348 49812
rect 5292 49758 5294 49810
rect 5294 49758 5346 49810
rect 5346 49758 5348 49810
rect 5292 49756 5348 49758
rect 4956 47234 5012 47236
rect 4956 47182 4958 47234
rect 4958 47182 5010 47234
rect 5010 47182 5012 47234
rect 4956 47180 5012 47182
rect 4844 46620 4900 46676
rect 4284 46508 4340 46564
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4396 46060 4452 46116
rect 4172 45500 4228 45556
rect 4060 43148 4116 43204
rect 4172 45276 4228 45332
rect 4620 44940 4676 44996
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 3276 42140 3332 42196
rect 3388 42364 3444 42420
rect 2604 41580 2660 41636
rect 2828 41970 2884 41972
rect 2828 41918 2830 41970
rect 2830 41918 2882 41970
rect 2882 41918 2884 41970
rect 2828 41916 2884 41918
rect 2940 41746 2996 41748
rect 2940 41694 2942 41746
rect 2942 41694 2994 41746
rect 2994 41694 2996 41746
rect 2940 41692 2996 41694
rect 1820 38050 1876 38052
rect 1820 37998 1822 38050
rect 1822 37998 1874 38050
rect 1874 37998 1876 38050
rect 1820 37996 1876 37998
rect 1932 37436 1988 37492
rect 2828 40572 2884 40628
rect 3164 41356 3220 41412
rect 2604 40460 2660 40516
rect 2492 40348 2548 40404
rect 2604 40290 2660 40292
rect 2604 40238 2606 40290
rect 2606 40238 2658 40290
rect 2658 40238 2660 40290
rect 2604 40236 2660 40238
rect 4172 42812 4228 42868
rect 4284 44044 4340 44100
rect 3948 42588 4004 42644
rect 3612 41916 3668 41972
rect 4172 42642 4228 42644
rect 4172 42590 4174 42642
rect 4174 42590 4226 42642
rect 4226 42590 4228 42642
rect 4172 42588 4228 42590
rect 3388 40236 3444 40292
rect 4732 44322 4788 44324
rect 4732 44270 4734 44322
rect 4734 44270 4786 44322
rect 4786 44270 4788 44322
rect 4732 44268 4788 44270
rect 4508 43372 4564 43428
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 5180 46732 5236 46788
rect 5068 45388 5124 45444
rect 5852 53564 5908 53620
rect 5740 53506 5796 53508
rect 5740 53454 5742 53506
rect 5742 53454 5794 53506
rect 5794 53454 5796 53506
rect 5740 53452 5796 53454
rect 6076 53340 6132 53396
rect 7084 56866 7140 56868
rect 7084 56814 7086 56866
rect 7086 56814 7138 56866
rect 7138 56814 7140 56866
rect 7084 56812 7140 56814
rect 6636 55298 6692 55300
rect 6636 55246 6638 55298
rect 6638 55246 6690 55298
rect 6690 55246 6692 55298
rect 6636 55244 6692 55246
rect 5628 52444 5684 52500
rect 5852 52722 5908 52724
rect 5852 52670 5854 52722
rect 5854 52670 5906 52722
rect 5906 52670 5908 52722
rect 5852 52668 5908 52670
rect 7196 55020 7252 55076
rect 6524 53618 6580 53620
rect 6524 53566 6526 53618
rect 6526 53566 6578 53618
rect 6578 53566 6580 53618
rect 6524 53564 6580 53566
rect 6748 53506 6804 53508
rect 6748 53454 6750 53506
rect 6750 53454 6802 53506
rect 6802 53454 6804 53506
rect 6748 53452 6804 53454
rect 6972 53340 7028 53396
rect 6860 52780 6916 52836
rect 6412 52108 6468 52164
rect 6300 51378 6356 51380
rect 6300 51326 6302 51378
rect 6302 51326 6354 51378
rect 6354 51326 6356 51378
rect 6300 51324 6356 51326
rect 6300 50540 6356 50596
rect 6076 50428 6132 50484
rect 6076 49756 6132 49812
rect 5964 49250 6020 49252
rect 5964 49198 5966 49250
rect 5966 49198 6018 49250
rect 6018 49198 6020 49250
rect 5964 49196 6020 49198
rect 6412 49138 6468 49140
rect 6412 49086 6414 49138
rect 6414 49086 6466 49138
rect 6466 49086 6468 49138
rect 6412 49084 6468 49086
rect 5852 47458 5908 47460
rect 5852 47406 5854 47458
rect 5854 47406 5906 47458
rect 5906 47406 5908 47458
rect 5852 47404 5908 47406
rect 5516 46786 5572 46788
rect 5516 46734 5518 46786
rect 5518 46734 5570 46786
rect 5570 46734 5572 46786
rect 5516 46732 5572 46734
rect 6188 46508 6244 46564
rect 6076 45666 6132 45668
rect 6076 45614 6078 45666
rect 6078 45614 6130 45666
rect 6130 45614 6132 45666
rect 6076 45612 6132 45614
rect 4060 42364 4116 42420
rect 2828 39730 2884 39732
rect 2828 39678 2830 39730
rect 2830 39678 2882 39730
rect 2882 39678 2884 39730
rect 2828 39676 2884 39678
rect 3052 39676 3108 39732
rect 2716 39340 2772 39396
rect 3612 41244 3668 41300
rect 3612 40460 3668 40516
rect 3724 40572 3780 40628
rect 3500 39676 3556 39732
rect 3836 39788 3892 39844
rect 3276 39564 3332 39620
rect 3276 39394 3332 39396
rect 3276 39342 3278 39394
rect 3278 39342 3330 39394
rect 3330 39342 3332 39394
rect 3276 39340 3332 39342
rect 2156 37938 2212 37940
rect 2156 37886 2158 37938
rect 2158 37886 2210 37938
rect 2210 37886 2212 37938
rect 2156 37884 2212 37886
rect 2268 37324 2324 37380
rect 2492 37996 2548 38052
rect 2716 38556 2772 38612
rect 2828 38050 2884 38052
rect 2828 37998 2830 38050
rect 2830 37998 2882 38050
rect 2882 37998 2884 38050
rect 2828 37996 2884 37998
rect 2940 37324 2996 37380
rect 2492 36988 2548 37044
rect 1932 36316 1988 36372
rect 2044 36204 2100 36260
rect 1932 33292 1988 33348
rect 2268 36764 2324 36820
rect 1708 32562 1764 32564
rect 1708 32510 1710 32562
rect 1710 32510 1762 32562
rect 1762 32510 1764 32562
rect 1708 32508 1764 32510
rect 1932 31276 1988 31332
rect 3500 37996 3556 38052
rect 3164 36764 3220 36820
rect 3276 37548 3332 37604
rect 2604 36370 2660 36372
rect 2604 36318 2606 36370
rect 2606 36318 2658 36370
rect 2658 36318 2660 36370
rect 2604 36316 2660 36318
rect 2492 36204 2548 36260
rect 2492 35922 2548 35924
rect 2492 35870 2494 35922
rect 2494 35870 2546 35922
rect 2546 35870 2548 35922
rect 2492 35868 2548 35870
rect 2492 33292 2548 33348
rect 3388 36988 3444 37044
rect 3724 37324 3780 37380
rect 3612 36482 3668 36484
rect 3612 36430 3614 36482
rect 3614 36430 3666 36482
rect 3666 36430 3668 36482
rect 3612 36428 3668 36430
rect 3500 35922 3556 35924
rect 3500 35870 3502 35922
rect 3502 35870 3554 35922
rect 3554 35870 3556 35922
rect 3500 35868 3556 35870
rect 3612 34188 3668 34244
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4620 41298 4676 41300
rect 4620 41246 4622 41298
rect 4622 41246 4674 41298
rect 4674 41246 4676 41298
rect 4620 41244 4676 41246
rect 4956 42028 5012 42084
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4508 39788 4564 39844
rect 4172 39340 4228 39396
rect 4284 39116 4340 39172
rect 4844 39564 4900 39620
rect 5068 41356 5124 41412
rect 5068 40962 5124 40964
rect 5068 40910 5070 40962
rect 5070 40910 5122 40962
rect 5122 40910 5124 40962
rect 5068 40908 5124 40910
rect 5628 40684 5684 40740
rect 5292 39676 5348 39732
rect 4732 38556 4788 38612
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4396 38050 4452 38052
rect 4396 37998 4398 38050
rect 4398 37998 4450 38050
rect 4450 37998 4452 38050
rect 4396 37996 4452 37998
rect 4284 37436 4340 37492
rect 4620 37938 4676 37940
rect 4620 37886 4622 37938
rect 4622 37886 4674 37938
rect 4674 37886 4676 37938
rect 4620 37884 4676 37886
rect 5180 38556 5236 38612
rect 4956 38050 5012 38052
rect 4956 37998 4958 38050
rect 4958 37998 5010 38050
rect 5010 37998 5012 38050
rect 4956 37996 5012 37998
rect 4396 37324 4452 37380
rect 4476 36874 4532 36876
rect 4284 36764 4340 36820
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 3836 36428 3892 36484
rect 4060 36652 4116 36708
rect 3948 34300 4004 34356
rect 3948 33516 4004 33572
rect 3948 32284 4004 32340
rect 3052 31276 3108 31332
rect 2828 30268 2884 30324
rect 3276 31778 3332 31780
rect 3276 31726 3278 31778
rect 3278 31726 3330 31778
rect 3330 31726 3332 31778
rect 3276 31724 3332 31726
rect 3164 31218 3220 31220
rect 3164 31166 3166 31218
rect 3166 31166 3218 31218
rect 3218 31166 3220 31218
rect 3164 31164 3220 31166
rect 1932 28700 1988 28756
rect 2940 29372 2996 29428
rect 2156 28364 2212 28420
rect 2716 27916 2772 27972
rect 2156 27858 2212 27860
rect 2156 27806 2158 27858
rect 2158 27806 2210 27858
rect 2210 27806 2212 27858
rect 2156 27804 2212 27806
rect 2604 27580 2660 27636
rect 2156 27468 2212 27524
rect 3388 30940 3444 30996
rect 3388 29708 3444 29764
rect 3164 28028 3220 28084
rect 3164 27804 3220 27860
rect 2268 26290 2324 26292
rect 2268 26238 2270 26290
rect 2270 26238 2322 26290
rect 2322 26238 2324 26290
rect 2268 26236 2324 26238
rect 1708 22652 1764 22708
rect 1820 22428 1876 22484
rect 3052 26236 3108 26292
rect 3276 26962 3332 26964
rect 3276 26910 3278 26962
rect 3278 26910 3330 26962
rect 3330 26910 3332 26962
rect 3276 26908 3332 26910
rect 2380 24892 2436 24948
rect 2268 23938 2324 23940
rect 2268 23886 2270 23938
rect 2270 23886 2322 23938
rect 2322 23886 2324 23938
rect 2268 23884 2324 23886
rect 2492 21532 2548 21588
rect 2940 24946 2996 24948
rect 2940 24894 2942 24946
rect 2942 24894 2994 24946
rect 2994 24894 2996 24946
rect 2940 24892 2996 24894
rect 4844 36540 4900 36596
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4172 34802 4228 34804
rect 4172 34750 4174 34802
rect 4174 34750 4226 34802
rect 4226 34750 4228 34802
rect 4172 34748 4228 34750
rect 5180 37490 5236 37492
rect 5180 37438 5182 37490
rect 5182 37438 5234 37490
rect 5234 37438 5236 37490
rect 5180 37436 5236 37438
rect 6188 44380 6244 44436
rect 6300 46620 6356 46676
rect 6972 49084 7028 49140
rect 6748 47964 6804 48020
rect 6748 47682 6804 47684
rect 6748 47630 6750 47682
rect 6750 47630 6802 47682
rect 6802 47630 6804 47682
rect 6748 47628 6804 47630
rect 7532 56866 7588 56868
rect 7532 56814 7534 56866
rect 7534 56814 7586 56866
rect 7586 56814 7588 56866
rect 7532 56812 7588 56814
rect 8316 61516 8372 61572
rect 8652 62524 8708 62580
rect 9436 62524 9492 62580
rect 9436 61570 9492 61572
rect 9436 61518 9438 61570
rect 9438 61518 9490 61570
rect 9490 61518 9492 61570
rect 9436 61516 9492 61518
rect 8876 61458 8932 61460
rect 8876 61406 8878 61458
rect 8878 61406 8930 61458
rect 8930 61406 8932 61458
rect 8876 61404 8932 61406
rect 9548 61404 9604 61460
rect 8764 60786 8820 60788
rect 8764 60734 8766 60786
rect 8766 60734 8818 60786
rect 8818 60734 8820 60786
rect 8764 60732 8820 60734
rect 8652 60674 8708 60676
rect 8652 60622 8654 60674
rect 8654 60622 8706 60674
rect 8706 60622 8708 60674
rect 8652 60620 8708 60622
rect 12012 64428 12068 64484
rect 12460 65436 12516 65492
rect 13020 65436 13076 65492
rect 12124 65324 12180 65380
rect 11452 63644 11508 63700
rect 10780 61458 10836 61460
rect 10780 61406 10782 61458
rect 10782 61406 10834 61458
rect 10834 61406 10836 61458
rect 10780 61404 10836 61406
rect 10668 60620 10724 60676
rect 12124 63922 12180 63924
rect 12124 63870 12126 63922
rect 12126 63870 12178 63922
rect 12178 63870 12180 63922
rect 12124 63868 12180 63870
rect 11788 63644 11844 63700
rect 14476 63868 14532 63924
rect 16380 63250 16436 63252
rect 16380 63198 16382 63250
rect 16382 63198 16434 63250
rect 16434 63198 16436 63250
rect 16380 63196 16436 63198
rect 11676 60620 11732 60676
rect 10668 59218 10724 59220
rect 10668 59166 10670 59218
rect 10670 59166 10722 59218
rect 10722 59166 10724 59218
rect 10668 59164 10724 59166
rect 12012 59330 12068 59332
rect 12012 59278 12014 59330
rect 12014 59278 12066 59330
rect 12066 59278 12068 59330
rect 12012 59276 12068 59278
rect 10892 58380 10948 58436
rect 7980 57820 8036 57876
rect 12012 58434 12068 58436
rect 12012 58382 12014 58434
rect 12014 58382 12066 58434
rect 12066 58382 12068 58434
rect 12012 58380 12068 58382
rect 12124 59164 12180 59220
rect 11900 57820 11956 57876
rect 7980 57036 8036 57092
rect 8316 57036 8372 57092
rect 9548 57090 9604 57092
rect 9548 57038 9550 57090
rect 9550 57038 9602 57090
rect 9602 57038 9604 57090
rect 9548 57036 9604 57038
rect 8988 56812 9044 56868
rect 7980 55468 8036 55524
rect 10780 57036 10836 57092
rect 12796 59218 12852 59220
rect 12796 59166 12798 59218
rect 12798 59166 12850 59218
rect 12850 59166 12852 59218
rect 12796 59164 12852 59166
rect 13244 59164 13300 59220
rect 15596 63138 15652 63140
rect 15596 63086 15598 63138
rect 15598 63086 15650 63138
rect 15650 63086 15652 63138
rect 15596 63084 15652 63086
rect 14252 59276 14308 59332
rect 14028 57874 14084 57876
rect 14028 57822 14030 57874
rect 14030 57822 14082 57874
rect 14082 57822 14084 57874
rect 14028 57820 14084 57822
rect 14812 59276 14868 59332
rect 15036 59052 15092 59108
rect 14700 57820 14756 57876
rect 12124 57090 12180 57092
rect 12124 57038 12126 57090
rect 12126 57038 12178 57090
rect 12178 57038 12180 57090
rect 12124 57036 12180 57038
rect 9996 56866 10052 56868
rect 9996 56814 9998 56866
rect 9998 56814 10050 56866
rect 10050 56814 10052 56866
rect 9996 56812 10052 56814
rect 7644 53842 7700 53844
rect 7644 53790 7646 53842
rect 7646 53790 7698 53842
rect 7698 53790 7700 53842
rect 7644 53788 7700 53790
rect 7532 53116 7588 53172
rect 13132 55020 13188 55076
rect 7980 53900 8036 53956
rect 9436 53900 9492 53956
rect 13804 54348 13860 54404
rect 8428 53506 8484 53508
rect 8428 53454 8430 53506
rect 8430 53454 8482 53506
rect 8482 53454 8484 53506
rect 8428 53452 8484 53454
rect 8876 53228 8932 53284
rect 7756 53116 7812 53172
rect 7644 53004 7700 53060
rect 7532 51324 7588 51380
rect 7308 51212 7364 51268
rect 7308 50594 7364 50596
rect 7308 50542 7310 50594
rect 7310 50542 7362 50594
rect 7362 50542 7364 50594
rect 7308 50540 7364 50542
rect 7644 50540 7700 50596
rect 7308 49084 7364 49140
rect 8428 53170 8484 53172
rect 8428 53118 8430 53170
rect 8430 53118 8482 53170
rect 8482 53118 8484 53170
rect 8428 53116 8484 53118
rect 8092 52834 8148 52836
rect 8092 52782 8094 52834
rect 8094 52782 8146 52834
rect 8146 52782 8148 52834
rect 8092 52780 8148 52782
rect 7868 50428 7924 50484
rect 12124 53506 12180 53508
rect 12124 53454 12126 53506
rect 12126 53454 12178 53506
rect 12178 53454 12180 53506
rect 12124 53452 12180 53454
rect 8988 51996 9044 52052
rect 9660 51996 9716 52052
rect 11116 51996 11172 52052
rect 10444 51884 10500 51940
rect 8540 51266 8596 51268
rect 8540 51214 8542 51266
rect 8542 51214 8594 51266
rect 8594 51214 8596 51266
rect 8540 51212 8596 51214
rect 8092 49644 8148 49700
rect 7532 48802 7588 48804
rect 7532 48750 7534 48802
rect 7534 48750 7586 48802
rect 7586 48750 7588 48802
rect 7532 48748 7588 48750
rect 7196 47964 7252 48020
rect 7196 46508 7252 46564
rect 6412 45666 6468 45668
rect 6412 45614 6414 45666
rect 6414 45614 6466 45666
rect 6466 45614 6468 45666
rect 6412 45612 6468 45614
rect 6860 45666 6916 45668
rect 6860 45614 6862 45666
rect 6862 45614 6914 45666
rect 6914 45614 6916 45666
rect 6860 45612 6916 45614
rect 7420 45612 7476 45668
rect 6748 44434 6804 44436
rect 6748 44382 6750 44434
rect 6750 44382 6802 44434
rect 6802 44382 6804 44434
rect 6748 44380 6804 44382
rect 7420 44380 7476 44436
rect 6524 44322 6580 44324
rect 6524 44270 6526 44322
rect 6526 44270 6578 44322
rect 6578 44270 6580 44322
rect 6524 44268 6580 44270
rect 6076 43932 6132 43988
rect 6412 43036 6468 43092
rect 6188 42754 6244 42756
rect 6188 42702 6190 42754
rect 6190 42702 6242 42754
rect 6242 42702 6244 42754
rect 6188 42700 6244 42702
rect 5852 39730 5908 39732
rect 5852 39678 5854 39730
rect 5854 39678 5906 39730
rect 5906 39678 5908 39730
rect 5852 39676 5908 39678
rect 6076 39116 6132 39172
rect 5740 38556 5796 38612
rect 5852 38220 5908 38276
rect 6860 43932 6916 43988
rect 6524 42364 6580 42420
rect 6748 42866 6804 42868
rect 6748 42814 6750 42866
rect 6750 42814 6802 42866
rect 6802 42814 6804 42866
rect 6748 42812 6804 42814
rect 6748 41804 6804 41860
rect 6300 38556 6356 38612
rect 6300 38220 6356 38276
rect 5516 36540 5572 36596
rect 5740 36540 5796 36596
rect 4956 34972 5012 35028
rect 4844 34242 4900 34244
rect 4844 34190 4846 34242
rect 4846 34190 4898 34242
rect 4898 34190 4900 34242
rect 4844 34188 4900 34190
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4508 33516 4564 33572
rect 4172 33346 4228 33348
rect 4172 33294 4174 33346
rect 4174 33294 4226 33346
rect 4226 33294 4228 33346
rect 4172 33292 4228 33294
rect 4172 30994 4228 30996
rect 4172 30942 4174 30994
rect 4174 30942 4226 30994
rect 4226 30942 4228 30994
rect 4172 30940 4228 30942
rect 3724 30156 3780 30212
rect 3836 28140 3892 28196
rect 4172 29932 4228 29988
rect 4060 28028 4116 28084
rect 4172 29426 4228 29428
rect 4172 29374 4174 29426
rect 4174 29374 4226 29426
rect 4226 29374 4228 29426
rect 4172 29372 4228 29374
rect 3724 27468 3780 27524
rect 4172 27244 4228 27300
rect 3724 26908 3780 26964
rect 4060 26514 4116 26516
rect 4060 26462 4062 26514
rect 4062 26462 4114 26514
rect 4114 26462 4116 26514
rect 4060 26460 4116 26462
rect 3388 24780 3444 24836
rect 3052 21586 3108 21588
rect 3052 21534 3054 21586
rect 3054 21534 3106 21586
rect 3106 21534 3108 21586
rect 3052 21532 3108 21534
rect 1932 18956 1988 19012
rect 2044 18620 2100 18676
rect 1708 17724 1764 17780
rect 1708 13468 1764 13524
rect 2044 17836 2100 17892
rect 2044 14642 2100 14644
rect 2044 14590 2046 14642
rect 2046 14590 2098 14642
rect 2098 14590 2100 14642
rect 2044 14588 2100 14590
rect 1820 14252 1876 14308
rect 1708 12850 1764 12852
rect 1708 12798 1710 12850
rect 1710 12798 1762 12850
rect 1762 12798 1764 12850
rect 1708 12796 1764 12798
rect 1932 12796 1988 12852
rect 2268 14140 2324 14196
rect 3052 20130 3108 20132
rect 3052 20078 3054 20130
rect 3054 20078 3106 20130
rect 3106 20078 3108 20130
rect 3052 20076 3108 20078
rect 3948 24556 4004 24612
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4844 32172 4900 32228
rect 4620 31948 4676 32004
rect 4396 31836 4452 31892
rect 4844 30994 4900 30996
rect 4844 30942 4846 30994
rect 4846 30942 4898 30994
rect 4898 30942 4900 30994
rect 4844 30940 4900 30942
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4732 29372 4788 29428
rect 5628 34748 5684 34804
rect 5628 34242 5684 34244
rect 5628 34190 5630 34242
rect 5630 34190 5682 34242
rect 5682 34190 5684 34242
rect 5628 34188 5684 34190
rect 5292 31164 5348 31220
rect 5068 31052 5124 31108
rect 4956 30268 5012 30324
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4732 28140 4788 28196
rect 4396 28082 4452 28084
rect 4396 28030 4398 28082
rect 4398 28030 4450 28082
rect 4450 28030 4452 28082
rect 4396 28028 4452 28030
rect 4396 27580 4452 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 5068 27356 5124 27412
rect 5292 27858 5348 27860
rect 5292 27806 5294 27858
rect 5294 27806 5346 27858
rect 5346 27806 5348 27858
rect 5292 27804 5348 27806
rect 5292 27634 5348 27636
rect 5292 27582 5294 27634
rect 5294 27582 5346 27634
rect 5346 27582 5348 27634
rect 5292 27580 5348 27582
rect 4844 26572 4900 26628
rect 5964 36652 6020 36708
rect 6188 37100 6244 37156
rect 6188 36540 6244 36596
rect 6188 36204 6244 36260
rect 6300 34242 6356 34244
rect 6300 34190 6302 34242
rect 6302 34190 6354 34242
rect 6354 34190 6356 34242
rect 6300 34188 6356 34190
rect 6076 34018 6132 34020
rect 6076 33966 6078 34018
rect 6078 33966 6130 34018
rect 6130 33966 6132 34018
rect 6076 33964 6132 33966
rect 6300 33628 6356 33684
rect 6300 33404 6356 33460
rect 5740 31948 5796 32004
rect 6300 31500 6356 31556
rect 6188 31276 6244 31332
rect 5516 31218 5572 31220
rect 5516 31166 5518 31218
rect 5518 31166 5570 31218
rect 5570 31166 5572 31218
rect 5516 31164 5572 31166
rect 5740 30994 5796 30996
rect 5740 30942 5742 30994
rect 5742 30942 5794 30994
rect 5794 30942 5796 30994
rect 5740 30940 5796 30942
rect 6524 36428 6580 36484
rect 9660 50428 9716 50484
rect 10556 50540 10612 50596
rect 9772 49644 9828 49700
rect 8540 48914 8596 48916
rect 8540 48862 8542 48914
rect 8542 48862 8594 48914
rect 8594 48862 8596 48914
rect 8540 48860 8596 48862
rect 9100 48860 9156 48916
rect 8876 48802 8932 48804
rect 8876 48750 8878 48802
rect 8878 48750 8930 48802
rect 8930 48750 8932 48802
rect 8876 48748 8932 48750
rect 8316 48076 8372 48132
rect 8876 48412 8932 48468
rect 9324 48412 9380 48468
rect 9660 48354 9716 48356
rect 9660 48302 9662 48354
rect 9662 48302 9714 48354
rect 9714 48302 9716 48354
rect 9660 48300 9716 48302
rect 8988 47404 9044 47460
rect 8316 46674 8372 46676
rect 8316 46622 8318 46674
rect 8318 46622 8370 46674
rect 8370 46622 8372 46674
rect 8316 46620 8372 46622
rect 7532 44268 7588 44324
rect 7196 43036 7252 43092
rect 7420 42700 7476 42756
rect 7084 42476 7140 42532
rect 7756 42924 7812 42980
rect 7532 41858 7588 41860
rect 7532 41806 7534 41858
rect 7534 41806 7586 41858
rect 7586 41806 7588 41858
rect 7532 41804 7588 41806
rect 7308 41692 7364 41748
rect 7084 40684 7140 40740
rect 6860 36988 6916 37044
rect 6748 36652 6804 36708
rect 6748 36482 6804 36484
rect 6748 36430 6750 36482
rect 6750 36430 6802 36482
rect 6802 36430 6804 36482
rect 6748 36428 6804 36430
rect 6972 35868 7028 35924
rect 7196 37996 7252 38052
rect 7308 37548 7364 37604
rect 7644 41132 7700 41188
rect 7868 40572 7924 40628
rect 7756 40460 7812 40516
rect 8428 45948 8484 46004
rect 9100 46002 9156 46004
rect 9100 45950 9102 46002
rect 9102 45950 9154 46002
rect 9154 45950 9156 46002
rect 9100 45948 9156 45950
rect 8652 43820 8708 43876
rect 8092 42364 8148 42420
rect 8092 38668 8148 38724
rect 7532 38220 7588 38276
rect 7644 38050 7700 38052
rect 7644 37998 7646 38050
rect 7646 37998 7698 38050
rect 7698 37998 7700 38050
rect 7644 37996 7700 37998
rect 7532 37884 7588 37940
rect 7532 37100 7588 37156
rect 7196 36370 7252 36372
rect 7196 36318 7198 36370
rect 7198 36318 7250 36370
rect 7250 36318 7252 36370
rect 7196 36316 7252 36318
rect 6636 34860 6692 34916
rect 6972 34802 7028 34804
rect 6972 34750 6974 34802
rect 6974 34750 7026 34802
rect 7026 34750 7028 34802
rect 6972 34748 7028 34750
rect 7196 34690 7252 34692
rect 7196 34638 7198 34690
rect 7198 34638 7250 34690
rect 7250 34638 7252 34690
rect 7196 34636 7252 34638
rect 6636 34188 6692 34244
rect 7084 33516 7140 33572
rect 7196 33964 7252 34020
rect 6972 33404 7028 33460
rect 6524 32562 6580 32564
rect 6524 32510 6526 32562
rect 6526 32510 6578 32562
rect 6578 32510 6580 32562
rect 6524 32508 6580 32510
rect 6636 32060 6692 32116
rect 6748 32732 6804 32788
rect 7084 32732 7140 32788
rect 8540 42812 8596 42868
rect 8428 42588 8484 42644
rect 9324 46956 9380 47012
rect 9996 48860 10052 48916
rect 9884 48412 9940 48468
rect 11452 51996 11508 52052
rect 11340 51772 11396 51828
rect 11564 51938 11620 51940
rect 11564 51886 11566 51938
rect 11566 51886 11618 51938
rect 11618 51886 11620 51938
rect 11564 51884 11620 51886
rect 11452 50706 11508 50708
rect 11452 50654 11454 50706
rect 11454 50654 11506 50706
rect 11506 50654 11508 50706
rect 11452 50652 11508 50654
rect 11340 50540 11396 50596
rect 11116 49698 11172 49700
rect 11116 49646 11118 49698
rect 11118 49646 11170 49698
rect 11170 49646 11172 49698
rect 11116 49644 11172 49646
rect 12572 53506 12628 53508
rect 12572 53454 12574 53506
rect 12574 53454 12626 53506
rect 12626 53454 12628 53506
rect 12572 53452 12628 53454
rect 12012 51772 12068 51828
rect 12684 50706 12740 50708
rect 12684 50654 12686 50706
rect 12686 50654 12738 50706
rect 12738 50654 12740 50706
rect 12684 50652 12740 50654
rect 12796 49698 12852 49700
rect 12796 49646 12798 49698
rect 12798 49646 12850 49698
rect 12850 49646 12852 49698
rect 12796 49644 12852 49646
rect 10332 48300 10388 48356
rect 10444 48130 10500 48132
rect 10444 48078 10446 48130
rect 10446 48078 10498 48130
rect 10498 48078 10500 48130
rect 10444 48076 10500 48078
rect 9772 46956 9828 47012
rect 10108 46786 10164 46788
rect 10108 46734 10110 46786
rect 10110 46734 10162 46786
rect 10162 46734 10164 46786
rect 10108 46732 10164 46734
rect 9212 42924 9268 42980
rect 8988 42194 9044 42196
rect 8988 42142 8990 42194
rect 8990 42142 9042 42194
rect 9042 42142 9044 42194
rect 8988 42140 9044 42142
rect 8540 40908 8596 40964
rect 8316 40348 8372 40404
rect 8428 37996 8484 38052
rect 10108 43708 10164 43764
rect 9660 42194 9716 42196
rect 9660 42142 9662 42194
rect 9662 42142 9714 42194
rect 9714 42142 9716 42194
rect 9660 42140 9716 42142
rect 10108 41970 10164 41972
rect 10108 41918 10110 41970
rect 10110 41918 10162 41970
rect 10162 41918 10164 41970
rect 10108 41916 10164 41918
rect 7532 36316 7588 36372
rect 7420 35868 7476 35924
rect 8204 37212 8260 37268
rect 8204 36988 8260 37044
rect 8540 37324 8596 37380
rect 8652 36988 8708 37044
rect 7756 34690 7812 34692
rect 7756 34638 7758 34690
rect 7758 34638 7810 34690
rect 7810 34638 7812 34690
rect 7756 34636 7812 34638
rect 8204 34860 8260 34916
rect 7532 33740 7588 33796
rect 7532 33516 7588 33572
rect 7084 32562 7140 32564
rect 7084 32510 7086 32562
rect 7086 32510 7138 32562
rect 7138 32510 7140 32562
rect 7084 32508 7140 32510
rect 6972 32172 7028 32228
rect 5964 30210 6020 30212
rect 5964 30158 5966 30210
rect 5966 30158 6018 30210
rect 6018 30158 6020 30210
rect 5964 30156 6020 30158
rect 5628 30044 5684 30100
rect 5740 29708 5796 29764
rect 4956 26460 5012 26516
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 6188 28642 6244 28644
rect 6188 28590 6190 28642
rect 6190 28590 6242 28642
rect 6242 28590 6244 28642
rect 6188 28588 6244 28590
rect 6076 28028 6132 28084
rect 4396 24834 4452 24836
rect 4396 24782 4398 24834
rect 4398 24782 4450 24834
rect 4450 24782 4452 24834
rect 4396 24780 4452 24782
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 3836 21084 3892 21140
rect 4284 23324 4340 23380
rect 3388 20018 3444 20020
rect 3388 19966 3390 20018
rect 3390 19966 3442 20018
rect 3442 19966 3444 20018
rect 3388 19964 3444 19966
rect 5740 27580 5796 27636
rect 6076 27298 6132 27300
rect 6076 27246 6078 27298
rect 6078 27246 6130 27298
rect 6130 27246 6132 27298
rect 6076 27244 6132 27246
rect 6412 29708 6468 29764
rect 6412 28812 6468 28868
rect 6412 27916 6468 27972
rect 5068 23996 5124 24052
rect 5628 25004 5684 25060
rect 5964 24834 6020 24836
rect 5964 24782 5966 24834
rect 5966 24782 6018 24834
rect 6018 24782 6020 24834
rect 5964 24780 6020 24782
rect 5628 23996 5684 24052
rect 5292 23660 5348 23716
rect 4956 23324 5012 23380
rect 5068 23436 5124 23492
rect 5740 23714 5796 23716
rect 5740 23662 5742 23714
rect 5742 23662 5794 23714
rect 5794 23662 5796 23714
rect 5740 23660 5796 23662
rect 5628 23436 5684 23492
rect 4844 23212 4900 23268
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4508 22594 4564 22596
rect 4508 22542 4510 22594
rect 4510 22542 4562 22594
rect 4562 22542 4564 22594
rect 4508 22540 4564 22542
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4284 20076 4340 20132
rect 2828 18620 2884 18676
rect 2716 18508 2772 18564
rect 2940 18396 2996 18452
rect 3500 19180 3556 19236
rect 3948 19234 4004 19236
rect 3948 19182 3950 19234
rect 3950 19182 4002 19234
rect 4002 19182 4004 19234
rect 3948 19180 4004 19182
rect 3724 18508 3780 18564
rect 3948 18620 4004 18676
rect 3500 18172 3556 18228
rect 2940 17276 2996 17332
rect 3388 17500 3444 17556
rect 4844 20076 4900 20132
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4844 18956 4900 19012
rect 4060 18172 4116 18228
rect 4508 18172 4564 18228
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 5852 23436 5908 23492
rect 5964 23660 6020 23716
rect 6188 26178 6244 26180
rect 6188 26126 6190 26178
rect 6190 26126 6242 26178
rect 6242 26126 6244 26178
rect 6188 26124 6244 26126
rect 6300 25004 6356 25060
rect 6860 31554 6916 31556
rect 6860 31502 6862 31554
rect 6862 31502 6914 31554
rect 6914 31502 6916 31554
rect 6860 31500 6916 31502
rect 7420 30716 7476 30772
rect 6860 29650 6916 29652
rect 6860 29598 6862 29650
rect 6862 29598 6914 29650
rect 6914 29598 6916 29650
rect 6860 29596 6916 29598
rect 7644 30098 7700 30100
rect 7644 30046 7646 30098
rect 7646 30046 7698 30098
rect 7698 30046 7700 30098
rect 7644 30044 7700 30046
rect 7532 29596 7588 29652
rect 7084 29426 7140 29428
rect 7084 29374 7086 29426
rect 7086 29374 7138 29426
rect 7138 29374 7140 29426
rect 7084 29372 7140 29374
rect 6636 28754 6692 28756
rect 6636 28702 6638 28754
rect 6638 28702 6690 28754
rect 6690 28702 6692 28754
rect 6636 28700 6692 28702
rect 6972 28642 7028 28644
rect 6972 28590 6974 28642
rect 6974 28590 7026 28642
rect 7026 28590 7028 28642
rect 6972 28588 7028 28590
rect 7980 33964 8036 34020
rect 8316 34130 8372 34132
rect 8316 34078 8318 34130
rect 8318 34078 8370 34130
rect 8370 34078 8372 34130
rect 8316 34076 8372 34078
rect 8092 33458 8148 33460
rect 8092 33406 8094 33458
rect 8094 33406 8146 33458
rect 8146 33406 8148 33458
rect 8092 33404 8148 33406
rect 9996 40402 10052 40404
rect 9996 40350 9998 40402
rect 9998 40350 10050 40402
rect 10050 40350 10052 40402
rect 9996 40348 10052 40350
rect 10108 40236 10164 40292
rect 9660 38834 9716 38836
rect 9660 38782 9662 38834
rect 9662 38782 9714 38834
rect 9714 38782 9716 38834
rect 9660 38780 9716 38782
rect 9436 38050 9492 38052
rect 9436 37998 9438 38050
rect 9438 37998 9490 38050
rect 9490 37998 9492 38050
rect 9436 37996 9492 37998
rect 9996 39564 10052 39620
rect 9996 39004 10052 39060
rect 9548 37548 9604 37604
rect 9884 37490 9940 37492
rect 9884 37438 9886 37490
rect 9886 37438 9938 37490
rect 9938 37438 9940 37490
rect 9884 37436 9940 37438
rect 8876 36652 8932 36708
rect 8652 34914 8708 34916
rect 8652 34862 8654 34914
rect 8654 34862 8706 34914
rect 8706 34862 8708 34914
rect 8652 34860 8708 34862
rect 9772 37378 9828 37380
rect 9772 37326 9774 37378
rect 9774 37326 9826 37378
rect 9826 37326 9828 37378
rect 9772 37324 9828 37326
rect 9996 36652 10052 36708
rect 9324 34860 9380 34916
rect 10332 43820 10388 43876
rect 10332 43596 10388 43652
rect 10556 43708 10612 43764
rect 10444 43372 10500 43428
rect 10332 42924 10388 42980
rect 10332 39564 10388 39620
rect 10892 43426 10948 43428
rect 10892 43374 10894 43426
rect 10894 43374 10946 43426
rect 10946 43374 10948 43426
rect 10892 43372 10948 43374
rect 11676 48412 11732 48468
rect 13580 53452 13636 53508
rect 14476 51996 14532 52052
rect 14924 52834 14980 52836
rect 14924 52782 14926 52834
rect 14926 52782 14978 52834
rect 14978 52782 14980 52834
rect 14924 52780 14980 52782
rect 12908 48412 12964 48468
rect 13244 50652 13300 50708
rect 14476 50706 14532 50708
rect 14476 50654 14478 50706
rect 14478 50654 14530 50706
rect 14530 50654 14532 50706
rect 14476 50652 14532 50654
rect 14252 50594 14308 50596
rect 14252 50542 14254 50594
rect 14254 50542 14306 50594
rect 14306 50542 14308 50594
rect 14252 50540 14308 50542
rect 13468 49756 13524 49812
rect 14028 48802 14084 48804
rect 14028 48750 14030 48802
rect 14030 48750 14082 48802
rect 14082 48750 14084 48802
rect 14028 48748 14084 48750
rect 11676 47346 11732 47348
rect 11676 47294 11678 47346
rect 11678 47294 11730 47346
rect 11730 47294 11732 47346
rect 11676 47292 11732 47294
rect 12236 47346 12292 47348
rect 12236 47294 12238 47346
rect 12238 47294 12290 47346
rect 12290 47294 12292 47346
rect 12236 47292 12292 47294
rect 10780 42924 10836 42980
rect 11116 46732 11172 46788
rect 10668 42812 10724 42868
rect 10556 42364 10612 42420
rect 13468 45836 13524 45892
rect 11340 43762 11396 43764
rect 11340 43710 11342 43762
rect 11342 43710 11394 43762
rect 11394 43710 11396 43762
rect 11340 43708 11396 43710
rect 11228 42476 11284 42532
rect 10332 38780 10388 38836
rect 10668 40908 10724 40964
rect 10668 39116 10724 39172
rect 10556 39058 10612 39060
rect 10556 39006 10558 39058
rect 10558 39006 10610 39058
rect 10610 39006 10612 39058
rect 10556 39004 10612 39006
rect 10444 38668 10500 38724
rect 10332 37996 10388 38052
rect 10556 37266 10612 37268
rect 10556 37214 10558 37266
rect 10558 37214 10610 37266
rect 10610 37214 10612 37266
rect 10556 37212 10612 37214
rect 10108 34748 10164 34804
rect 10220 35868 10276 35924
rect 8764 33404 8820 33460
rect 8988 32620 9044 32676
rect 8204 32450 8260 32452
rect 8204 32398 8206 32450
rect 8206 32398 8258 32450
rect 8258 32398 8260 32450
rect 8204 32396 8260 32398
rect 7980 30210 8036 30212
rect 7980 30158 7982 30210
rect 7982 30158 8034 30210
rect 8034 30158 8036 30210
rect 7980 30156 8036 30158
rect 11004 42140 11060 42196
rect 13580 43708 13636 43764
rect 13468 43036 13524 43092
rect 11788 42476 11844 42532
rect 12124 41916 12180 41972
rect 12572 42530 12628 42532
rect 12572 42478 12574 42530
rect 12574 42478 12626 42530
rect 12626 42478 12628 42530
rect 12572 42476 12628 42478
rect 11564 41186 11620 41188
rect 11564 41134 11566 41186
rect 11566 41134 11618 41186
rect 11618 41134 11620 41186
rect 11564 41132 11620 41134
rect 12684 41916 12740 41972
rect 12908 41916 12964 41972
rect 13916 43538 13972 43540
rect 13916 43486 13918 43538
rect 13918 43486 13970 43538
rect 13970 43486 13972 43538
rect 13916 43484 13972 43486
rect 14476 46508 14532 46564
rect 14476 42476 14532 42532
rect 14476 41970 14532 41972
rect 14476 41918 14478 41970
rect 14478 41918 14530 41970
rect 14530 41918 14532 41970
rect 14476 41916 14532 41918
rect 12684 41132 12740 41188
rect 13580 41132 13636 41188
rect 11340 40908 11396 40964
rect 12236 40962 12292 40964
rect 12236 40910 12238 40962
rect 12238 40910 12290 40962
rect 12290 40910 12292 40962
rect 12236 40908 12292 40910
rect 11004 40402 11060 40404
rect 11004 40350 11006 40402
rect 11006 40350 11058 40402
rect 11058 40350 11060 40402
rect 11004 40348 11060 40350
rect 12124 38780 12180 38836
rect 11116 37996 11172 38052
rect 14028 41186 14084 41188
rect 14028 41134 14030 41186
rect 14030 41134 14082 41186
rect 14082 41134 14084 41186
rect 14028 41132 14084 41134
rect 13580 40460 13636 40516
rect 12908 37996 12964 38052
rect 11004 37436 11060 37492
rect 11004 35868 11060 35924
rect 11564 37826 11620 37828
rect 11564 37774 11566 37826
rect 11566 37774 11618 37826
rect 11618 37774 11620 37826
rect 11564 37772 11620 37774
rect 12460 37772 12516 37828
rect 12908 36988 12964 37044
rect 14028 40348 14084 40404
rect 13916 39618 13972 39620
rect 13916 39566 13918 39618
rect 13918 39566 13970 39618
rect 13970 39566 13972 39618
rect 13916 39564 13972 39566
rect 13580 37996 13636 38052
rect 13692 38668 13748 38724
rect 11452 35756 11508 35812
rect 12684 35922 12740 35924
rect 12684 35870 12686 35922
rect 12686 35870 12738 35922
rect 12738 35870 12740 35922
rect 12684 35868 12740 35870
rect 12684 35644 12740 35700
rect 12908 35756 12964 35812
rect 10892 34972 10948 35028
rect 10556 34690 10612 34692
rect 10556 34638 10558 34690
rect 10558 34638 10610 34690
rect 10610 34638 10612 34690
rect 10556 34636 10612 34638
rect 10780 34914 10836 34916
rect 10780 34862 10782 34914
rect 10782 34862 10834 34914
rect 10834 34862 10836 34914
rect 10780 34860 10836 34862
rect 10780 34636 10836 34692
rect 9772 32620 9828 32676
rect 9548 32562 9604 32564
rect 9548 32510 9550 32562
rect 9550 32510 9602 32562
rect 9602 32510 9604 32562
rect 9548 32508 9604 32510
rect 10444 32562 10500 32564
rect 10444 32510 10446 32562
rect 10446 32510 10498 32562
rect 10498 32510 10500 32562
rect 10444 32508 10500 32510
rect 8204 30044 8260 30100
rect 8540 29596 8596 29652
rect 8092 28140 8148 28196
rect 7532 28028 7588 28084
rect 6636 27916 6692 27972
rect 6860 27858 6916 27860
rect 6860 27806 6862 27858
rect 6862 27806 6914 27858
rect 6914 27806 6916 27858
rect 6860 27804 6916 27806
rect 6636 27244 6692 27300
rect 7420 27858 7476 27860
rect 7420 27806 7422 27858
rect 7422 27806 7474 27858
rect 7474 27806 7476 27858
rect 7420 27804 7476 27806
rect 6860 27020 6916 27076
rect 6748 26514 6804 26516
rect 6748 26462 6750 26514
rect 6750 26462 6802 26514
rect 6802 26462 6804 26514
rect 6748 26460 6804 26462
rect 7196 26124 7252 26180
rect 7084 24780 7140 24836
rect 7196 25004 7252 25060
rect 6300 24668 6356 24724
rect 6972 24444 7028 24500
rect 5404 22988 5460 23044
rect 5740 22482 5796 22484
rect 5740 22430 5742 22482
rect 5742 22430 5794 22482
rect 5794 22430 5796 22482
rect 5740 22428 5796 22430
rect 5740 20130 5796 20132
rect 5740 20078 5742 20130
rect 5742 20078 5794 20130
rect 5794 20078 5796 20130
rect 5740 20076 5796 20078
rect 4956 18396 5012 18452
rect 5964 19628 6020 19684
rect 3724 17554 3780 17556
rect 3724 17502 3726 17554
rect 3726 17502 3778 17554
rect 3778 17502 3780 17554
rect 3724 17500 3780 17502
rect 3276 17276 3332 17332
rect 4844 17554 4900 17556
rect 4844 17502 4846 17554
rect 4846 17502 4898 17554
rect 4898 17502 4900 17554
rect 4844 17500 4900 17502
rect 4956 17442 5012 17444
rect 4956 17390 4958 17442
rect 4958 17390 5010 17442
rect 5010 17390 5012 17442
rect 4956 17388 5012 17390
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 2828 14642 2884 14644
rect 2828 14590 2830 14642
rect 2830 14590 2882 14642
rect 2882 14590 2884 14642
rect 2828 14588 2884 14590
rect 3164 14140 3220 14196
rect 5404 18562 5460 18564
rect 5404 18510 5406 18562
rect 5406 18510 5458 18562
rect 5458 18510 5460 18562
rect 5404 18508 5460 18510
rect 5180 18396 5236 18452
rect 5404 17724 5460 17780
rect 5068 17052 5124 17108
rect 5404 17276 5460 17332
rect 5852 18620 5908 18676
rect 6076 19010 6132 19012
rect 6076 18958 6078 19010
rect 6078 18958 6130 19010
rect 6130 18958 6132 19010
rect 6076 18956 6132 18958
rect 6524 23938 6580 23940
rect 6524 23886 6526 23938
rect 6526 23886 6578 23938
rect 6578 23886 6580 23938
rect 6524 23884 6580 23886
rect 6636 23826 6692 23828
rect 6636 23774 6638 23826
rect 6638 23774 6690 23826
rect 6690 23774 6692 23826
rect 6636 23772 6692 23774
rect 7196 24332 7252 24388
rect 7420 27186 7476 27188
rect 7420 27134 7422 27186
rect 7422 27134 7474 27186
rect 7474 27134 7476 27186
rect 7420 27132 7476 27134
rect 8092 27970 8148 27972
rect 8092 27918 8094 27970
rect 8094 27918 8146 27970
rect 8146 27918 8148 27970
rect 8092 27916 8148 27918
rect 7756 27132 7812 27188
rect 7644 27074 7700 27076
rect 7644 27022 7646 27074
rect 7646 27022 7698 27074
rect 7698 27022 7700 27074
rect 7644 27020 7700 27022
rect 8428 27020 8484 27076
rect 7532 26908 7588 26964
rect 7420 24722 7476 24724
rect 7420 24670 7422 24722
rect 7422 24670 7474 24722
rect 7474 24670 7476 24722
rect 7420 24668 7476 24670
rect 6860 23714 6916 23716
rect 6860 23662 6862 23714
rect 6862 23662 6914 23714
rect 6914 23662 6916 23714
rect 6860 23660 6916 23662
rect 7420 24220 7476 24276
rect 6524 23548 6580 23604
rect 6412 23436 6468 23492
rect 6300 22876 6356 22932
rect 6748 23436 6804 23492
rect 6748 22988 6804 23044
rect 6636 19628 6692 19684
rect 6300 18732 6356 18788
rect 6860 19010 6916 19012
rect 6860 18958 6862 19010
rect 6862 18958 6914 19010
rect 6914 18958 6916 19010
rect 6860 18956 6916 18958
rect 6524 18620 6580 18676
rect 6300 18450 6356 18452
rect 6300 18398 6302 18450
rect 6302 18398 6354 18450
rect 6354 18398 6356 18450
rect 6300 18396 6356 18398
rect 6524 18450 6580 18452
rect 6524 18398 6526 18450
rect 6526 18398 6578 18450
rect 6578 18398 6580 18450
rect 6524 18396 6580 18398
rect 6972 18450 7028 18452
rect 6972 18398 6974 18450
rect 6974 18398 7026 18450
rect 7026 18398 7028 18450
rect 6972 18396 7028 18398
rect 5852 17948 5908 18004
rect 6188 17948 6244 18004
rect 5740 17778 5796 17780
rect 5740 17726 5742 17778
rect 5742 17726 5794 17778
rect 5794 17726 5796 17778
rect 5740 17724 5796 17726
rect 5740 17052 5796 17108
rect 6076 17666 6132 17668
rect 6076 17614 6078 17666
rect 6078 17614 6130 17666
rect 6130 17614 6132 17666
rect 6076 17612 6132 17614
rect 6076 16994 6132 16996
rect 6076 16942 6078 16994
rect 6078 16942 6130 16994
rect 6130 16942 6132 16994
rect 6076 16940 6132 16942
rect 6076 16716 6132 16772
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 3724 14140 3780 14196
rect 3052 13468 3108 13524
rect 2492 13020 2548 13076
rect 2380 12908 2436 12964
rect 2828 12908 2884 12964
rect 2492 12850 2548 12852
rect 2492 12798 2494 12850
rect 2494 12798 2546 12850
rect 2546 12798 2548 12850
rect 2492 12796 2548 12798
rect 2716 10780 2772 10836
rect 3388 13074 3444 13076
rect 3388 13022 3390 13074
rect 3390 13022 3442 13074
rect 3442 13022 3444 13074
rect 3388 13020 3444 13022
rect 3388 10834 3444 10836
rect 3388 10782 3390 10834
rect 3390 10782 3442 10834
rect 3442 10782 3444 10834
rect 3388 10780 3444 10782
rect 4844 14306 4900 14308
rect 4844 14254 4846 14306
rect 4846 14254 4898 14306
rect 4898 14254 4900 14306
rect 4844 14252 4900 14254
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 6300 17554 6356 17556
rect 6300 17502 6302 17554
rect 6302 17502 6354 17554
rect 6354 17502 6356 17554
rect 6300 17500 6356 17502
rect 3724 12908 3780 12964
rect 4284 12962 4340 12964
rect 4284 12910 4286 12962
rect 4286 12910 4338 12962
rect 4338 12910 4340 12962
rect 4284 12908 4340 12910
rect 4956 12962 5012 12964
rect 4956 12910 4958 12962
rect 4958 12910 5010 12962
rect 5010 12910 5012 12962
rect 4956 12908 5012 12910
rect 5964 13804 6020 13860
rect 5180 12684 5236 12740
rect 4284 12290 4340 12292
rect 4284 12238 4286 12290
rect 4286 12238 4338 12290
rect 4338 12238 4340 12290
rect 4284 12236 4340 12238
rect 4732 12178 4788 12180
rect 4732 12126 4734 12178
rect 4734 12126 4786 12178
rect 4786 12126 4788 12178
rect 4732 12124 4788 12126
rect 4620 12066 4676 12068
rect 4620 12014 4622 12066
rect 4622 12014 4674 12066
rect 4674 12014 4676 12066
rect 4620 12012 4676 12014
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 3948 11564 4004 11620
rect 4844 11282 4900 11284
rect 4844 11230 4846 11282
rect 4846 11230 4898 11282
rect 4898 11230 4900 11282
rect 4844 11228 4900 11230
rect 3948 10834 4004 10836
rect 3948 10782 3950 10834
rect 3950 10782 4002 10834
rect 4002 10782 4004 10834
rect 3948 10780 4004 10782
rect 1932 7980 1988 8036
rect 1820 7868 1876 7924
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 5180 12236 5236 12292
rect 5068 12066 5124 12068
rect 5068 12014 5070 12066
rect 5070 12014 5122 12066
rect 5122 12014 5124 12066
rect 5068 12012 5124 12014
rect 5068 11506 5124 11508
rect 5068 11454 5070 11506
rect 5070 11454 5122 11506
rect 5122 11454 5124 11506
rect 5068 11452 5124 11454
rect 6188 13580 6244 13636
rect 5404 11900 5460 11956
rect 6748 17500 6804 17556
rect 6636 17388 6692 17444
rect 6636 16882 6692 16884
rect 6636 16830 6638 16882
rect 6638 16830 6690 16882
rect 6690 16830 6692 16882
rect 6636 16828 6692 16830
rect 6636 16604 6692 16660
rect 6860 14364 6916 14420
rect 6636 14252 6692 14308
rect 7308 23714 7364 23716
rect 7308 23662 7310 23714
rect 7310 23662 7362 23714
rect 7362 23662 7364 23714
rect 7308 23660 7364 23662
rect 7756 26850 7812 26852
rect 7756 26798 7758 26850
rect 7758 26798 7810 26850
rect 7810 26798 7812 26850
rect 7756 26796 7812 26798
rect 7644 26572 7700 26628
rect 7868 25676 7924 25732
rect 7756 25564 7812 25620
rect 8316 26850 8372 26852
rect 8316 26798 8318 26850
rect 8318 26798 8370 26850
rect 8370 26798 8372 26850
rect 8316 26796 8372 26798
rect 8316 26572 8372 26628
rect 7980 25506 8036 25508
rect 7980 25454 7982 25506
rect 7982 25454 8034 25506
rect 8034 25454 8036 25506
rect 7980 25452 8036 25454
rect 7868 25394 7924 25396
rect 7868 25342 7870 25394
rect 7870 25342 7922 25394
rect 7922 25342 7924 25394
rect 7868 25340 7924 25342
rect 8092 25282 8148 25284
rect 8092 25230 8094 25282
rect 8094 25230 8146 25282
rect 8146 25230 8148 25282
rect 8092 25228 8148 25230
rect 7644 24780 7700 24836
rect 7644 24444 7700 24500
rect 7756 24108 7812 24164
rect 7868 24332 7924 24388
rect 7868 23996 7924 24052
rect 7644 23436 7700 23492
rect 7756 23660 7812 23716
rect 7308 23266 7364 23268
rect 7308 23214 7310 23266
rect 7310 23214 7362 23266
rect 7362 23214 7364 23266
rect 7308 23212 7364 23214
rect 7420 23154 7476 23156
rect 7420 23102 7422 23154
rect 7422 23102 7474 23154
rect 7474 23102 7476 23154
rect 7420 23100 7476 23102
rect 7868 23436 7924 23492
rect 7196 22428 7252 22484
rect 8428 24332 8484 24388
rect 8316 24108 8372 24164
rect 8204 23996 8260 24052
rect 8092 23548 8148 23604
rect 8540 24108 8596 24164
rect 8428 23714 8484 23716
rect 8428 23662 8430 23714
rect 8430 23662 8482 23714
rect 8482 23662 8484 23714
rect 8428 23660 8484 23662
rect 8988 28812 9044 28868
rect 9212 27916 9268 27972
rect 8876 27132 8932 27188
rect 8764 27020 8820 27076
rect 8876 26514 8932 26516
rect 8876 26462 8878 26514
rect 8878 26462 8930 26514
rect 8930 26462 8932 26514
rect 8876 26460 8932 26462
rect 9100 25788 9156 25844
rect 8988 25618 9044 25620
rect 8988 25566 8990 25618
rect 8990 25566 9042 25618
rect 9042 25566 9044 25618
rect 8988 25564 9044 25566
rect 9884 29986 9940 29988
rect 9884 29934 9886 29986
rect 9886 29934 9938 29986
rect 9938 29934 9940 29986
rect 9884 29932 9940 29934
rect 9772 29426 9828 29428
rect 9772 29374 9774 29426
rect 9774 29374 9826 29426
rect 9826 29374 9828 29426
rect 9772 29372 9828 29374
rect 9884 28476 9940 28532
rect 9660 27916 9716 27972
rect 12796 35026 12852 35028
rect 12796 34974 12798 35026
rect 12798 34974 12850 35026
rect 12850 34974 12852 35026
rect 12796 34972 12852 34974
rect 10780 32508 10836 32564
rect 11788 34690 11844 34692
rect 11788 34638 11790 34690
rect 11790 34638 11842 34690
rect 11842 34638 11844 34690
rect 11788 34636 11844 34638
rect 12012 34690 12068 34692
rect 12012 34638 12014 34690
rect 12014 34638 12066 34690
rect 12066 34638 12068 34690
rect 12012 34636 12068 34638
rect 11116 32620 11172 32676
rect 11452 32396 11508 32452
rect 10556 30770 10612 30772
rect 10556 30718 10558 30770
rect 10558 30718 10610 30770
rect 10610 30718 10612 30770
rect 10556 30716 10612 30718
rect 10220 30098 10276 30100
rect 10220 30046 10222 30098
rect 10222 30046 10274 30098
rect 10274 30046 10276 30098
rect 10220 30044 10276 30046
rect 10668 30098 10724 30100
rect 10668 30046 10670 30098
rect 10670 30046 10722 30098
rect 10722 30046 10724 30098
rect 10668 30044 10724 30046
rect 11116 30098 11172 30100
rect 11116 30046 11118 30098
rect 11118 30046 11170 30098
rect 11170 30046 11172 30098
rect 11116 30044 11172 30046
rect 10556 29932 10612 29988
rect 10668 29650 10724 29652
rect 10668 29598 10670 29650
rect 10670 29598 10722 29650
rect 10722 29598 10724 29650
rect 10668 29596 10724 29598
rect 10332 29426 10388 29428
rect 10332 29374 10334 29426
rect 10334 29374 10386 29426
rect 10386 29374 10388 29426
rect 10332 29372 10388 29374
rect 11452 30604 11508 30660
rect 11452 29932 11508 29988
rect 11788 30044 11844 30100
rect 12012 33180 12068 33236
rect 12236 32674 12292 32676
rect 12236 32622 12238 32674
rect 12238 32622 12290 32674
rect 12290 32622 12292 32674
rect 12236 32620 12292 32622
rect 12124 30098 12180 30100
rect 12124 30046 12126 30098
rect 12126 30046 12178 30098
rect 12178 30046 12180 30098
rect 12124 30044 12180 30046
rect 12236 29986 12292 29988
rect 12236 29934 12238 29986
rect 12238 29934 12290 29986
rect 12290 29934 12292 29986
rect 12236 29932 12292 29934
rect 12348 29820 12404 29876
rect 10668 28812 10724 28868
rect 9660 26850 9716 26852
rect 9660 26798 9662 26850
rect 9662 26798 9714 26850
rect 9714 26798 9716 26850
rect 9660 26796 9716 26798
rect 8764 25340 8820 25396
rect 9212 24892 9268 24948
rect 8876 24834 8932 24836
rect 8876 24782 8878 24834
rect 8878 24782 8930 24834
rect 8930 24782 8932 24834
rect 8876 24780 8932 24782
rect 9548 24722 9604 24724
rect 9548 24670 9550 24722
rect 9550 24670 9602 24722
rect 9602 24670 9604 24722
rect 9548 24668 9604 24670
rect 9660 24610 9716 24612
rect 9660 24558 9662 24610
rect 9662 24558 9714 24610
rect 9714 24558 9716 24610
rect 9660 24556 9716 24558
rect 9100 24332 9156 24388
rect 8876 23996 8932 24052
rect 8316 23100 8372 23156
rect 8316 22540 8372 22596
rect 8876 23154 8932 23156
rect 8876 23102 8878 23154
rect 8878 23102 8930 23154
rect 8930 23102 8932 23154
rect 8876 23100 8932 23102
rect 7980 21756 8036 21812
rect 7980 21532 8036 21588
rect 9100 23436 9156 23492
rect 10220 27804 10276 27860
rect 10332 27356 10388 27412
rect 10556 27298 10612 27300
rect 10556 27246 10558 27298
rect 10558 27246 10610 27298
rect 10610 27246 10612 27298
rect 10556 27244 10612 27246
rect 11004 29036 11060 29092
rect 10108 27132 10164 27188
rect 10780 28700 10836 28756
rect 11788 28700 11844 28756
rect 10220 25788 10276 25844
rect 10108 25282 10164 25284
rect 10108 25230 10110 25282
rect 10110 25230 10162 25282
rect 10162 25230 10164 25282
rect 10108 25228 10164 25230
rect 10332 25506 10388 25508
rect 10332 25454 10334 25506
rect 10334 25454 10386 25506
rect 10386 25454 10388 25506
rect 10332 25452 10388 25454
rect 9884 24220 9940 24276
rect 10108 23884 10164 23940
rect 9772 23772 9828 23828
rect 10668 25116 10724 25172
rect 9212 23212 9268 23268
rect 9100 23100 9156 23156
rect 9772 22540 9828 22596
rect 9548 21810 9604 21812
rect 9548 21758 9550 21810
rect 9550 21758 9602 21810
rect 9602 21758 9604 21810
rect 9548 21756 9604 21758
rect 10444 23154 10500 23156
rect 10444 23102 10446 23154
rect 10446 23102 10498 23154
rect 10498 23102 10500 23154
rect 10444 23100 10500 23102
rect 10332 21644 10388 21700
rect 9772 21586 9828 21588
rect 9772 21534 9774 21586
rect 9774 21534 9826 21586
rect 9826 21534 9828 21586
rect 9772 21532 9828 21534
rect 9324 20914 9380 20916
rect 9324 20862 9326 20914
rect 9326 20862 9378 20914
rect 9378 20862 9380 20914
rect 9324 20860 9380 20862
rect 7196 18508 7252 18564
rect 7196 17948 7252 18004
rect 7308 18396 7364 18452
rect 9660 20524 9716 20580
rect 8092 18620 8148 18676
rect 8204 18732 8260 18788
rect 7756 18284 7812 18340
rect 7980 18508 8036 18564
rect 8092 18396 8148 18452
rect 7868 17724 7924 17780
rect 7532 17666 7588 17668
rect 7532 17614 7534 17666
rect 7534 17614 7586 17666
rect 7586 17614 7588 17666
rect 7532 17612 7588 17614
rect 7980 17948 8036 18004
rect 7308 17388 7364 17444
rect 8316 18284 8372 18340
rect 8652 18732 8708 18788
rect 8540 18396 8596 18452
rect 9436 18620 9492 18676
rect 9660 18562 9716 18564
rect 9660 18510 9662 18562
rect 9662 18510 9714 18562
rect 9714 18510 9716 18562
rect 9660 18508 9716 18510
rect 9436 17948 9492 18004
rect 8092 17500 8148 17556
rect 7756 17164 7812 17220
rect 8204 17164 8260 17220
rect 8428 17500 8484 17556
rect 8092 17052 8148 17108
rect 7532 16882 7588 16884
rect 7532 16830 7534 16882
rect 7534 16830 7586 16882
rect 7586 16830 7588 16882
rect 7532 16828 7588 16830
rect 8540 17666 8596 17668
rect 8540 17614 8542 17666
rect 8542 17614 8594 17666
rect 8594 17614 8596 17666
rect 8540 17612 8596 17614
rect 9324 17612 9380 17668
rect 9212 17554 9268 17556
rect 9212 17502 9214 17554
rect 9214 17502 9266 17554
rect 9266 17502 9268 17554
rect 9212 17500 9268 17502
rect 9772 17052 9828 17108
rect 8540 16940 8596 16996
rect 8428 16828 8484 16884
rect 10780 25340 10836 25396
rect 10892 24444 10948 24500
rect 10668 22540 10724 22596
rect 10892 22540 10948 22596
rect 10892 21644 10948 21700
rect 11116 28476 11172 28532
rect 11900 27916 11956 27972
rect 11788 27356 11844 27412
rect 11340 27186 11396 27188
rect 11340 27134 11342 27186
rect 11342 27134 11394 27186
rect 11394 27134 11396 27186
rect 11340 27132 11396 27134
rect 11676 26908 11732 26964
rect 11900 27244 11956 27300
rect 11676 25564 11732 25620
rect 11228 25394 11284 25396
rect 11228 25342 11230 25394
rect 11230 25342 11282 25394
rect 11282 25342 11284 25394
rect 11228 25340 11284 25342
rect 11340 25116 11396 25172
rect 11900 25116 11956 25172
rect 11228 24108 11284 24164
rect 11676 23548 11732 23604
rect 11676 22540 11732 22596
rect 11228 22428 11284 22484
rect 11004 20860 11060 20916
rect 10780 17836 10836 17892
rect 10556 16716 10612 16772
rect 10668 16044 10724 16100
rect 10556 15314 10612 15316
rect 10556 15262 10558 15314
rect 10558 15262 10610 15314
rect 10610 15262 10612 15314
rect 10556 15260 10612 15262
rect 9772 15148 9828 15204
rect 10444 14924 10500 14980
rect 9884 14530 9940 14532
rect 9884 14478 9886 14530
rect 9886 14478 9938 14530
rect 9938 14478 9940 14530
rect 9884 14476 9940 14478
rect 7420 14364 7476 14420
rect 6412 13244 6468 13300
rect 6524 13804 6580 13860
rect 5740 12124 5796 12180
rect 5628 11564 5684 11620
rect 5516 11452 5572 11508
rect 5852 12908 5908 12964
rect 6076 12962 6132 12964
rect 6076 12910 6078 12962
rect 6078 12910 6130 12962
rect 6130 12910 6132 12962
rect 6076 12908 6132 12910
rect 6748 13580 6804 13636
rect 6188 12460 6244 12516
rect 6076 12124 6132 12180
rect 5852 11900 5908 11956
rect 6188 11394 6244 11396
rect 6188 11342 6190 11394
rect 6190 11342 6242 11394
rect 6242 11342 6244 11394
rect 6188 11340 6244 11342
rect 6412 12460 6468 12516
rect 5852 11228 5908 11284
rect 5292 10556 5348 10612
rect 6076 10610 6132 10612
rect 6076 10558 6078 10610
rect 6078 10558 6130 10610
rect 6130 10558 6132 10610
rect 6076 10556 6132 10558
rect 3500 9436 3556 9492
rect 2716 9266 2772 9268
rect 2716 9214 2718 9266
rect 2718 9214 2770 9266
rect 2770 9214 2772 9266
rect 2716 9212 2772 9214
rect 2268 6860 2324 6916
rect 1708 6690 1764 6692
rect 1708 6638 1710 6690
rect 1710 6638 1762 6690
rect 1762 6638 1764 6690
rect 1708 6636 1764 6638
rect 2044 6636 2100 6692
rect 1820 6466 1876 6468
rect 1820 6414 1822 6466
rect 1822 6414 1874 6466
rect 1874 6414 1876 6466
rect 1820 6412 1876 6414
rect 2268 6412 2324 6468
rect 2716 8652 2772 8708
rect 2604 7980 2660 8036
rect 3052 7196 3108 7252
rect 2940 6524 2996 6580
rect 3612 8988 3668 9044
rect 3276 8652 3332 8708
rect 3388 6524 3444 6580
rect 4172 8204 4228 8260
rect 3836 6690 3892 6692
rect 3836 6638 3838 6690
rect 3838 6638 3890 6690
rect 3890 6638 3892 6690
rect 3836 6636 3892 6638
rect 6972 13522 7028 13524
rect 6972 13470 6974 13522
rect 6974 13470 7026 13522
rect 7026 13470 7028 13522
rect 6972 13468 7028 13470
rect 6748 12236 6804 12292
rect 6860 13074 6916 13076
rect 6860 13022 6862 13074
rect 6862 13022 6914 13074
rect 6914 13022 6916 13074
rect 6860 13020 6916 13022
rect 6524 12124 6580 12180
rect 6860 11788 6916 11844
rect 6524 11618 6580 11620
rect 6524 11566 6526 11618
rect 6526 11566 6578 11618
rect 6578 11566 6580 11618
rect 6524 11564 6580 11566
rect 6860 11506 6916 11508
rect 6860 11454 6862 11506
rect 6862 11454 6914 11506
rect 6914 11454 6916 11506
rect 6860 11452 6916 11454
rect 6636 11228 6692 11284
rect 6972 11394 7028 11396
rect 6972 11342 6974 11394
rect 6974 11342 7026 11394
rect 7026 11342 7028 11394
rect 6972 11340 7028 11342
rect 6972 10668 7028 10724
rect 6860 10556 6916 10612
rect 5852 9154 5908 9156
rect 5852 9102 5854 9154
rect 5854 9102 5906 9154
rect 5906 9102 5908 9154
rect 5852 9100 5908 9102
rect 6748 10108 6804 10164
rect 5964 9042 6020 9044
rect 5964 8990 5966 9042
rect 5966 8990 6018 9042
rect 6018 8990 6020 9042
rect 5964 8988 6020 8990
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4508 8370 4564 8372
rect 4508 8318 4510 8370
rect 4510 8318 4562 8370
rect 4562 8318 4564 8370
rect 4508 8316 4564 8318
rect 4956 8204 5012 8260
rect 4508 7474 4564 7476
rect 4508 7422 4510 7474
rect 4510 7422 4562 7474
rect 4562 7422 4564 7474
rect 4508 7420 4564 7422
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 5852 8258 5908 8260
rect 5852 8206 5854 8258
rect 5854 8206 5906 8258
rect 5906 8206 5908 8258
rect 5852 8204 5908 8206
rect 5404 7250 5460 7252
rect 5404 7198 5406 7250
rect 5406 7198 5458 7250
rect 5458 7198 5460 7250
rect 5404 7196 5460 7198
rect 4508 6578 4564 6580
rect 4508 6526 4510 6578
rect 4510 6526 4562 6578
rect 4562 6526 4564 6578
rect 4508 6524 4564 6526
rect 3948 6466 4004 6468
rect 3948 6414 3950 6466
rect 3950 6414 4002 6466
rect 4002 6414 4004 6466
rect 3948 6412 4004 6414
rect 3612 3612 3668 3668
rect 1708 3276 1764 3332
rect 3388 3276 3444 3332
rect 4284 6412 4340 6468
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 5068 6578 5124 6580
rect 5068 6526 5070 6578
rect 5070 6526 5122 6578
rect 5122 6526 5124 6578
rect 5068 6524 5124 6526
rect 5964 6578 6020 6580
rect 5964 6526 5966 6578
rect 5966 6526 6018 6578
rect 6018 6526 6020 6578
rect 5964 6524 6020 6526
rect 6076 4956 6132 5012
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 4620 3666 4676 3668
rect 4620 3614 4622 3666
rect 4622 3614 4674 3666
rect 4674 3614 4676 3666
rect 4620 3612 4676 3614
rect 6524 9042 6580 9044
rect 6524 8990 6526 9042
rect 6526 8990 6578 9042
rect 6578 8990 6580 9042
rect 6524 8988 6580 8990
rect 7308 12236 7364 12292
rect 7196 11900 7252 11956
rect 10444 14476 10500 14532
rect 10556 14140 10612 14196
rect 9660 13634 9716 13636
rect 9660 13582 9662 13634
rect 9662 13582 9714 13634
rect 9714 13582 9716 13634
rect 9660 13580 9716 13582
rect 8652 12962 8708 12964
rect 8652 12910 8654 12962
rect 8654 12910 8706 12962
rect 8706 12910 8708 12962
rect 8652 12908 8708 12910
rect 7420 10556 7476 10612
rect 7756 11676 7812 11732
rect 11004 18450 11060 18452
rect 11004 18398 11006 18450
rect 11006 18398 11058 18450
rect 11058 18398 11060 18450
rect 11004 18396 11060 18398
rect 11900 22428 11956 22484
rect 11564 21698 11620 21700
rect 11564 21646 11566 21698
rect 11566 21646 11618 21698
rect 11618 21646 11620 21698
rect 11564 21644 11620 21646
rect 11788 18450 11844 18452
rect 11788 18398 11790 18450
rect 11790 18398 11842 18450
rect 11842 18398 11844 18450
rect 11788 18396 11844 18398
rect 11004 16210 11060 16212
rect 11004 16158 11006 16210
rect 11006 16158 11058 16210
rect 11058 16158 11060 16210
rect 11004 16156 11060 16158
rect 12124 26908 12180 26964
rect 12908 30716 12964 30772
rect 12796 29820 12852 29876
rect 12684 28754 12740 28756
rect 12684 28702 12686 28754
rect 12686 28702 12738 28754
rect 12738 28702 12740 28754
rect 12684 28700 12740 28702
rect 12796 28588 12852 28644
rect 13580 35196 13636 35252
rect 13580 34690 13636 34692
rect 13580 34638 13582 34690
rect 13582 34638 13634 34690
rect 13634 34638 13636 34690
rect 13580 34636 13636 34638
rect 13244 29932 13300 29988
rect 13244 29426 13300 29428
rect 13244 29374 13246 29426
rect 13246 29374 13298 29426
rect 13298 29374 13300 29426
rect 13244 29372 13300 29374
rect 13020 29036 13076 29092
rect 13356 28700 13412 28756
rect 13580 28642 13636 28644
rect 13580 28590 13582 28642
rect 13582 28590 13634 28642
rect 13634 28590 13636 28642
rect 13580 28588 13636 28590
rect 14476 40236 14532 40292
rect 14924 50540 14980 50596
rect 15596 60396 15652 60452
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 19180 73052 19236 73108
rect 17724 71596 17780 71652
rect 17724 70588 17780 70644
rect 19180 71148 19236 71204
rect 18508 69298 18564 69300
rect 18508 69246 18510 69298
rect 18510 69246 18562 69298
rect 18562 69246 18564 69298
rect 18508 69244 18564 69246
rect 19068 69298 19124 69300
rect 19068 69246 19070 69298
rect 19070 69246 19122 69298
rect 19122 69246 19124 69298
rect 19068 69244 19124 69246
rect 18956 68796 19012 68852
rect 18284 67058 18340 67060
rect 18284 67006 18286 67058
rect 18286 67006 18338 67058
rect 18338 67006 18340 67058
rect 18284 67004 18340 67006
rect 18732 65378 18788 65380
rect 18732 65326 18734 65378
rect 18734 65326 18786 65378
rect 18786 65326 18788 65378
rect 18732 65324 18788 65326
rect 16828 63084 16884 63140
rect 17724 62466 17780 62468
rect 17724 62414 17726 62466
rect 17726 62414 17778 62466
rect 17778 62414 17780 62466
rect 17724 62412 17780 62414
rect 17948 62188 18004 62244
rect 21644 75682 21700 75684
rect 21644 75630 21646 75682
rect 21646 75630 21698 75682
rect 21698 75630 21700 75682
rect 21644 75628 21700 75630
rect 22428 75682 22484 75684
rect 22428 75630 22430 75682
rect 22430 75630 22482 75682
rect 22482 75630 22484 75682
rect 22428 75628 22484 75630
rect 20636 73052 20692 73108
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 20300 71596 20356 71652
rect 20748 71148 20804 71204
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20860 70588 20916 70644
rect 20044 70532 20100 70534
rect 21644 71202 21700 71204
rect 21644 71150 21646 71202
rect 21646 71150 21698 71202
rect 21698 71150 21700 71202
rect 21644 71148 21700 71150
rect 22428 70588 22484 70644
rect 22876 70588 22932 70644
rect 21532 69356 21588 69412
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 19740 68850 19796 68852
rect 19740 68798 19742 68850
rect 19742 68798 19794 68850
rect 19794 68798 19796 68850
rect 19740 68796 19796 68798
rect 20860 68626 20916 68628
rect 20860 68574 20862 68626
rect 20862 68574 20914 68626
rect 20914 68574 20916 68626
rect 20860 68572 20916 68574
rect 19516 68012 19572 68068
rect 20300 68066 20356 68068
rect 20300 68014 20302 68066
rect 20302 68014 20354 68066
rect 20354 68014 20356 68066
rect 20300 68012 20356 68014
rect 22540 69410 22596 69412
rect 22540 69358 22542 69410
rect 22542 69358 22594 69410
rect 22594 69358 22596 69410
rect 22540 69356 22596 69358
rect 24220 75682 24276 75684
rect 24220 75630 24222 75682
rect 24222 75630 24274 75682
rect 24274 75630 24276 75682
rect 24220 75628 24276 75630
rect 26796 75740 26852 75796
rect 24108 74844 24164 74900
rect 25228 75628 25284 75684
rect 28140 75794 28196 75796
rect 28140 75742 28142 75794
rect 28142 75742 28194 75794
rect 28194 75742 28196 75794
rect 28140 75740 28196 75742
rect 29372 75740 29428 75796
rect 25228 74898 25284 74900
rect 25228 74846 25230 74898
rect 25230 74846 25282 74898
rect 25282 74846 25284 74898
rect 25228 74844 25284 74846
rect 24220 73164 24276 73220
rect 25228 73164 25284 73220
rect 23660 71596 23716 71652
rect 21868 68572 21924 68628
rect 21980 68796 22036 68852
rect 21868 68402 21924 68404
rect 21868 68350 21870 68402
rect 21870 68350 21922 68402
rect 21922 68350 21924 68402
rect 21868 68348 21924 68350
rect 21420 68012 21476 68068
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 18956 63250 19012 63252
rect 18956 63198 18958 63250
rect 18958 63198 19010 63250
rect 19010 63198 19012 63250
rect 18956 63196 19012 63198
rect 18508 62466 18564 62468
rect 18508 62414 18510 62466
rect 18510 62414 18562 62466
rect 18562 62414 18564 62466
rect 18508 62412 18564 62414
rect 18508 62188 18564 62244
rect 15708 59890 15764 59892
rect 15708 59838 15710 59890
rect 15710 59838 15762 59890
rect 15762 59838 15764 59890
rect 15708 59836 15764 59838
rect 17500 60396 17556 60452
rect 18284 60396 18340 60452
rect 15596 59052 15652 59108
rect 16268 59276 16324 59332
rect 17388 59330 17444 59332
rect 17388 59278 17390 59330
rect 17390 59278 17442 59330
rect 17442 59278 17444 59330
rect 17388 59276 17444 59278
rect 18060 59836 18116 59892
rect 18620 61458 18676 61460
rect 18620 61406 18622 61458
rect 18622 61406 18674 61458
rect 18674 61406 18676 61458
rect 18620 61404 18676 61406
rect 18508 59500 18564 59556
rect 19628 63138 19684 63140
rect 19628 63086 19630 63138
rect 19630 63086 19682 63138
rect 19682 63086 19684 63138
rect 19628 63084 19684 63086
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 18956 62466 19012 62468
rect 18956 62414 18958 62466
rect 18958 62414 19010 62466
rect 19010 62414 19012 62466
rect 18956 62412 19012 62414
rect 19628 62466 19684 62468
rect 19628 62414 19630 62466
rect 19630 62414 19682 62466
rect 19682 62414 19684 62466
rect 19628 62412 19684 62414
rect 20300 62412 20356 62468
rect 20412 62860 20468 62916
rect 19516 61404 19572 61460
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 19740 59948 19796 60004
rect 19516 59500 19572 59556
rect 18396 59218 18452 59220
rect 18396 59166 18398 59218
rect 18398 59166 18450 59218
rect 18450 59166 18452 59218
rect 18396 59164 18452 59166
rect 18284 59052 18340 59108
rect 17948 57596 18004 57652
rect 18284 58268 18340 58324
rect 17052 56812 17108 56868
rect 18284 57148 18340 57204
rect 18396 58156 18452 58212
rect 17724 56588 17780 56644
rect 18172 56642 18228 56644
rect 18172 56590 18174 56642
rect 18174 56590 18226 56642
rect 18226 56590 18228 56642
rect 18172 56588 18228 56590
rect 18508 57650 18564 57652
rect 18508 57598 18510 57650
rect 18510 57598 18562 57650
rect 18562 57598 18564 57650
rect 18508 57596 18564 57598
rect 18844 59106 18900 59108
rect 18844 59054 18846 59106
rect 18846 59054 18898 59106
rect 18898 59054 18900 59106
rect 18844 59052 18900 59054
rect 19292 59052 19348 59108
rect 18844 58322 18900 58324
rect 18844 58270 18846 58322
rect 18846 58270 18898 58322
rect 18898 58270 18900 58322
rect 18844 58268 18900 58270
rect 19068 58210 19124 58212
rect 19068 58158 19070 58210
rect 19070 58158 19122 58210
rect 19122 58158 19124 58210
rect 19068 58156 19124 58158
rect 18620 56812 18676 56868
rect 18508 56588 18564 56644
rect 16380 54236 16436 54292
rect 17836 55020 17892 55076
rect 18508 55074 18564 55076
rect 18508 55022 18510 55074
rect 18510 55022 18562 55074
rect 18562 55022 18564 55074
rect 18508 55020 18564 55022
rect 18732 54684 18788 54740
rect 18844 57148 18900 57204
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 19628 59106 19684 59108
rect 19628 59054 19630 59106
rect 19630 59054 19682 59106
rect 19682 59054 19684 59106
rect 19628 59052 19684 59054
rect 19852 58322 19908 58324
rect 19852 58270 19854 58322
rect 19854 58270 19906 58322
rect 19906 58270 19908 58322
rect 19852 58268 19908 58270
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 19740 57036 19796 57092
rect 19852 57708 19908 57764
rect 19852 56812 19908 56868
rect 20076 56700 20132 56756
rect 19068 56588 19124 56644
rect 18172 54236 18228 54292
rect 18956 53676 19012 53732
rect 15372 52780 15428 52836
rect 18284 53564 18340 53620
rect 17948 51436 18004 51492
rect 15820 50706 15876 50708
rect 15820 50654 15822 50706
rect 15822 50654 15874 50706
rect 15874 50654 15876 50706
rect 15820 50652 15876 50654
rect 16156 50540 16212 50596
rect 14924 49644 14980 49700
rect 14924 48860 14980 48916
rect 14700 48524 14756 48580
rect 15596 49644 15652 49700
rect 17724 50428 17780 50484
rect 16156 49698 16212 49700
rect 16156 49646 16158 49698
rect 16158 49646 16210 49698
rect 16210 49646 16212 49698
rect 16156 49644 16212 49646
rect 16604 49756 16660 49812
rect 15484 48748 15540 48804
rect 16156 48466 16212 48468
rect 16156 48414 16158 48466
rect 16158 48414 16210 48466
rect 16210 48414 16212 48466
rect 16156 48412 16212 48414
rect 15372 46562 15428 46564
rect 15372 46510 15374 46562
rect 15374 46510 15426 46562
rect 15426 46510 15428 46562
rect 15372 46508 15428 46510
rect 16156 46620 16212 46676
rect 14924 45836 14980 45892
rect 14812 43484 14868 43540
rect 15708 45666 15764 45668
rect 15708 45614 15710 45666
rect 15710 45614 15762 45666
rect 15762 45614 15764 45666
rect 15708 45612 15764 45614
rect 16156 45612 16212 45668
rect 17612 48748 17668 48804
rect 16716 48412 16772 48468
rect 16828 47234 16884 47236
rect 16828 47182 16830 47234
rect 16830 47182 16882 47234
rect 16882 47182 16884 47234
rect 16828 47180 16884 47182
rect 16604 45724 16660 45780
rect 16268 44380 16324 44436
rect 15372 41916 15428 41972
rect 16380 44044 16436 44100
rect 16044 43596 16100 43652
rect 14812 39564 14868 39620
rect 14924 40236 14980 40292
rect 14700 39506 14756 39508
rect 14700 39454 14702 39506
rect 14702 39454 14754 39506
rect 14754 39454 14756 39506
rect 14700 39452 14756 39454
rect 14364 37154 14420 37156
rect 14364 37102 14366 37154
rect 14366 37102 14418 37154
rect 14418 37102 14420 37154
rect 14364 37100 14420 37102
rect 13804 33234 13860 33236
rect 13804 33182 13806 33234
rect 13806 33182 13858 33234
rect 13858 33182 13860 33234
rect 13804 33180 13860 33182
rect 14700 37996 14756 38052
rect 14700 36876 14756 36932
rect 14700 36482 14756 36484
rect 14700 36430 14702 36482
rect 14702 36430 14754 36482
rect 14754 36430 14756 36482
rect 14700 36428 14756 36430
rect 14700 32396 14756 32452
rect 13804 30210 13860 30212
rect 13804 30158 13806 30210
rect 13806 30158 13858 30210
rect 13858 30158 13860 30210
rect 13804 30156 13860 30158
rect 14476 30156 14532 30212
rect 14028 30098 14084 30100
rect 14028 30046 14030 30098
rect 14030 30046 14082 30098
rect 14082 30046 14084 30098
rect 14028 30044 14084 30046
rect 14476 28812 14532 28868
rect 14140 27970 14196 27972
rect 14140 27918 14142 27970
rect 14142 27918 14194 27970
rect 14194 27918 14196 27970
rect 14140 27916 14196 27918
rect 12572 25618 12628 25620
rect 12572 25566 12574 25618
rect 12574 25566 12626 25618
rect 12626 25566 12628 25618
rect 12572 25564 12628 25566
rect 12796 24444 12852 24500
rect 13244 24892 13300 24948
rect 13468 24108 13524 24164
rect 14812 30994 14868 30996
rect 14812 30942 14814 30994
rect 14814 30942 14866 30994
rect 14866 30942 14868 30994
rect 14812 30940 14868 30942
rect 14476 24892 14532 24948
rect 13916 24108 13972 24164
rect 13804 23996 13860 24052
rect 12572 23660 12628 23716
rect 12124 23212 12180 23268
rect 12124 22764 12180 22820
rect 12572 22428 12628 22484
rect 12908 23714 12964 23716
rect 12908 23662 12910 23714
rect 12910 23662 12962 23714
rect 12962 23662 12964 23714
rect 12908 23660 12964 23662
rect 13580 23660 13636 23716
rect 12572 20018 12628 20020
rect 12572 19966 12574 20018
rect 12574 19966 12626 20018
rect 12626 19966 12628 20018
rect 12572 19964 12628 19966
rect 13020 20018 13076 20020
rect 13020 19966 13022 20018
rect 13022 19966 13074 20018
rect 13074 19966 13076 20018
rect 13020 19964 13076 19966
rect 11564 16156 11620 16212
rect 11116 16098 11172 16100
rect 11116 16046 11118 16098
rect 11118 16046 11170 16098
rect 11170 16046 11172 16098
rect 11116 16044 11172 16046
rect 11340 15484 11396 15540
rect 11116 15314 11172 15316
rect 11116 15262 11118 15314
rect 11118 15262 11170 15314
rect 11170 15262 11172 15314
rect 11116 15260 11172 15262
rect 11452 15148 11508 15204
rect 11228 14140 11284 14196
rect 11116 13580 11172 13636
rect 9548 12908 9604 12964
rect 10444 12962 10500 12964
rect 10444 12910 10446 12962
rect 10446 12910 10498 12962
rect 10498 12910 10500 12962
rect 10444 12908 10500 12910
rect 9436 12850 9492 12852
rect 9436 12798 9438 12850
rect 9438 12798 9490 12850
rect 9490 12798 9492 12850
rect 9436 12796 9492 12798
rect 9996 12796 10052 12852
rect 8540 11900 8596 11956
rect 8092 11676 8148 11732
rect 7868 11452 7924 11508
rect 8316 11394 8372 11396
rect 8316 11342 8318 11394
rect 8318 11342 8370 11394
rect 8370 11342 8372 11394
rect 8316 11340 8372 11342
rect 8652 11506 8708 11508
rect 8652 11454 8654 11506
rect 8654 11454 8706 11506
rect 8706 11454 8708 11506
rect 8652 11452 8708 11454
rect 8764 11282 8820 11284
rect 8764 11230 8766 11282
rect 8766 11230 8818 11282
rect 8818 11230 8820 11282
rect 8764 11228 8820 11230
rect 7756 10108 7812 10164
rect 7084 9100 7140 9156
rect 7420 8988 7476 9044
rect 6748 8204 6804 8260
rect 7196 8204 7252 8260
rect 6524 7586 6580 7588
rect 6524 7534 6526 7586
rect 6526 7534 6578 7586
rect 6578 7534 6580 7586
rect 6524 7532 6580 7534
rect 6412 7420 6468 7476
rect 6636 7474 6692 7476
rect 6636 7422 6638 7474
rect 6638 7422 6690 7474
rect 6690 7422 6692 7474
rect 6636 7420 6692 7422
rect 8204 9042 8260 9044
rect 8204 8990 8206 9042
rect 8206 8990 8258 9042
rect 8258 8990 8260 9042
rect 8204 8988 8260 8990
rect 7868 7756 7924 7812
rect 7196 7698 7252 7700
rect 7196 7646 7198 7698
rect 7198 7646 7250 7698
rect 7250 7646 7252 7698
rect 7196 7644 7252 7646
rect 7756 7586 7812 7588
rect 7756 7534 7758 7586
rect 7758 7534 7810 7586
rect 7810 7534 7812 7586
rect 7756 7532 7812 7534
rect 6412 5122 6468 5124
rect 6412 5070 6414 5122
rect 6414 5070 6466 5122
rect 6466 5070 6468 5122
rect 6412 5068 6468 5070
rect 7308 6466 7364 6468
rect 7308 6414 7310 6466
rect 7310 6414 7362 6466
rect 7362 6414 7364 6466
rect 7308 6412 7364 6414
rect 6636 5852 6692 5908
rect 8428 7644 8484 7700
rect 8428 7474 8484 7476
rect 8428 7422 8430 7474
rect 8430 7422 8482 7474
rect 8482 7422 8484 7474
rect 8428 7420 8484 7422
rect 8316 7308 8372 7364
rect 7756 6524 7812 6580
rect 7532 6130 7588 6132
rect 7532 6078 7534 6130
rect 7534 6078 7586 6130
rect 7586 6078 7588 6130
rect 7532 6076 7588 6078
rect 8092 6076 8148 6132
rect 4956 3276 5012 3332
rect 5852 2940 5908 2996
rect 7420 5180 7476 5236
rect 7196 4620 7252 4676
rect 7532 4844 7588 4900
rect 7644 5852 7700 5908
rect 7980 5906 8036 5908
rect 7980 5854 7982 5906
rect 7982 5854 8034 5906
rect 8034 5854 8036 5906
rect 7980 5852 8036 5854
rect 7756 4508 7812 4564
rect 6748 3276 6804 3332
rect 4476 2378 4532 2380
rect 4476 2326 4478 2378
rect 4478 2326 4530 2378
rect 4530 2326 4532 2378
rect 4476 2324 4532 2326
rect 4580 2378 4636 2380
rect 4580 2326 4582 2378
rect 4582 2326 4634 2378
rect 4634 2326 4636 2378
rect 4580 2324 4636 2326
rect 4684 2378 4740 2380
rect 4684 2326 4686 2378
rect 4686 2326 4738 2378
rect 4738 2326 4740 2378
rect 4684 2324 4740 2326
rect 7420 3778 7476 3780
rect 7420 3726 7422 3778
rect 7422 3726 7474 3778
rect 7474 3726 7476 3778
rect 7420 3724 7476 3726
rect 8540 6578 8596 6580
rect 8540 6526 8542 6578
rect 8542 6526 8594 6578
rect 8594 6526 8596 6578
rect 8540 6524 8596 6526
rect 8204 4620 8260 4676
rect 8876 6018 8932 6020
rect 8876 5966 8878 6018
rect 8878 5966 8930 6018
rect 8930 5966 8932 6018
rect 8876 5964 8932 5966
rect 8316 5068 8372 5124
rect 8876 5180 8932 5236
rect 9324 11676 9380 11732
rect 10220 11228 10276 11284
rect 10668 12402 10724 12404
rect 10668 12350 10670 12402
rect 10670 12350 10722 12402
rect 10722 12350 10724 12402
rect 10668 12348 10724 12350
rect 9548 9938 9604 9940
rect 9548 9886 9550 9938
rect 9550 9886 9602 9938
rect 9602 9886 9604 9938
rect 9548 9884 9604 9886
rect 9100 7756 9156 7812
rect 9100 6412 9156 6468
rect 9324 7644 9380 7700
rect 11340 12348 11396 12404
rect 11340 11506 11396 11508
rect 11340 11454 11342 11506
rect 11342 11454 11394 11506
rect 11394 11454 11396 11506
rect 11340 11452 11396 11454
rect 11676 13468 11732 13524
rect 11900 15090 11956 15092
rect 11900 15038 11902 15090
rect 11902 15038 11954 15090
rect 11954 15038 11956 15090
rect 11900 15036 11956 15038
rect 12012 14476 12068 14532
rect 12460 18396 12516 18452
rect 12796 16716 12852 16772
rect 12572 15484 12628 15540
rect 12796 15260 12852 15316
rect 13020 15036 13076 15092
rect 12796 14476 12852 14532
rect 12460 14252 12516 14308
rect 11900 13468 11956 13524
rect 12236 13858 12292 13860
rect 12236 13806 12238 13858
rect 12238 13806 12290 13858
rect 12290 13806 12292 13858
rect 12236 13804 12292 13806
rect 12908 13468 12964 13524
rect 11788 12572 11844 12628
rect 11564 12236 11620 12292
rect 11564 11900 11620 11956
rect 12236 12572 12292 12628
rect 12124 12460 12180 12516
rect 12012 11788 12068 11844
rect 11900 11676 11956 11732
rect 10892 11228 10948 11284
rect 10668 10668 10724 10724
rect 10108 9548 10164 9604
rect 10108 9100 10164 9156
rect 9772 7756 9828 7812
rect 9884 7586 9940 7588
rect 9884 7534 9886 7586
rect 9886 7534 9938 7586
rect 9938 7534 9940 7586
rect 9884 7532 9940 7534
rect 9996 6636 10052 6692
rect 10556 8876 10612 8932
rect 10780 9548 10836 9604
rect 11564 9826 11620 9828
rect 11564 9774 11566 9826
rect 11566 9774 11618 9826
rect 11618 9774 11620 9826
rect 11564 9772 11620 9774
rect 11004 9042 11060 9044
rect 11004 8990 11006 9042
rect 11006 8990 11058 9042
rect 11058 8990 11060 9042
rect 11004 8988 11060 8990
rect 10444 7644 10500 7700
rect 11340 7532 11396 7588
rect 12572 12290 12628 12292
rect 12572 12238 12574 12290
rect 12574 12238 12626 12290
rect 12626 12238 12628 12290
rect 12572 12236 12628 12238
rect 12348 11676 12404 11732
rect 11900 9884 11956 9940
rect 11676 8876 11732 8932
rect 10220 7308 10276 7364
rect 10108 6748 10164 6804
rect 9548 6578 9604 6580
rect 9548 6526 9550 6578
rect 9550 6526 9602 6578
rect 9602 6526 9604 6578
rect 9548 6524 9604 6526
rect 9324 5852 9380 5908
rect 9884 5906 9940 5908
rect 9884 5854 9886 5906
rect 9886 5854 9938 5906
rect 9938 5854 9940 5906
rect 9884 5852 9940 5854
rect 10220 5964 10276 6020
rect 10892 6690 10948 6692
rect 10892 6638 10894 6690
rect 10894 6638 10946 6690
rect 10946 6638 10948 6690
rect 10892 6636 10948 6638
rect 10332 5292 10388 5348
rect 8764 4844 8820 4900
rect 8428 3724 8484 3780
rect 9660 4620 9716 4676
rect 8876 4562 8932 4564
rect 8876 4510 8878 4562
rect 8878 4510 8930 4562
rect 8930 4510 8932 4562
rect 8876 4508 8932 4510
rect 8876 4060 8932 4116
rect 10332 5010 10388 5012
rect 10332 4958 10334 5010
rect 10334 4958 10386 5010
rect 10386 4958 10388 5010
rect 10332 4956 10388 4958
rect 10332 4562 10388 4564
rect 10332 4510 10334 4562
rect 10334 4510 10386 4562
rect 10386 4510 10388 4562
rect 10332 4508 10388 4510
rect 10444 4450 10500 4452
rect 10444 4398 10446 4450
rect 10446 4398 10498 4450
rect 10498 4398 10500 4450
rect 10444 4396 10500 4398
rect 10892 5852 10948 5908
rect 10668 4508 10724 4564
rect 12124 9660 12180 9716
rect 12572 11452 12628 11508
rect 12572 10610 12628 10612
rect 12572 10558 12574 10610
rect 12574 10558 12626 10610
rect 12626 10558 12628 10610
rect 12572 10556 12628 10558
rect 12908 11452 12964 11508
rect 12908 9884 12964 9940
rect 12796 9660 12852 9716
rect 12012 8428 12068 8484
rect 12908 8428 12964 8484
rect 12684 7420 12740 7476
rect 12236 6748 12292 6804
rect 11788 6300 11844 6356
rect 11116 5740 11172 5796
rect 12684 6802 12740 6804
rect 12684 6750 12686 6802
rect 12686 6750 12738 6802
rect 12738 6750 12740 6802
rect 12684 6748 12740 6750
rect 11228 6076 11284 6132
rect 10444 4060 10500 4116
rect 7308 2546 7364 2548
rect 7308 2494 7310 2546
rect 7310 2494 7362 2546
rect 7362 2494 7364 2546
rect 7308 2492 7364 2494
rect 10108 2546 10164 2548
rect 10108 2494 10110 2546
rect 10110 2494 10162 2546
rect 10162 2494 10164 2546
rect 10108 2492 10164 2494
rect 11788 4508 11844 4564
rect 11340 3778 11396 3780
rect 11340 3726 11342 3778
rect 11342 3726 11394 3778
rect 11394 3726 11396 3778
rect 11340 3724 11396 3726
rect 12460 5964 12516 6020
rect 12572 6412 12628 6468
rect 12124 4396 12180 4452
rect 12460 5292 12516 5348
rect 12236 5068 12292 5124
rect 12348 5180 12404 5236
rect 13692 21420 13748 21476
rect 13468 21084 13524 21140
rect 14252 21474 14308 21476
rect 14252 21422 14254 21474
rect 14254 21422 14306 21474
rect 14306 21422 14308 21474
rect 14252 21420 14308 21422
rect 14476 21420 14532 21476
rect 14700 23996 14756 24052
rect 14700 23324 14756 23380
rect 14700 21532 14756 21588
rect 13468 20524 13524 20580
rect 14588 18396 14644 18452
rect 14812 18620 14868 18676
rect 13580 17388 13636 17444
rect 14700 17442 14756 17444
rect 14700 17390 14702 17442
rect 14702 17390 14754 17442
rect 14754 17390 14756 17442
rect 14700 17388 14756 17390
rect 14140 16882 14196 16884
rect 14140 16830 14142 16882
rect 14142 16830 14194 16882
rect 14194 16830 14196 16882
rect 14140 16828 14196 16830
rect 13468 14476 13524 14532
rect 13580 13804 13636 13860
rect 13132 12460 13188 12516
rect 13916 13468 13972 13524
rect 14028 14642 14084 14644
rect 14028 14590 14030 14642
rect 14030 14590 14082 14642
rect 14082 14590 14084 14642
rect 14028 14588 14084 14590
rect 15372 39452 15428 39508
rect 15372 38050 15428 38052
rect 15372 37998 15374 38050
rect 15374 37998 15426 38050
rect 15426 37998 15428 38050
rect 15372 37996 15428 37998
rect 15036 37100 15092 37156
rect 16604 43372 16660 43428
rect 16156 42476 16212 42532
rect 16828 46620 16884 46676
rect 17052 45612 17108 45668
rect 17500 44098 17556 44100
rect 17500 44046 17502 44098
rect 17502 44046 17554 44098
rect 17554 44046 17556 44098
rect 17500 44044 17556 44046
rect 17052 43708 17108 43764
rect 17612 43372 17668 43428
rect 16828 42588 16884 42644
rect 17500 42588 17556 42644
rect 16156 41970 16212 41972
rect 16156 41918 16158 41970
rect 16158 41918 16210 41970
rect 16210 41918 16212 41970
rect 16156 41916 16212 41918
rect 18060 48130 18116 48132
rect 18060 48078 18062 48130
rect 18062 48078 18114 48130
rect 18114 48078 18116 48130
rect 18060 48076 18116 48078
rect 18060 47180 18116 47236
rect 18732 50594 18788 50596
rect 18732 50542 18734 50594
rect 18734 50542 18786 50594
rect 18786 50542 18788 50594
rect 18732 50540 18788 50542
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 20412 60956 20468 61012
rect 20300 58322 20356 58324
rect 20300 58270 20302 58322
rect 20302 58270 20354 58322
rect 20354 58270 20356 58322
rect 20300 58268 20356 58270
rect 23324 68796 23380 68852
rect 22428 68684 22484 68740
rect 23100 68626 23156 68628
rect 23100 68574 23102 68626
rect 23102 68574 23154 68626
rect 23154 68574 23156 68626
rect 23100 68572 23156 68574
rect 22988 68348 23044 68404
rect 22428 67564 22484 67620
rect 22876 67618 22932 67620
rect 22876 67566 22878 67618
rect 22878 67566 22930 67618
rect 22930 67566 22932 67618
rect 22876 67564 22932 67566
rect 21420 66050 21476 66052
rect 21420 65998 21422 66050
rect 21422 65998 21474 66050
rect 21474 65998 21476 66050
rect 21420 65996 21476 65998
rect 21420 65324 21476 65380
rect 22316 65996 22372 66052
rect 21980 64146 22036 64148
rect 21980 64094 21982 64146
rect 21982 64094 22034 64146
rect 22034 64094 22036 64146
rect 21980 64092 22036 64094
rect 21532 63868 21588 63924
rect 22092 63868 22148 63924
rect 20748 62860 20804 62916
rect 20972 61292 21028 61348
rect 20636 61010 20692 61012
rect 20636 60958 20638 61010
rect 20638 60958 20690 61010
rect 20690 60958 20692 61010
rect 20636 60956 20692 60958
rect 21420 59948 21476 60004
rect 20188 55298 20244 55300
rect 20188 55246 20190 55298
rect 20190 55246 20242 55298
rect 20242 55246 20244 55298
rect 20188 55244 20244 55246
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19628 54738 19684 54740
rect 19628 54686 19630 54738
rect 19630 54686 19682 54738
rect 19682 54686 19684 54738
rect 19628 54684 19684 54686
rect 19516 54236 19572 54292
rect 18956 49308 19012 49364
rect 19180 52668 19236 52724
rect 18732 48860 18788 48916
rect 18844 48802 18900 48804
rect 18844 48750 18846 48802
rect 18846 48750 18898 48802
rect 18898 48750 18900 48802
rect 18844 48748 18900 48750
rect 18620 48242 18676 48244
rect 18620 48190 18622 48242
rect 18622 48190 18674 48242
rect 18674 48190 18676 48242
rect 18620 48188 18676 48190
rect 18844 47180 18900 47236
rect 18844 46562 18900 46564
rect 18844 46510 18846 46562
rect 18846 46510 18898 46562
rect 18898 46510 18900 46562
rect 18844 46508 18900 46510
rect 17836 43762 17892 43764
rect 17836 43710 17838 43762
rect 17838 43710 17890 43762
rect 17890 43710 17892 43762
rect 17836 43708 17892 43710
rect 17724 41970 17780 41972
rect 17724 41918 17726 41970
rect 17726 41918 17778 41970
rect 17778 41918 17780 41970
rect 17724 41916 17780 41918
rect 17164 41804 17220 41860
rect 20524 54236 20580 54292
rect 20748 55186 20804 55188
rect 20748 55134 20750 55186
rect 20750 55134 20802 55186
rect 20802 55134 20804 55186
rect 20748 55132 20804 55134
rect 20636 53788 20692 53844
rect 20076 53676 20132 53732
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 20524 53004 20580 53060
rect 19628 52722 19684 52724
rect 19628 52670 19630 52722
rect 19630 52670 19682 52722
rect 19682 52670 19684 52722
rect 19628 52668 19684 52670
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19852 50540 19908 50596
rect 21308 56588 21364 56644
rect 21756 59778 21812 59780
rect 21756 59726 21758 59778
rect 21758 59726 21810 59778
rect 21810 59726 21812 59778
rect 21756 59724 21812 59726
rect 21644 59388 21700 59444
rect 22428 64428 22484 64484
rect 22428 64092 22484 64148
rect 22316 62412 22372 62468
rect 22316 59388 22372 59444
rect 21980 59052 22036 59108
rect 22204 58828 22260 58884
rect 22876 64482 22932 64484
rect 22876 64430 22878 64482
rect 22878 64430 22930 64482
rect 22930 64430 22932 64482
rect 22876 64428 22932 64430
rect 22876 64034 22932 64036
rect 22876 63982 22878 64034
rect 22878 63982 22930 64034
rect 22930 63982 22932 64034
rect 22876 63980 22932 63982
rect 22764 63922 22820 63924
rect 22764 63870 22766 63922
rect 22766 63870 22818 63922
rect 22818 63870 22820 63922
rect 22764 63868 22820 63870
rect 24556 71650 24612 71652
rect 24556 71598 24558 71650
rect 24558 71598 24610 71650
rect 24610 71598 24612 71650
rect 24556 71596 24612 71598
rect 24108 70588 24164 70644
rect 23660 69244 23716 69300
rect 23996 70028 24052 70084
rect 23548 68684 23604 68740
rect 23324 64428 23380 64484
rect 23548 64540 23604 64596
rect 23324 62466 23380 62468
rect 23324 62414 23326 62466
rect 23326 62414 23378 62466
rect 23378 62414 23380 62466
rect 23324 62412 23380 62414
rect 23772 68850 23828 68852
rect 23772 68798 23774 68850
rect 23774 68798 23826 68850
rect 23826 68798 23828 68850
rect 23772 68796 23828 68798
rect 23996 68572 24052 68628
rect 24108 68460 24164 68516
rect 24220 68572 24276 68628
rect 24668 68738 24724 68740
rect 24668 68686 24670 68738
rect 24670 68686 24722 68738
rect 24722 68686 24724 68738
rect 24668 68684 24724 68686
rect 25004 68460 25060 68516
rect 23660 62466 23716 62468
rect 23660 62414 23662 62466
rect 23662 62414 23714 62466
rect 23714 62414 23716 62466
rect 23660 62412 23716 62414
rect 22652 61346 22708 61348
rect 22652 61294 22654 61346
rect 22654 61294 22706 61346
rect 22706 61294 22708 61346
rect 22652 61292 22708 61294
rect 22988 61292 23044 61348
rect 22876 59724 22932 59780
rect 21980 58380 22036 58436
rect 22652 59052 22708 59108
rect 21420 55244 21476 55300
rect 21644 53564 21700 53620
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19628 49810 19684 49812
rect 19628 49758 19630 49810
rect 19630 49758 19682 49810
rect 19682 49758 19684 49810
rect 19628 49756 19684 49758
rect 19516 49308 19572 49364
rect 19516 46844 19572 46900
rect 19292 46508 19348 46564
rect 18620 44434 18676 44436
rect 18620 44382 18622 44434
rect 18622 44382 18674 44434
rect 18674 44382 18676 44434
rect 18620 44380 18676 44382
rect 18284 43708 18340 43764
rect 18060 42530 18116 42532
rect 18060 42478 18062 42530
rect 18062 42478 18114 42530
rect 18114 42478 18116 42530
rect 18060 42476 18116 42478
rect 19292 45612 19348 45668
rect 19516 45778 19572 45780
rect 19516 45726 19518 45778
rect 19518 45726 19570 45778
rect 19570 45726 19572 45778
rect 19516 45724 19572 45726
rect 20076 48748 20132 48804
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 20300 48972 20356 49028
rect 19964 47234 20020 47236
rect 19964 47182 19966 47234
rect 19966 47182 20018 47234
rect 20018 47182 20020 47234
rect 19964 47180 20020 47182
rect 20300 48242 20356 48244
rect 20300 48190 20302 48242
rect 20302 48190 20354 48242
rect 20354 48190 20356 48242
rect 20300 48188 20356 48190
rect 20636 48076 20692 48132
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 20300 46620 20356 46676
rect 20076 46562 20132 46564
rect 20076 46510 20078 46562
rect 20078 46510 20130 46562
rect 20130 46510 20132 46562
rect 20076 46508 20132 46510
rect 19852 45724 19908 45780
rect 20188 46060 20244 46116
rect 20300 45836 20356 45892
rect 20636 46956 20692 47012
rect 20636 46060 20692 46116
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19180 44380 19236 44436
rect 18956 43372 19012 43428
rect 19180 43148 19236 43204
rect 18060 41746 18116 41748
rect 18060 41694 18062 41746
rect 18062 41694 18114 41746
rect 18114 41694 18116 41746
rect 18060 41692 18116 41694
rect 18396 40572 18452 40628
rect 16156 40348 16212 40404
rect 17500 40514 17556 40516
rect 17500 40462 17502 40514
rect 17502 40462 17554 40514
rect 17554 40462 17556 40514
rect 17500 40460 17556 40462
rect 18172 40402 18228 40404
rect 18172 40350 18174 40402
rect 18174 40350 18226 40402
rect 18226 40350 18228 40402
rect 18172 40348 18228 40350
rect 17948 39730 18004 39732
rect 17948 39678 17950 39730
rect 17950 39678 18002 39730
rect 18002 39678 18004 39730
rect 17948 39676 18004 39678
rect 16268 39564 16324 39620
rect 16604 38834 16660 38836
rect 16604 38782 16606 38834
rect 16606 38782 16658 38834
rect 16658 38782 16660 38834
rect 16604 38780 16660 38782
rect 15260 35532 15316 35588
rect 15932 36428 15988 36484
rect 15932 34972 15988 35028
rect 15932 34412 15988 34468
rect 15708 34188 15764 34244
rect 16828 37324 16884 37380
rect 16716 37154 16772 37156
rect 16716 37102 16718 37154
rect 16718 37102 16770 37154
rect 16770 37102 16772 37154
rect 16716 37100 16772 37102
rect 16492 37042 16548 37044
rect 16492 36990 16494 37042
rect 16494 36990 16546 37042
rect 16546 36990 16548 37042
rect 16492 36988 16548 36990
rect 17948 38834 18004 38836
rect 17948 38782 17950 38834
rect 17950 38782 18002 38834
rect 18002 38782 18004 38834
rect 17948 38780 18004 38782
rect 16828 36988 16884 37044
rect 16380 35586 16436 35588
rect 16380 35534 16382 35586
rect 16382 35534 16434 35586
rect 16434 35534 16436 35586
rect 16380 35532 16436 35534
rect 15820 33852 15876 33908
rect 15260 30940 15316 30996
rect 15484 32508 15540 32564
rect 16380 34018 16436 34020
rect 16380 33966 16382 34018
rect 16382 33966 16434 34018
rect 16434 33966 16436 34018
rect 16380 33964 16436 33966
rect 16380 33628 16436 33684
rect 15820 32508 15876 32564
rect 15260 30156 15316 30212
rect 18172 35810 18228 35812
rect 18172 35758 18174 35810
rect 18174 35758 18226 35810
rect 18226 35758 18228 35810
rect 18172 35756 18228 35758
rect 18060 35644 18116 35700
rect 17836 35532 17892 35588
rect 18396 35532 18452 35588
rect 19292 42754 19348 42756
rect 19292 42702 19294 42754
rect 19294 42702 19346 42754
rect 19346 42702 19348 42754
rect 19292 42700 19348 42702
rect 19404 42642 19460 42644
rect 19404 42590 19406 42642
rect 19406 42590 19458 42642
rect 19458 42590 19460 42642
rect 19404 42588 19460 42590
rect 19068 42476 19124 42532
rect 21084 49698 21140 49700
rect 21084 49646 21086 49698
rect 21086 49646 21138 49698
rect 21138 49646 21140 49698
rect 21084 49644 21140 49646
rect 21308 49026 21364 49028
rect 21308 48974 21310 49026
rect 21310 48974 21362 49026
rect 21362 48974 21364 49026
rect 21308 48972 21364 48974
rect 21308 48748 21364 48804
rect 21756 49644 21812 49700
rect 21420 48130 21476 48132
rect 21420 48078 21422 48130
rect 21422 48078 21474 48130
rect 21474 48078 21476 48130
rect 21420 48076 21476 48078
rect 21420 46732 21476 46788
rect 21308 46620 21364 46676
rect 20748 45164 20804 45220
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20636 43484 20692 43540
rect 19628 43372 19684 43428
rect 20076 43372 20132 43428
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 18732 41804 18788 41860
rect 19180 41692 19236 41748
rect 18732 40514 18788 40516
rect 18732 40462 18734 40514
rect 18734 40462 18786 40514
rect 18786 40462 18788 40514
rect 18732 40460 18788 40462
rect 18844 40348 18900 40404
rect 18956 39676 19012 39732
rect 19292 40460 19348 40516
rect 19068 38780 19124 38836
rect 19180 40124 19236 40180
rect 19180 37324 19236 37380
rect 19292 38892 19348 38948
rect 18956 36876 19012 36932
rect 19068 36764 19124 36820
rect 17388 35084 17444 35140
rect 17948 35026 18004 35028
rect 17948 34974 17950 35026
rect 17950 34974 18002 35026
rect 18002 34974 18004 35026
rect 17948 34972 18004 34974
rect 17052 33852 17108 33908
rect 17612 33628 17668 33684
rect 18508 35138 18564 35140
rect 18508 35086 18510 35138
rect 18510 35086 18562 35138
rect 18562 35086 18564 35138
rect 18508 35084 18564 35086
rect 19964 41298 20020 41300
rect 19964 41246 19966 41298
rect 19966 41246 20018 41298
rect 20018 41246 20020 41298
rect 19964 41244 20020 41246
rect 20860 42476 20916 42532
rect 20636 41804 20692 41860
rect 20748 41580 20804 41636
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19964 40402 20020 40404
rect 19964 40350 19966 40402
rect 19966 40350 20018 40402
rect 20018 40350 20020 40402
rect 19964 40348 20020 40350
rect 20524 40514 20580 40516
rect 20524 40462 20526 40514
rect 20526 40462 20578 40514
rect 20578 40462 20580 40514
rect 20524 40460 20580 40462
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 20188 39004 20244 39060
rect 20860 39564 20916 39620
rect 20412 39116 20468 39172
rect 19964 38892 20020 38948
rect 20636 38556 20692 38612
rect 21532 47068 21588 47124
rect 21756 46956 21812 47012
rect 21532 46620 21588 46676
rect 21644 46844 21700 46900
rect 21420 45666 21476 45668
rect 21420 45614 21422 45666
rect 21422 45614 21474 45666
rect 21474 45614 21476 45666
rect 21420 45612 21476 45614
rect 21308 43596 21364 43652
rect 21420 43538 21476 43540
rect 21420 43486 21422 43538
rect 21422 43486 21474 43538
rect 21474 43486 21476 43538
rect 21420 43484 21476 43486
rect 21868 46620 21924 46676
rect 21644 43484 21700 43540
rect 21756 45724 21812 45780
rect 21868 45164 21924 45220
rect 22204 52108 22260 52164
rect 22092 48076 22148 48132
rect 23212 59388 23268 59444
rect 23100 57036 23156 57092
rect 22764 55916 22820 55972
rect 22764 53676 22820 53732
rect 22764 53170 22820 53172
rect 22764 53118 22766 53170
rect 22766 53118 22818 53170
rect 22818 53118 22820 53170
rect 22764 53116 22820 53118
rect 22764 52050 22820 52052
rect 22764 51998 22766 52050
rect 22766 51998 22818 52050
rect 22818 51998 22820 52050
rect 22764 51996 22820 51998
rect 22764 51324 22820 51380
rect 22652 50988 22708 51044
rect 23324 57762 23380 57764
rect 23324 57710 23326 57762
rect 23326 57710 23378 57762
rect 23378 57710 23380 57762
rect 23324 57708 23380 57710
rect 24220 64540 24276 64596
rect 24108 64482 24164 64484
rect 24108 64430 24110 64482
rect 24110 64430 24162 64482
rect 24162 64430 24164 64482
rect 24108 64428 24164 64430
rect 24108 63868 24164 63924
rect 24332 60002 24388 60004
rect 24332 59950 24334 60002
rect 24334 59950 24386 60002
rect 24386 59950 24388 60002
rect 24332 59948 24388 59950
rect 24332 58828 24388 58884
rect 24332 58492 24388 58548
rect 23548 57148 23604 57204
rect 23884 56754 23940 56756
rect 23884 56702 23886 56754
rect 23886 56702 23938 56754
rect 23938 56702 23940 56754
rect 23884 56700 23940 56702
rect 25340 70252 25396 70308
rect 25900 74898 25956 74900
rect 25900 74846 25902 74898
rect 25902 74846 25954 74898
rect 25954 74846 25956 74898
rect 25900 74844 25956 74846
rect 31276 76188 31332 76244
rect 30156 75794 30212 75796
rect 30156 75742 30158 75794
rect 30158 75742 30210 75794
rect 30210 75742 30212 75794
rect 30156 75740 30212 75742
rect 30940 75794 30996 75796
rect 30940 75742 30942 75794
rect 30942 75742 30994 75794
rect 30994 75742 30996 75794
rect 30940 75740 30996 75742
rect 29932 75682 29988 75684
rect 29932 75630 29934 75682
rect 29934 75630 29986 75682
rect 29986 75630 29988 75682
rect 29932 75628 29988 75630
rect 30828 75628 30884 75684
rect 29820 74844 29876 74900
rect 25564 73218 25620 73220
rect 25564 73166 25566 73218
rect 25566 73166 25618 73218
rect 25618 73166 25620 73218
rect 25564 73164 25620 73166
rect 26684 73218 26740 73220
rect 26684 73166 26686 73218
rect 26686 73166 26738 73218
rect 26738 73166 26740 73218
rect 26684 73164 26740 73166
rect 26124 71650 26180 71652
rect 26124 71598 26126 71650
rect 26126 71598 26178 71650
rect 26178 71598 26180 71650
rect 26124 71596 26180 71598
rect 26348 71202 26404 71204
rect 26348 71150 26350 71202
rect 26350 71150 26402 71202
rect 26402 71150 26404 71202
rect 26348 71148 26404 71150
rect 26012 70252 26068 70308
rect 25788 70194 25844 70196
rect 25788 70142 25790 70194
rect 25790 70142 25842 70194
rect 25842 70142 25844 70194
rect 25788 70140 25844 70142
rect 25340 68684 25396 68740
rect 26908 70476 26964 70532
rect 26908 70028 26964 70084
rect 25788 68796 25844 68852
rect 25340 64988 25396 65044
rect 24780 61180 24836 61236
rect 25004 61292 25060 61348
rect 24556 61010 24612 61012
rect 24556 60958 24558 61010
rect 24558 60958 24610 61010
rect 24610 60958 24612 61010
rect 24556 60956 24612 60958
rect 24668 60674 24724 60676
rect 24668 60622 24670 60674
rect 24670 60622 24722 60674
rect 24722 60622 24724 60674
rect 24668 60620 24724 60622
rect 25340 63868 25396 63924
rect 24892 60114 24948 60116
rect 24892 60062 24894 60114
rect 24894 60062 24946 60114
rect 24946 60062 24948 60114
rect 24892 60060 24948 60062
rect 25004 59948 25060 60004
rect 24556 58434 24612 58436
rect 24556 58382 24558 58434
rect 24558 58382 24610 58434
rect 24610 58382 24612 58434
rect 24556 58380 24612 58382
rect 24556 57484 24612 57540
rect 24556 55916 24612 55972
rect 23212 54460 23268 54516
rect 23324 54572 23380 54628
rect 24108 54626 24164 54628
rect 24108 54574 24110 54626
rect 24110 54574 24162 54626
rect 24162 54574 24164 54626
rect 24108 54572 24164 54574
rect 24780 58546 24836 58548
rect 24780 58494 24782 58546
rect 24782 58494 24834 58546
rect 24834 58494 24836 58546
rect 24780 58492 24836 58494
rect 25004 58044 25060 58100
rect 25788 65212 25844 65268
rect 25676 64988 25732 65044
rect 25676 63980 25732 64036
rect 26348 61346 26404 61348
rect 26348 61294 26350 61346
rect 26350 61294 26402 61346
rect 26402 61294 26404 61346
rect 26348 61292 26404 61294
rect 25900 61180 25956 61236
rect 25676 58546 25732 58548
rect 25676 58494 25678 58546
rect 25678 58494 25730 58546
rect 25730 58494 25732 58546
rect 25676 58492 25732 58494
rect 25564 58268 25620 58324
rect 26348 60956 26404 61012
rect 26012 60674 26068 60676
rect 26012 60622 26014 60674
rect 26014 60622 26066 60674
rect 26066 60622 26068 60674
rect 26012 60620 26068 60622
rect 26572 65212 26628 65268
rect 26012 60060 26068 60116
rect 26348 59724 26404 59780
rect 26908 68514 26964 68516
rect 26908 68462 26910 68514
rect 26910 68462 26962 68514
rect 26962 68462 26964 68514
rect 26908 68460 26964 68462
rect 27356 72268 27412 72324
rect 28028 70194 28084 70196
rect 28028 70142 28030 70194
rect 28030 70142 28082 70194
rect 28082 70142 28084 70194
rect 28028 70140 28084 70142
rect 28364 70082 28420 70084
rect 28364 70030 28366 70082
rect 28366 70030 28418 70082
rect 28418 70030 28420 70082
rect 28364 70028 28420 70030
rect 27356 68460 27412 68516
rect 27356 67564 27412 67620
rect 27468 67058 27524 67060
rect 27468 67006 27470 67058
rect 27470 67006 27522 67058
rect 27522 67006 27524 67058
rect 27468 67004 27524 67006
rect 27804 65436 27860 65492
rect 26124 58434 26180 58436
rect 26124 58382 26126 58434
rect 26126 58382 26178 58434
rect 26178 58382 26180 58434
rect 26124 58380 26180 58382
rect 24780 57484 24836 57540
rect 25564 57596 25620 57652
rect 25340 57538 25396 57540
rect 25340 57486 25342 57538
rect 25342 57486 25394 57538
rect 25394 57486 25396 57538
rect 25340 57484 25396 57486
rect 25452 57090 25508 57092
rect 25452 57038 25454 57090
rect 25454 57038 25506 57090
rect 25506 57038 25508 57090
rect 25452 57036 25508 57038
rect 25676 56924 25732 56980
rect 23436 53842 23492 53844
rect 23436 53790 23438 53842
rect 23438 53790 23490 53842
rect 23490 53790 23492 53842
rect 23436 53788 23492 53790
rect 23212 53618 23268 53620
rect 23212 53566 23214 53618
rect 23214 53566 23266 53618
rect 23266 53566 23268 53618
rect 23212 53564 23268 53566
rect 23324 53452 23380 53508
rect 23212 53058 23268 53060
rect 23212 53006 23214 53058
rect 23214 53006 23266 53058
rect 23266 53006 23268 53058
rect 23212 53004 23268 53006
rect 23436 53116 23492 53172
rect 23212 52668 23268 52724
rect 23548 51996 23604 52052
rect 22652 50652 22708 50708
rect 22540 50594 22596 50596
rect 22540 50542 22542 50594
rect 22542 50542 22594 50594
rect 22594 50542 22596 50594
rect 22540 50540 22596 50542
rect 22540 48748 22596 48804
rect 22316 47180 22372 47236
rect 22316 46786 22372 46788
rect 22316 46734 22318 46786
rect 22318 46734 22370 46786
rect 22370 46734 22372 46786
rect 22316 46732 22372 46734
rect 22988 50594 23044 50596
rect 22988 50542 22990 50594
rect 22990 50542 23042 50594
rect 23042 50542 23044 50594
rect 22988 50540 23044 50542
rect 23436 50988 23492 51044
rect 22876 48972 22932 49028
rect 22764 46508 22820 46564
rect 23100 48748 23156 48804
rect 22316 45890 22372 45892
rect 22316 45838 22318 45890
rect 22318 45838 22370 45890
rect 22370 45838 22372 45890
rect 22316 45836 22372 45838
rect 23324 48802 23380 48804
rect 23324 48750 23326 48802
rect 23326 48750 23378 48802
rect 23378 48750 23380 48802
rect 23324 48748 23380 48750
rect 23660 51378 23716 51380
rect 23660 51326 23662 51378
rect 23662 51326 23714 51378
rect 23714 51326 23716 51378
rect 23660 51324 23716 51326
rect 23996 53170 24052 53172
rect 23996 53118 23998 53170
rect 23998 53118 24050 53170
rect 24050 53118 24052 53170
rect 23996 53116 24052 53118
rect 23548 47404 23604 47460
rect 23548 46844 23604 46900
rect 23436 46562 23492 46564
rect 23436 46510 23438 46562
rect 23438 46510 23490 46562
rect 23490 46510 23492 46562
rect 23436 46508 23492 46510
rect 22988 45890 23044 45892
rect 22988 45838 22990 45890
rect 22990 45838 23042 45890
rect 23042 45838 23044 45890
rect 22988 45836 23044 45838
rect 22316 45164 22372 45220
rect 21980 44716 22036 44772
rect 21532 42700 21588 42756
rect 21420 42140 21476 42196
rect 21420 41580 21476 41636
rect 21308 39116 21364 39172
rect 21084 39058 21140 39060
rect 21084 39006 21086 39058
rect 21086 39006 21138 39058
rect 21138 39006 21140 39058
rect 21084 39004 21140 39006
rect 21420 38892 21476 38948
rect 22988 44940 23044 44996
rect 22316 43820 22372 43876
rect 22428 44098 22484 44100
rect 22428 44046 22430 44098
rect 22430 44046 22482 44098
rect 22482 44046 22484 44098
rect 22428 44044 22484 44046
rect 22428 43708 22484 43764
rect 22764 44044 22820 44100
rect 23660 45890 23716 45892
rect 23660 45838 23662 45890
rect 23662 45838 23714 45890
rect 23714 45838 23716 45890
rect 23660 45836 23716 45838
rect 23212 44604 23268 44660
rect 23660 44994 23716 44996
rect 23660 44942 23662 44994
rect 23662 44942 23714 44994
rect 23714 44942 23716 44994
rect 23660 44940 23716 44942
rect 23212 43932 23268 43988
rect 22316 42530 22372 42532
rect 22316 42478 22318 42530
rect 22318 42478 22370 42530
rect 22370 42478 22372 42530
rect 22316 42476 22372 42478
rect 22092 42140 22148 42196
rect 21756 41244 21812 41300
rect 22652 41746 22708 41748
rect 22652 41694 22654 41746
rect 22654 41694 22706 41746
rect 22706 41694 22708 41746
rect 22652 41692 22708 41694
rect 21644 38834 21700 38836
rect 21644 38782 21646 38834
rect 21646 38782 21698 38834
rect 21698 38782 21700 38834
rect 21644 38780 21700 38782
rect 23548 43596 23604 43652
rect 23436 43148 23492 43204
rect 23436 42252 23492 42308
rect 23324 42194 23380 42196
rect 23324 42142 23326 42194
rect 23326 42142 23378 42194
rect 23378 42142 23380 42194
rect 23324 42140 23380 42142
rect 24444 52108 24500 52164
rect 24108 48860 24164 48916
rect 23884 48300 23940 48356
rect 23884 47404 23940 47460
rect 24444 48748 24500 48804
rect 24444 47458 24500 47460
rect 24444 47406 24446 47458
rect 24446 47406 24498 47458
rect 24498 47406 24500 47458
rect 24444 47404 24500 47406
rect 23996 46732 24052 46788
rect 24220 44994 24276 44996
rect 24220 44942 24222 44994
rect 24222 44942 24274 44994
rect 24274 44942 24276 44994
rect 24220 44940 24276 44942
rect 23996 43932 24052 43988
rect 23884 42028 23940 42084
rect 23996 43372 24052 43428
rect 23884 41356 23940 41412
rect 23212 40124 23268 40180
rect 21980 39618 22036 39620
rect 21980 39566 21982 39618
rect 21982 39566 22034 39618
rect 22034 39566 22036 39618
rect 21980 39564 22036 39566
rect 23436 39618 23492 39620
rect 23436 39566 23438 39618
rect 23438 39566 23490 39618
rect 23490 39566 23492 39618
rect 23436 39564 23492 39566
rect 23548 39506 23604 39508
rect 23548 39454 23550 39506
rect 23550 39454 23602 39506
rect 23602 39454 23604 39506
rect 23548 39452 23604 39454
rect 23660 39394 23716 39396
rect 23660 39342 23662 39394
rect 23662 39342 23714 39394
rect 23714 39342 23716 39394
rect 23660 39340 23716 39342
rect 21532 38556 21588 38612
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19740 36876 19796 36932
rect 20076 36204 20132 36260
rect 18396 33740 18452 33796
rect 16828 31948 16884 32004
rect 16268 30268 16324 30324
rect 15596 30210 15652 30212
rect 15596 30158 15598 30210
rect 15598 30158 15650 30210
rect 15650 30158 15652 30210
rect 15596 30156 15652 30158
rect 16940 30268 16996 30324
rect 17052 30156 17108 30212
rect 16044 29538 16100 29540
rect 16044 29486 16046 29538
rect 16046 29486 16098 29538
rect 16098 29486 16100 29538
rect 16044 29484 16100 29486
rect 16604 29372 16660 29428
rect 16268 28866 16324 28868
rect 16268 28814 16270 28866
rect 16270 28814 16322 28866
rect 16322 28814 16324 28866
rect 16268 28812 16324 28814
rect 15596 28028 15652 28084
rect 15596 27356 15652 27412
rect 15484 23938 15540 23940
rect 15484 23886 15486 23938
rect 15486 23886 15538 23938
rect 15538 23886 15540 23938
rect 15484 23884 15540 23886
rect 15036 23772 15092 23828
rect 16268 28082 16324 28084
rect 16268 28030 16270 28082
rect 16270 28030 16322 28082
rect 16322 28030 16324 28082
rect 16268 28028 16324 28030
rect 16940 28588 16996 28644
rect 16044 26572 16100 26628
rect 16492 24946 16548 24948
rect 16492 24894 16494 24946
rect 16494 24894 16546 24946
rect 16546 24894 16548 24946
rect 16492 24892 16548 24894
rect 15708 24556 15764 24612
rect 16044 24610 16100 24612
rect 16044 24558 16046 24610
rect 16046 24558 16098 24610
rect 16098 24558 16100 24610
rect 16044 24556 16100 24558
rect 16044 24108 16100 24164
rect 16716 23884 16772 23940
rect 16380 23826 16436 23828
rect 16380 23774 16382 23826
rect 16382 23774 16434 23826
rect 16434 23774 16436 23826
rect 16380 23772 16436 23774
rect 17052 26012 17108 26068
rect 15484 23378 15540 23380
rect 15484 23326 15486 23378
rect 15486 23326 15538 23378
rect 15538 23326 15540 23378
rect 15484 23324 15540 23326
rect 15596 19964 15652 20020
rect 15148 17388 15204 17444
rect 15036 16828 15092 16884
rect 14924 14588 14980 14644
rect 14140 13804 14196 13860
rect 14588 14252 14644 14308
rect 14028 13020 14084 13076
rect 14252 12348 14308 12404
rect 13468 10556 13524 10612
rect 14476 11676 14532 11732
rect 14364 11564 14420 11620
rect 14140 11506 14196 11508
rect 14140 11454 14142 11506
rect 14142 11454 14194 11506
rect 14194 11454 14196 11506
rect 14140 11452 14196 11454
rect 13356 8876 13412 8932
rect 13356 6690 13412 6692
rect 13356 6638 13358 6690
rect 13358 6638 13410 6690
rect 13410 6638 13412 6690
rect 13356 6636 13412 6638
rect 13020 6524 13076 6580
rect 14252 10610 14308 10612
rect 14252 10558 14254 10610
rect 14254 10558 14306 10610
rect 14306 10558 14308 10610
rect 14252 10556 14308 10558
rect 13916 8370 13972 8372
rect 13916 8318 13918 8370
rect 13918 8318 13970 8370
rect 13970 8318 13972 8370
rect 13916 8316 13972 8318
rect 14028 9714 14084 9716
rect 14028 9662 14030 9714
rect 14030 9662 14082 9714
rect 14082 9662 14084 9714
rect 14028 9660 14084 9662
rect 13804 6636 13860 6692
rect 13692 6578 13748 6580
rect 13692 6526 13694 6578
rect 13694 6526 13746 6578
rect 13746 6526 13748 6578
rect 13692 6524 13748 6526
rect 13804 6300 13860 6356
rect 13132 6018 13188 6020
rect 13132 5966 13134 6018
rect 13134 5966 13186 6018
rect 13186 5966 13188 6018
rect 13132 5964 13188 5966
rect 13692 5852 13748 5908
rect 14700 13356 14756 13412
rect 15372 13468 15428 13524
rect 15260 12348 15316 12404
rect 16940 23548 16996 23604
rect 16828 22316 16884 22372
rect 16380 21644 16436 21700
rect 15820 21420 15876 21476
rect 16380 20018 16436 20020
rect 16380 19966 16382 20018
rect 16382 19966 16434 20018
rect 16434 19966 16436 20018
rect 16380 19964 16436 19966
rect 16604 17388 16660 17444
rect 16268 16770 16324 16772
rect 16268 16718 16270 16770
rect 16270 16718 16322 16770
rect 16322 16718 16324 16770
rect 16268 16716 16324 16718
rect 16380 16044 16436 16100
rect 17052 16716 17108 16772
rect 17500 32172 17556 32228
rect 17948 32172 18004 32228
rect 18172 31948 18228 32004
rect 17388 29538 17444 29540
rect 17388 29486 17390 29538
rect 17390 29486 17442 29538
rect 17442 29486 17444 29538
rect 17388 29484 17444 29486
rect 17612 29426 17668 29428
rect 17612 29374 17614 29426
rect 17614 29374 17666 29426
rect 17666 29374 17668 29426
rect 17612 29372 17668 29374
rect 17500 28812 17556 28868
rect 17612 26796 17668 26852
rect 17276 26572 17332 26628
rect 17276 25618 17332 25620
rect 17276 25566 17278 25618
rect 17278 25566 17330 25618
rect 17330 25566 17332 25618
rect 17276 25564 17332 25566
rect 18284 31890 18340 31892
rect 18284 31838 18286 31890
rect 18286 31838 18338 31890
rect 18338 31838 18340 31890
rect 18284 31836 18340 31838
rect 18508 33964 18564 34020
rect 19068 33628 19124 33684
rect 19292 33852 19348 33908
rect 18732 32172 18788 32228
rect 18060 26066 18116 26068
rect 18060 26014 18062 26066
rect 18062 26014 18114 26066
rect 18114 26014 18116 26066
rect 18060 26012 18116 26014
rect 17500 24946 17556 24948
rect 17500 24894 17502 24946
rect 17502 24894 17554 24946
rect 17554 24894 17556 24946
rect 17500 24892 17556 24894
rect 17948 23154 18004 23156
rect 17948 23102 17950 23154
rect 17950 23102 18002 23154
rect 18002 23102 18004 23154
rect 17948 23100 18004 23102
rect 17836 22876 17892 22932
rect 17388 21698 17444 21700
rect 17388 21646 17390 21698
rect 17390 21646 17442 21698
rect 17442 21646 17444 21698
rect 17388 21644 17444 21646
rect 17612 22370 17668 22372
rect 17612 22318 17614 22370
rect 17614 22318 17666 22370
rect 17666 22318 17668 22370
rect 17612 22316 17668 22318
rect 17500 21084 17556 21140
rect 17724 18674 17780 18676
rect 17724 18622 17726 18674
rect 17726 18622 17778 18674
rect 17778 18622 17780 18674
rect 17724 18620 17780 18622
rect 18060 18450 18116 18452
rect 18060 18398 18062 18450
rect 18062 18398 18114 18450
rect 18114 18398 18116 18450
rect 18060 18396 18116 18398
rect 17500 17500 17556 17556
rect 15596 11676 15652 11732
rect 14588 10668 14644 10724
rect 16604 14252 16660 14308
rect 17388 14476 17444 14532
rect 16940 13132 16996 13188
rect 15932 12348 15988 12404
rect 15820 10556 15876 10612
rect 16604 10668 16660 10724
rect 17388 14306 17444 14308
rect 17388 14254 17390 14306
rect 17390 14254 17442 14306
rect 17442 14254 17444 14306
rect 17388 14252 17444 14254
rect 17388 13522 17444 13524
rect 17388 13470 17390 13522
rect 17390 13470 17442 13522
rect 17442 13470 17444 13522
rect 17388 13468 17444 13470
rect 17948 18172 18004 18228
rect 19292 32172 19348 32228
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19964 35532 20020 35588
rect 20412 35586 20468 35588
rect 20412 35534 20414 35586
rect 20414 35534 20466 35586
rect 20466 35534 20468 35586
rect 20412 35532 20468 35534
rect 19628 34972 19684 35028
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19628 34188 19684 34244
rect 19516 33292 19572 33348
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 21196 37490 21252 37492
rect 21196 37438 21198 37490
rect 21198 37438 21250 37490
rect 21250 37438 21252 37490
rect 21196 37436 21252 37438
rect 21532 37436 21588 37492
rect 23996 39452 24052 39508
rect 25340 55186 25396 55188
rect 25340 55134 25342 55186
rect 25342 55134 25394 55186
rect 25394 55134 25396 55186
rect 25340 55132 25396 55134
rect 25340 54626 25396 54628
rect 25340 54574 25342 54626
rect 25342 54574 25394 54626
rect 25394 54574 25396 54626
rect 25340 54572 25396 54574
rect 25228 54514 25284 54516
rect 25228 54462 25230 54514
rect 25230 54462 25282 54514
rect 25282 54462 25284 54514
rect 25228 54460 25284 54462
rect 25676 53788 25732 53844
rect 24668 50540 24724 50596
rect 24668 48130 24724 48132
rect 24668 48078 24670 48130
rect 24670 48078 24722 48130
rect 24722 48078 24724 48130
rect 24668 48076 24724 48078
rect 25004 48076 25060 48132
rect 24668 47068 24724 47124
rect 25340 50540 25396 50596
rect 25900 54514 25956 54516
rect 25900 54462 25902 54514
rect 25902 54462 25954 54514
rect 25954 54462 25956 54514
rect 25900 54460 25956 54462
rect 26012 53730 26068 53732
rect 26012 53678 26014 53730
rect 26014 53678 26066 53730
rect 26066 53678 26068 53730
rect 26012 53676 26068 53678
rect 25676 48914 25732 48916
rect 25676 48862 25678 48914
rect 25678 48862 25730 48914
rect 25730 48862 25732 48914
rect 25676 48860 25732 48862
rect 25228 48300 25284 48356
rect 25900 48300 25956 48356
rect 25676 47346 25732 47348
rect 25676 47294 25678 47346
rect 25678 47294 25730 47346
rect 25730 47294 25732 47346
rect 25676 47292 25732 47294
rect 24668 45052 24724 45108
rect 25452 45106 25508 45108
rect 25452 45054 25454 45106
rect 25454 45054 25506 45106
rect 25506 45054 25508 45106
rect 25452 45052 25508 45054
rect 25900 46620 25956 46676
rect 26236 57036 26292 57092
rect 26236 54572 26292 54628
rect 26572 58380 26628 58436
rect 26572 57372 26628 57428
rect 26908 61292 26964 61348
rect 26796 59724 26852 59780
rect 26796 58380 26852 58436
rect 26684 53676 26740 53732
rect 27020 59890 27076 59892
rect 27020 59838 27022 59890
rect 27022 59838 27074 59890
rect 27074 59838 27076 59890
rect 27020 59836 27076 59838
rect 26796 57148 26852 57204
rect 27132 58434 27188 58436
rect 27132 58382 27134 58434
rect 27134 58382 27186 58434
rect 27186 58382 27188 58434
rect 27132 58380 27188 58382
rect 27132 57260 27188 57316
rect 26908 53618 26964 53620
rect 26908 53566 26910 53618
rect 26910 53566 26962 53618
rect 26962 53566 26964 53618
rect 26908 53564 26964 53566
rect 26460 52220 26516 52276
rect 26572 51490 26628 51492
rect 26572 51438 26574 51490
rect 26574 51438 26626 51490
rect 26626 51438 26628 51490
rect 26572 51436 26628 51438
rect 26236 50482 26292 50484
rect 26236 50430 26238 50482
rect 26238 50430 26290 50482
rect 26290 50430 26292 50482
rect 26236 50428 26292 50430
rect 27020 50540 27076 50596
rect 27580 50818 27636 50820
rect 27580 50766 27582 50818
rect 27582 50766 27634 50818
rect 27634 50766 27636 50818
rect 27580 50764 27636 50766
rect 27244 50540 27300 50596
rect 27804 58434 27860 58436
rect 27804 58382 27806 58434
rect 27806 58382 27858 58434
rect 27858 58382 27860 58434
rect 27804 58380 27860 58382
rect 28252 63922 28308 63924
rect 28252 63870 28254 63922
rect 28254 63870 28306 63922
rect 28306 63870 28308 63922
rect 28252 63868 28308 63870
rect 28364 62354 28420 62356
rect 28364 62302 28366 62354
rect 28366 62302 28418 62354
rect 28418 62302 28420 62354
rect 28364 62300 28420 62302
rect 28588 64988 28644 65044
rect 28700 63922 28756 63924
rect 28700 63870 28702 63922
rect 28702 63870 28754 63922
rect 28754 63870 28756 63922
rect 28700 63868 28756 63870
rect 28140 59836 28196 59892
rect 28028 58156 28084 58212
rect 27916 57650 27972 57652
rect 27916 57598 27918 57650
rect 27918 57598 27970 57650
rect 27970 57598 27972 57650
rect 27916 57596 27972 57598
rect 27804 53788 27860 53844
rect 27804 50706 27860 50708
rect 27804 50654 27806 50706
rect 27806 50654 27858 50706
rect 27858 50654 27860 50706
rect 27804 50652 27860 50654
rect 28028 54684 28084 54740
rect 28140 54460 28196 54516
rect 28252 53788 28308 53844
rect 28140 52834 28196 52836
rect 28140 52782 28142 52834
rect 28142 52782 28194 52834
rect 28194 52782 28196 52834
rect 28140 52780 28196 52782
rect 26796 49196 26852 49252
rect 28140 51996 28196 52052
rect 28028 50764 28084 50820
rect 26796 48860 26852 48916
rect 26124 47458 26180 47460
rect 26124 47406 26126 47458
rect 26126 47406 26178 47458
rect 26178 47406 26180 47458
rect 26124 47404 26180 47406
rect 26572 47068 26628 47124
rect 26236 46674 26292 46676
rect 26236 46622 26238 46674
rect 26238 46622 26290 46674
rect 26290 46622 26292 46674
rect 26236 46620 26292 46622
rect 26236 46284 26292 46340
rect 27692 49250 27748 49252
rect 27692 49198 27694 49250
rect 27694 49198 27746 49250
rect 27746 49198 27748 49250
rect 27692 49196 27748 49198
rect 27356 47068 27412 47124
rect 27244 45724 27300 45780
rect 25676 45106 25732 45108
rect 25676 45054 25678 45106
rect 25678 45054 25730 45106
rect 25730 45054 25732 45106
rect 25676 45052 25732 45054
rect 25676 44604 25732 44660
rect 24668 43820 24724 43876
rect 25340 43426 25396 43428
rect 25340 43374 25342 43426
rect 25342 43374 25394 43426
rect 25394 43374 25396 43426
rect 25340 43372 25396 43374
rect 24668 41580 24724 41636
rect 24220 41298 24276 41300
rect 24220 41246 24222 41298
rect 24222 41246 24274 41298
rect 24274 41246 24276 41298
rect 24220 41244 24276 41246
rect 24220 39506 24276 39508
rect 24220 39454 24222 39506
rect 24222 39454 24274 39506
rect 24274 39454 24276 39506
rect 24220 39452 24276 39454
rect 20748 36764 20804 36820
rect 21420 36258 21476 36260
rect 21420 36206 21422 36258
rect 21422 36206 21474 36258
rect 21474 36206 21476 36258
rect 21420 36204 21476 36206
rect 21756 37154 21812 37156
rect 21756 37102 21758 37154
rect 21758 37102 21810 37154
rect 21810 37102 21812 37154
rect 21756 37100 21812 37102
rect 21644 35532 21700 35588
rect 22540 37772 22596 37828
rect 20636 33852 20692 33908
rect 20748 33740 20804 33796
rect 21756 34018 21812 34020
rect 21756 33966 21758 34018
rect 21758 33966 21810 34018
rect 21810 33966 21812 34018
rect 21756 33964 21812 33966
rect 21420 33852 21476 33908
rect 21644 33740 21700 33796
rect 23548 36204 23604 36260
rect 19516 31836 19572 31892
rect 19964 31890 20020 31892
rect 19964 31838 19966 31890
rect 19966 31838 20018 31890
rect 20018 31838 20020 31890
rect 19964 31836 20020 31838
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19628 30882 19684 30884
rect 19628 30830 19630 30882
rect 19630 30830 19682 30882
rect 19682 30830 19684 30882
rect 19628 30828 19684 30830
rect 18732 30156 18788 30212
rect 20076 30156 20132 30212
rect 19852 30044 19908 30100
rect 20636 30044 20692 30100
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20636 29484 20692 29540
rect 21420 29538 21476 29540
rect 21420 29486 21422 29538
rect 21422 29486 21474 29538
rect 21474 29486 21476 29538
rect 21420 29484 21476 29486
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19404 27020 19460 27076
rect 18732 26012 18788 26068
rect 18508 23100 18564 23156
rect 18956 23212 19012 23268
rect 18620 22930 18676 22932
rect 18620 22878 18622 22930
rect 18622 22878 18674 22930
rect 18674 22878 18676 22930
rect 18620 22876 18676 22878
rect 18508 22764 18564 22820
rect 18620 21474 18676 21476
rect 18620 21422 18622 21474
rect 18622 21422 18674 21474
rect 18674 21422 18676 21474
rect 18620 21420 18676 21422
rect 18284 18338 18340 18340
rect 18284 18286 18286 18338
rect 18286 18286 18338 18338
rect 18338 18286 18340 18338
rect 18284 18284 18340 18286
rect 17948 17612 18004 17668
rect 20524 27746 20580 27748
rect 20524 27694 20526 27746
rect 20526 27694 20578 27746
rect 20578 27694 20580 27746
rect 20524 27692 20580 27694
rect 22764 33346 22820 33348
rect 22764 33294 22766 33346
rect 22766 33294 22818 33346
rect 22818 33294 22820 33346
rect 22764 33292 22820 33294
rect 23548 32396 23604 32452
rect 22316 30210 22372 30212
rect 22316 30158 22318 30210
rect 22318 30158 22370 30210
rect 22370 30158 22372 30210
rect 22316 30156 22372 30158
rect 21868 27692 21924 27748
rect 21308 27074 21364 27076
rect 21308 27022 21310 27074
rect 21310 27022 21362 27074
rect 21362 27022 21364 27074
rect 21308 27020 21364 27022
rect 23884 29484 23940 29540
rect 23436 28700 23492 28756
rect 23212 28364 23268 28420
rect 22316 28252 22372 28308
rect 22764 27970 22820 27972
rect 22764 27918 22766 27970
rect 22766 27918 22818 27970
rect 22818 27918 22820 27970
rect 22764 27916 22820 27918
rect 21980 27132 22036 27188
rect 22316 27020 22372 27076
rect 24892 40962 24948 40964
rect 24892 40910 24894 40962
rect 24894 40910 24946 40962
rect 24946 40910 24948 40962
rect 24892 40908 24948 40910
rect 24668 40684 24724 40740
rect 24780 39340 24836 39396
rect 24780 39004 24836 39060
rect 24444 37212 24500 37268
rect 24668 36204 24724 36260
rect 24556 33852 24612 33908
rect 24220 33346 24276 33348
rect 24220 33294 24222 33346
rect 24222 33294 24274 33346
rect 24274 33294 24276 33346
rect 24220 33292 24276 33294
rect 24668 32450 24724 32452
rect 24668 32398 24670 32450
rect 24670 32398 24722 32450
rect 24722 32398 24724 32450
rect 24668 32396 24724 32398
rect 24556 31500 24612 31556
rect 24444 29708 24500 29764
rect 24444 28754 24500 28756
rect 24444 28702 24446 28754
rect 24446 28702 24498 28754
rect 24498 28702 24500 28754
rect 24444 28700 24500 28702
rect 23996 28476 24052 28532
rect 22540 26962 22596 26964
rect 22540 26910 22542 26962
rect 22542 26910 22594 26962
rect 22594 26910 22596 26962
rect 22540 26908 22596 26910
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20972 26796 21028 26852
rect 20972 26178 21028 26180
rect 20972 26126 20974 26178
rect 20974 26126 21026 26178
rect 21026 26126 21028 26178
rect 20972 26124 21028 26126
rect 21420 26124 21476 26180
rect 22092 25564 22148 25620
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19740 24610 19796 24612
rect 19740 24558 19742 24610
rect 19742 24558 19794 24610
rect 19794 24558 19796 24610
rect 19740 24556 19796 24558
rect 20188 24498 20244 24500
rect 20188 24446 20190 24498
rect 20190 24446 20242 24498
rect 20242 24446 20244 24498
rect 20188 24444 20244 24446
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19628 23266 19684 23268
rect 19628 23214 19630 23266
rect 19630 23214 19682 23266
rect 19682 23214 19684 23266
rect 19628 23212 19684 23214
rect 19180 22652 19236 22708
rect 19516 22316 19572 22372
rect 18956 20636 19012 20692
rect 19516 20188 19572 20244
rect 19068 20018 19124 20020
rect 19068 19966 19070 20018
rect 19070 19966 19122 20018
rect 19122 19966 19124 20018
rect 19068 19964 19124 19966
rect 18732 18450 18788 18452
rect 18732 18398 18734 18450
rect 18734 18398 18786 18450
rect 18786 18398 18788 18450
rect 18732 18396 18788 18398
rect 18956 18284 19012 18340
rect 18844 17836 18900 17892
rect 18732 17554 18788 17556
rect 18732 17502 18734 17554
rect 18734 17502 18786 17554
rect 18786 17502 18788 17554
rect 18732 17500 18788 17502
rect 17836 16882 17892 16884
rect 17836 16830 17838 16882
rect 17838 16830 17890 16882
rect 17890 16830 17892 16882
rect 17836 16828 17892 16830
rect 18620 16882 18676 16884
rect 18620 16830 18622 16882
rect 18622 16830 18674 16882
rect 18674 16830 18676 16882
rect 18620 16828 18676 16830
rect 19180 17666 19236 17668
rect 19180 17614 19182 17666
rect 19182 17614 19234 17666
rect 19234 17614 19236 17666
rect 19180 17612 19236 17614
rect 20524 22428 20580 22484
rect 21420 22482 21476 22484
rect 21420 22430 21422 22482
rect 21422 22430 21474 22482
rect 21474 22430 21476 22482
rect 21420 22428 21476 22430
rect 22092 23938 22148 23940
rect 22092 23886 22094 23938
rect 22094 23886 22146 23938
rect 22146 23886 22148 23938
rect 22092 23884 22148 23886
rect 22316 24722 22372 24724
rect 22316 24670 22318 24722
rect 22318 24670 22370 24722
rect 22370 24670 22372 24722
rect 22316 24668 22372 24670
rect 22204 22594 22260 22596
rect 22204 22542 22206 22594
rect 22206 22542 22258 22594
rect 22258 22542 22260 22594
rect 22204 22540 22260 22542
rect 20972 22316 21028 22372
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20860 21586 20916 21588
rect 20860 21534 20862 21586
rect 20862 21534 20914 21586
rect 20914 21534 20916 21586
rect 20860 21532 20916 21534
rect 21644 20188 21700 20244
rect 22428 21420 22484 21476
rect 23212 26908 23268 26964
rect 24108 27804 24164 27860
rect 23884 26796 23940 26852
rect 23212 26236 23268 26292
rect 22988 24556 23044 24612
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 17836 19684 17892
rect 20412 18172 20468 18228
rect 18172 16098 18228 16100
rect 18172 16046 18174 16098
rect 18174 16046 18226 16098
rect 18226 16046 18228 16098
rect 18172 16044 18228 16046
rect 18060 14476 18116 14532
rect 19180 16716 19236 16772
rect 19292 17106 19348 17108
rect 19292 17054 19294 17106
rect 19294 17054 19346 17106
rect 19346 17054 19348 17106
rect 19292 17052 19348 17054
rect 19516 17052 19572 17108
rect 19404 15372 19460 15428
rect 19068 14530 19124 14532
rect 19068 14478 19070 14530
rect 19070 14478 19122 14530
rect 19122 14478 19124 14530
rect 19068 14476 19124 14478
rect 18396 13916 18452 13972
rect 18844 14418 18900 14420
rect 18844 14366 18846 14418
rect 18846 14366 18898 14418
rect 18898 14366 18900 14418
rect 18844 14364 18900 14366
rect 17724 13132 17780 13188
rect 17612 12348 17668 12404
rect 15260 9938 15316 9940
rect 15260 9886 15262 9938
rect 15262 9886 15314 9938
rect 15314 9886 15316 9938
rect 15260 9884 15316 9886
rect 14924 8988 14980 9044
rect 14588 8316 14644 8372
rect 14364 7474 14420 7476
rect 14364 7422 14366 7474
rect 14366 7422 14418 7474
rect 14418 7422 14420 7474
rect 14364 7420 14420 7422
rect 14252 6636 14308 6692
rect 15372 9548 15428 9604
rect 15148 8930 15204 8932
rect 15148 8878 15150 8930
rect 15150 8878 15202 8930
rect 15202 8878 15204 8930
rect 15148 8876 15204 8878
rect 15148 7756 15204 7812
rect 14588 6188 14644 6244
rect 15372 7756 15428 7812
rect 16604 9042 16660 9044
rect 16604 8990 16606 9042
rect 16606 8990 16658 9042
rect 16658 8990 16660 9042
rect 16604 8988 16660 8990
rect 17836 11676 17892 11732
rect 16044 7474 16100 7476
rect 16044 7422 16046 7474
rect 16046 7422 16098 7474
rect 16098 7422 16100 7474
rect 16044 7420 16100 7422
rect 17948 8988 18004 9044
rect 17948 8316 18004 8372
rect 17500 6524 17556 6580
rect 15484 6188 15540 6244
rect 14476 6018 14532 6020
rect 14476 5966 14478 6018
rect 14478 5966 14530 6018
rect 14530 5966 14532 6018
rect 14476 5964 14532 5966
rect 14700 5906 14756 5908
rect 14700 5854 14702 5906
rect 14702 5854 14754 5906
rect 14754 5854 14756 5906
rect 14700 5852 14756 5854
rect 13468 5068 13524 5124
rect 14924 5794 14980 5796
rect 14924 5742 14926 5794
rect 14926 5742 14978 5794
rect 14978 5742 14980 5794
rect 14924 5740 14980 5742
rect 13804 5180 13860 5236
rect 14812 5292 14868 5348
rect 13244 4338 13300 4340
rect 13244 4286 13246 4338
rect 13246 4286 13298 4338
rect 13298 4286 13300 4338
rect 13244 4284 13300 4286
rect 14700 4172 14756 4228
rect 15708 5346 15764 5348
rect 15708 5294 15710 5346
rect 15710 5294 15762 5346
rect 15762 5294 15764 5346
rect 15708 5292 15764 5294
rect 15484 5234 15540 5236
rect 15484 5182 15486 5234
rect 15486 5182 15538 5234
rect 15538 5182 15540 5234
rect 15484 5180 15540 5182
rect 15820 5180 15876 5236
rect 15148 4844 15204 4900
rect 15148 4284 15204 4340
rect 16492 4898 16548 4900
rect 16492 4846 16494 4898
rect 16494 4846 16546 4898
rect 16546 4846 16548 4898
rect 16492 4844 16548 4846
rect 17052 4898 17108 4900
rect 17052 4846 17054 4898
rect 17054 4846 17106 4898
rect 17106 4846 17108 4898
rect 17052 4844 17108 4846
rect 18284 6412 18340 6468
rect 19516 13804 19572 13860
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20412 17276 20468 17332
rect 20044 17220 20100 17222
rect 20188 17106 20244 17108
rect 20188 17054 20190 17106
rect 20190 17054 20242 17106
rect 20242 17054 20244 17106
rect 20188 17052 20244 17054
rect 20412 16156 20468 16212
rect 20188 16044 20244 16100
rect 19740 15820 19796 15876
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20188 15484 20244 15540
rect 19740 14642 19796 14644
rect 19740 14590 19742 14642
rect 19742 14590 19794 14642
rect 19794 14590 19796 14642
rect 19740 14588 19796 14590
rect 20188 14642 20244 14644
rect 20188 14590 20190 14642
rect 20190 14590 20242 14642
rect 20242 14590 20244 14642
rect 20188 14588 20244 14590
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 18620 12178 18676 12180
rect 18620 12126 18622 12178
rect 18622 12126 18674 12178
rect 18674 12126 18676 12178
rect 18620 12124 18676 12126
rect 19068 12012 19124 12068
rect 18732 11676 18788 11732
rect 19068 11676 19124 11732
rect 19180 12124 19236 12180
rect 18844 8370 18900 8372
rect 18844 8318 18846 8370
rect 18846 8318 18898 8370
rect 18898 8318 18900 8370
rect 18844 8316 18900 8318
rect 19852 13916 19908 13972
rect 20076 13916 20132 13972
rect 20188 13858 20244 13860
rect 20188 13806 20190 13858
rect 20190 13806 20242 13858
rect 20242 13806 20244 13858
rect 20188 13804 20244 13806
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20412 14364 20468 14420
rect 22540 20524 22596 20580
rect 21308 17500 21364 17556
rect 22092 17276 22148 17332
rect 21308 16828 21364 16884
rect 20636 16044 20692 16100
rect 21084 16716 21140 16772
rect 22316 17052 22372 17108
rect 22540 19964 22596 20020
rect 21868 15426 21924 15428
rect 21868 15374 21870 15426
rect 21870 15374 21922 15426
rect 21922 15374 21924 15426
rect 21868 15372 21924 15374
rect 22540 15820 22596 15876
rect 22764 23884 22820 23940
rect 23884 26236 23940 26292
rect 23996 27132 24052 27188
rect 23996 26124 24052 26180
rect 22764 20972 22820 21028
rect 23100 22370 23156 22372
rect 23100 22318 23102 22370
rect 23102 22318 23154 22370
rect 23154 22318 23156 22370
rect 23100 22316 23156 22318
rect 22764 20132 22820 20188
rect 22876 20524 22932 20580
rect 23436 21474 23492 21476
rect 23436 21422 23438 21474
rect 23438 21422 23490 21474
rect 23490 21422 23492 21474
rect 23436 21420 23492 21422
rect 24332 23996 24388 24052
rect 24332 23826 24388 23828
rect 24332 23774 24334 23826
rect 24334 23774 24386 23826
rect 24386 23774 24388 23826
rect 24332 23772 24388 23774
rect 24332 22316 24388 22372
rect 23996 21756 24052 21812
rect 23884 21532 23940 21588
rect 23436 20300 23492 20356
rect 23548 20748 23604 20804
rect 23212 19234 23268 19236
rect 23212 19182 23214 19234
rect 23214 19182 23266 19234
rect 23266 19182 23268 19234
rect 23212 19180 23268 19182
rect 23100 18508 23156 18564
rect 23212 18674 23268 18676
rect 23212 18622 23214 18674
rect 23214 18622 23266 18674
rect 23266 18622 23268 18674
rect 23212 18620 23268 18622
rect 22764 16156 22820 16212
rect 22540 14588 22596 14644
rect 21756 13132 21812 13188
rect 21868 12460 21924 12516
rect 21420 12124 21476 12180
rect 21868 12124 21924 12180
rect 20188 8540 20244 8596
rect 19068 6636 19124 6692
rect 18620 6466 18676 6468
rect 18620 6414 18622 6466
rect 18622 6414 18674 6466
rect 18674 6414 18676 6466
rect 18620 6412 18676 6414
rect 17724 5180 17780 5236
rect 18620 5906 18676 5908
rect 18620 5854 18622 5906
rect 18622 5854 18674 5906
rect 18674 5854 18676 5906
rect 18620 5852 18676 5854
rect 18732 5292 18788 5348
rect 17500 4844 17556 4900
rect 18396 4508 18452 4564
rect 17500 4338 17556 4340
rect 17500 4286 17502 4338
rect 17502 4286 17554 4338
rect 17554 4286 17556 4338
rect 17500 4284 17556 4286
rect 18284 4284 18340 4340
rect 18060 3666 18116 3668
rect 18060 3614 18062 3666
rect 18062 3614 18114 3666
rect 18114 3614 18116 3666
rect 18060 3612 18116 3614
rect 20076 8316 20132 8372
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20300 6690 20356 6692
rect 20300 6638 20302 6690
rect 20302 6638 20354 6690
rect 20354 6638 20356 6690
rect 20300 6636 20356 6638
rect 19404 6524 19460 6580
rect 19516 6466 19572 6468
rect 19516 6414 19518 6466
rect 19518 6414 19570 6466
rect 19570 6414 19572 6466
rect 19516 6412 19572 6414
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 23548 18450 23604 18452
rect 23548 18398 23550 18450
rect 23550 18398 23602 18450
rect 23602 18398 23604 18450
rect 23548 18396 23604 18398
rect 23772 20972 23828 21028
rect 23884 20914 23940 20916
rect 23884 20862 23886 20914
rect 23886 20862 23938 20914
rect 23938 20862 23940 20914
rect 23884 20860 23940 20862
rect 24108 20860 24164 20916
rect 23996 20524 24052 20580
rect 23996 20018 24052 20020
rect 23996 19966 23998 20018
rect 23998 19966 24050 20018
rect 24050 19966 24052 20018
rect 23996 19964 24052 19966
rect 24668 27916 24724 27972
rect 24668 27132 24724 27188
rect 25452 38444 25508 38500
rect 25788 41298 25844 41300
rect 25788 41246 25790 41298
rect 25790 41246 25842 41298
rect 25842 41246 25844 41298
rect 25788 41244 25844 41246
rect 26684 44940 26740 44996
rect 26236 44604 26292 44660
rect 26124 44210 26180 44212
rect 26124 44158 26126 44210
rect 26126 44158 26178 44210
rect 26178 44158 26180 44210
rect 26124 44156 26180 44158
rect 26684 44156 26740 44212
rect 26460 44098 26516 44100
rect 26460 44046 26462 44098
rect 26462 44046 26514 44098
rect 26514 44046 26516 44098
rect 26460 44044 26516 44046
rect 27132 44940 27188 44996
rect 26012 42140 26068 42196
rect 26012 40908 26068 40964
rect 26460 40796 26516 40852
rect 26124 39618 26180 39620
rect 26124 39566 26126 39618
rect 26126 39566 26178 39618
rect 26178 39566 26180 39618
rect 26124 39564 26180 39566
rect 26236 39506 26292 39508
rect 26236 39454 26238 39506
rect 26238 39454 26290 39506
rect 26290 39454 26292 39506
rect 26236 39452 26292 39454
rect 25564 37324 25620 37380
rect 25564 37100 25620 37156
rect 25116 36316 25172 36372
rect 25004 33292 25060 33348
rect 24556 26796 24612 26852
rect 25228 32396 25284 32452
rect 25004 31948 25060 32004
rect 24556 26012 24612 26068
rect 26460 39116 26516 39172
rect 26460 38780 26516 38836
rect 26572 37884 26628 37940
rect 25900 36876 25956 36932
rect 25788 36482 25844 36484
rect 25788 36430 25790 36482
rect 25790 36430 25842 36482
rect 25842 36430 25844 36482
rect 25788 36428 25844 36430
rect 26348 36876 26404 36932
rect 26460 36652 26516 36708
rect 26124 36594 26180 36596
rect 26124 36542 26126 36594
rect 26126 36542 26178 36594
rect 26178 36542 26180 36594
rect 26124 36540 26180 36542
rect 26460 36428 26516 36484
rect 25900 36316 25956 36372
rect 26124 36370 26180 36372
rect 26124 36318 26126 36370
rect 26126 36318 26178 36370
rect 26178 36318 26180 36370
rect 26124 36316 26180 36318
rect 27020 44828 27076 44884
rect 27020 43932 27076 43988
rect 27020 43372 27076 43428
rect 26796 41186 26852 41188
rect 26796 41134 26798 41186
rect 26798 41134 26850 41186
rect 26850 41134 26852 41186
rect 26796 41132 26852 41134
rect 27356 45164 27412 45220
rect 27356 44492 27412 44548
rect 27580 47292 27636 47348
rect 27692 45612 27748 45668
rect 27692 44994 27748 44996
rect 27692 44942 27694 44994
rect 27694 44942 27746 44994
rect 27746 44942 27748 44994
rect 27692 44940 27748 44942
rect 28252 51548 28308 51604
rect 28252 50706 28308 50708
rect 28252 50654 28254 50706
rect 28254 50654 28306 50706
rect 28306 50654 28308 50706
rect 28252 50652 28308 50654
rect 28476 58210 28532 58212
rect 28476 58158 28478 58210
rect 28478 58158 28530 58210
rect 28530 58158 28532 58210
rect 28476 58156 28532 58158
rect 28476 57148 28532 57204
rect 29036 70194 29092 70196
rect 29036 70142 29038 70194
rect 29038 70142 29090 70194
rect 29090 70142 29092 70194
rect 29036 70140 29092 70142
rect 29260 72322 29316 72324
rect 29260 72270 29262 72322
rect 29262 72270 29314 72322
rect 29314 72270 29316 72322
rect 29260 72268 29316 72270
rect 33180 76188 33236 76244
rect 33964 76188 34020 76244
rect 32060 75682 32116 75684
rect 32060 75630 32062 75682
rect 32062 75630 32114 75682
rect 32114 75630 32116 75682
rect 32060 75628 32116 75630
rect 30380 74002 30436 74004
rect 30380 73950 30382 74002
rect 30382 73950 30434 74002
rect 30434 73950 30436 74002
rect 30380 73948 30436 73950
rect 32508 74786 32564 74788
rect 32508 74734 32510 74786
rect 32510 74734 32562 74786
rect 32562 74734 32564 74786
rect 32508 74732 32564 74734
rect 33404 74786 33460 74788
rect 33404 74734 33406 74786
rect 33406 74734 33458 74786
rect 33458 74734 33460 74786
rect 33404 74732 33460 74734
rect 33628 75516 33684 75572
rect 33628 75010 33684 75012
rect 33628 74958 33630 75010
rect 33630 74958 33682 75010
rect 33682 74958 33684 75010
rect 33628 74956 33684 74958
rect 34188 74786 34244 74788
rect 34188 74734 34190 74786
rect 34190 74734 34242 74786
rect 34242 74734 34244 74786
rect 34188 74732 34244 74734
rect 30044 73164 30100 73220
rect 30828 72546 30884 72548
rect 30828 72494 30830 72546
rect 30830 72494 30882 72546
rect 30882 72494 30884 72546
rect 30828 72492 30884 72494
rect 30268 72322 30324 72324
rect 30268 72270 30270 72322
rect 30270 72270 30322 72322
rect 30322 72270 30324 72322
rect 30268 72268 30324 72270
rect 29484 70140 29540 70196
rect 29932 70194 29988 70196
rect 29932 70142 29934 70194
rect 29934 70142 29986 70194
rect 29986 70142 29988 70194
rect 29932 70140 29988 70142
rect 29260 69916 29316 69972
rect 29708 70082 29764 70084
rect 29708 70030 29710 70082
rect 29710 70030 29762 70082
rect 29762 70030 29764 70082
rect 29708 70028 29764 70030
rect 29596 69132 29652 69188
rect 30716 69916 30772 69972
rect 30828 69132 30884 69188
rect 31164 70194 31220 70196
rect 31164 70142 31166 70194
rect 31166 70142 31218 70194
rect 31218 70142 31220 70194
rect 31164 70140 31220 70142
rect 29372 62300 29428 62356
rect 29148 59164 29204 59220
rect 29484 58156 29540 58212
rect 28812 54460 28868 54516
rect 28588 54402 28644 54404
rect 28588 54350 28590 54402
rect 28590 54350 28642 54402
rect 28642 54350 28644 54402
rect 28588 54348 28644 54350
rect 28924 54348 28980 54404
rect 28588 53730 28644 53732
rect 28588 53678 28590 53730
rect 28590 53678 28642 53730
rect 28642 53678 28644 53730
rect 28588 53676 28644 53678
rect 28588 52946 28644 52948
rect 28588 52894 28590 52946
rect 28590 52894 28642 52946
rect 28642 52894 28644 52946
rect 28588 52892 28644 52894
rect 29036 53452 29092 53508
rect 29372 53730 29428 53732
rect 29372 53678 29374 53730
rect 29374 53678 29426 53730
rect 29426 53678 29428 53730
rect 29372 53676 29428 53678
rect 29148 52780 29204 52836
rect 28924 52220 28980 52276
rect 28924 50428 28980 50484
rect 28028 49250 28084 49252
rect 28028 49198 28030 49250
rect 28030 49198 28082 49250
rect 28082 49198 28084 49250
rect 28028 49196 28084 49198
rect 28252 49868 28308 49924
rect 28364 48242 28420 48244
rect 28364 48190 28366 48242
rect 28366 48190 28418 48242
rect 28418 48190 28420 48242
rect 28364 48188 28420 48190
rect 27916 47068 27972 47124
rect 27916 44828 27972 44884
rect 28140 47404 28196 47460
rect 28140 46786 28196 46788
rect 28140 46734 28142 46786
rect 28142 46734 28194 46786
rect 28194 46734 28196 46786
rect 28140 46732 28196 46734
rect 28028 44604 28084 44660
rect 28140 45388 28196 45444
rect 27468 44380 27524 44436
rect 27356 43484 27412 43540
rect 27580 43932 27636 43988
rect 27244 43372 27300 43428
rect 27132 42028 27188 42084
rect 27020 41804 27076 41860
rect 27468 41410 27524 41412
rect 27468 41358 27470 41410
rect 27470 41358 27522 41410
rect 27522 41358 27524 41410
rect 27468 41356 27524 41358
rect 27804 43820 27860 43876
rect 27580 41580 27636 41636
rect 26908 40684 26964 40740
rect 26908 39452 26964 39508
rect 27468 40460 27524 40516
rect 27356 40402 27412 40404
rect 27356 40350 27358 40402
rect 27358 40350 27410 40402
rect 27410 40350 27412 40402
rect 27356 40348 27412 40350
rect 27244 39618 27300 39620
rect 27244 39566 27246 39618
rect 27246 39566 27298 39618
rect 27298 39566 27300 39618
rect 27244 39564 27300 39566
rect 27580 39506 27636 39508
rect 27580 39454 27582 39506
rect 27582 39454 27634 39506
rect 27634 39454 27636 39506
rect 27580 39452 27636 39454
rect 27804 41410 27860 41412
rect 27804 41358 27806 41410
rect 27806 41358 27858 41410
rect 27858 41358 27860 41410
rect 27804 41356 27860 41358
rect 27804 40572 27860 40628
rect 27356 38834 27412 38836
rect 27356 38782 27358 38834
rect 27358 38782 27410 38834
rect 27410 38782 27412 38834
rect 27356 38780 27412 38782
rect 26796 38108 26852 38164
rect 27356 38444 27412 38500
rect 27020 37490 27076 37492
rect 27020 37438 27022 37490
rect 27022 37438 27074 37490
rect 27074 37438 27076 37490
rect 27020 37436 27076 37438
rect 26908 36540 26964 36596
rect 26572 36316 26628 36372
rect 25788 36092 25844 36148
rect 25788 35308 25844 35364
rect 25900 35532 25956 35588
rect 26236 35980 26292 36036
rect 26012 33964 26068 34020
rect 25564 33292 25620 33348
rect 26124 32844 26180 32900
rect 25900 32508 25956 32564
rect 25564 31276 25620 31332
rect 25228 30828 25284 30884
rect 25676 30492 25732 30548
rect 25900 31554 25956 31556
rect 25900 31502 25902 31554
rect 25902 31502 25954 31554
rect 25954 31502 25956 31554
rect 25900 31500 25956 31502
rect 26236 31890 26292 31892
rect 26236 31838 26238 31890
rect 26238 31838 26290 31890
rect 26290 31838 26292 31890
rect 26236 31836 26292 31838
rect 26124 31778 26180 31780
rect 26124 31726 26126 31778
rect 26126 31726 26178 31778
rect 26178 31726 26180 31778
rect 26124 31724 26180 31726
rect 26460 35308 26516 35364
rect 26684 33852 26740 33908
rect 26572 33458 26628 33460
rect 26572 33406 26574 33458
rect 26574 33406 26626 33458
rect 26626 33406 26628 33458
rect 26572 33404 26628 33406
rect 27020 35756 27076 35812
rect 27020 34412 27076 34468
rect 27244 38162 27300 38164
rect 27244 38110 27246 38162
rect 27246 38110 27298 38162
rect 27298 38110 27300 38162
rect 27244 38108 27300 38110
rect 28028 44434 28084 44436
rect 28028 44382 28030 44434
rect 28030 44382 28082 44434
rect 28082 44382 28084 44434
rect 28028 44380 28084 44382
rect 28028 43484 28084 43540
rect 28252 45276 28308 45332
rect 28364 45164 28420 45220
rect 28364 44940 28420 44996
rect 28588 49868 28644 49924
rect 28588 48188 28644 48244
rect 28588 47458 28644 47460
rect 28588 47406 28590 47458
rect 28590 47406 28642 47458
rect 28642 47406 28644 47458
rect 28588 47404 28644 47406
rect 28588 45948 28644 46004
rect 28924 48300 28980 48356
rect 29036 50204 29092 50260
rect 28812 45500 28868 45556
rect 28924 48130 28980 48132
rect 28924 48078 28926 48130
rect 28926 48078 28978 48130
rect 28978 48078 28980 48130
rect 28924 48076 28980 48078
rect 29484 50706 29540 50708
rect 29484 50654 29486 50706
rect 29486 50654 29538 50706
rect 29538 50654 29540 50706
rect 29484 50652 29540 50654
rect 29260 49196 29316 49252
rect 30604 65436 30660 65492
rect 30604 64146 30660 64148
rect 30604 64094 30606 64146
rect 30606 64094 30658 64146
rect 30658 64094 30660 64146
rect 30604 64092 30660 64094
rect 30604 63250 30660 63252
rect 30604 63198 30606 63250
rect 30606 63198 30658 63250
rect 30658 63198 30660 63250
rect 30604 63196 30660 63198
rect 31276 64092 31332 64148
rect 30156 58210 30212 58212
rect 30156 58158 30158 58210
rect 30158 58158 30210 58210
rect 30210 58158 30212 58210
rect 30156 58156 30212 58158
rect 33404 74002 33460 74004
rect 33404 73950 33406 74002
rect 33406 73950 33458 74002
rect 33458 73950 33460 74002
rect 33404 73948 33460 73950
rect 34300 73948 34356 74004
rect 31948 72380 32004 72436
rect 31500 71932 31556 71988
rect 32956 72268 33012 72324
rect 32844 71708 32900 71764
rect 32508 71650 32564 71652
rect 32508 71598 32510 71650
rect 32510 71598 32562 71650
rect 32562 71598 32564 71650
rect 32508 71596 32564 71598
rect 33180 71986 33236 71988
rect 33180 71934 33182 71986
rect 33182 71934 33234 71986
rect 33234 71934 33236 71986
rect 33180 71932 33236 71934
rect 33068 71650 33124 71652
rect 33068 71598 33070 71650
rect 33070 71598 33122 71650
rect 33122 71598 33124 71650
rect 33068 71596 33124 71598
rect 33404 71596 33460 71652
rect 34972 76188 35028 76244
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 34524 74732 34580 74788
rect 35196 74956 35252 75012
rect 33852 72492 33908 72548
rect 34412 71708 34468 71764
rect 31612 70082 31668 70084
rect 31612 70030 31614 70082
rect 31614 70030 31666 70082
rect 31666 70030 31668 70082
rect 31612 70028 31668 70030
rect 32396 69132 32452 69188
rect 31500 67618 31556 67620
rect 31500 67566 31502 67618
rect 31502 67566 31554 67618
rect 31554 67566 31556 67618
rect 31500 67564 31556 67566
rect 31500 63922 31556 63924
rect 31500 63870 31502 63922
rect 31502 63870 31554 63922
rect 31554 63870 31556 63922
rect 31500 63868 31556 63870
rect 30716 60114 30772 60116
rect 30716 60062 30718 60114
rect 30718 60062 30770 60114
rect 30770 60062 30772 60114
rect 30716 60060 30772 60062
rect 30940 59724 30996 59780
rect 30604 58268 30660 58324
rect 30156 57484 30212 57540
rect 30268 57148 30324 57204
rect 29708 54738 29764 54740
rect 29708 54686 29710 54738
rect 29710 54686 29762 54738
rect 29762 54686 29764 54738
rect 29708 54684 29764 54686
rect 29708 53954 29764 53956
rect 29708 53902 29710 53954
rect 29710 53902 29762 53954
rect 29762 53902 29764 53954
rect 29708 53900 29764 53902
rect 29820 53676 29876 53732
rect 29708 53116 29764 53172
rect 29820 52668 29876 52724
rect 29820 51996 29876 52052
rect 29708 51884 29764 51940
rect 29708 50034 29764 50036
rect 29708 49982 29710 50034
rect 29710 49982 29762 50034
rect 29762 49982 29764 50034
rect 29708 49980 29764 49982
rect 29820 50428 29876 50484
rect 29708 49810 29764 49812
rect 29708 49758 29710 49810
rect 29710 49758 29762 49810
rect 29762 49758 29764 49810
rect 29708 49756 29764 49758
rect 29820 49250 29876 49252
rect 29820 49198 29822 49250
rect 29822 49198 29874 49250
rect 29874 49198 29876 49250
rect 29820 49196 29876 49198
rect 29596 47628 29652 47684
rect 29484 47404 29540 47460
rect 29036 46620 29092 46676
rect 29036 45612 29092 45668
rect 28924 45276 28980 45332
rect 29036 45388 29092 45444
rect 29148 44604 29204 44660
rect 29372 45948 29428 46004
rect 29372 45778 29428 45780
rect 29372 45726 29374 45778
rect 29374 45726 29426 45778
rect 29426 45726 29428 45778
rect 29372 45724 29428 45726
rect 29372 44994 29428 44996
rect 29372 44942 29374 44994
rect 29374 44942 29426 44994
rect 29426 44942 29428 44994
rect 29372 44940 29428 44942
rect 28252 43372 28308 43428
rect 28364 44044 28420 44100
rect 28140 42140 28196 42196
rect 28252 42028 28308 42084
rect 28028 41356 28084 41412
rect 28028 40684 28084 40740
rect 28252 41356 28308 41412
rect 28140 40460 28196 40516
rect 28252 40348 28308 40404
rect 28028 38834 28084 38836
rect 28028 38782 28030 38834
rect 28030 38782 28082 38834
rect 28082 38782 28084 38834
rect 28028 38780 28084 38782
rect 27804 38108 27860 38164
rect 27244 37938 27300 37940
rect 27244 37886 27246 37938
rect 27246 37886 27298 37938
rect 27298 37886 27300 37938
rect 27244 37884 27300 37886
rect 27356 37826 27412 37828
rect 27356 37774 27358 37826
rect 27358 37774 27410 37826
rect 27410 37774 27412 37826
rect 27356 37772 27412 37774
rect 27244 37660 27300 37716
rect 27356 37378 27412 37380
rect 27356 37326 27358 37378
rect 27358 37326 27410 37378
rect 27410 37326 27412 37378
rect 27356 37324 27412 37326
rect 27580 37212 27636 37268
rect 27468 36988 27524 37044
rect 27916 36764 27972 36820
rect 27804 36706 27860 36708
rect 27804 36654 27806 36706
rect 27806 36654 27858 36706
rect 27858 36654 27860 36706
rect 27804 36652 27860 36654
rect 27356 36204 27412 36260
rect 27916 35980 27972 36036
rect 26796 32508 26852 32564
rect 27244 35196 27300 35252
rect 26348 30828 26404 30884
rect 26684 31836 26740 31892
rect 27020 33964 27076 34020
rect 26572 31500 26628 31556
rect 26796 31276 26852 31332
rect 26236 30434 26292 30436
rect 26236 30382 26238 30434
rect 26238 30382 26290 30434
rect 26290 30382 26292 30434
rect 26236 30380 26292 30382
rect 25676 29484 25732 29540
rect 25116 28476 25172 28532
rect 26684 30492 26740 30548
rect 26012 29426 26068 29428
rect 26012 29374 26014 29426
rect 26014 29374 26066 29426
rect 26066 29374 26068 29426
rect 26012 29372 26068 29374
rect 26460 29650 26516 29652
rect 26460 29598 26462 29650
rect 26462 29598 26514 29650
rect 26514 29598 26516 29650
rect 26460 29596 26516 29598
rect 25788 28364 25844 28420
rect 25900 28140 25956 28196
rect 26684 28754 26740 28756
rect 26684 28702 26686 28754
rect 26686 28702 26738 28754
rect 26738 28702 26740 28754
rect 26684 28700 26740 28702
rect 25452 27858 25508 27860
rect 25452 27806 25454 27858
rect 25454 27806 25506 27858
rect 25506 27806 25508 27858
rect 25452 27804 25508 27806
rect 25228 27692 25284 27748
rect 25900 27692 25956 27748
rect 25676 27468 25732 27524
rect 26124 27186 26180 27188
rect 26124 27134 26126 27186
rect 26126 27134 26178 27186
rect 26178 27134 26180 27186
rect 26124 27132 26180 27134
rect 25564 26908 25620 26964
rect 25004 26684 25060 26740
rect 24556 23772 24612 23828
rect 24668 24668 24724 24724
rect 25452 26514 25508 26516
rect 25452 26462 25454 26514
rect 25454 26462 25506 26514
rect 25506 26462 25508 26514
rect 25452 26460 25508 26462
rect 25452 26066 25508 26068
rect 25452 26014 25454 26066
rect 25454 26014 25506 26066
rect 25506 26014 25508 26066
rect 25452 26012 25508 26014
rect 25452 24610 25508 24612
rect 25452 24558 25454 24610
rect 25454 24558 25506 24610
rect 25506 24558 25508 24610
rect 25452 24556 25508 24558
rect 24668 23660 24724 23716
rect 26012 26908 26068 26964
rect 26012 23996 26068 24052
rect 24556 22930 24612 22932
rect 24556 22878 24558 22930
rect 24558 22878 24610 22930
rect 24610 22878 24612 22930
rect 24556 22876 24612 22878
rect 23884 19234 23940 19236
rect 23884 19182 23886 19234
rect 23886 19182 23938 19234
rect 23938 19182 23940 19234
rect 23884 19180 23940 19182
rect 23660 17052 23716 17108
rect 24668 21810 24724 21812
rect 24668 21758 24670 21810
rect 24670 21758 24722 21810
rect 24722 21758 24724 21810
rect 24668 21756 24724 21758
rect 25340 22876 25396 22932
rect 25676 22876 25732 22932
rect 25228 21756 25284 21812
rect 25340 20076 25396 20132
rect 24668 19180 24724 19236
rect 24220 18396 24276 18452
rect 23212 14588 23268 14644
rect 22652 13970 22708 13972
rect 22652 13918 22654 13970
rect 22654 13918 22706 13970
rect 22706 13918 22708 13970
rect 22652 13916 22708 13918
rect 22988 13804 23044 13860
rect 22540 13468 22596 13524
rect 21644 11116 21700 11172
rect 20748 8540 20804 8596
rect 21868 8540 21924 8596
rect 21420 6636 21476 6692
rect 22652 12460 22708 12516
rect 22652 11452 22708 11508
rect 22764 11170 22820 11172
rect 22764 11118 22766 11170
rect 22766 11118 22818 11170
rect 22818 11118 22820 11170
rect 22764 11116 22820 11118
rect 23324 15036 23380 15092
rect 23996 15036 24052 15092
rect 25004 18396 25060 18452
rect 24780 17890 24836 17892
rect 24780 17838 24782 17890
rect 24782 17838 24834 17890
rect 24834 17838 24836 17890
rect 24780 17836 24836 17838
rect 23436 13916 23492 13972
rect 23324 13858 23380 13860
rect 23324 13806 23326 13858
rect 23326 13806 23378 13858
rect 23378 13806 23380 13858
rect 23324 13804 23380 13806
rect 23100 12178 23156 12180
rect 23100 12126 23102 12178
rect 23102 12126 23154 12178
rect 23154 12126 23156 12178
rect 23100 12124 23156 12126
rect 23324 11676 23380 11732
rect 23324 11394 23380 11396
rect 23324 11342 23326 11394
rect 23326 11342 23378 11394
rect 23378 11342 23380 11394
rect 23324 11340 23380 11342
rect 24220 14252 24276 14308
rect 24108 13468 24164 13524
rect 23996 13132 24052 13188
rect 24668 16882 24724 16884
rect 24668 16830 24670 16882
rect 24670 16830 24722 16882
rect 24722 16830 24724 16882
rect 24668 16828 24724 16830
rect 25116 16828 25172 16884
rect 25452 18620 25508 18676
rect 25564 16828 25620 16884
rect 26012 22876 26068 22932
rect 26124 22540 26180 22596
rect 25900 21420 25956 21476
rect 26012 20748 26068 20804
rect 26348 19964 26404 20020
rect 26572 27298 26628 27300
rect 26572 27246 26574 27298
rect 26574 27246 26626 27298
rect 26626 27246 26628 27298
rect 26572 27244 26628 27246
rect 26684 27132 26740 27188
rect 26012 18450 26068 18452
rect 26012 18398 26014 18450
rect 26014 18398 26066 18450
rect 26066 18398 26068 18450
rect 26012 18396 26068 18398
rect 26236 17890 26292 17892
rect 26236 17838 26238 17890
rect 26238 17838 26290 17890
rect 26290 17838 26292 17890
rect 26236 17836 26292 17838
rect 27916 34690 27972 34692
rect 27916 34638 27918 34690
rect 27918 34638 27970 34690
rect 27970 34638 27972 34690
rect 27916 34636 27972 34638
rect 27468 34188 27524 34244
rect 27132 33852 27188 33908
rect 27356 33234 27412 33236
rect 27356 33182 27358 33234
rect 27358 33182 27410 33234
rect 27410 33182 27412 33234
rect 27356 33180 27412 33182
rect 27356 32060 27412 32116
rect 26908 29596 26964 29652
rect 27132 29650 27188 29652
rect 27132 29598 27134 29650
rect 27134 29598 27186 29650
rect 27186 29598 27188 29650
rect 27132 29596 27188 29598
rect 26908 28140 26964 28196
rect 27020 27244 27076 27300
rect 27692 31836 27748 31892
rect 27468 30380 27524 30436
rect 27916 29484 27972 29540
rect 27356 29260 27412 29316
rect 28252 38556 28308 38612
rect 28700 44098 28756 44100
rect 28700 44046 28702 44098
rect 28702 44046 28754 44098
rect 28754 44046 28756 44098
rect 28700 44044 28756 44046
rect 29484 44268 29540 44324
rect 29484 44098 29540 44100
rect 29484 44046 29486 44098
rect 29486 44046 29538 44098
rect 29538 44046 29540 44098
rect 29484 44044 29540 44046
rect 28812 42194 28868 42196
rect 28812 42142 28814 42194
rect 28814 42142 28866 42194
rect 28866 42142 28868 42194
rect 28812 42140 28868 42142
rect 28924 40908 28980 40964
rect 28476 40572 28532 40628
rect 28924 40012 28980 40068
rect 28588 39730 28644 39732
rect 28588 39678 28590 39730
rect 28590 39678 28642 39730
rect 28642 39678 28644 39730
rect 28588 39676 28644 39678
rect 28588 39340 28644 39396
rect 28364 38444 28420 38500
rect 28252 37884 28308 37940
rect 28476 37436 28532 37492
rect 28588 37324 28644 37380
rect 28252 36428 28308 36484
rect 28588 36652 28644 36708
rect 28364 36258 28420 36260
rect 28364 36206 28366 36258
rect 28366 36206 28418 36258
rect 28418 36206 28420 36258
rect 28364 36204 28420 36206
rect 28140 35980 28196 36036
rect 28252 32844 28308 32900
rect 28252 32620 28308 32676
rect 28140 31724 28196 31780
rect 28140 30940 28196 30996
rect 27692 27858 27748 27860
rect 27692 27806 27694 27858
rect 27694 27806 27746 27858
rect 27746 27806 27748 27858
rect 27692 27804 27748 27806
rect 27244 27132 27300 27188
rect 27692 27580 27748 27636
rect 26908 26572 26964 26628
rect 27132 26852 27188 26908
rect 27020 24050 27076 24052
rect 27020 23998 27022 24050
rect 27022 23998 27074 24050
rect 27074 23998 27076 24050
rect 27020 23996 27076 23998
rect 26796 23772 26852 23828
rect 26684 23042 26740 23044
rect 26684 22990 26686 23042
rect 26686 22990 26738 23042
rect 26738 22990 26740 23042
rect 26684 22988 26740 22990
rect 27020 23154 27076 23156
rect 27020 23102 27022 23154
rect 27022 23102 27074 23154
rect 27074 23102 27076 23154
rect 27020 23100 27076 23102
rect 27020 22652 27076 22708
rect 26908 22540 26964 22596
rect 26908 22204 26964 22260
rect 26684 21756 26740 21812
rect 26572 20076 26628 20132
rect 25788 16156 25844 16212
rect 24892 14642 24948 14644
rect 24892 14590 24894 14642
rect 24894 14590 24946 14642
rect 24946 14590 24948 14642
rect 24892 14588 24948 14590
rect 24668 13970 24724 13972
rect 24668 13918 24670 13970
rect 24670 13918 24722 13970
rect 24722 13918 24724 13970
rect 24668 13916 24724 13918
rect 24108 11394 24164 11396
rect 24108 11342 24110 11394
rect 24110 11342 24162 11394
rect 24162 11342 24164 11394
rect 24108 11340 24164 11342
rect 23324 10892 23380 10948
rect 23548 9938 23604 9940
rect 23548 9886 23550 9938
rect 23550 9886 23602 9938
rect 23602 9886 23604 9938
rect 23548 9884 23604 9886
rect 20748 6524 20804 6580
rect 19964 5906 20020 5908
rect 19964 5854 19966 5906
rect 19966 5854 20018 5906
rect 20018 5854 20020 5906
rect 19964 5852 20020 5854
rect 19628 5068 19684 5124
rect 23100 5964 23156 6020
rect 21532 5292 21588 5348
rect 20412 5234 20468 5236
rect 20412 5182 20414 5234
rect 20414 5182 20466 5234
rect 20466 5182 20468 5234
rect 20412 5180 20468 5182
rect 22652 5180 22708 5236
rect 21868 5122 21924 5124
rect 21868 5070 21870 5122
rect 21870 5070 21922 5122
rect 21922 5070 21924 5122
rect 21868 5068 21924 5070
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19068 4172 19124 4228
rect 20300 4226 20356 4228
rect 20300 4174 20302 4226
rect 20302 4174 20354 4226
rect 20354 4174 20356 4226
rect 20300 4172 20356 4174
rect 18956 3666 19012 3668
rect 18956 3614 18958 3666
rect 18958 3614 19010 3666
rect 19010 3614 19012 3666
rect 18956 3612 19012 3614
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 18284 2994 18340 2996
rect 18284 2942 18286 2994
rect 18286 2942 18338 2994
rect 18338 2942 18340 2994
rect 18284 2940 18340 2942
rect 19180 2994 19236 2996
rect 19180 2942 19182 2994
rect 19182 2942 19234 2994
rect 19234 2942 19236 2994
rect 19180 2940 19236 2942
rect 19628 2940 19684 2996
rect 24220 9938 24276 9940
rect 24220 9886 24222 9938
rect 24222 9886 24274 9938
rect 24274 9886 24276 9938
rect 24220 9884 24276 9886
rect 25116 13580 25172 13636
rect 27244 26460 27300 26516
rect 27580 26402 27636 26404
rect 27580 26350 27582 26402
rect 27582 26350 27634 26402
rect 27634 26350 27636 26402
rect 27580 26348 27636 26350
rect 27580 23996 27636 24052
rect 28252 26796 28308 26852
rect 28252 26348 28308 26404
rect 27804 23996 27860 24052
rect 27916 23938 27972 23940
rect 27916 23886 27918 23938
rect 27918 23886 27970 23938
rect 27970 23886 27972 23938
rect 27916 23884 27972 23886
rect 28252 23996 28308 24052
rect 27356 22652 27412 22708
rect 27244 22258 27300 22260
rect 27244 22206 27246 22258
rect 27246 22206 27298 22258
rect 27298 22206 27300 22258
rect 27244 22204 27300 22206
rect 28028 22092 28084 22148
rect 28140 21474 28196 21476
rect 28140 21422 28142 21474
rect 28142 21422 28194 21474
rect 28194 21422 28196 21474
rect 28140 21420 28196 21422
rect 26908 17442 26964 17444
rect 26908 17390 26910 17442
rect 26910 17390 26962 17442
rect 26962 17390 26964 17442
rect 26908 17388 26964 17390
rect 26684 16828 26740 16884
rect 27356 17442 27412 17444
rect 27356 17390 27358 17442
rect 27358 17390 27410 17442
rect 27410 17390 27412 17442
rect 27356 17388 27412 17390
rect 28028 16882 28084 16884
rect 28028 16830 28030 16882
rect 28030 16830 28082 16882
rect 28082 16830 28084 16882
rect 28028 16828 28084 16830
rect 27356 16770 27412 16772
rect 27356 16718 27358 16770
rect 27358 16718 27410 16770
rect 27410 16718 27412 16770
rect 27356 16716 27412 16718
rect 26684 13634 26740 13636
rect 26684 13582 26686 13634
rect 26686 13582 26738 13634
rect 26738 13582 26740 13634
rect 26684 13580 26740 13582
rect 27132 14028 27188 14084
rect 26012 12738 26068 12740
rect 26012 12686 26014 12738
rect 26014 12686 26066 12738
rect 26066 12686 26068 12738
rect 26012 12684 26068 12686
rect 25228 12124 25284 12180
rect 24444 11452 24500 11508
rect 25116 11676 25172 11732
rect 25452 11506 25508 11508
rect 25452 11454 25454 11506
rect 25454 11454 25506 11506
rect 25506 11454 25508 11506
rect 25452 11452 25508 11454
rect 25900 11340 25956 11396
rect 23884 5852 23940 5908
rect 23100 5068 23156 5124
rect 23324 5292 23380 5348
rect 23436 5010 23492 5012
rect 23436 4958 23438 5010
rect 23438 4958 23490 5010
rect 23490 4958 23492 5010
rect 23436 4956 23492 4958
rect 26572 9660 26628 9716
rect 26908 9042 26964 9044
rect 26908 8990 26910 9042
rect 26910 8990 26962 9042
rect 26962 8990 26964 9042
rect 26908 8988 26964 8990
rect 27132 13580 27188 13636
rect 27132 8876 27188 8932
rect 28588 32844 28644 32900
rect 28588 32674 28644 32676
rect 28588 32622 28590 32674
rect 28590 32622 28642 32674
rect 28642 32622 28644 32674
rect 28588 32620 28644 32622
rect 28924 38220 28980 38276
rect 28924 37996 28980 38052
rect 28812 37100 28868 37156
rect 29372 43596 29428 43652
rect 29260 43426 29316 43428
rect 29260 43374 29262 43426
rect 29262 43374 29314 43426
rect 29314 43374 29316 43426
rect 29260 43372 29316 43374
rect 29260 42364 29316 42420
rect 29596 41244 29652 41300
rect 29260 41132 29316 41188
rect 29820 47570 29876 47572
rect 29820 47518 29822 47570
rect 29822 47518 29874 47570
rect 29874 47518 29876 47570
rect 29820 47516 29876 47518
rect 30044 54684 30100 54740
rect 30156 53900 30212 53956
rect 30156 52892 30212 52948
rect 30268 51266 30324 51268
rect 30268 51214 30270 51266
rect 30270 51214 30322 51266
rect 30322 51214 30324 51266
rect 30268 51212 30324 51214
rect 30716 57538 30772 57540
rect 30716 57486 30718 57538
rect 30718 57486 30770 57538
rect 30770 57486 30772 57538
rect 30716 57484 30772 57486
rect 30716 56978 30772 56980
rect 30716 56926 30718 56978
rect 30718 56926 30770 56978
rect 30770 56926 30772 56978
rect 30716 56924 30772 56926
rect 32060 65490 32116 65492
rect 32060 65438 32062 65490
rect 32062 65438 32114 65490
rect 32114 65438 32116 65490
rect 32060 65436 32116 65438
rect 32956 69186 33012 69188
rect 32956 69134 32958 69186
rect 32958 69134 33010 69186
rect 33010 69134 33012 69186
rect 32956 69132 33012 69134
rect 33628 70140 33684 70196
rect 33964 71372 34020 71428
rect 33628 69132 33684 69188
rect 33852 69356 33908 69412
rect 32620 66780 32676 66836
rect 32620 65436 32676 65492
rect 33292 66834 33348 66836
rect 33292 66782 33294 66834
rect 33294 66782 33346 66834
rect 33346 66782 33348 66834
rect 33292 66780 33348 66782
rect 33068 65436 33124 65492
rect 33740 67004 33796 67060
rect 31948 63980 32004 64036
rect 31724 62354 31780 62356
rect 31724 62302 31726 62354
rect 31726 62302 31778 62354
rect 31778 62302 31780 62354
rect 31724 62300 31780 62302
rect 32396 63196 32452 63252
rect 32844 64092 32900 64148
rect 32956 63980 33012 64036
rect 33516 65266 33572 65268
rect 33516 65214 33518 65266
rect 33518 65214 33570 65266
rect 33570 65214 33572 65266
rect 33516 65212 33572 65214
rect 34972 73052 35028 73108
rect 34748 71708 34804 71764
rect 34636 70306 34692 70308
rect 34636 70254 34638 70306
rect 34638 70254 34690 70306
rect 34690 70254 34692 70306
rect 34636 70252 34692 70254
rect 34748 70082 34804 70084
rect 34748 70030 34750 70082
rect 34750 70030 34802 70082
rect 34802 70030 34804 70082
rect 34748 70028 34804 70030
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 35308 74002 35364 74004
rect 35308 73950 35310 74002
rect 35310 73950 35362 74002
rect 35362 73950 35364 74002
rect 35308 73948 35364 73950
rect 35980 74002 36036 74004
rect 35980 73950 35982 74002
rect 35982 73950 36034 74002
rect 36034 73950 36036 74002
rect 35980 73948 36036 73950
rect 35644 73836 35700 73892
rect 36988 74956 37044 75012
rect 36316 73836 36372 73892
rect 37436 73948 37492 74004
rect 35644 73052 35700 73108
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 37100 71820 37156 71876
rect 35980 71708 36036 71764
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 36428 71708 36484 71764
rect 35084 70588 35140 70644
rect 35084 70194 35140 70196
rect 35084 70142 35086 70194
rect 35086 70142 35138 70194
rect 35138 70142 35140 70194
rect 35084 70140 35140 70142
rect 35644 70252 35700 70308
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 35868 70082 35924 70084
rect 35868 70030 35870 70082
rect 35870 70030 35922 70082
rect 35922 70030 35924 70082
rect 35868 70028 35924 70030
rect 33964 66892 34020 66948
rect 35868 69410 35924 69412
rect 35868 69358 35870 69410
rect 35870 69358 35922 69410
rect 35922 69358 35924 69410
rect 35868 69356 35924 69358
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 34748 67004 34804 67060
rect 34188 66946 34244 66948
rect 34188 66894 34190 66946
rect 34190 66894 34242 66946
rect 34242 66894 34244 66946
rect 34188 66892 34244 66894
rect 35308 67058 35364 67060
rect 35308 67006 35310 67058
rect 35310 67006 35362 67058
rect 35362 67006 35364 67058
rect 35308 67004 35364 67006
rect 34188 65490 34244 65492
rect 34188 65438 34190 65490
rect 34190 65438 34242 65490
rect 34242 65438 34244 65490
rect 34188 65436 34244 65438
rect 33180 63196 33236 63252
rect 34076 63196 34132 63252
rect 33180 62972 33236 63028
rect 32508 62300 32564 62356
rect 31276 60060 31332 60116
rect 31836 59724 31892 59780
rect 32956 62076 33012 62132
rect 33628 62076 33684 62132
rect 31612 58268 31668 58324
rect 32732 59778 32788 59780
rect 32732 59726 32734 59778
rect 32734 59726 32786 59778
rect 32786 59726 32788 59778
rect 32732 59724 32788 59726
rect 33180 59724 33236 59780
rect 32284 58492 32340 58548
rect 32396 57874 32452 57876
rect 32396 57822 32398 57874
rect 32398 57822 32450 57874
rect 32450 57822 32452 57874
rect 32396 57820 32452 57822
rect 31500 57148 31556 57204
rect 32060 57650 32116 57652
rect 32060 57598 32062 57650
rect 32062 57598 32114 57650
rect 32114 57598 32116 57650
rect 32060 57596 32116 57598
rect 30716 52274 30772 52276
rect 30716 52222 30718 52274
rect 30718 52222 30770 52274
rect 30770 52222 30772 52274
rect 30716 52220 30772 52222
rect 30716 51602 30772 51604
rect 30716 51550 30718 51602
rect 30718 51550 30770 51602
rect 30770 51550 30772 51602
rect 30716 51548 30772 51550
rect 31052 51212 31108 51268
rect 30156 50652 30212 50708
rect 30492 49868 30548 49924
rect 30380 49756 30436 49812
rect 30380 49196 30436 49252
rect 30492 49644 30548 49700
rect 30268 48914 30324 48916
rect 30268 48862 30270 48914
rect 30270 48862 30322 48914
rect 30322 48862 30324 48914
rect 30268 48860 30324 48862
rect 30044 47404 30100 47460
rect 29932 46956 29988 47012
rect 29820 46562 29876 46564
rect 29820 46510 29822 46562
rect 29822 46510 29874 46562
rect 29874 46510 29876 46562
rect 29820 46508 29876 46510
rect 29820 43708 29876 43764
rect 29932 44604 29988 44660
rect 29820 42924 29876 42980
rect 30156 45836 30212 45892
rect 30156 43708 30212 43764
rect 30044 43596 30100 43652
rect 30044 42476 30100 42532
rect 30044 41970 30100 41972
rect 30044 41918 30046 41970
rect 30046 41918 30098 41970
rect 30098 41918 30100 41970
rect 30044 41916 30100 41918
rect 29932 41298 29988 41300
rect 29932 41246 29934 41298
rect 29934 41246 29986 41298
rect 29986 41246 29988 41298
rect 29932 41244 29988 41246
rect 30380 48076 30436 48132
rect 30604 48076 30660 48132
rect 30716 50540 30772 50596
rect 30492 46620 30548 46676
rect 30828 49980 30884 50036
rect 31164 50652 31220 50708
rect 31164 50204 31220 50260
rect 31388 51548 31444 51604
rect 31276 50092 31332 50148
rect 31276 49922 31332 49924
rect 31276 49870 31278 49922
rect 31278 49870 31330 49922
rect 31330 49870 31332 49922
rect 31276 49868 31332 49870
rect 31500 50652 31556 50708
rect 31052 49532 31108 49588
rect 31052 47292 31108 47348
rect 31276 49532 31332 49588
rect 30716 46396 30772 46452
rect 30716 45778 30772 45780
rect 30716 45726 30718 45778
rect 30718 45726 30770 45778
rect 30770 45726 30772 45778
rect 30716 45724 30772 45726
rect 30380 45388 30436 45444
rect 30492 45218 30548 45220
rect 30492 45166 30494 45218
rect 30494 45166 30546 45218
rect 30546 45166 30548 45218
rect 30492 45164 30548 45166
rect 30380 44380 30436 44436
rect 31500 48188 31556 48244
rect 31388 48130 31444 48132
rect 31388 48078 31390 48130
rect 31390 48078 31442 48130
rect 31442 48078 31444 48130
rect 31388 48076 31444 48078
rect 31388 47516 31444 47572
rect 31276 45890 31332 45892
rect 31276 45838 31278 45890
rect 31278 45838 31330 45890
rect 31330 45838 31332 45890
rect 31276 45836 31332 45838
rect 31164 45330 31220 45332
rect 31164 45278 31166 45330
rect 31166 45278 31218 45330
rect 31218 45278 31220 45330
rect 31164 45276 31220 45278
rect 31500 45724 31556 45780
rect 30828 43708 30884 43764
rect 30380 43538 30436 43540
rect 30380 43486 30382 43538
rect 30382 43486 30434 43538
rect 30434 43486 30436 43538
rect 30380 43484 30436 43486
rect 30716 43484 30772 43540
rect 30268 42530 30324 42532
rect 30268 42478 30270 42530
rect 30270 42478 30322 42530
rect 30322 42478 30324 42530
rect 30268 42476 30324 42478
rect 30268 42140 30324 42196
rect 29820 40962 29876 40964
rect 29820 40910 29822 40962
rect 29822 40910 29874 40962
rect 29874 40910 29876 40962
rect 29820 40908 29876 40910
rect 29260 40796 29316 40852
rect 30156 40962 30212 40964
rect 30156 40910 30158 40962
rect 30158 40910 30210 40962
rect 30210 40910 30212 40962
rect 30156 40908 30212 40910
rect 29820 40684 29876 40740
rect 29484 39676 29540 39732
rect 29596 40012 29652 40068
rect 30156 40402 30212 40404
rect 30156 40350 30158 40402
rect 30158 40350 30210 40402
rect 30210 40350 30212 40402
rect 30156 40348 30212 40350
rect 30156 39842 30212 39844
rect 30156 39790 30158 39842
rect 30158 39790 30210 39842
rect 30210 39790 30212 39842
rect 30156 39788 30212 39790
rect 30156 39564 30212 39620
rect 29260 38780 29316 38836
rect 30044 39394 30100 39396
rect 30044 39342 30046 39394
rect 30046 39342 30098 39394
rect 30098 39342 30100 39394
rect 30044 39340 30100 39342
rect 29932 39116 29988 39172
rect 29932 38780 29988 38836
rect 29260 38274 29316 38276
rect 29260 38222 29262 38274
rect 29262 38222 29314 38274
rect 29314 38222 29316 38274
rect 29260 38220 29316 38222
rect 28924 35084 28980 35140
rect 29708 38162 29764 38164
rect 29708 38110 29710 38162
rect 29710 38110 29762 38162
rect 29762 38110 29764 38162
rect 29708 38108 29764 38110
rect 29484 37436 29540 37492
rect 29820 37266 29876 37268
rect 29820 37214 29822 37266
rect 29822 37214 29874 37266
rect 29874 37214 29876 37266
rect 29820 37212 29876 37214
rect 29596 35810 29652 35812
rect 29596 35758 29598 35810
rect 29598 35758 29650 35810
rect 29650 35758 29652 35810
rect 29596 35756 29652 35758
rect 28812 32060 28868 32116
rect 29484 35084 29540 35140
rect 28700 31276 28756 31332
rect 28812 30716 28868 30772
rect 28588 29986 28644 29988
rect 28588 29934 28590 29986
rect 28590 29934 28642 29986
rect 28642 29934 28644 29986
rect 28588 29932 28644 29934
rect 28812 29708 28868 29764
rect 28476 27580 28532 27636
rect 28588 29596 28644 29652
rect 28476 26908 28532 26964
rect 28476 26572 28532 26628
rect 28476 26348 28532 26404
rect 28812 29148 28868 29204
rect 29148 34636 29204 34692
rect 29036 34412 29092 34468
rect 29036 34076 29092 34132
rect 29372 34636 29428 34692
rect 29148 34188 29204 34244
rect 29260 34300 29316 34356
rect 29372 33740 29428 33796
rect 29260 31890 29316 31892
rect 29260 31838 29262 31890
rect 29262 31838 29314 31890
rect 29314 31838 29316 31890
rect 29260 31836 29316 31838
rect 29148 30994 29204 30996
rect 29148 30942 29150 30994
rect 29150 30942 29202 30994
rect 29202 30942 29204 30994
rect 29148 30940 29204 30942
rect 29148 29426 29204 29428
rect 29148 29374 29150 29426
rect 29150 29374 29202 29426
rect 29202 29374 29204 29426
rect 29148 29372 29204 29374
rect 29372 31500 29428 31556
rect 29372 30770 29428 30772
rect 29372 30718 29374 30770
rect 29374 30718 29426 30770
rect 29426 30718 29428 30770
rect 29372 30716 29428 30718
rect 29260 28700 29316 28756
rect 29372 29484 29428 29540
rect 28924 28028 28980 28084
rect 28812 27132 28868 27188
rect 29260 27132 29316 27188
rect 29932 36764 29988 36820
rect 29820 36482 29876 36484
rect 29820 36430 29822 36482
rect 29822 36430 29874 36482
rect 29874 36430 29876 36482
rect 29820 36428 29876 36430
rect 30156 36652 30212 36708
rect 30716 41916 30772 41972
rect 30716 40348 30772 40404
rect 30604 39788 30660 39844
rect 30492 38220 30548 38276
rect 30940 43650 30996 43652
rect 30940 43598 30942 43650
rect 30942 43598 30994 43650
rect 30994 43598 30996 43650
rect 30940 43596 30996 43598
rect 31164 43372 31220 43428
rect 31164 43148 31220 43204
rect 31836 51938 31892 51940
rect 31836 51886 31838 51938
rect 31838 51886 31890 51938
rect 31890 51886 31892 51938
rect 31836 51884 31892 51886
rect 32060 57372 32116 57428
rect 33740 58546 33796 58548
rect 33740 58494 33742 58546
rect 33742 58494 33794 58546
rect 33794 58494 33796 58546
rect 33740 58492 33796 58494
rect 34076 57874 34132 57876
rect 34076 57822 34078 57874
rect 34078 57822 34130 57874
rect 34130 57822 34132 57874
rect 34076 57820 34132 57822
rect 33068 57596 33124 57652
rect 33740 57148 33796 57204
rect 32060 52722 32116 52724
rect 32060 52670 32062 52722
rect 32062 52670 32114 52722
rect 32114 52670 32116 52722
rect 32060 52668 32116 52670
rect 31724 48972 31780 49028
rect 32284 51938 32340 51940
rect 32284 51886 32286 51938
rect 32286 51886 32338 51938
rect 32338 51886 32340 51938
rect 32284 51884 32340 51886
rect 31948 49698 32004 49700
rect 31948 49646 31950 49698
rect 31950 49646 32002 49698
rect 32002 49646 32004 49698
rect 31948 49644 32004 49646
rect 32396 50594 32452 50596
rect 32396 50542 32398 50594
rect 32398 50542 32450 50594
rect 32450 50542 32452 50594
rect 32396 50540 32452 50542
rect 32508 49756 32564 49812
rect 32396 49698 32452 49700
rect 32396 49646 32398 49698
rect 32398 49646 32450 49698
rect 32450 49646 32452 49698
rect 32396 49644 32452 49646
rect 32172 47628 32228 47684
rect 32060 47346 32116 47348
rect 32060 47294 32062 47346
rect 32062 47294 32114 47346
rect 32114 47294 32116 47346
rect 32060 47292 32116 47294
rect 31388 43820 31444 43876
rect 31276 42812 31332 42868
rect 31164 41916 31220 41972
rect 31500 43036 31556 43092
rect 31500 42476 31556 42532
rect 31276 40908 31332 40964
rect 31388 42140 31444 42196
rect 30940 40012 30996 40068
rect 30716 38556 30772 38612
rect 30716 37772 30772 37828
rect 30604 37490 30660 37492
rect 30604 37438 30606 37490
rect 30606 37438 30658 37490
rect 30658 37438 30660 37490
rect 30604 37436 30660 37438
rect 31500 41804 31556 41860
rect 31276 39564 31332 39620
rect 31836 46898 31892 46900
rect 31836 46846 31838 46898
rect 31838 46846 31890 46898
rect 31890 46846 31892 46898
rect 31836 46844 31892 46846
rect 32732 52050 32788 52052
rect 32732 51998 32734 52050
rect 32734 51998 32786 52050
rect 32786 51998 32788 52050
rect 32732 51996 32788 51998
rect 32844 51884 32900 51940
rect 32732 50540 32788 50596
rect 33628 52946 33684 52948
rect 33628 52894 33630 52946
rect 33630 52894 33682 52946
rect 33682 52894 33684 52946
rect 33628 52892 33684 52894
rect 33292 52668 33348 52724
rect 33180 52220 33236 52276
rect 33068 51884 33124 51940
rect 33068 50764 33124 50820
rect 32620 46956 32676 47012
rect 32508 46844 32564 46900
rect 32396 46786 32452 46788
rect 32396 46734 32398 46786
rect 32398 46734 32450 46786
rect 32450 46734 32452 46786
rect 32396 46732 32452 46734
rect 32284 46508 32340 46564
rect 32508 45330 32564 45332
rect 32508 45278 32510 45330
rect 32510 45278 32562 45330
rect 32562 45278 32564 45330
rect 32508 45276 32564 45278
rect 32060 44492 32116 44548
rect 31836 43426 31892 43428
rect 31836 43374 31838 43426
rect 31838 43374 31890 43426
rect 31890 43374 31892 43426
rect 31836 43372 31892 43374
rect 31724 43148 31780 43204
rect 31836 42700 31892 42756
rect 31948 42140 32004 42196
rect 33068 49810 33124 49812
rect 33068 49758 33070 49810
rect 33070 49758 33122 49810
rect 33122 49758 33124 49810
rect 33068 49756 33124 49758
rect 32956 49644 33012 49700
rect 32956 48914 33012 48916
rect 32956 48862 32958 48914
rect 32958 48862 33010 48914
rect 33010 48862 33012 48914
rect 32956 48860 33012 48862
rect 33068 48242 33124 48244
rect 33068 48190 33070 48242
rect 33070 48190 33122 48242
rect 33122 48190 33124 48242
rect 33068 48188 33124 48190
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 35756 66050 35812 66052
rect 35756 65998 35758 66050
rect 35758 65998 35810 66050
rect 35810 65998 35812 66050
rect 35756 65996 35812 65998
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 35644 64092 35700 64148
rect 34524 63980 34580 64036
rect 35196 64034 35252 64036
rect 35196 63982 35198 64034
rect 35198 63982 35250 64034
rect 35250 63982 35252 64034
rect 35196 63980 35252 63982
rect 35308 63922 35364 63924
rect 35308 63870 35310 63922
rect 35310 63870 35362 63922
rect 35362 63870 35364 63922
rect 35308 63868 35364 63870
rect 35756 63868 35812 63924
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 35644 63026 35700 63028
rect 35644 62974 35646 63026
rect 35646 62974 35698 63026
rect 35698 62974 35700 63026
rect 35644 62972 35700 62974
rect 34860 62914 34916 62916
rect 34860 62862 34862 62914
rect 34862 62862 34914 62914
rect 34914 62862 34916 62914
rect 34860 62860 34916 62862
rect 36092 69020 36148 69076
rect 36540 71596 36596 71652
rect 37548 71762 37604 71764
rect 37548 71710 37550 71762
rect 37550 71710 37602 71762
rect 37602 71710 37604 71762
rect 37548 71708 37604 71710
rect 38332 71708 38388 71764
rect 37212 71538 37268 71540
rect 37212 71486 37214 71538
rect 37214 71486 37266 71538
rect 37266 71486 37268 71538
rect 37212 71484 37268 71486
rect 36988 70588 37044 70644
rect 37996 70588 38052 70644
rect 38780 71596 38836 71652
rect 37100 69410 37156 69412
rect 37100 69358 37102 69410
rect 37102 69358 37154 69410
rect 37154 69358 37156 69410
rect 37100 69356 37156 69358
rect 36204 68908 36260 68964
rect 36988 69020 37044 69076
rect 37100 68908 37156 68964
rect 36428 66162 36484 66164
rect 36428 66110 36430 66162
rect 36430 66110 36482 66162
rect 36482 66110 36484 66162
rect 36428 66108 36484 66110
rect 36988 65996 37044 66052
rect 36204 64876 36260 64932
rect 36988 64930 37044 64932
rect 36988 64878 36990 64930
rect 36990 64878 37042 64930
rect 37042 64878 37044 64930
rect 36988 64876 37044 64878
rect 35980 64092 36036 64148
rect 36428 63196 36484 63252
rect 36316 62972 36372 63028
rect 36092 62188 36148 62244
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 34636 59724 34692 59780
rect 34300 58434 34356 58436
rect 34300 58382 34302 58434
rect 34302 58382 34354 58434
rect 34354 58382 34356 58434
rect 34300 58380 34356 58382
rect 34300 56978 34356 56980
rect 34300 56926 34302 56978
rect 34302 56926 34354 56978
rect 34354 56926 34356 56978
rect 34300 56924 34356 56926
rect 33516 52162 33572 52164
rect 33516 52110 33518 52162
rect 33518 52110 33570 52162
rect 33570 52110 33572 52162
rect 33516 52108 33572 52110
rect 33964 51884 34020 51940
rect 33628 50876 33684 50932
rect 33628 50652 33684 50708
rect 33292 46732 33348 46788
rect 33292 46562 33348 46564
rect 33292 46510 33294 46562
rect 33294 46510 33346 46562
rect 33346 46510 33348 46562
rect 33292 46508 33348 46510
rect 33292 45836 33348 45892
rect 33068 44492 33124 44548
rect 33740 50540 33796 50596
rect 33740 49756 33796 49812
rect 33964 49644 34020 49700
rect 34188 54460 34244 54516
rect 34188 52108 34244 52164
rect 34188 51100 34244 51156
rect 33628 45276 33684 45332
rect 33740 49026 33796 49028
rect 33740 48974 33742 49026
rect 33742 48974 33794 49026
rect 33794 48974 33796 49026
rect 33740 48972 33796 48974
rect 33628 45106 33684 45108
rect 33628 45054 33630 45106
rect 33630 45054 33682 45106
rect 33682 45054 33684 45106
rect 33628 45052 33684 45054
rect 33628 44492 33684 44548
rect 32172 43484 32228 43540
rect 32060 42924 32116 42980
rect 31276 37938 31332 37940
rect 31276 37886 31278 37938
rect 31278 37886 31330 37938
rect 31330 37886 31332 37938
rect 31276 37884 31332 37886
rect 30940 37100 30996 37156
rect 31388 37266 31444 37268
rect 31388 37214 31390 37266
rect 31390 37214 31442 37266
rect 31442 37214 31444 37266
rect 31388 37212 31444 37214
rect 30156 36482 30212 36484
rect 30156 36430 30158 36482
rect 30158 36430 30210 36482
rect 30210 36430 30212 36482
rect 30156 36428 30212 36430
rect 30044 35868 30100 35924
rect 30156 35308 30212 35364
rect 29932 34690 29988 34692
rect 29932 34638 29934 34690
rect 29934 34638 29986 34690
rect 29986 34638 29988 34690
rect 29932 34636 29988 34638
rect 29820 34524 29876 34580
rect 29708 34130 29764 34132
rect 29708 34078 29710 34130
rect 29710 34078 29762 34130
rect 29762 34078 29764 34130
rect 29708 34076 29764 34078
rect 29708 32508 29764 32564
rect 30156 34242 30212 34244
rect 30156 34190 30158 34242
rect 30158 34190 30210 34242
rect 30210 34190 30212 34242
rect 30156 34188 30212 34190
rect 30380 33740 30436 33796
rect 30268 33458 30324 33460
rect 30268 33406 30270 33458
rect 30270 33406 30322 33458
rect 30322 33406 30324 33458
rect 30268 33404 30324 33406
rect 30828 36316 30884 36372
rect 30716 35810 30772 35812
rect 30716 35758 30718 35810
rect 30718 35758 30770 35810
rect 30770 35758 30772 35810
rect 30716 35756 30772 35758
rect 30604 33516 30660 33572
rect 30604 33346 30660 33348
rect 30604 33294 30606 33346
rect 30606 33294 30658 33346
rect 30658 33294 30660 33346
rect 30604 33292 30660 33294
rect 30156 31836 30212 31892
rect 30940 35868 30996 35924
rect 31052 36316 31108 36372
rect 30940 35698 30996 35700
rect 30940 35646 30942 35698
rect 30942 35646 30994 35698
rect 30994 35646 30996 35698
rect 30940 35644 30996 35646
rect 30940 35420 30996 35476
rect 31164 35420 31220 35476
rect 31388 35868 31444 35924
rect 31052 34188 31108 34244
rect 30492 31218 30548 31220
rect 30492 31166 30494 31218
rect 30494 31166 30546 31218
rect 30546 31166 30548 31218
rect 30492 31164 30548 31166
rect 29932 29708 29988 29764
rect 30044 29820 30100 29876
rect 30044 29372 30100 29428
rect 30604 28924 30660 28980
rect 29708 28700 29764 28756
rect 29932 28754 29988 28756
rect 29932 28702 29934 28754
rect 29934 28702 29986 28754
rect 29986 28702 29988 28754
rect 29932 28700 29988 28702
rect 30380 28588 30436 28644
rect 30156 28082 30212 28084
rect 30156 28030 30158 28082
rect 30158 28030 30210 28082
rect 30210 28030 30212 28082
rect 30156 28028 30212 28030
rect 29932 27858 29988 27860
rect 29932 27806 29934 27858
rect 29934 27806 29986 27858
rect 29986 27806 29988 27858
rect 29932 27804 29988 27806
rect 29484 27074 29540 27076
rect 29484 27022 29486 27074
rect 29486 27022 29538 27074
rect 29538 27022 29540 27074
rect 29484 27020 29540 27022
rect 29820 27020 29876 27076
rect 29036 26572 29092 26628
rect 29036 26402 29092 26404
rect 29036 26350 29038 26402
rect 29038 26350 29090 26402
rect 29090 26350 29092 26402
rect 29036 26348 29092 26350
rect 29708 25618 29764 25620
rect 29708 25566 29710 25618
rect 29710 25566 29762 25618
rect 29762 25566 29764 25618
rect 29708 25564 29764 25566
rect 29708 25228 29764 25284
rect 30604 27356 30660 27412
rect 30268 27298 30324 27300
rect 30268 27246 30270 27298
rect 30270 27246 30322 27298
rect 30322 27246 30324 27298
rect 30268 27244 30324 27246
rect 30940 31666 30996 31668
rect 30940 31614 30942 31666
rect 30942 31614 30994 31666
rect 30994 31614 30996 31666
rect 30940 31612 30996 31614
rect 31052 31164 31108 31220
rect 30828 29820 30884 29876
rect 31612 37100 31668 37156
rect 31612 36370 31668 36372
rect 31612 36318 31614 36370
rect 31614 36318 31666 36370
rect 31666 36318 31668 36370
rect 31612 36316 31668 36318
rect 32620 42028 32676 42084
rect 32284 41020 32340 41076
rect 32060 40684 32116 40740
rect 31948 40514 32004 40516
rect 31948 40462 31950 40514
rect 31950 40462 32002 40514
rect 32002 40462 32004 40514
rect 31948 40460 32004 40462
rect 31948 39116 32004 39172
rect 32284 40348 32340 40404
rect 32172 40178 32228 40180
rect 32172 40126 32174 40178
rect 32174 40126 32226 40178
rect 32226 40126 32228 40178
rect 32172 40124 32228 40126
rect 32172 39340 32228 39396
rect 32060 37996 32116 38052
rect 32508 39506 32564 39508
rect 32508 39454 32510 39506
rect 32510 39454 32562 39506
rect 32562 39454 32564 39506
rect 32508 39452 32564 39454
rect 32508 38668 32564 38724
rect 31948 37884 32004 37940
rect 31836 37378 31892 37380
rect 31836 37326 31838 37378
rect 31838 37326 31890 37378
rect 31890 37326 31892 37378
rect 31836 37324 31892 37326
rect 31948 37212 32004 37268
rect 31724 36540 31780 36596
rect 31724 35420 31780 35476
rect 31612 31778 31668 31780
rect 31612 31726 31614 31778
rect 31614 31726 31666 31778
rect 31666 31726 31668 31778
rect 31612 31724 31668 31726
rect 32060 36988 32116 37044
rect 31836 34636 31892 34692
rect 31836 33404 31892 33460
rect 31388 31388 31444 31444
rect 31500 30492 31556 30548
rect 31164 30380 31220 30436
rect 31500 30044 31556 30100
rect 31500 29820 31556 29876
rect 31836 31106 31892 31108
rect 31836 31054 31838 31106
rect 31838 31054 31890 31106
rect 31890 31054 31892 31106
rect 31836 31052 31892 31054
rect 32060 34636 32116 34692
rect 32060 31500 32116 31556
rect 32060 30604 32116 30660
rect 32284 38444 32340 38500
rect 32508 38332 32564 38388
rect 32956 43708 33012 43764
rect 33180 43036 33236 43092
rect 33068 42588 33124 42644
rect 33180 42140 33236 42196
rect 33292 41580 33348 41636
rect 33068 41074 33124 41076
rect 33068 41022 33070 41074
rect 33070 41022 33122 41074
rect 33122 41022 33124 41074
rect 33068 41020 33124 41022
rect 33516 44268 33572 44324
rect 33516 42588 33572 42644
rect 33516 41580 33572 41636
rect 33852 45052 33908 45108
rect 33964 43314 34020 43316
rect 33964 43262 33966 43314
rect 33966 43262 34018 43314
rect 34018 43262 34020 43314
rect 33964 43260 34020 43262
rect 33964 42642 34020 42644
rect 33964 42590 33966 42642
rect 33966 42590 34018 42642
rect 34018 42590 34020 42642
rect 33964 42588 34020 42590
rect 33852 41804 33908 41860
rect 33740 41132 33796 41188
rect 33628 40514 33684 40516
rect 33628 40462 33630 40514
rect 33630 40462 33682 40514
rect 33682 40462 33684 40514
rect 33628 40460 33684 40462
rect 33964 40572 34020 40628
rect 33516 40012 33572 40068
rect 33852 40348 33908 40404
rect 33068 39116 33124 39172
rect 33180 39340 33236 39396
rect 33740 39340 33796 39396
rect 32732 37436 32788 37492
rect 32956 36988 33012 37044
rect 32620 36764 32676 36820
rect 32284 36594 32340 36596
rect 32284 36542 32286 36594
rect 32286 36542 32338 36594
rect 32338 36542 32340 36594
rect 32284 36540 32340 36542
rect 33292 38050 33348 38052
rect 33292 37998 33294 38050
rect 33294 37998 33346 38050
rect 33346 37998 33348 38050
rect 33292 37996 33348 37998
rect 32732 35756 32788 35812
rect 32508 35586 32564 35588
rect 32508 35534 32510 35586
rect 32510 35534 32562 35586
rect 32562 35534 32564 35586
rect 32508 35532 32564 35534
rect 32844 35420 32900 35476
rect 32508 35308 32564 35364
rect 32620 34636 32676 34692
rect 32508 33516 32564 33572
rect 32620 32956 32676 33012
rect 32620 32732 32676 32788
rect 32284 31612 32340 31668
rect 32284 31218 32340 31220
rect 32284 31166 32286 31218
rect 32286 31166 32338 31218
rect 32338 31166 32340 31218
rect 32284 31164 32340 31166
rect 32732 31164 32788 31220
rect 32396 30770 32452 30772
rect 32396 30718 32398 30770
rect 32398 30718 32450 30770
rect 32450 30718 32452 30770
rect 32396 30716 32452 30718
rect 31724 29932 31780 29988
rect 31948 29820 32004 29876
rect 32060 30044 32116 30100
rect 31052 28700 31108 28756
rect 30828 27580 30884 27636
rect 30716 27244 30772 27300
rect 30380 25564 30436 25620
rect 29932 23100 29988 23156
rect 28700 22092 28756 22148
rect 29260 22146 29316 22148
rect 29260 22094 29262 22146
rect 29262 22094 29314 22146
rect 29314 22094 29316 22146
rect 29260 22092 29316 22094
rect 29148 17554 29204 17556
rect 29148 17502 29150 17554
rect 29150 17502 29202 17554
rect 29202 17502 29204 17554
rect 29148 17500 29204 17502
rect 28588 15314 28644 15316
rect 28588 15262 28590 15314
rect 28590 15262 28642 15314
rect 28642 15262 28644 15314
rect 28588 15260 28644 15262
rect 28812 16994 28868 16996
rect 28812 16942 28814 16994
rect 28814 16942 28866 16994
rect 28866 16942 28868 16994
rect 28812 16940 28868 16942
rect 28364 14028 28420 14084
rect 28028 13580 28084 13636
rect 27356 12684 27412 12740
rect 28700 14642 28756 14644
rect 28700 14590 28702 14642
rect 28702 14590 28754 14642
rect 28754 14590 28756 14642
rect 28700 14588 28756 14590
rect 28588 12348 28644 12404
rect 28252 11394 28308 11396
rect 28252 11342 28254 11394
rect 28254 11342 28306 11394
rect 28306 11342 28308 11394
rect 28252 11340 28308 11342
rect 27916 9884 27972 9940
rect 27356 9548 27412 9604
rect 27804 9042 27860 9044
rect 27804 8990 27806 9042
rect 27806 8990 27858 9042
rect 27858 8990 27860 9042
rect 27804 8988 27860 8990
rect 27468 8876 27524 8932
rect 25788 6018 25844 6020
rect 25788 5966 25790 6018
rect 25790 5966 25842 6018
rect 25842 5966 25844 6018
rect 25788 5964 25844 5966
rect 25228 5740 25284 5796
rect 24220 4956 24276 5012
rect 24444 5068 24500 5124
rect 26012 5740 26068 5796
rect 24668 4450 24724 4452
rect 24668 4398 24670 4450
rect 24670 4398 24722 4450
rect 24722 4398 24724 4450
rect 24668 4396 24724 4398
rect 25452 5122 25508 5124
rect 25452 5070 25454 5122
rect 25454 5070 25506 5122
rect 25506 5070 25508 5122
rect 25452 5068 25508 5070
rect 26908 6914 26964 6916
rect 26908 6862 26910 6914
rect 26910 6862 26962 6914
rect 26962 6862 26964 6914
rect 26908 6860 26964 6862
rect 27580 6860 27636 6916
rect 27244 6690 27300 6692
rect 27244 6638 27246 6690
rect 27246 6638 27298 6690
rect 27298 6638 27300 6690
rect 27244 6636 27300 6638
rect 26684 6018 26740 6020
rect 26684 5966 26686 6018
rect 26686 5966 26738 6018
rect 26738 5966 26740 6018
rect 26684 5964 26740 5966
rect 25788 5122 25844 5124
rect 25788 5070 25790 5122
rect 25790 5070 25842 5122
rect 25842 5070 25844 5122
rect 25788 5068 25844 5070
rect 23436 2770 23492 2772
rect 23436 2718 23438 2770
rect 23438 2718 23490 2770
rect 23490 2718 23492 2770
rect 23436 2716 23492 2718
rect 24220 2770 24276 2772
rect 24220 2718 24222 2770
rect 24222 2718 24274 2770
rect 24274 2718 24276 2770
rect 24220 2716 24276 2718
rect 26460 5122 26516 5124
rect 26460 5070 26462 5122
rect 26462 5070 26514 5122
rect 26514 5070 26516 5122
rect 26460 5068 26516 5070
rect 27244 6076 27300 6132
rect 27132 5068 27188 5124
rect 26012 4450 26068 4452
rect 26012 4398 26014 4450
rect 26014 4398 26066 4450
rect 26066 4398 26068 4450
rect 26012 4396 26068 4398
rect 28588 9602 28644 9604
rect 28588 9550 28590 9602
rect 28590 9550 28642 9602
rect 28642 9550 28644 9602
rect 28588 9548 28644 9550
rect 29148 15260 29204 15316
rect 29484 20690 29540 20692
rect 29484 20638 29486 20690
rect 29486 20638 29538 20690
rect 29538 20638 29540 20690
rect 29484 20636 29540 20638
rect 30604 23324 30660 23380
rect 30380 23154 30436 23156
rect 30380 23102 30382 23154
rect 30382 23102 30434 23154
rect 30434 23102 30436 23154
rect 30380 23100 30436 23102
rect 31052 27132 31108 27188
rect 31948 29426 32004 29428
rect 31948 29374 31950 29426
rect 31950 29374 32002 29426
rect 32002 29374 32004 29426
rect 31948 29372 32004 29374
rect 30828 27074 30884 27076
rect 30828 27022 30830 27074
rect 30830 27022 30882 27074
rect 30882 27022 30884 27074
rect 30828 27020 30884 27022
rect 31276 26962 31332 26964
rect 31276 26910 31278 26962
rect 31278 26910 31330 26962
rect 31330 26910 31332 26962
rect 31276 26908 31332 26910
rect 32172 29650 32228 29652
rect 32172 29598 32174 29650
rect 32174 29598 32226 29650
rect 32226 29598 32228 29650
rect 32172 29596 32228 29598
rect 32396 29538 32452 29540
rect 32396 29486 32398 29538
rect 32398 29486 32450 29538
rect 32450 29486 32452 29538
rect 32396 29484 32452 29486
rect 32508 29372 32564 29428
rect 32172 28812 32228 28868
rect 32284 28924 32340 28980
rect 32620 30604 32676 30660
rect 32620 29148 32676 29204
rect 32620 28252 32676 28308
rect 31500 26796 31556 26852
rect 31388 26460 31444 26516
rect 31612 25788 31668 25844
rect 31164 25004 31220 25060
rect 31164 23660 31220 23716
rect 31612 23714 31668 23716
rect 31612 23662 31614 23714
rect 31614 23662 31666 23714
rect 31666 23662 31668 23714
rect 31612 23660 31668 23662
rect 31612 23100 31668 23156
rect 30828 21644 30884 21700
rect 30492 21586 30548 21588
rect 30492 21534 30494 21586
rect 30494 21534 30546 21586
rect 30546 21534 30548 21586
rect 30492 21532 30548 21534
rect 30380 20524 30436 20580
rect 29708 16994 29764 16996
rect 29708 16942 29710 16994
rect 29710 16942 29762 16994
rect 29762 16942 29764 16994
rect 29708 16940 29764 16942
rect 29484 16658 29540 16660
rect 29484 16606 29486 16658
rect 29486 16606 29538 16658
rect 29538 16606 29540 16658
rect 29484 16604 29540 16606
rect 29932 17388 29988 17444
rect 30268 17106 30324 17108
rect 30268 17054 30270 17106
rect 30270 17054 30322 17106
rect 30322 17054 30324 17106
rect 30268 17052 30324 17054
rect 29932 16604 29988 16660
rect 30268 16604 30324 16660
rect 29820 14700 29876 14756
rect 29260 14588 29316 14644
rect 29372 14476 29428 14532
rect 29932 14476 29988 14532
rect 29596 14306 29652 14308
rect 29596 14254 29598 14306
rect 29598 14254 29650 14306
rect 29650 14254 29652 14306
rect 29596 14252 29652 14254
rect 29932 13132 29988 13188
rect 29596 12738 29652 12740
rect 29596 12686 29598 12738
rect 29598 12686 29650 12738
rect 29650 12686 29652 12738
rect 29596 12684 29652 12686
rect 29932 12348 29988 12404
rect 29708 12236 29764 12292
rect 28924 9884 28980 9940
rect 29932 11564 29988 11620
rect 28924 9548 28980 9604
rect 30604 20412 30660 20468
rect 30156 14700 30212 14756
rect 30380 14530 30436 14532
rect 30380 14478 30382 14530
rect 30382 14478 30434 14530
rect 30434 14478 30436 14530
rect 30380 14476 30436 14478
rect 30156 14364 30212 14420
rect 30492 14252 30548 14308
rect 30380 12684 30436 12740
rect 30268 11564 30324 11620
rect 29372 9826 29428 9828
rect 29372 9774 29374 9826
rect 29374 9774 29426 9826
rect 29426 9774 29428 9826
rect 29372 9772 29428 9774
rect 31164 21532 31220 21588
rect 31052 17724 31108 17780
rect 30828 15874 30884 15876
rect 30828 15822 30830 15874
rect 30830 15822 30882 15874
rect 30882 15822 30884 15874
rect 30828 15820 30884 15822
rect 31948 27580 32004 27636
rect 31948 27356 32004 27412
rect 32172 27244 32228 27300
rect 31948 24780 32004 24836
rect 32060 27132 32116 27188
rect 33068 35644 33124 35700
rect 33628 39058 33684 39060
rect 33628 39006 33630 39058
rect 33630 39006 33682 39058
rect 33682 39006 33684 39058
rect 33628 39004 33684 39006
rect 34076 41692 34132 41748
rect 34524 58492 34580 58548
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 35084 58380 35140 58436
rect 34972 56978 35028 56980
rect 34972 56926 34974 56978
rect 34974 56926 35026 56978
rect 35026 56926 35028 56978
rect 34972 56924 35028 56926
rect 34860 54514 34916 54516
rect 34860 54462 34862 54514
rect 34862 54462 34914 54514
rect 34914 54462 34916 54514
rect 34860 54460 34916 54462
rect 34636 52892 34692 52948
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 35420 57036 35476 57092
rect 35420 56252 35476 56308
rect 35532 56924 35588 56980
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 35196 55468 35252 55524
rect 36092 55468 36148 55524
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35532 53116 35588 53172
rect 35532 52946 35588 52948
rect 35532 52894 35534 52946
rect 35534 52894 35586 52946
rect 35586 52894 35588 52946
rect 35532 52892 35588 52894
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35644 52444 35700 52500
rect 34524 51938 34580 51940
rect 34524 51886 34526 51938
rect 34526 51886 34578 51938
rect 34578 51886 34580 51938
rect 34524 51884 34580 51886
rect 34972 51212 35028 51268
rect 34860 50876 34916 50932
rect 34860 50594 34916 50596
rect 34860 50542 34862 50594
rect 34862 50542 34914 50594
rect 34914 50542 34916 50594
rect 34860 50540 34916 50542
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 34748 50428 34804 50484
rect 35756 50706 35812 50708
rect 35756 50654 35758 50706
rect 35758 50654 35810 50706
rect 35810 50654 35812 50706
rect 35756 50652 35812 50654
rect 34748 49810 34804 49812
rect 34748 49758 34750 49810
rect 34750 49758 34802 49810
rect 34802 49758 34804 49810
rect 34748 49756 34804 49758
rect 34972 48748 35028 48804
rect 36204 52444 36260 52500
rect 35980 51266 36036 51268
rect 35980 51214 35982 51266
rect 35982 51214 36034 51266
rect 36034 51214 36036 51266
rect 35980 51212 36036 51214
rect 36204 50594 36260 50596
rect 36204 50542 36206 50594
rect 36206 50542 36258 50594
rect 36258 50542 36260 50594
rect 36204 50540 36260 50542
rect 35868 50428 35924 50484
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35644 48748 35700 48804
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 34412 47458 34468 47460
rect 34412 47406 34414 47458
rect 34414 47406 34466 47458
rect 34466 47406 34468 47458
rect 34412 47404 34468 47406
rect 34636 47068 34692 47124
rect 34636 46786 34692 46788
rect 34636 46734 34638 46786
rect 34638 46734 34690 46786
rect 34690 46734 34692 46786
rect 34636 46732 34692 46734
rect 34300 45330 34356 45332
rect 34300 45278 34302 45330
rect 34302 45278 34354 45330
rect 34354 45278 34356 45330
rect 34300 45276 34356 45278
rect 34636 45276 34692 45332
rect 34636 44716 34692 44772
rect 35084 47516 35140 47572
rect 35532 47234 35588 47236
rect 35532 47182 35534 47234
rect 35534 47182 35586 47234
rect 35586 47182 35588 47234
rect 35532 47180 35588 47182
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35196 45890 35252 45892
rect 35196 45838 35198 45890
rect 35198 45838 35250 45890
rect 35250 45838 35252 45890
rect 35196 45836 35252 45838
rect 35532 45836 35588 45892
rect 35084 45612 35140 45668
rect 35084 45330 35140 45332
rect 35084 45278 35086 45330
rect 35086 45278 35138 45330
rect 35138 45278 35140 45330
rect 35084 45276 35140 45278
rect 34972 44940 35028 44996
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35196 44098 35252 44100
rect 35196 44046 35198 44098
rect 35198 44046 35250 44098
rect 35250 44046 35252 44098
rect 35196 44044 35252 44046
rect 34748 42476 34804 42532
rect 34972 42364 35028 42420
rect 34524 41580 34580 41636
rect 34860 42140 34916 42196
rect 34300 40012 34356 40068
rect 34076 39676 34132 39732
rect 34188 39900 34244 39956
rect 33964 39506 34020 39508
rect 33964 39454 33966 39506
rect 33966 39454 34018 39506
rect 34018 39454 34020 39506
rect 33964 39452 34020 39454
rect 33740 37884 33796 37940
rect 33628 37324 33684 37380
rect 33740 37212 33796 37268
rect 33404 35980 33460 36036
rect 33404 35420 33460 35476
rect 33180 34412 33236 34468
rect 33628 34354 33684 34356
rect 33628 34302 33630 34354
rect 33630 34302 33682 34354
rect 33682 34302 33684 34354
rect 33628 34300 33684 34302
rect 33068 33740 33124 33796
rect 33292 33516 33348 33572
rect 33180 32956 33236 33012
rect 33180 31500 33236 31556
rect 33068 30604 33124 30660
rect 33404 32396 33460 32452
rect 33628 31948 33684 32004
rect 33740 31724 33796 31780
rect 33628 31612 33684 31668
rect 32956 29596 33012 29652
rect 33404 30716 33460 30772
rect 33740 30604 33796 30660
rect 32956 27692 33012 27748
rect 32620 27244 32676 27300
rect 32620 26572 32676 26628
rect 32396 26236 32452 26292
rect 32284 25228 32340 25284
rect 32060 23660 32116 23716
rect 31500 21586 31556 21588
rect 31500 21534 31502 21586
rect 31502 21534 31554 21586
rect 31554 21534 31556 21586
rect 31500 21532 31556 21534
rect 31388 20860 31444 20916
rect 31612 18508 31668 18564
rect 32172 23100 32228 23156
rect 32396 24444 32452 24500
rect 33292 29986 33348 29988
rect 33292 29934 33294 29986
rect 33294 29934 33346 29986
rect 33346 29934 33348 29986
rect 33292 29932 33348 29934
rect 33180 29820 33236 29876
rect 33740 30322 33796 30324
rect 33740 30270 33742 30322
rect 33742 30270 33794 30322
rect 33794 30270 33796 30322
rect 33740 30268 33796 30270
rect 33964 37436 34020 37492
rect 33964 33964 34020 34020
rect 33964 33292 34020 33348
rect 34300 39116 34356 39172
rect 34636 41132 34692 41188
rect 34524 40962 34580 40964
rect 34524 40910 34526 40962
rect 34526 40910 34578 40962
rect 34578 40910 34580 40962
rect 34524 40908 34580 40910
rect 34412 38556 34468 38612
rect 34300 37938 34356 37940
rect 34300 37886 34302 37938
rect 34302 37886 34354 37938
rect 34354 37886 34356 37938
rect 34300 37884 34356 37886
rect 34188 36988 34244 37044
rect 34188 35756 34244 35812
rect 35420 43596 35476 43652
rect 35532 43484 35588 43540
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35196 42866 35252 42868
rect 35196 42814 35198 42866
rect 35198 42814 35250 42866
rect 35250 42814 35252 42866
rect 35196 42812 35252 42814
rect 35756 45388 35812 45444
rect 38332 66892 38388 66948
rect 37772 66162 37828 66164
rect 37772 66110 37774 66162
rect 37774 66110 37826 66162
rect 37826 66110 37828 66162
rect 37772 66108 37828 66110
rect 37324 63138 37380 63140
rect 37324 63086 37326 63138
rect 37326 63086 37378 63138
rect 37378 63086 37380 63138
rect 37324 63084 37380 63086
rect 37324 62188 37380 62244
rect 37996 63250 38052 63252
rect 37996 63198 37998 63250
rect 37998 63198 38050 63250
rect 38050 63198 38052 63250
rect 37996 63196 38052 63198
rect 37548 61404 37604 61460
rect 37548 58434 37604 58436
rect 37548 58382 37550 58434
rect 37550 58382 37602 58434
rect 37602 58382 37604 58434
rect 37548 58380 37604 58382
rect 37884 58156 37940 58212
rect 37660 57932 37716 57988
rect 37324 54572 37380 54628
rect 37436 51938 37492 51940
rect 37436 51886 37438 51938
rect 37438 51886 37490 51938
rect 37490 51886 37492 51938
rect 37436 51884 37492 51886
rect 36540 49698 36596 49700
rect 36540 49646 36542 49698
rect 36542 49646 36594 49698
rect 36594 49646 36596 49698
rect 36540 49644 36596 49646
rect 36540 48748 36596 48804
rect 36092 47458 36148 47460
rect 36092 47406 36094 47458
rect 36094 47406 36146 47458
rect 36146 47406 36148 47458
rect 36092 47404 36148 47406
rect 36764 48354 36820 48356
rect 36764 48302 36766 48354
rect 36766 48302 36818 48354
rect 36818 48302 36820 48354
rect 36764 48300 36820 48302
rect 37100 48802 37156 48804
rect 37100 48750 37102 48802
rect 37102 48750 37154 48802
rect 37154 48750 37156 48802
rect 37100 48748 37156 48750
rect 37100 48412 37156 48468
rect 37324 47516 37380 47572
rect 37212 47404 37268 47460
rect 36540 47068 36596 47124
rect 36204 46844 36260 46900
rect 35980 46060 36036 46116
rect 36092 45890 36148 45892
rect 36092 45838 36094 45890
rect 36094 45838 36146 45890
rect 36146 45838 36148 45890
rect 36092 45836 36148 45838
rect 35980 44380 36036 44436
rect 35868 43596 35924 43652
rect 35644 42140 35700 42196
rect 34860 40684 34916 40740
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 34636 39004 34692 39060
rect 34748 40012 34804 40068
rect 34524 37212 34580 37268
rect 34300 34972 34356 35028
rect 34412 34300 34468 34356
rect 34300 34018 34356 34020
rect 34300 33966 34302 34018
rect 34302 33966 34354 34018
rect 34354 33966 34356 34018
rect 34300 33964 34356 33966
rect 35532 41356 35588 41412
rect 35532 41074 35588 41076
rect 35532 41022 35534 41074
rect 35534 41022 35586 41074
rect 35586 41022 35588 41074
rect 35532 41020 35588 41022
rect 34972 39394 35028 39396
rect 34972 39342 34974 39394
rect 34974 39342 35026 39394
rect 35026 39342 35028 39394
rect 34972 39340 35028 39342
rect 35084 40908 35140 40964
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 39730 35252 39732
rect 35196 39678 35198 39730
rect 35198 39678 35250 39730
rect 35250 39678 35252 39730
rect 35196 39676 35252 39678
rect 35868 42140 35924 42196
rect 35980 42028 36036 42084
rect 36204 43708 36260 43764
rect 36316 43596 36372 43652
rect 35868 40460 35924 40516
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 34748 37100 34804 37156
rect 34636 36652 34692 36708
rect 34860 36988 34916 37044
rect 34748 36204 34804 36260
rect 34748 34188 34804 34244
rect 34748 33964 34804 34020
rect 34636 33628 34692 33684
rect 34076 32450 34132 32452
rect 34076 32398 34078 32450
rect 34078 32398 34130 32450
rect 34130 32398 34132 32450
rect 34076 32396 34132 32398
rect 34300 33068 34356 33124
rect 34636 32844 34692 32900
rect 34412 32732 34468 32788
rect 34300 32396 34356 32452
rect 33964 31052 34020 31108
rect 33964 30492 34020 30548
rect 34188 31388 34244 31444
rect 34300 31052 34356 31108
rect 34300 30268 34356 30324
rect 33740 29820 33796 29876
rect 34076 29820 34132 29876
rect 33516 28866 33572 28868
rect 33516 28814 33518 28866
rect 33518 28814 33570 28866
rect 33570 28814 33572 28866
rect 33516 28812 33572 28814
rect 33740 28754 33796 28756
rect 33740 28702 33742 28754
rect 33742 28702 33794 28754
rect 33794 28702 33796 28754
rect 33740 28700 33796 28702
rect 33628 28252 33684 28308
rect 33068 26290 33124 26292
rect 33068 26238 33070 26290
rect 33070 26238 33122 26290
rect 33122 26238 33124 26290
rect 33068 26236 33124 26238
rect 32508 23884 32564 23940
rect 32396 23772 32452 23828
rect 32508 23660 32564 23716
rect 32844 24444 32900 24500
rect 32956 24892 33012 24948
rect 32844 23714 32900 23716
rect 32844 23662 32846 23714
rect 32846 23662 32898 23714
rect 32898 23662 32900 23714
rect 32844 23660 32900 23662
rect 31948 21810 32004 21812
rect 31948 21758 31950 21810
rect 31950 21758 32002 21810
rect 32002 21758 32004 21810
rect 31948 21756 32004 21758
rect 32284 20914 32340 20916
rect 32284 20862 32286 20914
rect 32286 20862 32338 20914
rect 32338 20862 32340 20914
rect 32284 20860 32340 20862
rect 32060 20076 32116 20132
rect 31388 16658 31444 16660
rect 31388 16606 31390 16658
rect 31390 16606 31442 16658
rect 31442 16606 31444 16658
rect 31388 16604 31444 16606
rect 31164 15202 31220 15204
rect 31164 15150 31166 15202
rect 31166 15150 31218 15202
rect 31218 15150 31220 15202
rect 31164 15148 31220 15150
rect 30828 14588 30884 14644
rect 30828 14418 30884 14420
rect 30828 14366 30830 14418
rect 30830 14366 30882 14418
rect 30882 14366 30884 14418
rect 30828 14364 30884 14366
rect 30940 12236 30996 12292
rect 31612 15820 31668 15876
rect 32060 16604 32116 16660
rect 31724 14588 31780 14644
rect 32060 14364 32116 14420
rect 32060 13692 32116 13748
rect 32396 18284 32452 18340
rect 33180 24780 33236 24836
rect 33068 23938 33124 23940
rect 33068 23886 33070 23938
rect 33070 23886 33122 23938
rect 33122 23886 33124 23938
rect 33068 23884 33124 23886
rect 32956 20860 33012 20916
rect 33180 23378 33236 23380
rect 33180 23326 33182 23378
rect 33182 23326 33234 23378
rect 33234 23326 33236 23378
rect 33180 23324 33236 23326
rect 33180 20076 33236 20132
rect 32620 17500 32676 17556
rect 33068 18284 33124 18340
rect 33180 17778 33236 17780
rect 33180 17726 33182 17778
rect 33182 17726 33234 17778
rect 33234 17726 33236 17778
rect 33180 17724 33236 17726
rect 33404 25282 33460 25284
rect 33404 25230 33406 25282
rect 33406 25230 33458 25282
rect 33458 25230 33460 25282
rect 33404 25228 33460 25230
rect 33404 23100 33460 23156
rect 33516 21756 33572 21812
rect 33740 19852 33796 19908
rect 33516 17724 33572 17780
rect 33628 17164 33684 17220
rect 33516 16994 33572 16996
rect 33516 16942 33518 16994
rect 33518 16942 33570 16994
rect 33570 16942 33572 16994
rect 33516 16940 33572 16942
rect 33964 29148 34020 29204
rect 34748 31164 34804 31220
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35308 36652 35364 36708
rect 35868 38556 35924 38612
rect 35868 38162 35924 38164
rect 35868 38110 35870 38162
rect 35870 38110 35922 38162
rect 35922 38110 35924 38162
rect 35868 38108 35924 38110
rect 35644 37996 35700 38052
rect 35532 36258 35588 36260
rect 35532 36206 35534 36258
rect 35534 36206 35586 36258
rect 35586 36206 35588 36258
rect 35532 36204 35588 36206
rect 35196 35698 35252 35700
rect 35196 35646 35198 35698
rect 35198 35646 35250 35698
rect 35250 35646 35252 35698
rect 35196 35644 35252 35646
rect 36092 41468 36148 41524
rect 36092 38050 36148 38052
rect 36092 37998 36094 38050
rect 36094 37998 36146 38050
rect 36146 37998 36148 38050
rect 36092 37996 36148 37998
rect 36316 41132 36372 41188
rect 36540 41020 36596 41076
rect 36652 44940 36708 44996
rect 36316 40796 36372 40852
rect 37100 46786 37156 46788
rect 37100 46734 37102 46786
rect 37102 46734 37154 46786
rect 37154 46734 37156 46786
rect 37100 46732 37156 46734
rect 39228 66332 39284 66388
rect 39900 66386 39956 66388
rect 39900 66334 39902 66386
rect 39902 66334 39954 66386
rect 39954 66334 39956 66386
rect 39900 66332 39956 66334
rect 39004 65378 39060 65380
rect 39004 65326 39006 65378
rect 39006 65326 39058 65378
rect 39058 65326 39060 65378
rect 39004 65324 39060 65326
rect 39676 65378 39732 65380
rect 39676 65326 39678 65378
rect 39678 65326 39730 65378
rect 39730 65326 39732 65378
rect 39676 65324 39732 65326
rect 38444 63196 38500 63252
rect 39228 63250 39284 63252
rect 39228 63198 39230 63250
rect 39230 63198 39282 63250
rect 39282 63198 39284 63250
rect 39228 63196 39284 63198
rect 38444 61404 38500 61460
rect 38108 57932 38164 57988
rect 37660 52162 37716 52164
rect 37660 52110 37662 52162
rect 37662 52110 37714 52162
rect 37714 52110 37716 52162
rect 37660 52108 37716 52110
rect 37660 51548 37716 51604
rect 37660 50706 37716 50708
rect 37660 50654 37662 50706
rect 37662 50654 37714 50706
rect 37714 50654 37716 50706
rect 37660 50652 37716 50654
rect 38220 58044 38276 58100
rect 40124 61516 40180 61572
rect 39116 58156 39172 58212
rect 40796 61516 40852 61572
rect 39676 59724 39732 59780
rect 38780 57762 38836 57764
rect 38780 57710 38782 57762
rect 38782 57710 38834 57762
rect 38834 57710 38836 57762
rect 38780 57708 38836 57710
rect 42812 60620 42868 60676
rect 43820 60674 43876 60676
rect 43820 60622 43822 60674
rect 43822 60622 43874 60674
rect 43874 60622 43876 60674
rect 43820 60620 43876 60622
rect 40572 59778 40628 59780
rect 40572 59726 40574 59778
rect 40574 59726 40626 59778
rect 40626 59726 40628 59778
rect 40572 59724 40628 59726
rect 41468 59724 41524 59780
rect 39676 57708 39732 57764
rect 38668 56306 38724 56308
rect 38668 56254 38670 56306
rect 38670 56254 38722 56306
rect 38722 56254 38724 56306
rect 38668 56252 38724 56254
rect 41020 56252 41076 56308
rect 40684 56028 40740 56084
rect 38332 54626 38388 54628
rect 38332 54574 38334 54626
rect 38334 54574 38386 54626
rect 38386 54574 38388 54626
rect 38332 54572 38388 54574
rect 38668 54402 38724 54404
rect 38668 54350 38670 54402
rect 38670 54350 38722 54402
rect 38722 54350 38724 54402
rect 38668 54348 38724 54350
rect 38892 53170 38948 53172
rect 38892 53118 38894 53170
rect 38894 53118 38946 53170
rect 38946 53118 38948 53170
rect 38892 53116 38948 53118
rect 38332 52220 38388 52276
rect 38668 51884 38724 51940
rect 40236 52780 40292 52836
rect 39900 51996 39956 52052
rect 39228 51548 39284 51604
rect 38332 51324 38388 51380
rect 37660 48972 37716 49028
rect 37660 48466 37716 48468
rect 37660 48414 37662 48466
rect 37662 48414 37714 48466
rect 37714 48414 37716 48466
rect 37660 48412 37716 48414
rect 37772 48300 37828 48356
rect 37100 44994 37156 44996
rect 37100 44942 37102 44994
rect 37102 44942 37154 44994
rect 37154 44942 37156 44994
rect 37100 44940 37156 44942
rect 37212 44098 37268 44100
rect 37212 44046 37214 44098
rect 37214 44046 37266 44098
rect 37266 44046 37268 44098
rect 37212 44044 37268 44046
rect 37772 45612 37828 45668
rect 37548 45388 37604 45444
rect 37548 44268 37604 44324
rect 37660 44156 37716 44212
rect 37212 43484 37268 43540
rect 36764 42700 36820 42756
rect 36988 42140 37044 42196
rect 37100 41356 37156 41412
rect 36764 40684 36820 40740
rect 36428 40124 36484 40180
rect 37548 42754 37604 42756
rect 37548 42702 37550 42754
rect 37550 42702 37602 42754
rect 37602 42702 37604 42754
rect 37548 42700 37604 42702
rect 37436 42642 37492 42644
rect 37436 42590 37438 42642
rect 37438 42590 37490 42642
rect 37490 42590 37492 42642
rect 37436 42588 37492 42590
rect 37324 42082 37380 42084
rect 37324 42030 37326 42082
rect 37326 42030 37378 42082
rect 37378 42030 37380 42082
rect 37324 42028 37380 42030
rect 36764 40124 36820 40180
rect 37100 39730 37156 39732
rect 37100 39678 37102 39730
rect 37102 39678 37154 39730
rect 37154 39678 37156 39730
rect 37100 39676 37156 39678
rect 37660 41020 37716 41076
rect 37548 39788 37604 39844
rect 37772 40236 37828 40292
rect 36652 39116 36708 39172
rect 36204 37266 36260 37268
rect 36204 37214 36206 37266
rect 36206 37214 36258 37266
rect 36258 37214 36260 37266
rect 36204 37212 36260 37214
rect 36092 36428 36148 36484
rect 35644 35532 35700 35588
rect 35084 35420 35140 35476
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 35084 35252 35140
rect 34972 34636 35028 34692
rect 34972 33628 35028 33684
rect 35420 34242 35476 34244
rect 35420 34190 35422 34242
rect 35422 34190 35474 34242
rect 35474 34190 35476 34242
rect 35420 34188 35476 34190
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 34636 30492 34692 30548
rect 34412 30044 34468 30100
rect 34412 28924 34468 28980
rect 34860 30716 34916 30772
rect 34972 31388 35028 31444
rect 34972 30940 35028 30996
rect 34860 30434 34916 30436
rect 34860 30382 34862 30434
rect 34862 30382 34914 30434
rect 34914 30382 34916 30434
rect 34860 30380 34916 30382
rect 34636 29986 34692 29988
rect 34636 29934 34638 29986
rect 34638 29934 34690 29986
rect 34690 29934 34692 29986
rect 34636 29932 34692 29934
rect 34524 29484 34580 29540
rect 34636 29426 34692 29428
rect 34636 29374 34638 29426
rect 34638 29374 34690 29426
rect 34690 29374 34692 29426
rect 34636 29372 34692 29374
rect 34860 29484 34916 29540
rect 34860 28812 34916 28868
rect 34412 28642 34468 28644
rect 34412 28590 34414 28642
rect 34414 28590 34466 28642
rect 34466 28590 34468 28642
rect 34412 28588 34468 28590
rect 35532 32562 35588 32564
rect 35532 32510 35534 32562
rect 35534 32510 35586 32562
rect 35586 32510 35588 32562
rect 35532 32508 35588 32510
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35532 31836 35588 31892
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35308 30098 35364 30100
rect 35308 30046 35310 30098
rect 35310 30046 35362 30098
rect 35362 30046 35364 30098
rect 35308 30044 35364 30046
rect 35532 29650 35588 29652
rect 35532 29598 35534 29650
rect 35534 29598 35586 29650
rect 35586 29598 35588 29650
rect 35532 29596 35588 29598
rect 35868 31052 35924 31108
rect 35756 30828 35812 30884
rect 36204 35420 36260 35476
rect 36092 33180 36148 33236
rect 36764 37996 36820 38052
rect 36428 37938 36484 37940
rect 36428 37886 36430 37938
rect 36430 37886 36482 37938
rect 36482 37886 36484 37938
rect 36428 37884 36484 37886
rect 37436 38556 37492 38612
rect 37212 37884 37268 37940
rect 37212 37154 37268 37156
rect 37212 37102 37214 37154
rect 37214 37102 37266 37154
rect 37266 37102 37268 37154
rect 37212 37100 37268 37102
rect 36988 36652 37044 36708
rect 36652 35586 36708 35588
rect 36652 35534 36654 35586
rect 36654 35534 36706 35586
rect 36706 35534 36708 35586
rect 36652 35532 36708 35534
rect 36540 34860 36596 34916
rect 37212 36876 37268 36932
rect 37212 35532 37268 35588
rect 37212 34914 37268 34916
rect 37212 34862 37214 34914
rect 37214 34862 37266 34914
rect 37266 34862 37268 34914
rect 37212 34860 37268 34862
rect 36540 33964 36596 34020
rect 36428 32396 36484 32452
rect 35756 30268 35812 30324
rect 36204 30210 36260 30212
rect 36204 30158 36206 30210
rect 36206 30158 36258 30210
rect 36258 30158 36260 30210
rect 36204 30156 36260 30158
rect 36428 30156 36484 30212
rect 36204 29708 36260 29764
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35420 28642 35476 28644
rect 35420 28590 35422 28642
rect 35422 28590 35474 28642
rect 35474 28590 35476 28642
rect 35420 28588 35476 28590
rect 34076 22204 34132 22260
rect 33852 17052 33908 17108
rect 35084 27858 35140 27860
rect 35084 27806 35086 27858
rect 35086 27806 35138 27858
rect 35138 27806 35140 27858
rect 35084 27804 35140 27806
rect 35420 27804 35476 27860
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 26796 35252 26852
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35980 28642 36036 28644
rect 35980 28590 35982 28642
rect 35982 28590 36034 28642
rect 36034 28590 36036 28642
rect 35980 28588 36036 28590
rect 35644 26796 35700 26852
rect 34300 23154 34356 23156
rect 34300 23102 34302 23154
rect 34302 23102 34354 23154
rect 34354 23102 34356 23154
rect 34300 23100 34356 23102
rect 33964 21756 34020 21812
rect 34076 19964 34132 20020
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35084 22370 35140 22372
rect 35084 22318 35086 22370
rect 35086 22318 35138 22370
rect 35138 22318 35140 22370
rect 35084 22316 35140 22318
rect 35196 21756 35252 21812
rect 35868 21644 35924 21700
rect 33964 17164 34020 17220
rect 33740 16716 33796 16772
rect 33516 16210 33572 16212
rect 33516 16158 33518 16210
rect 33518 16158 33570 16210
rect 33570 16158 33572 16210
rect 33516 16156 33572 16158
rect 34076 16156 34132 16212
rect 33964 16044 34020 16100
rect 34076 15538 34132 15540
rect 34076 15486 34078 15538
rect 34078 15486 34130 15538
rect 34130 15486 34132 15538
rect 34076 15484 34132 15486
rect 33068 15148 33124 15204
rect 32284 13020 32340 13076
rect 31612 12850 31668 12852
rect 31612 12798 31614 12850
rect 31614 12798 31666 12850
rect 31666 12798 31668 12850
rect 31612 12796 31668 12798
rect 32508 12796 32564 12852
rect 33068 13020 33124 13076
rect 30492 9826 30548 9828
rect 30492 9774 30494 9826
rect 30494 9774 30546 9826
rect 30546 9774 30548 9826
rect 30492 9772 30548 9774
rect 31388 9884 31444 9940
rect 29596 8092 29652 8148
rect 27916 6636 27972 6692
rect 27692 6130 27748 6132
rect 27692 6078 27694 6130
rect 27694 6078 27746 6130
rect 27746 6078 27748 6130
rect 27692 6076 27748 6078
rect 28140 5404 28196 5460
rect 28812 6076 28868 6132
rect 29596 5964 29652 6020
rect 27468 4172 27524 4228
rect 28140 4226 28196 4228
rect 28140 4174 28142 4226
rect 28142 4174 28194 4226
rect 28194 4174 28196 4226
rect 28140 4172 28196 4174
rect 30044 9548 30100 9604
rect 30380 6130 30436 6132
rect 30380 6078 30382 6130
rect 30382 6078 30434 6130
rect 30434 6078 30436 6130
rect 30380 6076 30436 6078
rect 30940 9602 30996 9604
rect 30940 9550 30942 9602
rect 30942 9550 30994 9602
rect 30994 9550 30996 9602
rect 30940 9548 30996 9550
rect 31724 9826 31780 9828
rect 31724 9774 31726 9826
rect 31726 9774 31778 9826
rect 31778 9774 31780 9826
rect 31724 9772 31780 9774
rect 31500 8988 31556 9044
rect 32060 9042 32116 9044
rect 32060 8990 32062 9042
rect 32062 8990 32114 9042
rect 32114 8990 32116 9042
rect 32060 8988 32116 8990
rect 31164 8146 31220 8148
rect 31164 8094 31166 8146
rect 31166 8094 31218 8146
rect 31218 8094 31220 8146
rect 31164 8092 31220 8094
rect 31612 8092 31668 8148
rect 32060 8204 32116 8260
rect 32732 8092 32788 8148
rect 30716 6018 30772 6020
rect 30716 5966 30718 6018
rect 30718 5966 30770 6018
rect 30770 5966 30772 6018
rect 30716 5964 30772 5966
rect 30940 6076 30996 6132
rect 33292 13746 33348 13748
rect 33292 13694 33294 13746
rect 33294 13694 33346 13746
rect 33346 13694 33348 13746
rect 33292 13692 33348 13694
rect 34076 13746 34132 13748
rect 34076 13694 34078 13746
rect 34078 13694 34130 13746
rect 34130 13694 34132 13746
rect 34076 13692 34132 13694
rect 33404 13074 33460 13076
rect 33404 13022 33406 13074
rect 33406 13022 33458 13074
rect 33458 13022 33460 13074
rect 33404 13020 33460 13022
rect 34076 13074 34132 13076
rect 34076 13022 34078 13074
rect 34078 13022 34130 13074
rect 34130 13022 34132 13074
rect 34076 13020 34132 13022
rect 34412 21308 34468 21364
rect 35084 21308 35140 21364
rect 34860 20076 34916 20132
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 36428 29372 36484 29428
rect 36764 30828 36820 30884
rect 36540 29932 36596 29988
rect 36092 21532 36148 21588
rect 36204 27804 36260 27860
rect 36428 27580 36484 27636
rect 36652 30044 36708 30100
rect 36652 28924 36708 28980
rect 37212 30268 37268 30324
rect 37100 29986 37156 29988
rect 37100 29934 37102 29986
rect 37102 29934 37154 29986
rect 37154 29934 37156 29986
rect 37100 29932 37156 29934
rect 36876 28642 36932 28644
rect 36876 28590 36878 28642
rect 36878 28590 36930 28642
rect 36930 28590 36932 28642
rect 36876 28588 36932 28590
rect 37100 28588 37156 28644
rect 36876 28082 36932 28084
rect 36876 28030 36878 28082
rect 36878 28030 36930 28082
rect 36930 28030 36932 28082
rect 36876 28028 36932 28030
rect 36988 27186 37044 27188
rect 36988 27134 36990 27186
rect 36990 27134 37042 27186
rect 37042 27134 37044 27186
rect 36988 27132 37044 27134
rect 37212 28418 37268 28420
rect 37212 28366 37214 28418
rect 37214 28366 37266 28418
rect 37266 28366 37268 28418
rect 37212 28364 37268 28366
rect 39452 51378 39508 51380
rect 39452 51326 39454 51378
rect 39454 51326 39506 51378
rect 39506 51326 39508 51378
rect 39452 51324 39508 51326
rect 38332 49026 38388 49028
rect 38332 48974 38334 49026
rect 38334 48974 38386 49026
rect 38386 48974 38388 49026
rect 38332 48972 38388 48974
rect 38668 50428 38724 50484
rect 38108 46396 38164 46452
rect 38556 47516 38612 47572
rect 38220 46060 38276 46116
rect 39116 47180 39172 47236
rect 39900 47180 39956 47236
rect 40348 51602 40404 51604
rect 40348 51550 40350 51602
rect 40350 51550 40402 51602
rect 40402 51550 40404 51602
rect 40348 51548 40404 51550
rect 40124 48972 40180 49028
rect 40348 47570 40404 47572
rect 40348 47518 40350 47570
rect 40350 47518 40402 47570
rect 40402 47518 40404 47570
rect 40348 47516 40404 47518
rect 39564 46732 39620 46788
rect 38780 46396 38836 46452
rect 38332 45948 38388 46004
rect 38220 45666 38276 45668
rect 38220 45614 38222 45666
rect 38222 45614 38274 45666
rect 38274 45614 38276 45666
rect 38220 45612 38276 45614
rect 38668 45388 38724 45444
rect 37996 44380 38052 44436
rect 38444 44380 38500 44436
rect 38332 43820 38388 43876
rect 38220 43650 38276 43652
rect 38220 43598 38222 43650
rect 38222 43598 38274 43650
rect 38274 43598 38276 43650
rect 38220 43596 38276 43598
rect 38220 42530 38276 42532
rect 38220 42478 38222 42530
rect 38222 42478 38274 42530
rect 38274 42478 38276 42530
rect 38220 42476 38276 42478
rect 38780 42028 38836 42084
rect 39452 45724 39508 45780
rect 39004 44492 39060 44548
rect 39340 44994 39396 44996
rect 39340 44942 39342 44994
rect 39342 44942 39394 44994
rect 39394 44942 39396 44994
rect 39340 44940 39396 44942
rect 39452 44210 39508 44212
rect 39452 44158 39454 44210
rect 39454 44158 39506 44210
rect 39506 44158 39508 44210
rect 39452 44156 39508 44158
rect 39116 43820 39172 43876
rect 38332 41186 38388 41188
rect 38332 41134 38334 41186
rect 38334 41134 38386 41186
rect 38386 41134 38388 41186
rect 38332 41132 38388 41134
rect 38556 40796 38612 40852
rect 38332 40460 38388 40516
rect 38332 39842 38388 39844
rect 38332 39790 38334 39842
rect 38334 39790 38386 39842
rect 38386 39790 38388 39842
rect 38332 39788 38388 39790
rect 38444 39116 38500 39172
rect 38444 38780 38500 38836
rect 38108 38556 38164 38612
rect 37996 38162 38052 38164
rect 37996 38110 37998 38162
rect 37998 38110 38050 38162
rect 38050 38110 38052 38162
rect 37996 38108 38052 38110
rect 37660 37266 37716 37268
rect 37660 37214 37662 37266
rect 37662 37214 37714 37266
rect 37714 37214 37716 37266
rect 37660 37212 37716 37214
rect 38108 37154 38164 37156
rect 38108 37102 38110 37154
rect 38110 37102 38162 37154
rect 38162 37102 38164 37154
rect 38108 37100 38164 37102
rect 38892 40572 38948 40628
rect 37996 36594 38052 36596
rect 37996 36542 37998 36594
rect 37998 36542 38050 36594
rect 38050 36542 38052 36594
rect 37996 36540 38052 36542
rect 38332 36428 38388 36484
rect 37772 36204 37828 36260
rect 37996 36316 38052 36372
rect 38108 36204 38164 36260
rect 38108 31724 38164 31780
rect 37660 31666 37716 31668
rect 37660 31614 37662 31666
rect 37662 31614 37714 31666
rect 37714 31614 37716 31666
rect 37660 31612 37716 31614
rect 38108 31388 38164 31444
rect 38220 31500 38276 31556
rect 37436 31106 37492 31108
rect 37436 31054 37438 31106
rect 37438 31054 37490 31106
rect 37490 31054 37492 31106
rect 37436 31052 37492 31054
rect 37548 28476 37604 28532
rect 37548 28028 37604 28084
rect 37436 27580 37492 27636
rect 38220 30268 38276 30324
rect 38108 29932 38164 29988
rect 37772 28364 37828 28420
rect 37660 27356 37716 27412
rect 36652 25228 36708 25284
rect 36428 24892 36484 24948
rect 37772 26684 37828 26740
rect 37660 26514 37716 26516
rect 37660 26462 37662 26514
rect 37662 26462 37714 26514
rect 37714 26462 37716 26514
rect 37660 26460 37716 26462
rect 37212 24946 37268 24948
rect 37212 24894 37214 24946
rect 37214 24894 37266 24946
rect 37266 24894 37268 24946
rect 37212 24892 37268 24894
rect 36652 22428 36708 22484
rect 37100 22370 37156 22372
rect 37100 22318 37102 22370
rect 37102 22318 37154 22370
rect 37154 22318 37156 22370
rect 37100 22316 37156 22318
rect 36204 21420 36260 21476
rect 36876 21308 36932 21364
rect 36540 20972 36596 21028
rect 35532 20130 35588 20132
rect 35532 20078 35534 20130
rect 35534 20078 35586 20130
rect 35586 20078 35588 20130
rect 35532 20076 35588 20078
rect 36204 20076 36260 20132
rect 35196 19964 35252 20020
rect 34412 16940 34468 16996
rect 34300 15148 34356 15204
rect 34972 16716 35028 16772
rect 34524 16268 34580 16324
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 37772 22482 37828 22484
rect 37772 22430 37774 22482
rect 37774 22430 37826 22482
rect 37826 22430 37828 22482
rect 37772 22428 37828 22430
rect 38668 31164 38724 31220
rect 38444 28364 38500 28420
rect 38892 39676 38948 39732
rect 38892 38780 38948 38836
rect 39452 40348 39508 40404
rect 39340 39676 39396 39732
rect 38892 33122 38948 33124
rect 38892 33070 38894 33122
rect 38894 33070 38946 33122
rect 38946 33070 38948 33122
rect 38892 33068 38948 33070
rect 38892 31666 38948 31668
rect 38892 31614 38894 31666
rect 38894 31614 38946 31666
rect 38946 31614 38948 31666
rect 38892 31612 38948 31614
rect 38892 29148 38948 29204
rect 38780 24892 38836 24948
rect 38556 24050 38612 24052
rect 38556 23998 38558 24050
rect 38558 23998 38610 24050
rect 38610 23998 38612 24050
rect 38556 23996 38612 23998
rect 38220 23436 38276 23492
rect 38220 22316 38276 22372
rect 38892 21644 38948 21700
rect 38332 21420 38388 21476
rect 38780 21474 38836 21476
rect 38780 21422 38782 21474
rect 38782 21422 38834 21474
rect 38834 21422 38836 21474
rect 38780 21420 38836 21422
rect 37660 20524 37716 20580
rect 37548 20076 37604 20132
rect 36652 18338 36708 18340
rect 36652 18286 36654 18338
rect 36654 18286 36706 18338
rect 36706 18286 36708 18338
rect 36652 18284 36708 18286
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35644 17164 35700 17220
rect 35196 17106 35252 17108
rect 35196 17054 35198 17106
rect 35198 17054 35250 17106
rect 35250 17054 35252 17106
rect 35196 17052 35252 17054
rect 36204 17164 36260 17220
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35196 16098 35252 16100
rect 35196 16046 35198 16098
rect 35198 16046 35250 16098
rect 35250 16046 35252 16098
rect 35196 16044 35252 16046
rect 34748 15484 34804 15540
rect 34412 14530 34468 14532
rect 34412 14478 34414 14530
rect 34414 14478 34466 14530
rect 34466 14478 34468 14530
rect 34412 14476 34468 14478
rect 33180 12178 33236 12180
rect 33180 12126 33182 12178
rect 33182 12126 33234 12178
rect 33234 12126 33236 12178
rect 33180 12124 33236 12126
rect 33404 12124 33460 12180
rect 33740 12178 33796 12180
rect 33740 12126 33742 12178
rect 33742 12126 33794 12178
rect 33794 12126 33796 12178
rect 33740 12124 33796 12126
rect 33404 9042 33460 9044
rect 33404 8990 33406 9042
rect 33406 8990 33458 9042
rect 33458 8990 33460 9042
rect 33404 8988 33460 8990
rect 33628 8988 33684 9044
rect 33516 8316 33572 8372
rect 33404 8092 33460 8148
rect 35756 17052 35812 17108
rect 35308 15314 35364 15316
rect 35308 15262 35310 15314
rect 35310 15262 35362 15314
rect 35362 15262 35364 15314
rect 35308 15260 35364 15262
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 36204 16268 36260 16324
rect 35756 14812 35812 14868
rect 34972 14642 35028 14644
rect 34972 14590 34974 14642
rect 34974 14590 35026 14642
rect 35026 14590 35028 14642
rect 34972 14588 35028 14590
rect 35420 14700 35476 14756
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35644 13132 35700 13188
rect 35980 15986 36036 15988
rect 35980 15934 35982 15986
rect 35982 15934 36034 15986
rect 36034 15934 36036 15986
rect 35980 15932 36036 15934
rect 37324 18508 37380 18564
rect 36652 17724 36708 17780
rect 36764 17164 36820 17220
rect 36540 16882 36596 16884
rect 36540 16830 36542 16882
rect 36542 16830 36594 16882
rect 36594 16830 36596 16882
rect 36540 16828 36596 16830
rect 36428 15820 36484 15876
rect 35980 15708 36036 15764
rect 36652 15932 36708 15988
rect 37660 16940 37716 16996
rect 38220 20914 38276 20916
rect 38220 20862 38222 20914
rect 38222 20862 38274 20914
rect 38274 20862 38276 20914
rect 38220 20860 38276 20862
rect 38220 20300 38276 20356
rect 37884 18508 37940 18564
rect 36540 14642 36596 14644
rect 36540 14590 36542 14642
rect 36542 14590 36594 14642
rect 36594 14590 36596 14642
rect 36540 14588 36596 14590
rect 37212 14812 37268 14868
rect 39452 39394 39508 39396
rect 39452 39342 39454 39394
rect 39454 39342 39506 39394
rect 39506 39342 39508 39394
rect 39452 39340 39508 39342
rect 39340 38946 39396 38948
rect 39340 38894 39342 38946
rect 39342 38894 39394 38946
rect 39394 38894 39396 38946
rect 39340 38892 39396 38894
rect 39228 38780 39284 38836
rect 39452 34300 39508 34356
rect 39228 33068 39284 33124
rect 39340 32450 39396 32452
rect 39340 32398 39342 32450
rect 39342 32398 39394 32450
rect 39394 32398 39396 32450
rect 39340 32396 39396 32398
rect 40348 45724 40404 45780
rect 40012 44940 40068 44996
rect 39900 44434 39956 44436
rect 39900 44382 39902 44434
rect 39902 44382 39954 44434
rect 39954 44382 39956 44434
rect 39900 44380 39956 44382
rect 40348 44492 40404 44548
rect 41020 55468 41076 55524
rect 41020 54460 41076 54516
rect 41244 55410 41300 55412
rect 41244 55358 41246 55410
rect 41246 55358 41298 55410
rect 41298 55358 41300 55410
rect 41244 55356 41300 55358
rect 41356 54684 41412 54740
rect 41356 54514 41412 54516
rect 41356 54462 41358 54514
rect 41358 54462 41410 54514
rect 41410 54462 41412 54514
rect 41356 54460 41412 54462
rect 42252 59778 42308 59780
rect 42252 59726 42254 59778
rect 42254 59726 42306 59778
rect 42306 59726 42308 59778
rect 42252 59724 42308 59726
rect 41916 57148 41972 57204
rect 42700 57148 42756 57204
rect 41580 54348 41636 54404
rect 41804 56082 41860 56084
rect 41804 56030 41806 56082
rect 41806 56030 41858 56082
rect 41858 56030 41860 56082
rect 41804 56028 41860 56030
rect 42476 56082 42532 56084
rect 42476 56030 42478 56082
rect 42478 56030 42530 56082
rect 42530 56030 42532 56082
rect 42476 56028 42532 56030
rect 41916 55020 41972 55076
rect 42364 55410 42420 55412
rect 42364 55358 42366 55410
rect 42366 55358 42418 55410
rect 42418 55358 42420 55410
rect 42364 55356 42420 55358
rect 42812 55410 42868 55412
rect 42812 55358 42814 55410
rect 42814 55358 42866 55410
rect 42866 55358 42868 55410
rect 42812 55356 42868 55358
rect 44156 55356 44212 55412
rect 42252 55074 42308 55076
rect 42252 55022 42254 55074
rect 42254 55022 42306 55074
rect 42306 55022 42308 55074
rect 42252 55020 42308 55022
rect 41020 52834 41076 52836
rect 41020 52782 41022 52834
rect 41022 52782 41074 52834
rect 41074 52782 41076 52834
rect 41020 52780 41076 52782
rect 41132 52220 41188 52276
rect 41356 52220 41412 52276
rect 42364 54460 42420 54516
rect 42140 53452 42196 53508
rect 42812 54348 42868 54404
rect 42812 53788 42868 53844
rect 42364 53170 42420 53172
rect 42364 53118 42366 53170
rect 42366 53118 42418 53170
rect 42418 53118 42420 53170
rect 42364 53116 42420 53118
rect 42140 52780 42196 52836
rect 42476 52386 42532 52388
rect 42476 52334 42478 52386
rect 42478 52334 42530 52386
rect 42530 52334 42532 52386
rect 42476 52332 42532 52334
rect 41468 51548 41524 51604
rect 42028 51324 42084 51380
rect 42364 52162 42420 52164
rect 42364 52110 42366 52162
rect 42366 52110 42418 52162
rect 42418 52110 42420 52162
rect 42364 52108 42420 52110
rect 42140 51548 42196 51604
rect 42252 51378 42308 51380
rect 42252 51326 42254 51378
rect 42254 51326 42306 51378
rect 42306 51326 42308 51378
rect 42252 51324 42308 51326
rect 41356 51100 41412 51156
rect 41356 50482 41412 50484
rect 41356 50430 41358 50482
rect 41358 50430 41410 50482
rect 41410 50430 41412 50482
rect 41356 50428 41412 50430
rect 41020 48636 41076 48692
rect 41244 48354 41300 48356
rect 41244 48302 41246 48354
rect 41246 48302 41298 48354
rect 41298 48302 41300 48354
rect 41244 48300 41300 48302
rect 41580 48242 41636 48244
rect 41580 48190 41582 48242
rect 41582 48190 41634 48242
rect 41634 48190 41636 48242
rect 41580 48188 41636 48190
rect 41356 47068 41412 47124
rect 41244 46898 41300 46900
rect 41244 46846 41246 46898
rect 41246 46846 41298 46898
rect 41298 46846 41300 46898
rect 41244 46844 41300 46846
rect 41132 45724 41188 45780
rect 42028 50764 42084 50820
rect 42028 50428 42084 50484
rect 41916 49698 41972 49700
rect 41916 49646 41918 49698
rect 41918 49646 41970 49698
rect 41970 49646 41972 49698
rect 41916 49644 41972 49646
rect 41244 45276 41300 45332
rect 41916 46732 41972 46788
rect 41244 44994 41300 44996
rect 41244 44942 41246 44994
rect 41246 44942 41298 44994
rect 41298 44942 41300 44994
rect 41244 44940 41300 44942
rect 41692 45276 41748 45332
rect 41244 44604 41300 44660
rect 40796 44210 40852 44212
rect 40796 44158 40798 44210
rect 40798 44158 40850 44210
rect 40850 44158 40852 44210
rect 40796 44156 40852 44158
rect 40908 44044 40964 44100
rect 40348 43820 40404 43876
rect 40124 43596 40180 43652
rect 40124 42140 40180 42196
rect 40236 41916 40292 41972
rect 39676 40572 39732 40628
rect 39788 41468 39844 41524
rect 39676 39004 39732 39060
rect 39788 38780 39844 38836
rect 40012 39564 40068 39620
rect 40236 41746 40292 41748
rect 40236 41694 40238 41746
rect 40238 41694 40290 41746
rect 40290 41694 40292 41746
rect 40236 41692 40292 41694
rect 40348 40236 40404 40292
rect 40348 40012 40404 40068
rect 40124 39228 40180 39284
rect 41020 43650 41076 43652
rect 41020 43598 41022 43650
rect 41022 43598 41074 43650
rect 41074 43598 41076 43650
rect 41020 43596 41076 43598
rect 41132 44492 41188 44548
rect 40684 40348 40740 40404
rect 40796 40572 40852 40628
rect 40908 40908 40964 40964
rect 41020 40684 41076 40740
rect 40796 39788 40852 39844
rect 40684 39228 40740 39284
rect 41244 44098 41300 44100
rect 41244 44046 41246 44098
rect 41246 44046 41298 44098
rect 41298 44046 41300 44098
rect 41244 44044 41300 44046
rect 41244 41804 41300 41860
rect 41244 40460 41300 40516
rect 41692 44492 41748 44548
rect 41916 45500 41972 45556
rect 42140 48300 42196 48356
rect 42252 47852 42308 47908
rect 43596 53788 43652 53844
rect 43148 53506 43204 53508
rect 43148 53454 43150 53506
rect 43150 53454 43202 53506
rect 43202 53454 43204 53506
rect 43148 53452 43204 53454
rect 43148 53116 43204 53172
rect 43372 52332 43428 52388
rect 42812 52108 42868 52164
rect 42476 48636 42532 48692
rect 42252 47180 42308 47236
rect 42364 47068 42420 47124
rect 42028 44380 42084 44436
rect 42364 45500 42420 45556
rect 42700 48188 42756 48244
rect 42700 47404 42756 47460
rect 42588 47292 42644 47348
rect 43148 49698 43204 49700
rect 43148 49646 43150 49698
rect 43150 49646 43202 49698
rect 43202 49646 43204 49698
rect 43148 49644 43204 49646
rect 42924 48636 42980 48692
rect 43260 47292 43316 47348
rect 42588 45612 42644 45668
rect 42700 45500 42756 45556
rect 42924 45612 42980 45668
rect 42476 45276 42532 45332
rect 42364 45164 42420 45220
rect 43148 45500 43204 45556
rect 42700 44940 42756 44996
rect 42588 44322 42644 44324
rect 42588 44270 42590 44322
rect 42590 44270 42642 44322
rect 42642 44270 42644 44322
rect 42588 44268 42644 44270
rect 41804 43762 41860 43764
rect 41804 43710 41806 43762
rect 41806 43710 41858 43762
rect 41858 43710 41860 43762
rect 41804 43708 41860 43710
rect 41468 41970 41524 41972
rect 41468 41918 41470 41970
rect 41470 41918 41522 41970
rect 41522 41918 41524 41970
rect 41468 41916 41524 41918
rect 41692 41692 41748 41748
rect 41692 40684 41748 40740
rect 41356 39900 41412 39956
rect 41468 40348 41524 40404
rect 41244 39788 41300 39844
rect 41132 39340 41188 39396
rect 41468 39004 41524 39060
rect 41468 38834 41524 38836
rect 41468 38782 41470 38834
rect 41470 38782 41522 38834
rect 41522 38782 41524 38834
rect 41468 38780 41524 38782
rect 41356 38556 41412 38612
rect 42252 41970 42308 41972
rect 42252 41918 42254 41970
rect 42254 41918 42306 41970
rect 42306 41918 42308 41970
rect 42252 41916 42308 41918
rect 42028 40012 42084 40068
rect 42140 40460 42196 40516
rect 42252 40348 42308 40404
rect 42588 39618 42644 39620
rect 42588 39566 42590 39618
rect 42590 39566 42642 39618
rect 42642 39566 42644 39618
rect 42588 39564 42644 39566
rect 42364 39340 42420 39396
rect 41916 39058 41972 39060
rect 41916 39006 41918 39058
rect 41918 39006 41970 39058
rect 41970 39006 41972 39058
rect 41916 39004 41972 39006
rect 41580 37490 41636 37492
rect 41580 37438 41582 37490
rect 41582 37438 41634 37490
rect 41634 37438 41636 37490
rect 41580 37436 41636 37438
rect 40908 37100 40964 37156
rect 41356 36594 41412 36596
rect 41356 36542 41358 36594
rect 41358 36542 41410 36594
rect 41410 36542 41412 36594
rect 41356 36540 41412 36542
rect 42924 44156 42980 44212
rect 43036 45276 43092 45332
rect 42812 41970 42868 41972
rect 42812 41918 42814 41970
rect 42814 41918 42866 41970
rect 42866 41918 42868 41970
rect 42812 41916 42868 41918
rect 42812 40684 42868 40740
rect 42140 38556 42196 38612
rect 42924 38332 42980 38388
rect 45164 52780 45220 52836
rect 45052 52274 45108 52276
rect 45052 52222 45054 52274
rect 45054 52222 45106 52274
rect 45106 52222 45108 52274
rect 45052 52220 45108 52222
rect 46060 52834 46116 52836
rect 46060 52782 46062 52834
rect 46062 52782 46114 52834
rect 46114 52782 46116 52834
rect 46060 52780 46116 52782
rect 43932 52162 43988 52164
rect 43932 52110 43934 52162
rect 43934 52110 43986 52162
rect 43986 52110 43988 52162
rect 43932 52108 43988 52110
rect 43708 51602 43764 51604
rect 43708 51550 43710 51602
rect 43710 51550 43762 51602
rect 43762 51550 43764 51602
rect 43708 51548 43764 51550
rect 44156 51602 44212 51604
rect 44156 51550 44158 51602
rect 44158 51550 44210 51602
rect 44210 51550 44212 51602
rect 44156 51548 44212 51550
rect 43820 47346 43876 47348
rect 43820 47294 43822 47346
rect 43822 47294 43874 47346
rect 43874 47294 43876 47346
rect 43820 47292 43876 47294
rect 43596 46786 43652 46788
rect 43596 46734 43598 46786
rect 43598 46734 43650 46786
rect 43650 46734 43652 46786
rect 43596 46732 43652 46734
rect 44156 46732 44212 46788
rect 43484 45276 43540 45332
rect 44044 45666 44100 45668
rect 44044 45614 44046 45666
rect 44046 45614 44098 45666
rect 44098 45614 44100 45666
rect 44044 45612 44100 45614
rect 43596 45500 43652 45556
rect 43372 45052 43428 45108
rect 43484 44604 43540 44660
rect 43372 44434 43428 44436
rect 43372 44382 43374 44434
rect 43374 44382 43426 44434
rect 43426 44382 43428 44434
rect 43372 44380 43428 44382
rect 43372 44156 43428 44212
rect 43372 41858 43428 41860
rect 43372 41806 43374 41858
rect 43374 41806 43426 41858
rect 43426 41806 43428 41858
rect 43372 41804 43428 41806
rect 43260 40290 43316 40292
rect 43260 40238 43262 40290
rect 43262 40238 43314 40290
rect 43314 40238 43316 40290
rect 43260 40236 43316 40238
rect 43148 38556 43204 38612
rect 42700 37826 42756 37828
rect 42700 37774 42702 37826
rect 42702 37774 42754 37826
rect 42754 37774 42756 37826
rect 42700 37772 42756 37774
rect 43148 37660 43204 37716
rect 44044 44322 44100 44324
rect 44044 44270 44046 44322
rect 44046 44270 44098 44322
rect 44098 44270 44100 44322
rect 44044 44268 44100 44270
rect 43596 43596 43652 43652
rect 44268 43650 44324 43652
rect 44268 43598 44270 43650
rect 44270 43598 44322 43650
rect 44322 43598 44324 43650
rect 44268 43596 44324 43598
rect 43596 40572 43652 40628
rect 43596 40402 43652 40404
rect 43596 40350 43598 40402
rect 43598 40350 43650 40402
rect 43650 40350 43652 40402
rect 43596 40348 43652 40350
rect 43484 38220 43540 38276
rect 43372 37826 43428 37828
rect 43372 37774 43374 37826
rect 43374 37774 43426 37826
rect 43426 37774 43428 37826
rect 43372 37772 43428 37774
rect 42364 36540 42420 36596
rect 40908 32396 40964 32452
rect 39452 29202 39508 29204
rect 39452 29150 39454 29202
rect 39454 29150 39506 29202
rect 39506 29150 39508 29202
rect 39452 29148 39508 29150
rect 40124 31500 40180 31556
rect 40572 31554 40628 31556
rect 40572 31502 40574 31554
rect 40574 31502 40626 31554
rect 40626 31502 40628 31554
rect 40572 31500 40628 31502
rect 40348 30210 40404 30212
rect 40348 30158 40350 30210
rect 40350 30158 40402 30210
rect 40402 30158 40404 30210
rect 40348 30156 40404 30158
rect 40796 31164 40852 31220
rect 40908 30828 40964 30884
rect 42028 35644 42084 35700
rect 43484 35644 43540 35700
rect 42700 34354 42756 34356
rect 42700 34302 42702 34354
rect 42702 34302 42754 34354
rect 42754 34302 42756 34354
rect 42700 34300 42756 34302
rect 42028 33068 42084 33124
rect 42476 32786 42532 32788
rect 42476 32734 42478 32786
rect 42478 32734 42530 32786
rect 42530 32734 42532 32786
rect 42476 32732 42532 32734
rect 43036 34300 43092 34356
rect 43036 33068 43092 33124
rect 43148 32732 43204 32788
rect 43036 32562 43092 32564
rect 43036 32510 43038 32562
rect 43038 32510 43090 32562
rect 43090 32510 43092 32562
rect 43036 32508 43092 32510
rect 44268 40908 44324 40964
rect 45948 46786 46004 46788
rect 45948 46734 45950 46786
rect 45950 46734 46002 46786
rect 46002 46734 46004 46786
rect 45948 46732 46004 46734
rect 44940 45500 44996 45556
rect 45164 45164 45220 45220
rect 44828 44268 44884 44324
rect 44604 41468 44660 41524
rect 45164 41468 45220 41524
rect 43820 38274 43876 38276
rect 43820 38222 43822 38274
rect 43822 38222 43874 38274
rect 43874 38222 43876 38274
rect 43820 38220 43876 38222
rect 44940 40962 44996 40964
rect 44940 40910 44942 40962
rect 44942 40910 44994 40962
rect 44994 40910 44996 40962
rect 44940 40908 44996 40910
rect 48076 45164 48132 45220
rect 44156 38556 44212 38612
rect 44044 37938 44100 37940
rect 44044 37886 44046 37938
rect 44046 37886 44098 37938
rect 44098 37886 44100 37938
rect 44044 37884 44100 37886
rect 44156 38332 44212 38388
rect 46396 39618 46452 39620
rect 46396 39566 46398 39618
rect 46398 39566 46450 39618
rect 46450 39566 46452 39618
rect 46396 39564 46452 39566
rect 45836 38556 45892 38612
rect 44268 36876 44324 36932
rect 44268 34300 44324 34356
rect 44268 33628 44324 33684
rect 43596 32060 43652 32116
rect 41356 31612 41412 31668
rect 41244 31164 41300 31220
rect 41804 31666 41860 31668
rect 41804 31614 41806 31666
rect 41806 31614 41858 31666
rect 41858 31614 41860 31666
rect 41804 31612 41860 31614
rect 41916 31500 41972 31556
rect 41692 30268 41748 30324
rect 41580 30210 41636 30212
rect 41580 30158 41582 30210
rect 41582 30158 41634 30210
rect 41634 30158 41636 30210
rect 41580 30156 41636 30158
rect 42028 31164 42084 31220
rect 41020 29314 41076 29316
rect 41020 29262 41022 29314
rect 41022 29262 41074 29314
rect 41074 29262 41076 29314
rect 41020 29260 41076 29262
rect 41020 28588 41076 28644
rect 39228 26796 39284 26852
rect 39116 26460 39172 26516
rect 39228 21810 39284 21812
rect 39228 21758 39230 21810
rect 39230 21758 39282 21810
rect 39282 21758 39284 21810
rect 39228 21756 39284 21758
rect 39228 21026 39284 21028
rect 39228 20974 39230 21026
rect 39230 20974 39282 21026
rect 39282 20974 39284 21026
rect 39228 20972 39284 20974
rect 38332 19010 38388 19012
rect 38332 18958 38334 19010
rect 38334 18958 38386 19010
rect 38386 18958 38388 19010
rect 38332 18956 38388 18958
rect 38332 18284 38388 18340
rect 38668 18956 38724 19012
rect 38668 17276 38724 17332
rect 38332 17164 38388 17220
rect 37996 16716 38052 16772
rect 37996 13692 38052 13748
rect 38108 16828 38164 16884
rect 36764 13132 36820 13188
rect 35868 13020 35924 13076
rect 35756 12572 35812 12628
rect 34524 11452 34580 11508
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35084 11506 35140 11508
rect 35084 11454 35086 11506
rect 35086 11454 35138 11506
rect 35138 11454 35140 11506
rect 35084 11452 35140 11454
rect 35308 11394 35364 11396
rect 35308 11342 35310 11394
rect 35310 11342 35362 11394
rect 35362 11342 35364 11394
rect 35308 11340 35364 11342
rect 36092 12572 36148 12628
rect 35756 11340 35812 11396
rect 35868 12460 35924 12516
rect 34636 10722 34692 10724
rect 34636 10670 34638 10722
rect 34638 10670 34690 10722
rect 34690 10670 34692 10722
rect 34636 10668 34692 10670
rect 34972 10668 35028 10724
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 34412 8370 34468 8372
rect 34412 8318 34414 8370
rect 34414 8318 34466 8370
rect 34466 8318 34468 8370
rect 34412 8316 34468 8318
rect 35756 8258 35812 8260
rect 35756 8206 35758 8258
rect 35758 8206 35810 8258
rect 35810 8206 35812 8258
rect 35756 8204 35812 8206
rect 35644 8092 35700 8148
rect 33068 5292 33124 5348
rect 33516 5292 33572 5348
rect 30156 4956 30212 5012
rect 25788 2828 25844 2884
rect 25340 2716 25396 2772
rect 26796 2770 26852 2772
rect 26796 2718 26798 2770
rect 26798 2718 26850 2770
rect 26850 2718 26852 2770
rect 26796 2716 26852 2718
rect 30940 4956 30996 5012
rect 32508 4450 32564 4452
rect 32508 4398 32510 4450
rect 32510 4398 32562 4450
rect 32562 4398 32564 4450
rect 32508 4396 32564 4398
rect 33628 4956 33684 5012
rect 33740 4508 33796 4564
rect 33852 4450 33908 4452
rect 33852 4398 33854 4450
rect 33854 4398 33906 4450
rect 33906 4398 33908 4450
rect 33852 4396 33908 4398
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 34076 5346 34132 5348
rect 34076 5294 34078 5346
rect 34078 5294 34130 5346
rect 34130 5294 34132 5346
rect 34076 5292 34132 5294
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 34972 5292 35028 5348
rect 35644 5346 35700 5348
rect 35644 5294 35646 5346
rect 35646 5294 35698 5346
rect 35698 5294 35700 5346
rect 35644 5292 35700 5294
rect 34300 5234 34356 5236
rect 34300 5182 34302 5234
rect 34302 5182 34354 5234
rect 34354 5182 34356 5234
rect 34300 5180 34356 5182
rect 34748 5234 34804 5236
rect 34748 5182 34750 5234
rect 34750 5182 34802 5234
rect 34802 5182 34804 5234
rect 34748 5180 34804 5182
rect 36316 8930 36372 8932
rect 36316 8878 36318 8930
rect 36318 8878 36370 8930
rect 36370 8878 36372 8930
rect 36316 8876 36372 8878
rect 37100 8876 37156 8932
rect 37324 9100 37380 9156
rect 35868 4956 35924 5012
rect 35980 8428 36036 8484
rect 35980 8092 36036 8148
rect 33964 4060 34020 4116
rect 33740 3778 33796 3780
rect 33740 3726 33742 3778
rect 33742 3726 33794 3778
rect 33794 3726 33796 3778
rect 33740 3724 33796 3726
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 34412 3724 34468 3780
rect 35980 4396 36036 4452
rect 37324 8428 37380 8484
rect 37548 8876 37604 8932
rect 36204 8092 36260 8148
rect 36316 8204 36372 8260
rect 36092 5180 36148 5236
rect 37324 8258 37380 8260
rect 37324 8206 37326 8258
rect 37326 8206 37378 8258
rect 37378 8206 37380 8258
rect 37324 8204 37380 8206
rect 36988 8146 37044 8148
rect 36988 8094 36990 8146
rect 36990 8094 37042 8146
rect 37042 8094 37044 8146
rect 36988 8092 37044 8094
rect 37212 6972 37268 7028
rect 35756 4172 35812 4228
rect 38332 16268 38388 16324
rect 38444 17052 38500 17108
rect 38892 20018 38948 20020
rect 38892 19966 38894 20018
rect 38894 19966 38946 20018
rect 38946 19966 38948 20018
rect 38892 19964 38948 19966
rect 39900 27804 39956 27860
rect 40348 27580 40404 27636
rect 41020 27858 41076 27860
rect 41020 27806 41022 27858
rect 41022 27806 41074 27858
rect 41074 27806 41076 27858
rect 41020 27804 41076 27806
rect 40460 26962 40516 26964
rect 40460 26910 40462 26962
rect 40462 26910 40514 26962
rect 40514 26910 40516 26962
rect 40460 26908 40516 26910
rect 39900 26796 39956 26852
rect 41244 29148 41300 29204
rect 41580 29148 41636 29204
rect 41356 28642 41412 28644
rect 41356 28590 41358 28642
rect 41358 28590 41410 28642
rect 41410 28590 41412 28642
rect 41356 28588 41412 28590
rect 42028 29596 42084 29652
rect 42252 30268 42308 30324
rect 42252 28700 42308 28756
rect 42364 29650 42420 29652
rect 42364 29598 42366 29650
rect 42366 29598 42418 29650
rect 42418 29598 42420 29650
rect 42364 29596 42420 29598
rect 41692 27580 41748 27636
rect 41132 26908 41188 26964
rect 41020 24892 41076 24948
rect 41468 24892 41524 24948
rect 40348 23548 40404 23604
rect 40908 23042 40964 23044
rect 40908 22990 40910 23042
rect 40910 22990 40962 23042
rect 40962 22990 40964 23042
rect 40908 22988 40964 22990
rect 41916 28252 41972 28308
rect 41916 24108 41972 24164
rect 43148 31164 43204 31220
rect 42812 29596 42868 29652
rect 43372 30882 43428 30884
rect 43372 30830 43374 30882
rect 43374 30830 43426 30882
rect 43426 30830 43428 30882
rect 43372 30828 43428 30830
rect 43148 30434 43204 30436
rect 43148 30382 43150 30434
rect 43150 30382 43202 30434
rect 43202 30382 43204 30434
rect 43148 30380 43204 30382
rect 42924 28754 42980 28756
rect 42924 28702 42926 28754
rect 42926 28702 42978 28754
rect 42978 28702 42980 28754
rect 42924 28700 42980 28702
rect 42700 27132 42756 27188
rect 43036 27692 43092 27748
rect 43372 27692 43428 27748
rect 44268 32508 44324 32564
rect 44268 31948 44324 32004
rect 45276 37100 45332 37156
rect 45612 37042 45668 37044
rect 45612 36990 45614 37042
rect 45614 36990 45666 37042
rect 45666 36990 45668 37042
rect 45612 36988 45668 36990
rect 48076 36594 48132 36596
rect 48076 36542 48078 36594
rect 48078 36542 48130 36594
rect 48130 36542 48132 36594
rect 48076 36540 48132 36542
rect 44828 33628 44884 33684
rect 44828 31948 44884 32004
rect 44380 30380 44436 30436
rect 45052 32060 45108 32116
rect 46284 32060 46340 32116
rect 46396 31836 46452 31892
rect 47740 31890 47796 31892
rect 47740 31838 47742 31890
rect 47742 31838 47794 31890
rect 47794 31838 47796 31890
rect 47740 31836 47796 31838
rect 45500 30994 45556 30996
rect 45500 30942 45502 30994
rect 45502 30942 45554 30994
rect 45554 30942 45556 30994
rect 45500 30940 45556 30942
rect 45052 30882 45108 30884
rect 45052 30830 45054 30882
rect 45054 30830 45106 30882
rect 45106 30830 45108 30882
rect 45052 30828 45108 30830
rect 46284 30994 46340 30996
rect 46284 30942 46286 30994
rect 46286 30942 46338 30994
rect 46338 30942 46340 30994
rect 46284 30940 46340 30942
rect 44268 28642 44324 28644
rect 44268 28590 44270 28642
rect 44270 28590 44322 28642
rect 44322 28590 44324 28642
rect 44268 28588 44324 28590
rect 44940 28642 44996 28644
rect 44940 28590 44942 28642
rect 44942 28590 44994 28642
rect 44994 28590 44996 28642
rect 44940 28588 44996 28590
rect 43820 28252 43876 28308
rect 43820 27746 43876 27748
rect 43820 27694 43822 27746
rect 43822 27694 43874 27746
rect 43874 27694 43876 27746
rect 43820 27692 43876 27694
rect 43596 27244 43652 27300
rect 45388 27244 45444 27300
rect 43372 27186 43428 27188
rect 43372 27134 43374 27186
rect 43374 27134 43426 27186
rect 43426 27134 43428 27186
rect 43372 27132 43428 27134
rect 43036 27020 43092 27076
rect 43596 27074 43652 27076
rect 43596 27022 43598 27074
rect 43598 27022 43650 27074
rect 43650 27022 43652 27074
rect 43596 27020 43652 27022
rect 44268 27020 44324 27076
rect 42812 24946 42868 24948
rect 42812 24894 42814 24946
rect 42814 24894 42866 24946
rect 42866 24894 42868 24946
rect 42812 24892 42868 24894
rect 43260 24892 43316 24948
rect 47180 26908 47236 26964
rect 44268 25116 44324 25172
rect 42588 24162 42644 24164
rect 42588 24110 42590 24162
rect 42590 24110 42642 24162
rect 42642 24110 42644 24162
rect 42588 24108 42644 24110
rect 42812 24050 42868 24052
rect 42812 23998 42814 24050
rect 42814 23998 42866 24050
rect 42866 23998 42868 24050
rect 42812 23996 42868 23998
rect 43932 24108 43988 24164
rect 43708 23884 43764 23940
rect 43708 23154 43764 23156
rect 43708 23102 43710 23154
rect 43710 23102 43762 23154
rect 43762 23102 43764 23154
rect 43708 23100 43764 23102
rect 42028 22988 42084 23044
rect 41916 21586 41972 21588
rect 41916 21534 41918 21586
rect 41918 21534 41970 21586
rect 41970 21534 41972 21586
rect 41916 21532 41972 21534
rect 42476 21586 42532 21588
rect 42476 21534 42478 21586
rect 42478 21534 42530 21586
rect 42530 21534 42532 21586
rect 42476 21532 42532 21534
rect 40012 21420 40068 21476
rect 39788 18284 39844 18340
rect 40124 20300 40180 20356
rect 38892 16882 38948 16884
rect 38892 16830 38894 16882
rect 38894 16830 38946 16882
rect 38946 16830 38948 16882
rect 38892 16828 38948 16830
rect 39340 17276 39396 17332
rect 39788 17052 39844 17108
rect 39564 16828 39620 16884
rect 38444 14812 38500 14868
rect 39004 14530 39060 14532
rect 39004 14478 39006 14530
rect 39006 14478 39058 14530
rect 39058 14478 39060 14530
rect 39004 14476 39060 14478
rect 39452 14530 39508 14532
rect 39452 14478 39454 14530
rect 39454 14478 39506 14530
rect 39506 14478 39508 14530
rect 39452 14476 39508 14478
rect 39788 16882 39844 16884
rect 39788 16830 39790 16882
rect 39790 16830 39842 16882
rect 39842 16830 39844 16882
rect 39788 16828 39844 16830
rect 39900 17666 39956 17668
rect 39900 17614 39902 17666
rect 39902 17614 39954 17666
rect 39954 17614 39956 17666
rect 39900 17612 39956 17614
rect 39788 16156 39844 16212
rect 39676 15932 39732 15988
rect 39788 15372 39844 15428
rect 40348 20300 40404 20356
rect 44268 23938 44324 23940
rect 44268 23886 44270 23938
rect 44270 23886 44322 23938
rect 44322 23886 44324 23938
rect 44268 23884 44324 23886
rect 45164 25116 45220 25172
rect 47740 24050 47796 24052
rect 47740 23998 47742 24050
rect 47742 23998 47794 24050
rect 47794 23998 47796 24050
rect 47740 23996 47796 23998
rect 43932 19292 43988 19348
rect 44604 19906 44660 19908
rect 44604 19854 44606 19906
rect 44606 19854 44658 19906
rect 44658 19854 44660 19906
rect 44604 19852 44660 19854
rect 44940 19292 44996 19348
rect 44492 18956 44548 19012
rect 41916 17836 41972 17892
rect 40908 17612 40964 17668
rect 40236 17052 40292 17108
rect 40460 16828 40516 16884
rect 40012 15426 40068 15428
rect 40012 15374 40014 15426
rect 40014 15374 40066 15426
rect 40066 15374 40068 15426
rect 40012 15372 40068 15374
rect 41468 17276 41524 17332
rect 41916 17106 41972 17108
rect 41916 17054 41918 17106
rect 41918 17054 41970 17106
rect 41970 17054 41972 17106
rect 41916 17052 41972 17054
rect 45388 19010 45444 19012
rect 45388 18958 45390 19010
rect 45390 18958 45442 19010
rect 45442 18958 45444 19010
rect 45388 18956 45444 18958
rect 45276 17890 45332 17892
rect 45276 17838 45278 17890
rect 45278 17838 45330 17890
rect 45330 17838 45332 17890
rect 45276 17836 45332 17838
rect 42028 16716 42084 16772
rect 41132 16268 41188 16324
rect 41468 16098 41524 16100
rect 41468 16046 41470 16098
rect 41470 16046 41522 16098
rect 41522 16046 41524 16098
rect 41468 16044 41524 16046
rect 39900 13746 39956 13748
rect 39900 13694 39902 13746
rect 39902 13694 39954 13746
rect 39954 13694 39956 13746
rect 39900 13692 39956 13694
rect 39452 11394 39508 11396
rect 39452 11342 39454 11394
rect 39454 11342 39506 11394
rect 39506 11342 39508 11394
rect 39452 11340 39508 11342
rect 38556 10668 38612 10724
rect 39116 10834 39172 10836
rect 39116 10782 39118 10834
rect 39118 10782 39170 10834
rect 39170 10782 39172 10834
rect 39116 10780 39172 10782
rect 38892 10722 38948 10724
rect 38892 10670 38894 10722
rect 38894 10670 38946 10722
rect 38946 10670 38948 10722
rect 38892 10668 38948 10670
rect 39788 10722 39844 10724
rect 39788 10670 39790 10722
rect 39790 10670 39842 10722
rect 39842 10670 39844 10722
rect 39788 10668 39844 10670
rect 41020 15426 41076 15428
rect 41020 15374 41022 15426
rect 41022 15374 41074 15426
rect 41074 15374 41076 15426
rect 41020 15372 41076 15374
rect 40236 14252 40292 14308
rect 40908 14476 40964 14532
rect 41580 15314 41636 15316
rect 41580 15262 41582 15314
rect 41582 15262 41634 15314
rect 41634 15262 41636 15314
rect 41580 15260 41636 15262
rect 43036 16770 43092 16772
rect 43036 16718 43038 16770
rect 43038 16718 43090 16770
rect 43090 16718 43092 16770
rect 43036 16716 43092 16718
rect 43484 16716 43540 16772
rect 43708 16322 43764 16324
rect 43708 16270 43710 16322
rect 43710 16270 43762 16322
rect 43762 16270 43764 16322
rect 43708 16268 43764 16270
rect 42028 15260 42084 15316
rect 41580 14476 41636 14532
rect 42924 14418 42980 14420
rect 42924 14366 42926 14418
rect 42926 14366 42978 14418
rect 42978 14366 42980 14418
rect 42924 14364 42980 14366
rect 43820 14364 43876 14420
rect 42812 14306 42868 14308
rect 42812 14254 42814 14306
rect 42814 14254 42866 14306
rect 42866 14254 42868 14306
rect 42812 14252 42868 14254
rect 40908 10834 40964 10836
rect 40908 10782 40910 10834
rect 40910 10782 40962 10834
rect 40962 10782 40964 10834
rect 40908 10780 40964 10782
rect 39564 9996 39620 10052
rect 40124 9884 40180 9940
rect 40572 9996 40628 10052
rect 43036 9938 43092 9940
rect 43036 9886 43038 9938
rect 43038 9886 43090 9938
rect 43090 9886 43092 9938
rect 43036 9884 43092 9886
rect 43708 9212 43764 9268
rect 41020 9154 41076 9156
rect 41020 9102 41022 9154
rect 41022 9102 41074 9154
rect 41074 9102 41076 9154
rect 41020 9100 41076 9102
rect 38108 6972 38164 7028
rect 38892 6972 38948 7028
rect 36988 4956 37044 5012
rect 36204 4396 36260 4452
rect 36764 4396 36820 4452
rect 36316 4060 36372 4116
rect 38444 4226 38500 4228
rect 38444 4174 38446 4226
rect 38446 4174 38498 4226
rect 38498 4174 38500 4226
rect 38444 4172 38500 4174
rect 39116 4338 39172 4340
rect 39116 4286 39118 4338
rect 39118 4286 39170 4338
rect 39170 4286 39172 4338
rect 39116 4284 39172 4286
rect 39788 4284 39844 4340
rect 35196 2378 35252 2380
rect 35196 2326 35198 2378
rect 35198 2326 35250 2378
rect 35250 2326 35252 2378
rect 35196 2324 35252 2326
rect 35300 2378 35356 2380
rect 35300 2326 35302 2378
rect 35302 2326 35354 2378
rect 35354 2326 35356 2378
rect 35300 2324 35356 2326
rect 35404 2378 35460 2380
rect 35404 2326 35406 2378
rect 35406 2326 35458 2378
rect 35458 2326 35460 2378
rect 35404 2324 35460 2326
rect 19836 1594 19892 1596
rect 19836 1542 19838 1594
rect 19838 1542 19890 1594
rect 19890 1542 19892 1594
rect 19836 1540 19892 1542
rect 19940 1594 19996 1596
rect 19940 1542 19942 1594
rect 19942 1542 19994 1594
rect 19994 1542 19996 1594
rect 19940 1540 19996 1542
rect 20044 1594 20100 1596
rect 20044 1542 20046 1594
rect 20046 1542 20098 1594
rect 20098 1542 20100 1594
rect 20044 1540 20100 1542
<< metal3 >>
rect 19826 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20110 78428
rect 4466 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4750 77644
rect 35186 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35470 77644
rect 30482 77196 30492 77252
rect 30548 77196 31276 77252
rect 31332 77196 31342 77252
rect 7522 76972 7532 77028
rect 7588 76972 8204 77028
rect 8260 76972 8876 77028
rect 8932 76972 10108 77028
rect 10164 76972 11228 77028
rect 11284 76972 11294 77028
rect 0 76916 400 76944
rect 0 76860 3388 76916
rect 3444 76860 3454 76916
rect 0 76832 400 76860
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 3042 76636 3052 76692
rect 3108 76636 3612 76692
rect 3668 76636 4284 76692
rect 4340 76636 4956 76692
rect 5012 76636 5022 76692
rect 10434 76412 10444 76468
rect 10500 76412 13020 76468
rect 13076 76412 13086 76468
rect 18498 76412 18508 76468
rect 18564 76412 21756 76468
rect 21812 76412 21822 76468
rect 21410 76300 21420 76356
rect 21476 76300 23548 76356
rect 23604 76300 23614 76356
rect 12562 76188 12572 76244
rect 12628 76188 13804 76244
rect 13860 76188 15148 76244
rect 15204 76188 15214 76244
rect 31266 76188 31276 76244
rect 31332 76188 33180 76244
rect 33236 76188 33964 76244
rect 34020 76188 34972 76244
rect 35028 76188 35038 76244
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 19282 75852 19292 75908
rect 19348 75852 21308 75908
rect 21364 75852 21374 75908
rect 24546 75740 24556 75796
rect 24612 75740 26796 75796
rect 26852 75740 26862 75796
rect 28130 75740 28140 75796
rect 28196 75740 29372 75796
rect 29428 75740 30156 75796
rect 30212 75740 30940 75796
rect 30996 75740 31006 75796
rect 3266 75628 3276 75684
rect 3332 75628 4396 75684
rect 4452 75628 4462 75684
rect 20738 75628 20748 75684
rect 20804 75628 21644 75684
rect 21700 75628 22428 75684
rect 22484 75628 22494 75684
rect 24210 75628 24220 75684
rect 24276 75628 25228 75684
rect 25284 75628 25294 75684
rect 29922 75628 29932 75684
rect 29988 75628 30828 75684
rect 30884 75628 30894 75684
rect 32050 75628 32060 75684
rect 32116 75628 33684 75684
rect 33628 75572 33684 75628
rect 33618 75516 33628 75572
rect 33684 75516 33694 75572
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 4274 75068 4284 75124
rect 4340 75068 4956 75124
rect 5012 75068 5740 75124
rect 5796 75068 5806 75124
rect 33618 74956 33628 75012
rect 33684 74956 35196 75012
rect 35252 74956 36988 75012
rect 37044 74956 37054 75012
rect 24098 74844 24108 74900
rect 24164 74844 25228 74900
rect 25284 74844 25900 74900
rect 25956 74844 29820 74900
rect 29876 74844 29886 74900
rect 32498 74732 32508 74788
rect 32564 74732 33404 74788
rect 33460 74732 34188 74788
rect 34244 74732 34524 74788
rect 34580 74732 34590 74788
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 9650 73948 9660 74004
rect 9716 73948 10668 74004
rect 10724 73948 12292 74004
rect 30370 73948 30380 74004
rect 30436 73948 33404 74004
rect 33460 73948 33470 74004
rect 34290 73948 34300 74004
rect 34356 73948 35308 74004
rect 35364 73948 35980 74004
rect 36036 73948 37436 74004
rect 37492 73948 37502 74004
rect 12236 73892 12292 73948
rect 12226 73836 12236 73892
rect 12292 73836 12302 73892
rect 35634 73836 35644 73892
rect 35700 73836 36316 73892
rect 36372 73836 36382 73892
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 24210 73164 24220 73220
rect 24276 73164 25228 73220
rect 25284 73164 25564 73220
rect 25620 73164 25630 73220
rect 26674 73164 26684 73220
rect 26740 73164 30044 73220
rect 30100 73164 30110 73220
rect 13010 73052 13020 73108
rect 13076 73052 14252 73108
rect 14308 73052 14318 73108
rect 19170 73052 19180 73108
rect 19236 73052 20636 73108
rect 20692 73052 20702 73108
rect 34962 73052 34972 73108
rect 35028 73052 35644 73108
rect 35700 73052 35710 73108
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 30818 72492 30828 72548
rect 30884 72492 33852 72548
rect 33908 72492 33918 72548
rect 3154 72380 3164 72436
rect 3220 72380 4060 72436
rect 4116 72380 4126 72436
rect 29260 72380 31948 72436
rect 32004 72380 32014 72436
rect 29260 72324 29316 72380
rect 27346 72268 27356 72324
rect 27412 72268 29260 72324
rect 29316 72268 29326 72324
rect 30258 72268 30268 72324
rect 30324 72268 32956 72324
rect 33012 72268 33022 72324
rect 2930 72156 2940 72212
rect 2996 72156 3500 72212
rect 3556 72156 4004 72212
rect 0 71988 400 72016
rect 3948 71988 4004 72156
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 0 71932 3724 71988
rect 3780 71932 3790 71988
rect 3938 71932 3948 71988
rect 4004 71932 5068 71988
rect 5124 71932 5134 71988
rect 31490 71932 31500 71988
rect 31556 71932 33180 71988
rect 33236 71932 33246 71988
rect 0 71904 400 71932
rect 35980 71820 37100 71876
rect 37156 71820 37166 71876
rect 35980 71764 36036 71820
rect 32834 71708 32844 71764
rect 32900 71708 34412 71764
rect 34468 71708 34748 71764
rect 34804 71708 35980 71764
rect 36036 71708 36046 71764
rect 36418 71708 36428 71764
rect 36484 71708 37548 71764
rect 37604 71708 38332 71764
rect 38388 71708 38398 71764
rect 17714 71596 17724 71652
rect 17780 71596 20300 71652
rect 20356 71596 20366 71652
rect 23650 71596 23660 71652
rect 23716 71596 24556 71652
rect 24612 71596 24622 71652
rect 26114 71596 26124 71652
rect 26180 71596 32508 71652
rect 32564 71596 33068 71652
rect 33124 71596 33134 71652
rect 33394 71596 33404 71652
rect 33460 71596 36540 71652
rect 36596 71596 38780 71652
rect 38836 71596 38846 71652
rect 33068 71428 33124 71596
rect 33964 71484 37212 71540
rect 37268 71484 37278 71540
rect 33964 71428 34020 71484
rect 33068 71372 33964 71428
rect 34020 71372 34030 71428
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 19170 71148 19180 71204
rect 19236 71148 20748 71204
rect 20804 71148 21644 71204
rect 21700 71148 26348 71204
rect 26404 71148 26414 71204
rect 1810 70924 1820 70980
rect 1876 70924 2380 70980
rect 2436 70924 2716 70980
rect 2772 70924 4172 70980
rect 4228 70924 4238 70980
rect 3602 70812 3612 70868
rect 3668 70812 4060 70868
rect 4116 70812 5628 70868
rect 5684 70812 5694 70868
rect 16818 70588 16828 70644
rect 16884 70588 17724 70644
rect 17780 70588 17790 70644
rect 20850 70588 20860 70644
rect 20916 70588 22428 70644
rect 22484 70588 22876 70644
rect 22932 70588 24108 70644
rect 24164 70588 24174 70644
rect 35074 70588 35084 70644
rect 35140 70588 36988 70644
rect 37044 70588 37996 70644
rect 38052 70588 38062 70644
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 26852 70308 26908 70532
rect 26964 70476 26974 70532
rect 25330 70252 25340 70308
rect 25396 70252 26012 70308
rect 26068 70252 26908 70308
rect 34626 70252 34636 70308
rect 34692 70252 35644 70308
rect 35700 70252 35710 70308
rect 6626 70140 6636 70196
rect 6692 70140 7532 70196
rect 7588 70140 7598 70196
rect 9874 70140 9884 70196
rect 9940 70140 10668 70196
rect 10724 70140 12348 70196
rect 12404 70140 12414 70196
rect 13346 70140 13356 70196
rect 13412 70140 14700 70196
rect 14756 70140 14766 70196
rect 25778 70140 25788 70196
rect 25844 70140 28028 70196
rect 28084 70140 28094 70196
rect 29026 70140 29036 70196
rect 29092 70140 29484 70196
rect 29540 70140 29932 70196
rect 29988 70140 31164 70196
rect 31220 70140 31230 70196
rect 33618 70140 33628 70196
rect 33684 70140 35084 70196
rect 35140 70140 35150 70196
rect 23986 70028 23996 70084
rect 24052 70028 26908 70084
rect 26964 70028 28364 70084
rect 28420 70028 28430 70084
rect 29698 70028 29708 70084
rect 29764 70028 31612 70084
rect 31668 70028 31678 70084
rect 34738 70028 34748 70084
rect 34804 70028 35868 70084
rect 35924 70028 35934 70084
rect 29250 69916 29260 69972
rect 29316 69916 30716 69972
rect 30772 69916 30782 69972
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 3826 69468 3836 69524
rect 3892 69468 4284 69524
rect 4340 69468 4620 69524
rect 4676 69468 5740 69524
rect 5796 69468 6188 69524
rect 6244 69468 6254 69524
rect 21522 69356 21532 69412
rect 21588 69356 22540 69412
rect 22596 69356 22606 69412
rect 33842 69356 33852 69412
rect 33908 69356 35868 69412
rect 35924 69356 37100 69412
rect 37156 69356 37166 69412
rect 18498 69244 18508 69300
rect 18564 69244 19068 69300
rect 19124 69244 23660 69300
rect 23716 69244 23726 69300
rect 10322 69132 10332 69188
rect 10388 69132 10780 69188
rect 10836 69132 11452 69188
rect 11508 69132 11900 69188
rect 11956 69132 11966 69188
rect 29586 69132 29596 69188
rect 29652 69132 30828 69188
rect 30884 69132 32396 69188
rect 32452 69132 32956 69188
rect 33012 69132 33628 69188
rect 33684 69132 33694 69188
rect 36082 69020 36092 69076
rect 36148 69020 36988 69076
rect 37044 69020 37054 69076
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 36194 68908 36204 68964
rect 36260 68908 37100 68964
rect 37156 68908 37166 68964
rect 18946 68796 18956 68852
rect 19012 68796 19740 68852
rect 19796 68796 19806 68852
rect 21970 68796 21980 68852
rect 22036 68796 23324 68852
rect 23380 68796 23772 68852
rect 23828 68796 25788 68852
rect 25844 68796 25854 68852
rect 22418 68684 22428 68740
rect 22484 68684 23548 68740
rect 23604 68684 24668 68740
rect 24724 68684 25340 68740
rect 25396 68684 25406 68740
rect 20850 68572 20860 68628
rect 20916 68572 21868 68628
rect 21924 68572 23100 68628
rect 23156 68572 23996 68628
rect 24052 68572 24220 68628
rect 24276 68572 24286 68628
rect 24098 68460 24108 68516
rect 24164 68460 25004 68516
rect 25060 68460 26908 68516
rect 26964 68460 27356 68516
rect 27412 68460 27422 68516
rect 21858 68348 21868 68404
rect 21924 68348 22988 68404
rect 23044 68348 23054 68404
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 4946 68012 4956 68068
rect 5012 68012 5740 68068
rect 5796 68012 5806 68068
rect 10322 68012 10332 68068
rect 10388 68012 10780 68068
rect 10836 68012 10846 68068
rect 19506 68012 19516 68068
rect 19572 68012 20300 68068
rect 20356 68012 21420 68068
rect 21476 68012 21486 68068
rect 8306 67900 8316 67956
rect 8372 67900 9436 67956
rect 9492 67900 9502 67956
rect 2930 67788 2940 67844
rect 2996 67788 3500 67844
rect 3556 67788 3566 67844
rect 6066 67788 6076 67844
rect 6132 67788 7644 67844
rect 7700 67788 7710 67844
rect 22418 67564 22428 67620
rect 22484 67564 22652 67620
rect 22708 67564 22876 67620
rect 22932 67564 22942 67620
rect 27346 67564 27356 67620
rect 27412 67564 31500 67620
rect 31556 67564 31566 67620
rect 2594 67452 2604 67508
rect 2660 67452 2940 67508
rect 2996 67452 3006 67508
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 6402 67228 6412 67284
rect 6468 67228 7196 67284
rect 7252 67228 7262 67284
rect 3154 67116 3164 67172
rect 3220 67116 3612 67172
rect 3668 67116 3678 67172
rect 0 67060 400 67088
rect 0 67004 532 67060
rect 2482 67004 2492 67060
rect 2548 67004 3052 67060
rect 3108 67004 3118 67060
rect 0 66976 400 67004
rect 476 66836 532 67004
rect 6748 66948 6804 67228
rect 8754 67004 8764 67060
rect 8820 67004 10668 67060
rect 10724 67004 11676 67060
rect 11732 67004 11742 67060
rect 18274 67004 18284 67060
rect 18340 67004 27468 67060
rect 27524 67004 27534 67060
rect 33730 67004 33740 67060
rect 33796 67004 34748 67060
rect 34804 67004 35308 67060
rect 35364 67004 35374 67060
rect 2930 66892 2940 66948
rect 2996 66892 4844 66948
rect 4900 66892 5516 66948
rect 5572 66892 6076 66948
rect 6132 66892 6142 66948
rect 6738 66892 6748 66948
rect 6804 66892 6814 66948
rect 33954 66892 33964 66948
rect 34020 66892 34188 66948
rect 34244 66892 38332 66948
rect 38388 66892 38398 66948
rect 252 66780 532 66836
rect 6962 66780 6972 66836
rect 7028 66780 7532 66836
rect 7588 66780 7598 66836
rect 32610 66780 32620 66836
rect 32676 66780 33292 66836
rect 33348 66780 33358 66836
rect 252 66052 308 66780
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 39218 66332 39228 66388
rect 39284 66332 39900 66388
rect 39956 66332 39966 66388
rect 6850 66220 6860 66276
rect 6916 66220 7308 66276
rect 7364 66220 7644 66276
rect 7700 66220 7710 66276
rect 36418 66108 36428 66164
rect 36484 66108 37772 66164
rect 37828 66108 37838 66164
rect 252 65996 3388 66052
rect 3714 65996 3724 66052
rect 3780 65996 4172 66052
rect 4228 65996 4238 66052
rect 9650 65996 9660 66052
rect 9716 65996 10220 66052
rect 10276 65996 10780 66052
rect 10836 65996 11340 66052
rect 11396 65996 11406 66052
rect 21410 65996 21420 66052
rect 21476 65996 22316 66052
rect 22372 65996 22382 66052
rect 35746 65996 35756 66052
rect 35812 65996 36988 66052
rect 37044 65996 37054 66052
rect 3332 65828 3388 65996
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 3332 65772 3500 65828
rect 3556 65772 3566 65828
rect 6412 65436 6748 65492
rect 6804 65436 7756 65492
rect 7812 65436 7822 65492
rect 9426 65436 9436 65492
rect 9492 65436 10780 65492
rect 10836 65436 12460 65492
rect 12516 65436 13020 65492
rect 13076 65436 13086 65492
rect 27794 65436 27804 65492
rect 27860 65436 30604 65492
rect 30660 65436 32060 65492
rect 32116 65436 32620 65492
rect 32676 65436 32686 65492
rect 33058 65436 33068 65492
rect 33124 65436 34188 65492
rect 34244 65436 34254 65492
rect 6412 65380 6468 65436
rect 3602 65324 3612 65380
rect 3668 65324 3948 65380
rect 4004 65324 6468 65380
rect 6626 65324 6636 65380
rect 6692 65324 8204 65380
rect 8260 65324 8988 65380
rect 9044 65324 9548 65380
rect 9604 65324 9614 65380
rect 11106 65324 11116 65380
rect 11172 65324 12124 65380
rect 12180 65324 12190 65380
rect 18722 65324 18732 65380
rect 18788 65324 21420 65380
rect 21476 65324 21486 65380
rect 32620 65268 32676 65436
rect 38994 65324 39004 65380
rect 39060 65324 39676 65380
rect 39732 65324 39742 65380
rect 25778 65212 25788 65268
rect 25844 65212 26572 65268
rect 26628 65212 26638 65268
rect 32620 65212 33516 65268
rect 33572 65212 33582 65268
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 25330 64988 25340 65044
rect 25396 64988 25676 65044
rect 25732 64988 28588 65044
rect 28644 64988 28654 65044
rect 36194 64876 36204 64932
rect 36260 64876 36988 64932
rect 37044 64876 37054 64932
rect 10098 64652 10108 64708
rect 10164 64652 10780 64708
rect 10836 64652 11116 64708
rect 11172 64652 11182 64708
rect 23538 64540 23548 64596
rect 23604 64540 24220 64596
rect 24276 64540 24286 64596
rect 10658 64428 10668 64484
rect 10724 64428 11452 64484
rect 11508 64428 12012 64484
rect 12068 64428 12078 64484
rect 22418 64428 22428 64484
rect 22484 64428 22876 64484
rect 22932 64428 23324 64484
rect 23380 64428 24108 64484
rect 24164 64428 24174 64484
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 21970 64092 21980 64148
rect 22036 64092 22428 64148
rect 22484 64092 22494 64148
rect 30594 64092 30604 64148
rect 30660 64092 31276 64148
rect 31332 64092 31342 64148
rect 32834 64092 32844 64148
rect 32900 64092 35644 64148
rect 35700 64092 35980 64148
rect 36036 64092 36046 64148
rect 22866 63980 22876 64036
rect 22932 63980 25676 64036
rect 25732 63980 25742 64036
rect 31938 63980 31948 64036
rect 32004 63980 32956 64036
rect 33012 63980 34524 64036
rect 34580 63980 35196 64036
rect 35252 63980 35262 64036
rect 12114 63868 12124 63924
rect 12180 63868 14476 63924
rect 14532 63868 14542 63924
rect 21522 63868 21532 63924
rect 21588 63868 22092 63924
rect 22148 63868 22764 63924
rect 22820 63868 22830 63924
rect 24098 63868 24108 63924
rect 24164 63868 25340 63924
rect 25396 63868 25406 63924
rect 28242 63868 28252 63924
rect 28308 63868 28700 63924
rect 28756 63868 28766 63924
rect 31490 63868 31500 63924
rect 31556 63868 35308 63924
rect 35364 63868 35756 63924
rect 35812 63868 35822 63924
rect 11442 63644 11452 63700
rect 11508 63644 11788 63700
rect 11844 63644 11854 63700
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 3042 63196 3052 63252
rect 3108 63196 4508 63252
rect 4564 63196 5292 63252
rect 5348 63196 6076 63252
rect 6132 63196 6412 63252
rect 6468 63196 7420 63252
rect 7476 63196 7486 63252
rect 16370 63196 16380 63252
rect 16436 63196 18956 63252
rect 19012 63196 19022 63252
rect 30594 63196 30604 63252
rect 30660 63196 32396 63252
rect 32452 63196 32462 63252
rect 33170 63196 33180 63252
rect 33236 63196 34076 63252
rect 34132 63196 36428 63252
rect 36484 63196 37996 63252
rect 38052 63196 38444 63252
rect 38500 63196 38510 63252
rect 38612 63196 39228 63252
rect 39284 63196 39294 63252
rect 38612 63140 38668 63196
rect 15586 63084 15596 63140
rect 15652 63084 16828 63140
rect 16884 63084 19628 63140
rect 19684 63084 20188 63140
rect 37314 63084 37324 63140
rect 37380 63084 38668 63140
rect 2706 62972 2716 63028
rect 2772 62972 3724 63028
rect 3780 62972 3790 63028
rect 20132 62916 20188 63084
rect 33170 62972 33180 63028
rect 33236 62972 35644 63028
rect 35700 62972 36316 63028
rect 36372 62972 36382 63028
rect 20132 62860 20412 62916
rect 20468 62860 20748 62916
rect 20804 62860 20814 62916
rect 34822 62860 34860 62916
rect 34916 62860 34926 62916
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 7410 62524 7420 62580
rect 7476 62524 8652 62580
rect 8708 62524 9436 62580
rect 9492 62524 9502 62580
rect 17714 62412 17724 62468
rect 17780 62412 18508 62468
rect 18564 62412 18956 62468
rect 19012 62412 19022 62468
rect 19618 62412 19628 62468
rect 19684 62412 20300 62468
rect 20356 62412 20366 62468
rect 22306 62412 22316 62468
rect 22372 62412 23324 62468
rect 23380 62412 23660 62468
rect 23716 62412 23726 62468
rect 28354 62300 28364 62356
rect 28420 62300 29372 62356
rect 29428 62300 31724 62356
rect 31780 62300 32508 62356
rect 32564 62300 32574 62356
rect 17938 62188 17948 62244
rect 18004 62188 18508 62244
rect 18564 62188 18574 62244
rect 35308 62188 36092 62244
rect 36148 62188 37324 62244
rect 37380 62188 37390 62244
rect 0 62132 400 62160
rect 35308 62132 35364 62188
rect 0 62076 4116 62132
rect 4722 62076 4732 62132
rect 4788 62076 5852 62132
rect 5908 62076 5918 62132
rect 32946 62076 32956 62132
rect 33012 62076 33628 62132
rect 33684 62076 35364 62132
rect 0 62048 400 62076
rect 4060 61908 4116 62076
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 4050 61852 4060 61908
rect 4116 61852 4126 61908
rect 3938 61740 3948 61796
rect 4004 61740 4620 61796
rect 4676 61740 4686 61796
rect 7634 61516 7644 61572
rect 7700 61516 8316 61572
rect 8372 61516 9436 61572
rect 9492 61516 9502 61572
rect 40114 61516 40124 61572
rect 40180 61516 40796 61572
rect 40852 61516 40862 61572
rect 4274 61404 4284 61460
rect 4340 61404 5628 61460
rect 5684 61404 5694 61460
rect 8866 61404 8876 61460
rect 8932 61404 9548 61460
rect 9604 61404 10780 61460
rect 10836 61404 10846 61460
rect 18610 61404 18620 61460
rect 18676 61404 19516 61460
rect 19572 61404 19582 61460
rect 37538 61404 37548 61460
rect 37604 61404 38444 61460
rect 38500 61404 38510 61460
rect 20962 61292 20972 61348
rect 21028 61292 22652 61348
rect 22708 61292 22988 61348
rect 23044 61292 25004 61348
rect 25060 61292 25070 61348
rect 26338 61292 26348 61348
rect 26404 61292 26908 61348
rect 26964 61292 26974 61348
rect 24770 61180 24780 61236
rect 24836 61180 25900 61236
rect 25956 61180 25966 61236
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 20402 60956 20412 61012
rect 20468 60956 20636 61012
rect 20692 60956 20702 61012
rect 24546 60956 24556 61012
rect 24612 60956 26348 61012
rect 26404 60956 26414 61012
rect 7634 60732 7644 60788
rect 7700 60732 8764 60788
rect 8820 60732 8830 60788
rect 3266 60620 3276 60676
rect 3332 60620 3724 60676
rect 3780 60620 3790 60676
rect 4162 60620 4172 60676
rect 4228 60620 4620 60676
rect 4676 60620 5068 60676
rect 5124 60620 5134 60676
rect 8642 60620 8652 60676
rect 8708 60620 10668 60676
rect 10724 60620 11676 60676
rect 11732 60620 11742 60676
rect 24658 60620 24668 60676
rect 24724 60620 26012 60676
rect 26068 60620 26078 60676
rect 42802 60620 42812 60676
rect 42868 60620 43820 60676
rect 43876 60620 43886 60676
rect 4946 60508 4956 60564
rect 5012 60508 5852 60564
rect 5908 60508 5918 60564
rect 15586 60396 15596 60452
rect 15652 60396 17500 60452
rect 17556 60396 18284 60452
rect 18340 60396 18350 60452
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 24882 60060 24892 60116
rect 24948 60060 26012 60116
rect 26068 60060 26078 60116
rect 30706 60060 30716 60116
rect 30772 60060 31276 60116
rect 31332 60060 31342 60116
rect 19730 59948 19740 60004
rect 19796 59948 21420 60004
rect 21476 59948 24332 60004
rect 24388 59948 25004 60004
rect 25060 59948 25070 60004
rect 6290 59836 6300 59892
rect 6356 59836 7532 59892
rect 7588 59836 7598 59892
rect 15698 59836 15708 59892
rect 15764 59836 18060 59892
rect 18116 59836 18126 59892
rect 27010 59836 27020 59892
rect 27076 59836 28140 59892
rect 28196 59836 28206 59892
rect 21746 59724 21756 59780
rect 21812 59724 22876 59780
rect 22932 59724 22942 59780
rect 26338 59724 26348 59780
rect 26404 59724 26796 59780
rect 26852 59724 26862 59780
rect 30930 59724 30940 59780
rect 30996 59724 31836 59780
rect 31892 59724 32732 59780
rect 32788 59724 33180 59780
rect 33236 59724 34636 59780
rect 34692 59724 34702 59780
rect 39666 59724 39676 59780
rect 39732 59724 40572 59780
rect 40628 59724 40638 59780
rect 41458 59724 41468 59780
rect 41524 59724 42252 59780
rect 42308 59724 42318 59780
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 18498 59500 18508 59556
rect 18564 59500 19516 59556
rect 19572 59500 19582 59556
rect 21634 59388 21644 59444
rect 21700 59388 22316 59444
rect 22372 59388 23212 59444
rect 23268 59388 23278 59444
rect 12002 59276 12012 59332
rect 12068 59276 14252 59332
rect 14308 59276 14812 59332
rect 14868 59276 14878 59332
rect 16258 59276 16268 59332
rect 16324 59276 17388 59332
rect 17444 59276 17454 59332
rect 10658 59164 10668 59220
rect 10724 59164 12124 59220
rect 12180 59164 12796 59220
rect 12852 59164 13244 59220
rect 13300 59164 13310 59220
rect 18386 59164 18396 59220
rect 18452 59164 29148 59220
rect 29204 59164 29214 59220
rect 15026 59052 15036 59108
rect 15092 59052 15596 59108
rect 15652 59052 15662 59108
rect 18274 59052 18284 59108
rect 18340 59052 18844 59108
rect 18900 59052 18910 59108
rect 19282 59052 19292 59108
rect 19348 59052 19628 59108
rect 19684 59052 21980 59108
rect 22036 59052 22046 59108
rect 22614 59052 22652 59108
rect 22708 59052 22718 59108
rect 5730 58940 5740 58996
rect 5796 58940 6300 58996
rect 6356 58940 6366 58996
rect 3490 58828 3500 58884
rect 3556 58828 3948 58884
rect 4004 58828 4014 58884
rect 22194 58828 22204 58884
rect 22260 58828 24332 58884
rect 24388 58828 24398 58884
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 24322 58492 24332 58548
rect 24388 58492 24780 58548
rect 24836 58492 25676 58548
rect 25732 58492 25742 58548
rect 32274 58492 32284 58548
rect 32340 58492 33740 58548
rect 33796 58492 34524 58548
rect 34580 58492 34590 58548
rect 2706 58380 2716 58436
rect 2772 58380 4060 58436
rect 4116 58380 4284 58436
rect 4340 58380 5292 58436
rect 5348 58380 5358 58436
rect 6514 58380 6524 58436
rect 6580 58380 7196 58436
rect 7252 58380 7262 58436
rect 10882 58380 10892 58436
rect 10948 58380 12012 58436
rect 12068 58380 12078 58436
rect 21970 58380 21980 58436
rect 22036 58380 24556 58436
rect 24612 58380 26124 58436
rect 26180 58380 26572 58436
rect 26628 58380 26638 58436
rect 26786 58380 26796 58436
rect 26852 58380 27132 58436
rect 27188 58380 27804 58436
rect 27860 58380 27870 58436
rect 34290 58380 34300 58436
rect 34356 58380 35084 58436
rect 35140 58380 37548 58436
rect 37604 58380 37614 58436
rect 18274 58268 18284 58324
rect 18340 58268 18844 58324
rect 18900 58268 19852 58324
rect 19908 58268 20300 58324
rect 20356 58268 20366 58324
rect 25526 58268 25564 58324
rect 25620 58268 25630 58324
rect 30594 58268 30604 58324
rect 30660 58268 31612 58324
rect 31668 58268 31678 58324
rect 18386 58156 18396 58212
rect 18452 58156 19068 58212
rect 19124 58156 19134 58212
rect 28018 58156 28028 58212
rect 28084 58156 28476 58212
rect 28532 58156 28542 58212
rect 29474 58156 29484 58212
rect 29540 58156 30156 58212
rect 30212 58156 30222 58212
rect 37874 58156 37884 58212
rect 37940 58156 39116 58212
rect 39172 58156 39182 58212
rect 24994 58044 25004 58100
rect 25060 58044 38220 58100
rect 38276 58044 38668 58100
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 37650 57932 37660 57988
rect 37716 57932 38108 57988
rect 38164 57932 38174 57988
rect 5282 57820 5292 57876
rect 5348 57820 6412 57876
rect 6468 57820 6748 57876
rect 6804 57820 7980 57876
rect 8036 57820 8046 57876
rect 11890 57820 11900 57876
rect 11956 57820 14028 57876
rect 14084 57820 14700 57876
rect 14756 57820 14766 57876
rect 32386 57820 32396 57876
rect 32452 57820 34076 57876
rect 34132 57820 34142 57876
rect 38612 57764 38668 58044
rect 19842 57708 19852 57764
rect 19908 57708 23324 57764
rect 23380 57708 23390 57764
rect 38612 57708 38780 57764
rect 38836 57708 39676 57764
rect 39732 57708 39742 57764
rect 1922 57596 1932 57652
rect 1988 57596 3276 57652
rect 3332 57596 5180 57652
rect 5236 57596 5246 57652
rect 17938 57596 17948 57652
rect 18004 57596 18508 57652
rect 18564 57596 18574 57652
rect 25526 57596 25564 57652
rect 25620 57596 25630 57652
rect 25788 57596 27916 57652
rect 27972 57596 27982 57652
rect 32050 57596 32060 57652
rect 32116 57596 33068 57652
rect 33124 57596 33134 57652
rect 25788 57540 25844 57596
rect 3042 57484 3052 57540
rect 3108 57484 4060 57540
rect 4116 57484 7308 57540
rect 7364 57484 7374 57540
rect 24546 57484 24556 57540
rect 24612 57484 24780 57540
rect 24836 57484 25340 57540
rect 25396 57484 25844 57540
rect 30146 57484 30156 57540
rect 30212 57484 30716 57540
rect 30772 57484 30782 57540
rect 3490 57372 3500 57428
rect 3556 57372 4508 57428
rect 4564 57372 4574 57428
rect 26562 57372 26572 57428
rect 26628 57372 32060 57428
rect 32116 57372 32126 57428
rect 23090 57260 23100 57316
rect 23156 57260 27132 57316
rect 27188 57260 27198 57316
rect 0 57204 400 57232
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 0 57148 3556 57204
rect 18274 57148 18284 57204
rect 18340 57148 18844 57204
rect 18900 57148 18910 57204
rect 23538 57148 23548 57204
rect 23604 57148 26796 57204
rect 26852 57148 26862 57204
rect 28466 57148 28476 57204
rect 28532 57148 30268 57204
rect 30324 57148 30334 57204
rect 31490 57148 31500 57204
rect 31556 57148 33740 57204
rect 33796 57148 35028 57204
rect 41906 57148 41916 57204
rect 41972 57148 42700 57204
rect 42756 57148 42766 57204
rect 0 57120 400 57148
rect 3500 57092 3556 57148
rect 34972 57092 35028 57148
rect 3500 57036 6804 57092
rect 7970 57036 7980 57092
rect 8036 57036 8316 57092
rect 8372 57036 9548 57092
rect 9604 57036 10780 57092
rect 10836 57036 12124 57092
rect 12180 57036 12190 57092
rect 19730 57036 19740 57092
rect 19796 57036 23100 57092
rect 23156 57036 23166 57092
rect 25442 57036 25452 57092
rect 25508 57036 26236 57092
rect 26292 57036 26302 57092
rect 34972 57036 35420 57092
rect 35476 57036 35486 57092
rect 6748 56980 6804 57036
rect 6738 56924 6748 56980
rect 6804 56924 6814 56980
rect 25638 56924 25676 56980
rect 25732 56924 30716 56980
rect 30772 56924 30782 56980
rect 34290 56924 34300 56980
rect 34356 56924 34972 56980
rect 35028 56924 35532 56980
rect 35588 56924 35598 56980
rect 2930 56812 2940 56868
rect 2996 56812 5852 56868
rect 5908 56812 5918 56868
rect 7074 56812 7084 56868
rect 7140 56812 7532 56868
rect 7588 56812 8988 56868
rect 9044 56812 9996 56868
rect 10052 56812 10062 56868
rect 17042 56812 17052 56868
rect 17108 56812 18620 56868
rect 18676 56812 19852 56868
rect 19908 56812 19918 56868
rect 20066 56700 20076 56756
rect 20132 56700 23884 56756
rect 23940 56700 23950 56756
rect 17714 56588 17724 56644
rect 17780 56588 18172 56644
rect 18228 56588 18508 56644
rect 18564 56588 18574 56644
rect 19058 56588 19068 56644
rect 19124 56588 21308 56644
rect 21364 56588 21374 56644
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 35410 56252 35420 56308
rect 35476 56252 38668 56308
rect 38724 56252 41020 56308
rect 41076 56252 41086 56308
rect 40674 56028 40684 56084
rect 40740 56028 41804 56084
rect 41860 56028 42476 56084
rect 42532 56028 42542 56084
rect 22754 55916 22764 55972
rect 22820 55916 24556 55972
rect 24612 55916 24622 55972
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 6636 55468 7980 55524
rect 8036 55468 8046 55524
rect 35186 55468 35196 55524
rect 35252 55468 36092 55524
rect 36148 55468 36158 55524
rect 41010 55468 41020 55524
rect 41076 55468 42868 55524
rect 3714 55356 3724 55412
rect 3780 55356 4172 55412
rect 4228 55356 4238 55412
rect 6636 55300 6692 55468
rect 42812 55412 42868 55468
rect 41234 55356 41244 55412
rect 41300 55356 42364 55412
rect 42420 55356 42430 55412
rect 42802 55356 42812 55412
rect 42868 55356 44156 55412
rect 44212 55356 44222 55412
rect 1922 55244 1932 55300
rect 1988 55244 4620 55300
rect 4676 55244 6636 55300
rect 6692 55244 6702 55300
rect 20178 55244 20188 55300
rect 20244 55244 21420 55300
rect 21476 55244 21486 55300
rect 3714 55132 3724 55188
rect 3780 55132 4060 55188
rect 4116 55132 6188 55188
rect 6244 55132 6254 55188
rect 20738 55132 20748 55188
rect 20804 55132 25340 55188
rect 25396 55132 25406 55188
rect 4162 55020 4172 55076
rect 4228 55020 4732 55076
rect 4788 55020 5740 55076
rect 5796 55020 5806 55076
rect 6066 55020 6076 55076
rect 6132 55020 7196 55076
rect 7252 55020 7262 55076
rect 13122 55020 13132 55076
rect 13188 55020 15148 55076
rect 17826 55020 17836 55076
rect 17892 55020 18508 55076
rect 18564 55020 23100 55076
rect 23156 55020 23166 55076
rect 41906 55020 41916 55076
rect 41972 55020 42252 55076
rect 42308 55020 42318 55076
rect 5170 54908 5180 54964
rect 5236 54908 5964 54964
rect 6020 54908 6030 54964
rect 2594 54684 2604 54740
rect 2660 54684 3612 54740
rect 3668 54684 3678 54740
rect 15092 54516 15148 55020
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 18722 54684 18732 54740
rect 18788 54684 19628 54740
rect 19684 54684 19694 54740
rect 28018 54684 28028 54740
rect 28084 54684 29708 54740
rect 29764 54684 30044 54740
rect 30100 54684 41356 54740
rect 41412 54684 41422 54740
rect 23314 54572 23324 54628
rect 23380 54572 24108 54628
rect 24164 54572 25340 54628
rect 25396 54572 25406 54628
rect 26226 54572 26236 54628
rect 26292 54572 37324 54628
rect 37380 54572 38332 54628
rect 38388 54572 38668 54628
rect 3266 54460 3276 54516
rect 3332 54460 3612 54516
rect 3668 54460 3678 54516
rect 15092 54460 23212 54516
rect 23268 54460 25228 54516
rect 25284 54460 25900 54516
rect 25956 54460 25966 54516
rect 28130 54460 28140 54516
rect 28196 54460 28812 54516
rect 28868 54460 28878 54516
rect 34178 54460 34188 54516
rect 34244 54460 34860 54516
rect 34916 54460 34926 54516
rect 1922 54348 1932 54404
rect 1988 54348 2492 54404
rect 2548 54348 2558 54404
rect 13794 54348 13804 54404
rect 13860 54348 15148 54404
rect 28578 54348 28588 54404
rect 28644 54348 28924 54404
rect 28980 54348 28990 54404
rect 38612 54348 38668 54572
rect 41010 54460 41020 54516
rect 41076 54460 41356 54516
rect 41412 54460 42364 54516
rect 42420 54460 42430 54516
rect 38724 54348 41580 54404
rect 41636 54348 42812 54404
rect 42868 54348 42878 54404
rect 15092 54292 15148 54348
rect 15092 54236 16380 54292
rect 16436 54236 18172 54292
rect 18228 54236 19516 54292
rect 19572 54236 20524 54292
rect 20580 54236 20590 54292
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 4162 53900 4172 53956
rect 4228 53900 4508 53956
rect 4564 53900 7980 53956
rect 8036 53900 9436 53956
rect 9492 53900 9502 53956
rect 29698 53900 29708 53956
rect 29764 53900 30156 53956
rect 30212 53900 30222 53956
rect 3602 53788 3612 53844
rect 3668 53788 7644 53844
rect 7700 53788 7710 53844
rect 20626 53788 20636 53844
rect 20692 53788 23436 53844
rect 23492 53788 25676 53844
rect 25732 53788 25742 53844
rect 27794 53788 27804 53844
rect 27860 53788 28252 53844
rect 28308 53788 28644 53844
rect 42802 53788 42812 53844
rect 42868 53788 43596 53844
rect 43652 53788 43662 53844
rect 28588 53732 28644 53788
rect 3154 53676 3164 53732
rect 3220 53676 4172 53732
rect 4228 53676 4238 53732
rect 18946 53676 18956 53732
rect 19012 53676 20076 53732
rect 20132 53676 22764 53732
rect 22820 53676 22830 53732
rect 26002 53676 26012 53732
rect 26068 53676 26684 53732
rect 26740 53676 26750 53732
rect 28578 53676 28588 53732
rect 28644 53676 29372 53732
rect 29428 53676 29820 53732
rect 29876 53676 29886 53732
rect 4274 53564 4284 53620
rect 4340 53564 5516 53620
rect 5572 53564 5852 53620
rect 5908 53564 6524 53620
rect 6580 53564 6590 53620
rect 18274 53564 18284 53620
rect 18340 53564 21644 53620
rect 21700 53564 21710 53620
rect 23202 53564 23212 53620
rect 23268 53564 26908 53620
rect 26964 53564 26974 53620
rect 3714 53452 3724 53508
rect 3780 53452 5740 53508
rect 5796 53452 5806 53508
rect 6738 53452 6748 53508
rect 6804 53452 8428 53508
rect 8484 53452 8494 53508
rect 12114 53452 12124 53508
rect 12180 53452 12572 53508
rect 12628 53452 13580 53508
rect 13636 53452 13646 53508
rect 23314 53452 23324 53508
rect 23380 53452 29036 53508
rect 29092 53452 29102 53508
rect 42130 53452 42140 53508
rect 42196 53452 43148 53508
rect 43204 53452 43214 53508
rect 4834 53340 4844 53396
rect 4900 53340 6076 53396
rect 6132 53340 6972 53396
rect 7028 53340 7038 53396
rect 7532 53340 8932 53396
rect 7532 53172 7588 53340
rect 8876 53284 8932 53340
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 8866 53228 8876 53284
rect 8932 53228 8942 53284
rect 4050 53116 4060 53172
rect 4116 53116 5292 53172
rect 5348 53116 7532 53172
rect 7588 53116 7598 53172
rect 7746 53116 7756 53172
rect 7812 53116 8428 53172
rect 8484 53116 8494 53172
rect 22754 53116 22764 53172
rect 22820 53116 23436 53172
rect 23492 53116 23502 53172
rect 23986 53116 23996 53172
rect 24052 53116 25676 53172
rect 25732 53116 29708 53172
rect 29764 53116 29774 53172
rect 35522 53116 35532 53172
rect 35588 53116 38892 53172
rect 38948 53116 39900 53172
rect 39956 53116 42364 53172
rect 42420 53116 43148 53172
rect 43204 53116 43214 53172
rect 23996 53060 24052 53116
rect 4274 53004 4284 53060
rect 4340 53004 7644 53060
rect 7700 53004 7710 53060
rect 20514 53004 20524 53060
rect 20580 53004 23212 53060
rect 23268 53004 24052 53060
rect 4274 52892 4284 52948
rect 4340 52892 4508 52948
rect 4564 52892 4574 52948
rect 28578 52892 28588 52948
rect 28644 52892 30156 52948
rect 30212 52892 33628 52948
rect 33684 52892 34636 52948
rect 34692 52892 35532 52948
rect 35588 52892 35598 52948
rect 2258 52780 2268 52836
rect 2324 52780 3276 52836
rect 3332 52780 4172 52836
rect 4228 52780 4238 52836
rect 6850 52780 6860 52836
rect 6916 52780 8092 52836
rect 8148 52780 8158 52836
rect 14914 52780 14924 52836
rect 14980 52780 15372 52836
rect 15428 52780 15438 52836
rect 28130 52780 28140 52836
rect 28196 52780 29148 52836
rect 29204 52780 29214 52836
rect 40226 52780 40236 52836
rect 40292 52780 41020 52836
rect 41076 52780 42140 52836
rect 42196 52780 42206 52836
rect 45154 52780 45164 52836
rect 45220 52780 46060 52836
rect 46116 52780 46126 52836
rect 2594 52668 2604 52724
rect 2660 52668 3500 52724
rect 3556 52668 5852 52724
rect 5908 52668 5918 52724
rect 19170 52668 19180 52724
rect 19236 52668 19628 52724
rect 19684 52668 23212 52724
rect 23268 52668 23278 52724
rect 29810 52668 29820 52724
rect 29876 52668 32060 52724
rect 32116 52668 33292 52724
rect 33348 52668 33358 52724
rect 2258 52556 2268 52612
rect 2324 52556 4060 52612
rect 4116 52556 4126 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 4834 52444 4844 52500
rect 4900 52444 5628 52500
rect 5684 52444 5694 52500
rect 35634 52444 35644 52500
rect 35700 52444 36204 52500
rect 36260 52444 36270 52500
rect 3714 52332 3724 52388
rect 3780 52332 4060 52388
rect 4116 52332 4126 52388
rect 42466 52332 42476 52388
rect 42532 52332 43372 52388
rect 43428 52332 43438 52388
rect 0 52276 400 52304
rect 0 52220 5292 52276
rect 5348 52220 5358 52276
rect 26450 52220 26460 52276
rect 26516 52220 28924 52276
rect 28980 52220 30716 52276
rect 30772 52220 30782 52276
rect 33170 52220 33180 52276
rect 33236 52220 38332 52276
rect 38388 52220 41132 52276
rect 41188 52220 41356 52276
rect 41412 52220 41422 52276
rect 42364 52220 45052 52276
rect 45108 52220 45118 52276
rect 0 52192 400 52220
rect 42364 52164 42420 52220
rect 3714 52108 3724 52164
rect 3780 52108 6412 52164
rect 6468 52108 6478 52164
rect 22194 52108 22204 52164
rect 22260 52108 24444 52164
rect 24500 52108 24510 52164
rect 33506 52108 33516 52164
rect 33572 52108 34188 52164
rect 34244 52108 34254 52164
rect 37650 52108 37660 52164
rect 37716 52108 42364 52164
rect 42420 52108 42430 52164
rect 42802 52108 42812 52164
rect 42868 52108 43932 52164
rect 43988 52108 43998 52164
rect 8978 51996 8988 52052
rect 9044 51996 9660 52052
rect 9716 51996 11116 52052
rect 11172 51996 11452 52052
rect 11508 51996 14476 52052
rect 14532 51996 14542 52052
rect 22754 51996 22764 52052
rect 22820 51996 23548 52052
rect 23604 51996 23614 52052
rect 28130 51996 28140 52052
rect 28196 51996 29820 52052
rect 29876 51996 29886 52052
rect 31836 51996 32732 52052
rect 32788 51996 32798 52052
rect 39862 51996 39900 52052
rect 39956 51996 39966 52052
rect 31836 51940 31892 51996
rect 2706 51884 2716 51940
rect 2772 51884 3276 51940
rect 3332 51884 4284 51940
rect 4340 51884 4396 51940
rect 4452 51884 4462 51940
rect 10434 51884 10444 51940
rect 10500 51884 11564 51940
rect 11620 51884 11630 51940
rect 29698 51884 29708 51940
rect 29764 51884 31052 51940
rect 31108 51884 31836 51940
rect 31892 51884 31902 51940
rect 32274 51884 32284 51940
rect 32340 51884 32844 51940
rect 32900 51884 33068 51940
rect 33124 51884 33134 51940
rect 33954 51884 33964 51940
rect 34020 51884 34524 51940
rect 34580 51884 34590 51940
rect 37426 51884 37436 51940
rect 37492 51884 38668 51940
rect 38724 51884 38734 51940
rect 11330 51772 11340 51828
rect 11396 51772 12012 51828
rect 12068 51772 12078 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 28242 51548 28252 51604
rect 28308 51548 30716 51604
rect 30772 51548 31388 51604
rect 31444 51548 31454 51604
rect 37650 51548 37660 51604
rect 37716 51548 39228 51604
rect 39284 51548 40348 51604
rect 40404 51548 41468 51604
rect 41524 51548 41534 51604
rect 42130 51548 42140 51604
rect 42196 51548 43708 51604
rect 43764 51548 44156 51604
rect 44212 51548 44222 51604
rect 17938 51436 17948 51492
rect 18004 51436 26572 51492
rect 26628 51436 26638 51492
rect 6290 51324 6300 51380
rect 6356 51324 7532 51380
rect 7588 51324 7598 51380
rect 22754 51324 22764 51380
rect 22820 51324 23660 51380
rect 23716 51324 23726 51380
rect 38322 51324 38332 51380
rect 38388 51324 39452 51380
rect 39508 51324 39518 51380
rect 42018 51324 42028 51380
rect 42084 51324 42252 51380
rect 42308 51324 42318 51380
rect 3154 51212 3164 51268
rect 3220 51212 3724 51268
rect 3780 51212 4172 51268
rect 4228 51212 4508 51268
rect 4564 51212 4574 51268
rect 7298 51212 7308 51268
rect 7364 51212 8540 51268
rect 8596 51212 8606 51268
rect 30258 51212 30268 51268
rect 30324 51212 31052 51268
rect 31108 51212 31118 51268
rect 34962 51212 34972 51268
rect 35028 51212 35980 51268
rect 36036 51212 36046 51268
rect 2034 50988 2044 51044
rect 2100 50988 3388 51044
rect 3444 50988 3454 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 8372 50596 8428 51212
rect 34178 51100 34188 51156
rect 34244 51100 41356 51156
rect 41412 51100 41422 51156
rect 22642 50988 22652 51044
rect 22708 50988 23436 51044
rect 23492 50988 23502 51044
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 33618 50876 33628 50932
rect 33684 50876 34860 50932
rect 34916 50876 34926 50932
rect 26852 50764 27580 50820
rect 27636 50764 28028 50820
rect 28084 50764 28094 50820
rect 33058 50764 33068 50820
rect 33124 50764 42028 50820
rect 42084 50764 42094 50820
rect 11442 50652 11452 50708
rect 11508 50652 12684 50708
rect 12740 50652 13244 50708
rect 13300 50652 13310 50708
rect 14466 50652 14476 50708
rect 14532 50652 15820 50708
rect 15876 50652 22652 50708
rect 22708 50652 22718 50708
rect 3490 50540 3500 50596
rect 3556 50540 3948 50596
rect 4004 50540 4844 50596
rect 4900 50540 4910 50596
rect 6290 50540 6300 50596
rect 6356 50540 7308 50596
rect 7364 50540 7374 50596
rect 7634 50540 7644 50596
rect 7700 50540 10556 50596
rect 10612 50540 10622 50596
rect 11330 50540 11340 50596
rect 11396 50540 14252 50596
rect 14308 50540 14924 50596
rect 14980 50540 14990 50596
rect 16146 50540 16156 50596
rect 16212 50540 18732 50596
rect 18788 50540 19852 50596
rect 19908 50540 22540 50596
rect 22596 50540 22988 50596
rect 23044 50540 24668 50596
rect 24724 50540 25340 50596
rect 25396 50540 25406 50596
rect 26852 50484 26908 50764
rect 27794 50652 27804 50708
rect 27860 50652 28252 50708
rect 28308 50652 28318 50708
rect 29446 50652 29484 50708
rect 29540 50652 29550 50708
rect 30146 50652 30156 50708
rect 30212 50652 31164 50708
rect 31220 50652 31500 50708
rect 31556 50652 33628 50708
rect 33684 50652 35756 50708
rect 35812 50652 37660 50708
rect 37716 50652 37726 50708
rect 27010 50540 27020 50596
rect 27076 50540 27244 50596
rect 27300 50540 27310 50596
rect 30146 50540 30156 50596
rect 30212 50540 30716 50596
rect 30772 50540 32396 50596
rect 32452 50540 32462 50596
rect 32722 50540 32732 50596
rect 32788 50540 33740 50596
rect 33796 50540 33806 50596
rect 34850 50540 34860 50596
rect 34916 50540 36204 50596
rect 36260 50540 36270 50596
rect 2706 50428 2716 50484
rect 2772 50428 3724 50484
rect 3780 50428 4732 50484
rect 4788 50428 4798 50484
rect 6066 50428 6076 50484
rect 6132 50428 7868 50484
rect 7924 50428 9660 50484
rect 9716 50428 9726 50484
rect 17714 50428 17724 50484
rect 17780 50428 26236 50484
rect 26292 50428 26908 50484
rect 28914 50428 28924 50484
rect 28980 50428 29820 50484
rect 29876 50428 29886 50484
rect 34738 50428 34748 50484
rect 34804 50428 35868 50484
rect 35924 50428 38668 50484
rect 38724 50428 38734 50484
rect 41346 50428 41356 50484
rect 41412 50428 42028 50484
rect 42084 50428 42094 50484
rect 3266 50316 3276 50372
rect 3332 50316 3500 50372
rect 3556 50316 3566 50372
rect 29026 50204 29036 50260
rect 29092 50204 31164 50260
rect 31220 50204 31230 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 31238 50092 31276 50148
rect 31332 50092 31342 50148
rect 29698 49980 29708 50036
rect 29764 49980 30828 50036
rect 30884 49980 30894 50036
rect 3938 49868 3948 49924
rect 4004 49868 4844 49924
rect 4900 49868 4910 49924
rect 28242 49868 28252 49924
rect 28308 49868 28588 49924
rect 28644 49868 30492 49924
rect 30548 49868 30558 49924
rect 31266 49868 31276 49924
rect 31332 49868 31342 49924
rect 31276 49812 31332 49868
rect 1810 49756 1820 49812
rect 1876 49756 5292 49812
rect 5348 49756 6076 49812
rect 6132 49756 6142 49812
rect 11116 49756 13468 49812
rect 13524 49756 13534 49812
rect 16594 49756 16604 49812
rect 16660 49756 19628 49812
rect 19684 49756 19694 49812
rect 29698 49756 29708 49812
rect 29764 49756 30156 49812
rect 30212 49756 30222 49812
rect 30370 49756 30380 49812
rect 30436 49756 31332 49812
rect 32498 49756 32508 49812
rect 32564 49756 33068 49812
rect 33124 49756 33134 49812
rect 33730 49756 33740 49812
rect 33796 49756 34748 49812
rect 34804 49756 34814 49812
rect 11116 49700 11172 49756
rect 3938 49644 3948 49700
rect 4004 49644 4396 49700
rect 4452 49644 4462 49700
rect 8082 49644 8092 49700
rect 8148 49644 9772 49700
rect 9828 49644 11116 49700
rect 11172 49644 11182 49700
rect 12786 49644 12796 49700
rect 12852 49644 14924 49700
rect 14980 49644 14990 49700
rect 15586 49644 15596 49700
rect 15652 49644 16156 49700
rect 16212 49644 16222 49700
rect 21074 49644 21084 49700
rect 21140 49644 21756 49700
rect 21812 49644 21822 49700
rect 30482 49644 30492 49700
rect 30548 49644 31948 49700
rect 32004 49644 32014 49700
rect 32386 49644 32396 49700
rect 32452 49644 32956 49700
rect 33012 49644 33964 49700
rect 34020 49644 36540 49700
rect 36596 49644 36606 49700
rect 41906 49644 41916 49700
rect 41972 49644 43148 49700
rect 43204 49644 43214 49700
rect 31014 49532 31052 49588
rect 31108 49532 31118 49588
rect 31238 49532 31276 49588
rect 31332 49532 31342 49588
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 18946 49308 18956 49364
rect 19012 49308 19516 49364
rect 19572 49308 19582 49364
rect 2930 49196 2940 49252
rect 2996 49196 3388 49252
rect 4274 49196 4284 49252
rect 4340 49196 5964 49252
rect 6020 49196 6030 49252
rect 26786 49196 26796 49252
rect 26852 49196 27692 49252
rect 27748 49196 27758 49252
rect 28018 49196 28028 49252
rect 28084 49196 29260 49252
rect 29316 49196 29326 49252
rect 29810 49196 29820 49252
rect 29876 49196 30380 49252
rect 30436 49196 30446 49252
rect 3332 49140 3388 49196
rect 3332 49084 4508 49140
rect 4564 49084 6412 49140
rect 6468 49084 6972 49140
rect 7028 49084 7308 49140
rect 7364 49084 7374 49140
rect 2146 48972 2156 49028
rect 2212 48972 3052 49028
rect 3108 48972 3118 49028
rect 3266 48972 3276 49028
rect 3332 48972 4284 49028
rect 4340 48972 4350 49028
rect 20290 48972 20300 49028
rect 20356 48972 21308 49028
rect 21364 48972 22876 49028
rect 22932 48972 22942 49028
rect 31714 48972 31724 49028
rect 31780 48972 33740 49028
rect 33796 48972 33806 49028
rect 37650 48972 37660 49028
rect 37716 48972 38332 49028
rect 38388 48972 40124 49028
rect 40180 48972 40190 49028
rect 1922 48860 1932 48916
rect 1988 48860 2268 48916
rect 2324 48860 3388 48916
rect 3444 48860 3454 48916
rect 8530 48860 8540 48916
rect 8596 48860 9100 48916
rect 9156 48860 9996 48916
rect 10052 48860 10062 48916
rect 14914 48860 14924 48916
rect 14980 48860 18732 48916
rect 18788 48860 18798 48916
rect 24098 48860 24108 48916
rect 24164 48860 25676 48916
rect 25732 48860 26796 48916
rect 26852 48860 26862 48916
rect 30258 48860 30268 48916
rect 30324 48860 32956 48916
rect 33012 48860 33022 48916
rect 7522 48748 7532 48804
rect 7588 48748 8876 48804
rect 8932 48748 8942 48804
rect 14018 48748 14028 48804
rect 14084 48748 15484 48804
rect 15540 48748 15550 48804
rect 17602 48748 17612 48804
rect 17668 48748 18844 48804
rect 18900 48748 20076 48804
rect 20132 48748 20142 48804
rect 21298 48748 21308 48804
rect 21364 48748 22540 48804
rect 22596 48748 22606 48804
rect 23062 48748 23100 48804
rect 23156 48748 23166 48804
rect 23314 48748 23324 48804
rect 23380 48748 24444 48804
rect 24500 48748 24510 48804
rect 34962 48748 34972 48804
rect 35028 48748 35644 48804
rect 35700 48748 35710 48804
rect 36530 48748 36540 48804
rect 36596 48748 37100 48804
rect 37156 48748 38668 48804
rect 38612 48692 38668 48748
rect 38612 48636 41020 48692
rect 41076 48636 42476 48692
rect 42532 48636 42924 48692
rect 42980 48636 42990 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 11676 48524 14700 48580
rect 14756 48524 14766 48580
rect 11676 48468 11732 48524
rect 2818 48412 2828 48468
rect 2884 48412 4060 48468
rect 4116 48412 4126 48468
rect 8866 48412 8876 48468
rect 8932 48412 9324 48468
rect 9380 48412 9884 48468
rect 9940 48412 11676 48468
rect 11732 48412 11742 48468
rect 12898 48412 12908 48468
rect 12964 48412 16156 48468
rect 16212 48412 16716 48468
rect 16772 48412 16782 48468
rect 35252 48412 37100 48468
rect 37156 48412 37660 48468
rect 37716 48412 37726 48468
rect 9650 48300 9660 48356
rect 9716 48300 10332 48356
rect 10388 48300 10398 48356
rect 23874 48300 23884 48356
rect 23940 48300 25228 48356
rect 25284 48300 25900 48356
rect 25956 48300 25966 48356
rect 28886 48300 28924 48356
rect 28980 48300 28990 48356
rect 35252 48244 35308 48412
rect 36754 48300 36764 48356
rect 36820 48300 37772 48356
rect 37828 48300 37838 48356
rect 41234 48300 41244 48356
rect 41300 48300 42140 48356
rect 42196 48300 42206 48356
rect 18610 48188 18620 48244
rect 18676 48188 20300 48244
rect 20356 48188 20366 48244
rect 24668 48188 28364 48244
rect 28420 48188 28588 48244
rect 28644 48188 31500 48244
rect 31556 48188 31566 48244
rect 33058 48188 33068 48244
rect 33124 48188 35308 48244
rect 41570 48188 41580 48244
rect 41636 48188 42700 48244
rect 42756 48188 42766 48244
rect 24668 48132 24724 48188
rect 2370 48076 2380 48132
rect 2436 48076 3276 48132
rect 3332 48076 3500 48132
rect 3556 48076 3566 48132
rect 8306 48076 8316 48132
rect 8372 48076 10444 48132
rect 10500 48076 10510 48132
rect 18050 48076 18060 48132
rect 18116 48076 20636 48132
rect 20692 48076 20702 48132
rect 21410 48076 21420 48132
rect 21476 48076 22092 48132
rect 22148 48076 22158 48132
rect 24658 48076 24668 48132
rect 24724 48076 24734 48132
rect 24994 48076 25004 48132
rect 25060 48076 28924 48132
rect 28980 48076 30380 48132
rect 30436 48076 30604 48132
rect 30660 48076 31388 48132
rect 31444 48076 31454 48132
rect 2482 47964 2492 48020
rect 2548 47964 3164 48020
rect 3220 47964 3230 48020
rect 6738 47964 6748 48020
rect 6804 47964 7196 48020
rect 7252 47964 7262 48020
rect 42242 47852 42252 47908
rect 42308 47852 42318 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 1922 47740 1932 47796
rect 1988 47740 2716 47796
rect 2772 47740 2782 47796
rect 4610 47628 4620 47684
rect 4676 47628 6748 47684
rect 6804 47628 6814 47684
rect 29586 47628 29596 47684
rect 29652 47628 32172 47684
rect 32228 47628 32238 47684
rect 28588 47516 29820 47572
rect 29876 47516 29886 47572
rect 31378 47516 31388 47572
rect 31444 47516 35084 47572
rect 35140 47516 35150 47572
rect 37314 47516 37324 47572
rect 37380 47516 38556 47572
rect 38612 47516 40348 47572
rect 40404 47516 40414 47572
rect 28588 47460 28644 47516
rect 2258 47404 2268 47460
rect 2324 47404 2884 47460
rect 3154 47404 3164 47460
rect 3220 47404 3500 47460
rect 3556 47404 3566 47460
rect 4050 47404 4060 47460
rect 4116 47404 4126 47460
rect 5842 47404 5852 47460
rect 5908 47404 8988 47460
rect 9044 47404 9054 47460
rect 23538 47404 23548 47460
rect 23604 47404 23884 47460
rect 23940 47404 23950 47460
rect 24434 47404 24444 47460
rect 24500 47404 26124 47460
rect 26180 47404 28140 47460
rect 28196 47404 28588 47460
rect 28644 47404 28654 47460
rect 29474 47404 29484 47460
rect 29540 47404 30044 47460
rect 30100 47404 30110 47460
rect 34402 47404 34412 47460
rect 34468 47404 36092 47460
rect 36148 47404 37212 47460
rect 37268 47404 37278 47460
rect 0 47348 400 47376
rect 0 47292 2380 47348
rect 2436 47292 2446 47348
rect 0 47264 400 47292
rect 2828 47236 2884 47404
rect 4060 47348 4116 47404
rect 42252 47348 42308 47852
rect 42690 47404 42700 47460
rect 42756 47404 42868 47460
rect 4060 47292 5012 47348
rect 11666 47292 11676 47348
rect 11732 47292 12236 47348
rect 12292 47292 12302 47348
rect 25666 47292 25676 47348
rect 25732 47292 27580 47348
rect 27636 47292 27646 47348
rect 31042 47292 31052 47348
rect 31108 47292 32060 47348
rect 32116 47292 32126 47348
rect 42252 47292 42588 47348
rect 42644 47292 42654 47348
rect 4956 47236 5012 47292
rect 42812 47236 42868 47404
rect 43250 47292 43260 47348
rect 43316 47292 43820 47348
rect 43876 47292 43886 47348
rect 2828 47180 4116 47236
rect 4946 47180 4956 47236
rect 5012 47180 5022 47236
rect 16818 47180 16828 47236
rect 16884 47180 18060 47236
rect 18116 47180 18126 47236
rect 18834 47180 18844 47236
rect 18900 47180 19964 47236
rect 20020 47180 20244 47236
rect 22306 47180 22316 47236
rect 22372 47180 35532 47236
rect 35588 47180 35598 47236
rect 39106 47180 39116 47236
rect 39172 47180 39900 47236
rect 39956 47180 39966 47236
rect 42242 47180 42252 47236
rect 42308 47180 42868 47236
rect 4060 47012 4116 47180
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 20188 47012 20244 47180
rect 21522 47068 21532 47124
rect 21588 47068 24668 47124
rect 24724 47068 24734 47124
rect 26562 47068 26572 47124
rect 26628 47068 27356 47124
rect 27412 47068 27916 47124
rect 27972 47068 27982 47124
rect 34626 47068 34636 47124
rect 34692 47068 36540 47124
rect 36596 47068 36606 47124
rect 41346 47068 41356 47124
rect 41412 47068 42364 47124
rect 42420 47068 42430 47124
rect 2930 46956 2940 47012
rect 2996 46956 3612 47012
rect 3668 46956 3678 47012
rect 4050 46956 4060 47012
rect 4116 46956 4126 47012
rect 9314 46956 9324 47012
rect 9380 46956 9772 47012
rect 9828 46956 9838 47012
rect 20188 46956 20636 47012
rect 20692 46956 21756 47012
rect 21812 46956 21822 47012
rect 29922 46956 29932 47012
rect 29988 46956 32620 47012
rect 32676 46956 32686 47012
rect 19506 46844 19516 46900
rect 19572 46844 21644 46900
rect 21700 46844 23548 46900
rect 23604 46844 23614 46900
rect 31826 46844 31836 46900
rect 31892 46844 32508 46900
rect 32564 46844 32574 46900
rect 36194 46844 36204 46900
rect 36260 46844 41244 46900
rect 41300 46844 41310 46900
rect 5142 46732 5180 46788
rect 5236 46732 5516 46788
rect 5572 46732 5582 46788
rect 10098 46732 10108 46788
rect 10164 46732 11116 46788
rect 11172 46732 11182 46788
rect 21410 46732 21420 46788
rect 21476 46732 22316 46788
rect 22372 46732 22382 46788
rect 23986 46732 23996 46788
rect 24052 46732 28140 46788
rect 28196 46732 32396 46788
rect 32452 46732 33292 46788
rect 33348 46732 34636 46788
rect 34692 46732 34702 46788
rect 37090 46732 37100 46788
rect 37156 46732 39564 46788
rect 39620 46732 39630 46788
rect 41906 46732 41916 46788
rect 41972 46732 43596 46788
rect 43652 46732 43662 46788
rect 44146 46732 44156 46788
rect 44212 46732 45948 46788
rect 46004 46732 46014 46788
rect 23996 46676 24052 46732
rect 3266 46620 3276 46676
rect 3332 46620 3612 46676
rect 3668 46620 4844 46676
rect 4900 46620 4910 46676
rect 6290 46620 6300 46676
rect 6356 46620 8316 46676
rect 8372 46620 8382 46676
rect 16146 46620 16156 46676
rect 16212 46620 16828 46676
rect 16884 46620 16894 46676
rect 20290 46620 20300 46676
rect 20356 46620 21308 46676
rect 21364 46620 21532 46676
rect 21588 46620 21598 46676
rect 21858 46620 21868 46676
rect 21924 46620 24052 46676
rect 25890 46620 25900 46676
rect 25956 46620 26236 46676
rect 26292 46620 26302 46676
rect 29026 46620 29036 46676
rect 29092 46620 30492 46676
rect 30548 46620 30558 46676
rect 2594 46508 2604 46564
rect 2660 46508 2670 46564
rect 3042 46508 3052 46564
rect 3108 46508 4284 46564
rect 4340 46508 4350 46564
rect 6178 46508 6188 46564
rect 6244 46508 7196 46564
rect 7252 46508 7262 46564
rect 14466 46508 14476 46564
rect 14532 46508 15372 46564
rect 15428 46508 15438 46564
rect 18834 46508 18844 46564
rect 18900 46508 19292 46564
rect 19348 46508 19358 46564
rect 20066 46508 20076 46564
rect 20132 46508 22764 46564
rect 22820 46508 22830 46564
rect 23426 46508 23436 46564
rect 23492 46508 29820 46564
rect 29876 46508 29886 46564
rect 32274 46508 32284 46564
rect 32340 46508 33292 46564
rect 33348 46508 33358 46564
rect 2604 46452 2660 46508
rect 2604 46396 3276 46452
rect 3332 46396 3342 46452
rect 30678 46396 30716 46452
rect 30772 46396 30782 46452
rect 38098 46396 38108 46452
rect 38164 46396 38780 46452
rect 38836 46396 38846 46452
rect 2146 46284 2156 46340
rect 2212 46284 2940 46340
rect 2996 46284 3006 46340
rect 26226 46284 26236 46340
rect 26292 46284 26908 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 2370 46060 2380 46116
rect 2436 46060 2940 46116
rect 2996 46060 3500 46116
rect 3556 46060 3566 46116
rect 3714 46060 3724 46116
rect 3780 46060 4396 46116
rect 4452 46060 4462 46116
rect 20178 46060 20188 46116
rect 20244 46060 20636 46116
rect 20692 46060 20702 46116
rect 26852 46004 26908 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 35970 46060 35980 46116
rect 36036 46060 38220 46116
rect 38276 46060 38286 46116
rect 8418 45948 8428 46004
rect 8484 45948 9100 46004
rect 9156 45948 9166 46004
rect 26852 45948 28588 46004
rect 28644 45948 29372 46004
rect 29428 45948 29438 46004
rect 38322 45948 38332 46004
rect 38388 45948 41972 46004
rect 3266 45836 3276 45892
rect 3332 45836 3612 45892
rect 3668 45836 3678 45892
rect 13458 45836 13468 45892
rect 13524 45836 14924 45892
rect 14980 45836 20300 45892
rect 20356 45836 20366 45892
rect 22306 45836 22316 45892
rect 22372 45836 22988 45892
rect 23044 45836 23660 45892
rect 23716 45836 23726 45892
rect 30146 45836 30156 45892
rect 30212 45836 31276 45892
rect 31332 45836 31342 45892
rect 33282 45836 33292 45892
rect 33348 45836 35196 45892
rect 35252 45836 35532 45892
rect 35588 45836 36092 45892
rect 36148 45836 36158 45892
rect 16594 45724 16604 45780
rect 16660 45724 19516 45780
rect 19572 45724 19582 45780
rect 19842 45724 19852 45780
rect 19908 45724 21756 45780
rect 21812 45724 21822 45780
rect 27234 45724 27244 45780
rect 27300 45724 29372 45780
rect 29428 45724 29438 45780
rect 30706 45724 30716 45780
rect 30772 45724 31500 45780
rect 31556 45724 31566 45780
rect 39442 45724 39452 45780
rect 39508 45724 40348 45780
rect 40404 45724 41132 45780
rect 41188 45724 41198 45780
rect 6066 45612 6076 45668
rect 6132 45612 6412 45668
rect 6468 45612 6860 45668
rect 6916 45612 7420 45668
rect 7476 45612 7486 45668
rect 15698 45612 15708 45668
rect 15764 45612 16156 45668
rect 16212 45612 17052 45668
rect 17108 45612 17118 45668
rect 19282 45612 19292 45668
rect 19348 45612 21420 45668
rect 21476 45612 21486 45668
rect 27682 45612 27692 45668
rect 27748 45612 29036 45668
rect 29092 45612 29102 45668
rect 35074 45612 35084 45668
rect 35140 45612 37772 45668
rect 37828 45612 38220 45668
rect 38276 45612 38286 45668
rect 41916 45556 41972 45948
rect 42578 45612 42588 45668
rect 42644 45612 42924 45668
rect 42980 45612 44044 45668
rect 44100 45612 44110 45668
rect 3042 45500 3052 45556
rect 3108 45500 4172 45556
rect 4228 45500 4238 45556
rect 28774 45500 28812 45556
rect 28868 45500 28878 45556
rect 41906 45500 41916 45556
rect 41972 45500 42364 45556
rect 42420 45500 42700 45556
rect 42756 45500 43148 45556
rect 43204 45500 43214 45556
rect 43586 45500 43596 45556
rect 43652 45500 44940 45556
rect 44996 45500 45006 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 4172 45388 5068 45444
rect 5124 45388 5134 45444
rect 28130 45388 28140 45444
rect 28196 45388 29036 45444
rect 29092 45388 30380 45444
rect 30436 45388 30446 45444
rect 35746 45388 35756 45444
rect 35812 45388 37548 45444
rect 37604 45388 38668 45444
rect 38724 45388 38734 45444
rect 4172 45332 4228 45388
rect 38668 45332 38724 45388
rect 4162 45276 4172 45332
rect 4228 45276 4238 45332
rect 28242 45276 28252 45332
rect 28308 45276 28924 45332
rect 28980 45276 28990 45332
rect 31154 45276 31164 45332
rect 31220 45276 32508 45332
rect 32564 45276 32574 45332
rect 33618 45276 33628 45332
rect 33684 45276 34300 45332
rect 34356 45276 34366 45332
rect 34626 45276 34636 45332
rect 34692 45276 35084 45332
rect 35140 45276 35150 45332
rect 38668 45276 41244 45332
rect 41300 45276 41310 45332
rect 41682 45276 41692 45332
rect 41748 45276 42476 45332
rect 42532 45276 42542 45332
rect 43026 45276 43036 45332
rect 43092 45276 43484 45332
rect 43540 45276 43550 45332
rect 33628 45220 33684 45276
rect 20738 45164 20748 45220
rect 20804 45164 21868 45220
rect 21924 45164 22316 45220
rect 22372 45164 22382 45220
rect 27346 45164 27356 45220
rect 27412 45164 28364 45220
rect 28420 45164 28430 45220
rect 30482 45164 30492 45220
rect 30548 45164 33684 45220
rect 42354 45164 42364 45220
rect 42420 45164 45164 45220
rect 45220 45164 48076 45220
rect 48132 45164 48142 45220
rect 24658 45052 24668 45108
rect 24724 45052 25452 45108
rect 25508 45052 25518 45108
rect 25666 45052 25676 45108
rect 25732 45052 33628 45108
rect 33684 45052 33852 45108
rect 33908 45052 33918 45108
rect 40012 45052 43372 45108
rect 43428 45052 43438 45108
rect 40012 44996 40068 45052
rect 2370 44940 2380 44996
rect 2436 44940 2940 44996
rect 2996 44940 3836 44996
rect 3892 44940 4620 44996
rect 4676 44940 4686 44996
rect 22978 44940 22988 44996
rect 23044 44940 23660 44996
rect 23716 44940 23726 44996
rect 24210 44940 24220 44996
rect 24276 44940 26684 44996
rect 26740 44940 26750 44996
rect 27122 44940 27132 44996
rect 27188 44940 27692 44996
rect 27748 44940 27758 44996
rect 28354 44940 28364 44996
rect 28420 44940 29372 44996
rect 29428 44940 29438 44996
rect 34962 44940 34972 44996
rect 35028 44940 36652 44996
rect 36708 44940 37100 44996
rect 37156 44940 37166 44996
rect 39330 44940 39340 44996
rect 39396 44940 40012 44996
rect 40068 44940 40078 44996
rect 41234 44940 41244 44996
rect 41300 44940 42700 44996
rect 42756 44940 42766 44996
rect 27010 44828 27020 44884
rect 27076 44828 27916 44884
rect 27972 44828 27982 44884
rect 21970 44716 21980 44772
rect 22036 44716 34636 44772
rect 34692 44716 34702 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 23202 44604 23212 44660
rect 23268 44604 25676 44660
rect 25732 44604 26236 44660
rect 26292 44604 26302 44660
rect 28018 44604 28028 44660
rect 28084 44604 28094 44660
rect 29138 44604 29148 44660
rect 29204 44604 29932 44660
rect 29988 44604 29998 44660
rect 41234 44604 41244 44660
rect 41300 44604 43484 44660
rect 43540 44604 43550 44660
rect 28028 44548 28084 44604
rect 2034 44492 2044 44548
rect 2100 44492 2268 44548
rect 2324 44492 2334 44548
rect 27346 44492 27356 44548
rect 27412 44492 28084 44548
rect 32050 44492 32060 44548
rect 32116 44492 33068 44548
rect 33124 44492 33134 44548
rect 33618 44492 33628 44548
rect 33684 44492 39004 44548
rect 39060 44492 40348 44548
rect 40404 44492 41132 44548
rect 41188 44492 41692 44548
rect 41748 44492 41758 44548
rect 6178 44380 6188 44436
rect 6244 44380 6748 44436
rect 6804 44380 7420 44436
rect 7476 44380 7486 44436
rect 16258 44380 16268 44436
rect 16324 44380 18620 44436
rect 18676 44380 19180 44436
rect 19236 44380 19246 44436
rect 27458 44380 27468 44436
rect 27524 44380 28028 44436
rect 28084 44380 30380 44436
rect 30436 44380 30446 44436
rect 35942 44380 35980 44436
rect 36036 44380 36046 44436
rect 37986 44380 37996 44436
rect 38052 44380 38444 44436
rect 38500 44380 39900 44436
rect 39956 44380 39966 44436
rect 42018 44380 42028 44436
rect 42084 44380 43372 44436
rect 43428 44380 43438 44436
rect 2482 44268 2492 44324
rect 2548 44268 2940 44324
rect 2996 44268 3388 44324
rect 3444 44268 3454 44324
rect 4722 44268 4732 44324
rect 4788 44268 6524 44324
rect 6580 44268 7532 44324
rect 7588 44268 7598 44324
rect 29362 44268 29372 44324
rect 29428 44268 29484 44324
rect 29540 44268 29550 44324
rect 33506 44268 33516 44324
rect 33572 44268 37548 44324
rect 37604 44268 37614 44324
rect 42578 44268 42588 44324
rect 42644 44268 44044 44324
rect 44100 44268 44828 44324
rect 44884 44268 44894 44324
rect 4732 44212 4788 44268
rect 2818 44156 2828 44212
rect 2884 44156 4788 44212
rect 26114 44156 26124 44212
rect 26180 44156 26684 44212
rect 26740 44156 26750 44212
rect 37650 44156 37660 44212
rect 37716 44156 39452 44212
rect 39508 44156 40796 44212
rect 40852 44156 42924 44212
rect 42980 44156 43372 44212
rect 43428 44156 43438 44212
rect 3500 44100 3556 44156
rect 3490 44044 3500 44100
rect 3556 44044 3566 44100
rect 3826 44044 3836 44100
rect 3892 44044 4284 44100
rect 4340 44044 4350 44100
rect 16370 44044 16380 44100
rect 16436 44044 17500 44100
rect 17556 44044 17566 44100
rect 22418 44044 22428 44100
rect 22484 44044 22764 44100
rect 22820 44044 22830 44100
rect 26450 44044 26460 44100
rect 26516 44044 28364 44100
rect 28420 44044 28430 44100
rect 28690 44044 28700 44100
rect 28756 44044 29036 44100
rect 29092 44044 29102 44100
rect 29474 44044 29484 44100
rect 29540 44044 29596 44100
rect 29652 44044 29662 44100
rect 35186 44044 35196 44100
rect 35252 44044 37212 44100
rect 37268 44044 37278 44100
rect 40898 44044 40908 44100
rect 40964 44044 41244 44100
rect 41300 44044 41310 44100
rect 2930 43932 2940 43988
rect 2996 43932 3388 43988
rect 3444 43932 3454 43988
rect 6066 43932 6076 43988
rect 6132 43932 6860 43988
rect 6916 43932 6926 43988
rect 23202 43932 23212 43988
rect 23268 43932 23996 43988
rect 24052 43932 24062 43988
rect 27010 43932 27020 43988
rect 27076 43932 27580 43988
rect 27636 43932 27646 43988
rect 3388 43876 3444 43932
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 3388 43820 8652 43876
rect 8708 43820 10332 43876
rect 10388 43820 10398 43876
rect 22306 43820 22316 43876
rect 22372 43820 24668 43876
rect 24724 43820 24734 43876
rect 27794 43820 27804 43876
rect 27860 43820 31388 43876
rect 31444 43820 31454 43876
rect 38322 43820 38332 43876
rect 38388 43820 39116 43876
rect 39172 43820 40348 43876
rect 40404 43820 40414 43876
rect 10098 43708 10108 43764
rect 10164 43708 10556 43764
rect 10612 43708 11340 43764
rect 11396 43708 13580 43764
rect 13636 43708 13646 43764
rect 17042 43708 17052 43764
rect 17108 43708 17836 43764
rect 17892 43708 18284 43764
rect 18340 43708 22428 43764
rect 22484 43708 22494 43764
rect 23548 43708 29820 43764
rect 29876 43708 29886 43764
rect 30146 43708 30156 43764
rect 30212 43708 30828 43764
rect 30884 43708 30894 43764
rect 32946 43708 32956 43764
rect 33012 43708 33124 43764
rect 36194 43708 36204 43764
rect 36260 43708 41804 43764
rect 41860 43708 41870 43764
rect 10322 43596 10332 43652
rect 10388 43596 16044 43652
rect 16100 43596 16110 43652
rect 17052 43540 17108 43708
rect 23548 43652 23604 43708
rect 21298 43596 21308 43652
rect 21364 43596 23548 43652
rect 23604 43596 23614 43652
rect 29362 43596 29372 43652
rect 29428 43596 30044 43652
rect 30100 43596 30940 43652
rect 30996 43596 31006 43652
rect 13906 43484 13916 43540
rect 13972 43484 14812 43540
rect 14868 43484 17108 43540
rect 20626 43484 20636 43540
rect 20692 43484 21420 43540
rect 21476 43484 21644 43540
rect 21700 43484 21710 43540
rect 27346 43484 27356 43540
rect 27412 43484 28028 43540
rect 28084 43484 30380 43540
rect 30436 43484 30716 43540
rect 30772 43484 32172 43540
rect 32228 43484 32238 43540
rect 33068 43428 33124 43708
rect 35410 43596 35420 43652
rect 35476 43596 35868 43652
rect 35924 43596 35934 43652
rect 36306 43596 36316 43652
rect 36372 43596 38220 43652
rect 38276 43596 38286 43652
rect 40114 43596 40124 43652
rect 40180 43596 41020 43652
rect 41076 43596 41086 43652
rect 43586 43596 43596 43652
rect 43652 43596 44268 43652
rect 44324 43596 44334 43652
rect 35522 43484 35532 43540
rect 35588 43484 37212 43540
rect 37268 43484 38332 43540
rect 38388 43484 38398 43540
rect 4498 43372 4508 43428
rect 4564 43372 4956 43428
rect 5012 43372 5022 43428
rect 10434 43372 10444 43428
rect 10500 43372 10892 43428
rect 10948 43372 15148 43428
rect 16594 43372 16604 43428
rect 16660 43372 17612 43428
rect 17668 43372 18956 43428
rect 19012 43372 19628 43428
rect 19684 43372 20076 43428
rect 20132 43372 20142 43428
rect 23986 43372 23996 43428
rect 24052 43372 25340 43428
rect 25396 43372 27020 43428
rect 27076 43372 27244 43428
rect 27300 43372 28252 43428
rect 28308 43372 29260 43428
rect 29316 43372 29326 43428
rect 31154 43372 31164 43428
rect 31220 43372 31836 43428
rect 31892 43372 33124 43428
rect 4022 43148 4060 43204
rect 4116 43148 4126 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 15092 43092 15148 43372
rect 16604 43092 16660 43372
rect 33926 43260 33964 43316
rect 34020 43260 34030 43316
rect 19170 43148 19180 43204
rect 19236 43148 23436 43204
rect 23492 43148 23502 43204
rect 31154 43148 31164 43204
rect 31220 43148 31724 43204
rect 31780 43148 31790 43204
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 6402 43036 6412 43092
rect 6468 43036 7196 43092
rect 7252 43036 13468 43092
rect 13524 43036 13534 43092
rect 15092 43036 16660 43092
rect 31490 43036 31500 43092
rect 31556 43036 33180 43092
rect 33236 43036 33246 43092
rect 7746 42924 7756 42980
rect 7812 42924 9212 42980
rect 9268 42924 9278 42980
rect 10322 42924 10332 42980
rect 10388 42924 10780 42980
rect 10836 42924 10846 42980
rect 29810 42924 29820 42980
rect 29876 42924 32060 42980
rect 32116 42924 32126 42980
rect 4162 42812 4172 42868
rect 4228 42812 4238 42868
rect 6738 42812 6748 42868
rect 6804 42812 8540 42868
rect 8596 42812 8606 42868
rect 10658 42812 10668 42868
rect 10724 42812 10734 42868
rect 31266 42812 31276 42868
rect 31332 42812 35196 42868
rect 35252 42812 35262 42868
rect 4172 42756 4228 42812
rect 3948 42700 4228 42756
rect 6178 42700 6188 42756
rect 6244 42700 7420 42756
rect 7476 42700 7486 42756
rect 3948 42644 4004 42700
rect 2370 42588 2380 42644
rect 2436 42588 2940 42644
rect 2996 42588 3006 42644
rect 3938 42588 3948 42644
rect 4004 42588 4014 42644
rect 4162 42588 4172 42644
rect 4228 42588 8428 42644
rect 8484 42588 8494 42644
rect 10668 42532 10724 42812
rect 19282 42700 19292 42756
rect 19348 42700 21532 42756
rect 21588 42700 21598 42756
rect 31826 42700 31836 42756
rect 31892 42700 36764 42756
rect 36820 42700 37548 42756
rect 37604 42700 37614 42756
rect 16818 42588 16828 42644
rect 16884 42588 17500 42644
rect 17556 42588 19404 42644
rect 19460 42588 19470 42644
rect 33058 42588 33068 42644
rect 33124 42588 33516 42644
rect 33572 42588 33582 42644
rect 33954 42588 33964 42644
rect 34020 42588 37436 42644
rect 37492 42588 37502 42644
rect 7074 42476 7084 42532
rect 7140 42476 11228 42532
rect 11284 42476 11788 42532
rect 11844 42476 11854 42532
rect 12562 42476 12572 42532
rect 12628 42476 14476 42532
rect 14532 42476 16156 42532
rect 16212 42476 18060 42532
rect 18116 42476 19068 42532
rect 19124 42476 19134 42532
rect 20850 42476 20860 42532
rect 20916 42476 22316 42532
rect 22372 42476 22382 42532
rect 30034 42476 30044 42532
rect 30100 42476 30268 42532
rect 30324 42476 31500 42532
rect 31556 42476 31566 42532
rect 0 42420 400 42448
rect 33516 42420 33572 42588
rect 34738 42476 34748 42532
rect 34804 42476 38220 42532
rect 38276 42476 38286 42532
rect 0 42364 3388 42420
rect 3444 42364 3454 42420
rect 4022 42364 4060 42420
rect 4116 42364 4126 42420
rect 6514 42364 6524 42420
rect 6580 42364 8092 42420
rect 8148 42364 8158 42420
rect 10546 42364 10556 42420
rect 10612 42364 10622 42420
rect 29222 42364 29260 42420
rect 29316 42364 29326 42420
rect 33516 42364 34972 42420
rect 35028 42364 35038 42420
rect 0 42336 400 42364
rect 10556 42196 10612 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 23426 42252 23436 42308
rect 23492 42252 38668 42308
rect 38612 42196 38668 42252
rect 2482 42140 2492 42196
rect 2548 42140 3052 42196
rect 3108 42140 3118 42196
rect 3266 42140 3276 42196
rect 3332 42140 3342 42196
rect 8978 42140 8988 42196
rect 9044 42140 9660 42196
rect 9716 42140 9726 42196
rect 10556 42140 11004 42196
rect 11060 42140 11070 42196
rect 21410 42140 21420 42196
rect 21476 42140 22092 42196
rect 22148 42140 23324 42196
rect 23380 42140 23390 42196
rect 26002 42140 26012 42196
rect 26068 42140 28140 42196
rect 28196 42140 28206 42196
rect 28774 42140 28812 42196
rect 28868 42140 29708 42196
rect 29764 42140 30268 42196
rect 30324 42140 30334 42196
rect 31378 42140 31388 42196
rect 31444 42140 31948 42196
rect 32004 42140 33180 42196
rect 33236 42140 34860 42196
rect 34916 42140 34926 42196
rect 35634 42140 35644 42196
rect 35700 42140 35868 42196
rect 35924 42140 36988 42196
rect 37044 42140 37054 42196
rect 38612 42140 40124 42196
rect 40180 42140 40190 42196
rect 3276 42084 3332 42140
rect 1586 42028 1596 42084
rect 1652 42028 3332 42084
rect 4918 42028 4956 42084
rect 5012 42028 5022 42084
rect 23874 42028 23884 42084
rect 23940 42028 23950 42084
rect 2818 41916 2828 41972
rect 2884 41916 3612 41972
rect 3668 41916 3678 41972
rect 10098 41916 10108 41972
rect 10164 41916 12124 41972
rect 12180 41916 12684 41972
rect 12740 41916 12750 41972
rect 12898 41916 12908 41972
rect 12964 41916 14476 41972
rect 14532 41916 15372 41972
rect 15428 41916 15438 41972
rect 16146 41916 16156 41972
rect 16212 41916 17724 41972
rect 17780 41916 17790 41972
rect 6738 41804 6748 41860
rect 6804 41804 7532 41860
rect 7588 41804 7598 41860
rect 17154 41804 17164 41860
rect 17220 41804 18732 41860
rect 18788 41804 20636 41860
rect 20692 41804 20702 41860
rect 23884 41748 23940 42028
rect 26684 41860 26740 42140
rect 27122 42028 27132 42084
rect 27188 42028 28252 42084
rect 28308 42028 31444 42084
rect 32610 42028 32620 42084
rect 32676 42028 35980 42084
rect 36036 42028 36046 42084
rect 37314 42028 37324 42084
rect 37380 42028 38780 42084
rect 38836 42028 38846 42084
rect 31388 41972 31444 42028
rect 30034 41916 30044 41972
rect 30100 41916 30716 41972
rect 30772 41916 31164 41972
rect 31220 41916 31230 41972
rect 31388 41916 34300 41972
rect 34356 41916 34366 41972
rect 40226 41916 40236 41972
rect 40292 41916 41468 41972
rect 41524 41916 41534 41972
rect 42242 41916 42252 41972
rect 42308 41916 42812 41972
rect 42868 41916 42878 41972
rect 26684 41804 27020 41860
rect 27076 41804 27086 41860
rect 31490 41804 31500 41860
rect 31556 41804 33852 41860
rect 33908 41804 33918 41860
rect 41234 41804 41244 41860
rect 41300 41804 43372 41860
rect 43428 41804 43438 41860
rect 2930 41692 2940 41748
rect 2996 41692 7308 41748
rect 7364 41692 7374 41748
rect 18050 41692 18060 41748
rect 18116 41692 19180 41748
rect 19236 41692 19246 41748
rect 22642 41692 22652 41748
rect 22708 41692 34076 41748
rect 34132 41692 34142 41748
rect 40226 41692 40236 41748
rect 40292 41692 41692 41748
rect 41748 41692 41758 41748
rect 2034 41580 2044 41636
rect 2100 41580 2604 41636
rect 2660 41580 2670 41636
rect 20738 41580 20748 41636
rect 20804 41580 21420 41636
rect 21476 41580 22428 41636
rect 22484 41580 24668 41636
rect 24724 41580 24734 41636
rect 27570 41580 27580 41636
rect 27636 41580 33292 41636
rect 33348 41580 33358 41636
rect 33506 41580 33516 41636
rect 33572 41580 34524 41636
rect 34580 41580 34590 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 26852 41468 35028 41524
rect 35970 41468 35980 41524
rect 36036 41468 36092 41524
rect 36148 41468 39788 41524
rect 39844 41468 44604 41524
rect 44660 41468 45164 41524
rect 45220 41468 45230 41524
rect 26852 41412 26908 41468
rect 34972 41412 35028 41468
rect 3154 41356 3164 41412
rect 3220 41356 5068 41412
rect 5124 41356 5134 41412
rect 23874 41356 23884 41412
rect 23940 41356 26908 41412
rect 27458 41356 27468 41412
rect 27524 41356 27534 41412
rect 27794 41356 27804 41412
rect 27860 41356 28028 41412
rect 28084 41356 28252 41412
rect 28308 41356 28318 41412
rect 34972 41356 35532 41412
rect 35588 41356 37100 41412
rect 37156 41356 37166 41412
rect 3602 41244 3612 41300
rect 3668 41244 4620 41300
rect 4676 41244 4686 41300
rect 19954 41244 19964 41300
rect 20020 41244 21756 41300
rect 21812 41244 21822 41300
rect 24210 41244 24220 41300
rect 24276 41244 25788 41300
rect 25844 41244 25854 41300
rect 27468 41188 27524 41356
rect 29586 41244 29596 41300
rect 29652 41244 29932 41300
rect 29988 41244 29998 41300
rect 1810 41132 1820 41188
rect 1876 41132 3388 41188
rect 7634 41132 7644 41188
rect 7700 41132 11564 41188
rect 11620 41132 11630 41188
rect 12674 41132 12684 41188
rect 12740 41132 13580 41188
rect 13636 41132 14028 41188
rect 14084 41132 14094 41188
rect 26786 41132 26796 41188
rect 26852 41132 27524 41188
rect 29250 41132 29260 41188
rect 29316 41132 29326 41188
rect 33730 41132 33740 41188
rect 33796 41132 34636 41188
rect 34692 41132 34702 41188
rect 36306 41132 36316 41188
rect 36372 41132 38332 41188
rect 38388 41132 38398 41188
rect 3332 40964 3388 41132
rect 29260 40964 29316 41132
rect 32274 41020 32284 41076
rect 32340 41020 33068 41076
rect 33124 41020 33134 41076
rect 35522 41020 35532 41076
rect 35588 41020 36540 41076
rect 36596 41020 36606 41076
rect 37650 41020 37660 41076
rect 37716 41020 38668 41076
rect 38612 40964 38668 41020
rect 3332 40908 5068 40964
rect 5124 40908 8540 40964
rect 8596 40908 8606 40964
rect 10658 40908 10668 40964
rect 10724 40908 11340 40964
rect 11396 40908 12236 40964
rect 12292 40908 12302 40964
rect 24882 40908 24892 40964
rect 24948 40908 26012 40964
rect 26068 40908 26078 40964
rect 28914 40908 28924 40964
rect 28980 40908 29820 40964
rect 29876 40908 29886 40964
rect 30146 40908 30156 40964
rect 30212 40908 30828 40964
rect 30884 40908 31276 40964
rect 31332 40908 31342 40964
rect 34514 40908 34524 40964
rect 34580 40908 35084 40964
rect 35140 40908 35150 40964
rect 38612 40908 40908 40964
rect 40964 40908 40974 40964
rect 44258 40908 44268 40964
rect 44324 40908 44940 40964
rect 44996 40908 45006 40964
rect 26450 40796 26460 40852
rect 26516 40796 28924 40852
rect 28980 40796 28990 40852
rect 29222 40796 29260 40852
rect 29316 40796 29326 40852
rect 36306 40796 36316 40852
rect 36372 40796 38556 40852
rect 38612 40796 38622 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 3332 40684 5628 40740
rect 5684 40684 7084 40740
rect 7140 40684 7150 40740
rect 23492 40684 24668 40740
rect 24724 40684 26908 40740
rect 26964 40684 28028 40740
rect 28084 40684 29820 40740
rect 29876 40684 32060 40740
rect 32116 40684 32126 40740
rect 34850 40684 34860 40740
rect 34916 40684 36764 40740
rect 36820 40684 41020 40740
rect 41076 40684 41692 40740
rect 41748 40684 42812 40740
rect 42868 40684 42878 40740
rect 3332 40628 3388 40684
rect 23492 40628 23548 40684
rect 2594 40572 2604 40628
rect 2660 40572 2828 40628
rect 2884 40572 3388 40628
rect 3714 40572 3724 40628
rect 3780 40572 7868 40628
rect 7924 40572 7934 40628
rect 18386 40572 18396 40628
rect 18452 40572 23548 40628
rect 26852 40572 27804 40628
rect 27860 40572 27870 40628
rect 28466 40572 28476 40628
rect 28532 40572 33964 40628
rect 34020 40572 34030 40628
rect 38882 40572 38892 40628
rect 38948 40572 39676 40628
rect 39732 40572 39742 40628
rect 40786 40572 40796 40628
rect 40852 40572 43596 40628
rect 43652 40572 43662 40628
rect 26852 40516 26908 40572
rect 2594 40460 2604 40516
rect 2660 40460 3612 40516
rect 3668 40460 3678 40516
rect 7746 40460 7756 40516
rect 7812 40460 10052 40516
rect 13570 40460 13580 40516
rect 13636 40460 17500 40516
rect 17556 40460 17566 40516
rect 18722 40460 18732 40516
rect 18788 40460 19292 40516
rect 19348 40460 20524 40516
rect 20580 40460 26908 40516
rect 27458 40460 27468 40516
rect 27524 40460 28140 40516
rect 28196 40460 31948 40516
rect 32004 40460 32014 40516
rect 33618 40460 33628 40516
rect 33684 40460 33908 40516
rect 35858 40460 35868 40516
rect 35924 40460 38332 40516
rect 38388 40460 41244 40516
rect 41300 40460 42140 40516
rect 42196 40460 42206 40516
rect 9996 40404 10052 40460
rect 33852 40404 33908 40460
rect 2454 40348 2492 40404
rect 2548 40348 2558 40404
rect 8306 40348 8316 40404
rect 8372 40292 8428 40404
rect 9986 40348 9996 40404
rect 10052 40348 11004 40404
rect 11060 40348 11070 40404
rect 14018 40348 14028 40404
rect 14084 40348 16156 40404
rect 16212 40348 16222 40404
rect 18162 40348 18172 40404
rect 18228 40348 18844 40404
rect 18900 40348 19964 40404
rect 20020 40348 20030 40404
rect 27346 40348 27356 40404
rect 27412 40348 28252 40404
rect 28308 40348 30156 40404
rect 30212 40348 30716 40404
rect 30772 40348 32284 40404
rect 32340 40348 32350 40404
rect 33842 40348 33852 40404
rect 33908 40348 33918 40404
rect 39442 40348 39452 40404
rect 39508 40348 40684 40404
rect 40740 40348 40750 40404
rect 41458 40348 41468 40404
rect 41524 40348 42252 40404
rect 42308 40348 42318 40404
rect 43260 40348 43596 40404
rect 43652 40348 43662 40404
rect 43260 40292 43316 40348
rect 2594 40236 2604 40292
rect 2660 40236 3388 40292
rect 3444 40236 3454 40292
rect 8372 40236 10108 40292
rect 10164 40236 10174 40292
rect 14466 40236 14476 40292
rect 14532 40236 14924 40292
rect 14980 40236 37772 40292
rect 37828 40236 40348 40292
rect 40404 40236 40414 40292
rect 43250 40236 43260 40292
rect 43316 40236 43326 40292
rect 19170 40124 19180 40180
rect 19236 40124 23212 40180
rect 23268 40124 32172 40180
rect 32228 40124 32238 40180
rect 36418 40124 36428 40180
rect 36484 40124 36764 40180
rect 36820 40124 36830 40180
rect 28886 40012 28924 40068
rect 28980 40012 28990 40068
rect 29558 40012 29596 40068
rect 29652 40012 29662 40068
rect 29810 40012 29820 40068
rect 29876 40012 30940 40068
rect 30996 40012 31006 40068
rect 33506 40012 33516 40068
rect 33572 40012 33582 40068
rect 34290 40012 34300 40068
rect 34356 40012 34748 40068
rect 34804 40012 34814 40068
rect 40338 40012 40348 40068
rect 40404 40012 42028 40068
rect 42084 40012 42094 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 33516 39956 33572 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 33516 39900 34188 39956
rect 34244 39900 34254 39956
rect 35532 39900 41356 39956
rect 41412 39900 41422 39956
rect 35532 39844 35588 39900
rect 3826 39788 3836 39844
rect 3892 39788 4508 39844
rect 4564 39788 5180 39844
rect 5236 39788 5246 39844
rect 30146 39788 30156 39844
rect 30212 39788 30604 39844
rect 30660 39788 35588 39844
rect 37538 39788 37548 39844
rect 37604 39788 38332 39844
rect 38388 39788 40796 39844
rect 40852 39788 41244 39844
rect 41300 39788 41310 39844
rect 2818 39676 2828 39732
rect 2884 39676 3052 39732
rect 3108 39676 3500 39732
rect 3556 39676 5124 39732
rect 5282 39676 5292 39732
rect 5348 39676 5852 39732
rect 5908 39676 5918 39732
rect 17938 39676 17948 39732
rect 18004 39676 18956 39732
rect 19012 39676 19022 39732
rect 28578 39676 28588 39732
rect 28644 39676 29484 39732
rect 29540 39676 29550 39732
rect 34066 39676 34076 39732
rect 34132 39676 35196 39732
rect 35252 39676 37100 39732
rect 37156 39676 37166 39732
rect 38882 39676 38892 39732
rect 38948 39676 39340 39732
rect 39396 39676 39406 39732
rect 5068 39620 5124 39676
rect 3266 39564 3276 39620
rect 3332 39564 4844 39620
rect 4900 39564 4910 39620
rect 5068 39564 9996 39620
rect 10052 39564 10332 39620
rect 10388 39564 10398 39620
rect 13906 39564 13916 39620
rect 13972 39564 14812 39620
rect 14868 39564 16268 39620
rect 16324 39564 16334 39620
rect 20850 39564 20860 39620
rect 20916 39564 21980 39620
rect 22036 39564 23436 39620
rect 23492 39564 25060 39620
rect 26114 39564 26124 39620
rect 26180 39564 27244 39620
rect 27300 39564 27310 39620
rect 30146 39564 30156 39620
rect 30212 39564 31276 39620
rect 31332 39564 31342 39620
rect 40002 39564 40012 39620
rect 40068 39564 42588 39620
rect 42644 39564 46396 39620
rect 46452 39564 46462 39620
rect 14690 39452 14700 39508
rect 14756 39452 15372 39508
rect 15428 39452 15438 39508
rect 23538 39452 23548 39508
rect 23604 39452 23996 39508
rect 24052 39452 24220 39508
rect 24276 39452 24286 39508
rect 25004 39396 25060 39564
rect 26226 39452 26236 39508
rect 26292 39452 26908 39508
rect 26964 39452 26974 39508
rect 27542 39452 27580 39508
rect 27636 39452 27646 39508
rect 32498 39452 32508 39508
rect 32564 39452 33964 39508
rect 34020 39452 34030 39508
rect 2706 39340 2716 39396
rect 2772 39340 3276 39396
rect 3332 39340 4172 39396
rect 4228 39340 4238 39396
rect 23650 39340 23660 39396
rect 23716 39340 24780 39396
rect 24836 39340 24846 39396
rect 25004 39340 28588 39396
rect 28644 39340 28654 39396
rect 29586 39340 29596 39396
rect 29652 39340 30044 39396
rect 30100 39340 30110 39396
rect 32162 39340 32172 39396
rect 32228 39340 33180 39396
rect 33236 39340 33246 39396
rect 33730 39340 33740 39396
rect 33796 39340 34972 39396
rect 35028 39340 35038 39396
rect 39442 39340 39452 39396
rect 39508 39340 41132 39396
rect 41188 39340 42364 39396
rect 42420 39340 42430 39396
rect 33180 39284 33236 39340
rect 33180 39228 40124 39284
rect 40180 39228 40684 39284
rect 40740 39228 40750 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 4274 39116 4284 39172
rect 4340 39116 6076 39172
rect 6132 39116 10668 39172
rect 10724 39116 10734 39172
rect 20402 39116 20412 39172
rect 20468 39116 21308 39172
rect 21364 39116 21374 39172
rect 26422 39116 26460 39172
rect 26516 39116 26526 39172
rect 29922 39116 29932 39172
rect 29988 39116 31948 39172
rect 32004 39116 33068 39172
rect 33124 39116 33134 39172
rect 34290 39116 34300 39172
rect 34356 39116 36652 39172
rect 36708 39116 38444 39172
rect 38500 39116 38510 39172
rect 9986 39004 9996 39060
rect 10052 39004 10556 39060
rect 10612 39004 10622 39060
rect 20178 39004 20188 39060
rect 20244 39004 21084 39060
rect 21140 39004 21150 39060
rect 24770 39004 24780 39060
rect 24836 39004 26908 39060
rect 33618 39004 33628 39060
rect 33684 39004 34636 39060
rect 34692 39004 34702 39060
rect 39666 39004 39676 39060
rect 39732 39004 41468 39060
rect 41524 39004 41916 39060
rect 41972 39004 41982 39060
rect 26852 38948 26908 39004
rect 39676 38948 39732 39004
rect 19282 38892 19292 38948
rect 19348 38892 19964 38948
rect 20020 38892 21420 38948
rect 21476 38892 21486 38948
rect 26852 38892 39340 38948
rect 39396 38892 39732 38948
rect 9650 38780 9660 38836
rect 9716 38780 10332 38836
rect 10388 38780 12124 38836
rect 12180 38780 12190 38836
rect 16594 38780 16604 38836
rect 16660 38780 17948 38836
rect 18004 38780 19068 38836
rect 19124 38780 19134 38836
rect 21634 38780 21644 38836
rect 21700 38780 26460 38836
rect 26516 38780 26526 38836
rect 27346 38780 27356 38836
rect 27412 38780 28028 38836
rect 28084 38780 28094 38836
rect 29250 38780 29260 38836
rect 29316 38780 29932 38836
rect 29988 38780 29998 38836
rect 38434 38780 38444 38836
rect 38500 38780 38892 38836
rect 38948 38780 38958 38836
rect 39218 38780 39228 38836
rect 39284 38780 39788 38836
rect 39844 38780 41468 38836
rect 41524 38780 41534 38836
rect 8082 38668 8092 38724
rect 8148 38668 10444 38724
rect 10500 38668 13692 38724
rect 13748 38668 13758 38724
rect 32284 38668 32508 38724
rect 32564 38668 32574 38724
rect 2594 38556 2604 38612
rect 2660 38556 2716 38612
rect 2772 38556 4732 38612
rect 4788 38556 4798 38612
rect 5170 38556 5180 38612
rect 5236 38556 5740 38612
rect 5796 38556 6300 38612
rect 6356 38556 6366 38612
rect 20626 38556 20636 38612
rect 20692 38556 21532 38612
rect 21588 38556 21598 38612
rect 28242 38556 28252 38612
rect 28308 38556 30716 38612
rect 30772 38556 30782 38612
rect 32284 38500 32340 38668
rect 34402 38556 34412 38612
rect 34468 38556 35868 38612
rect 35924 38556 35934 38612
rect 37426 38556 37436 38612
rect 37492 38556 38108 38612
rect 38164 38556 38174 38612
rect 41346 38556 41356 38612
rect 41412 38556 42140 38612
rect 42196 38556 43148 38612
rect 43204 38556 43214 38612
rect 44146 38556 44156 38612
rect 44212 38556 45836 38612
rect 45892 38556 45902 38612
rect 25442 38444 25452 38500
rect 25508 38444 26908 38500
rect 27346 38444 27356 38500
rect 27412 38444 28364 38500
rect 28420 38444 28430 38500
rect 32274 38444 32284 38500
rect 32340 38444 32350 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 26852 38388 26908 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 26852 38332 32508 38388
rect 32564 38332 32574 38388
rect 42914 38332 42924 38388
rect 42980 38332 44156 38388
rect 44212 38332 44222 38388
rect 2258 38220 2268 38276
rect 2324 38220 5852 38276
rect 5908 38220 5918 38276
rect 6290 38220 6300 38276
rect 6356 38220 7532 38276
rect 7588 38220 7598 38276
rect 28914 38220 28924 38276
rect 28980 38220 29260 38276
rect 29316 38220 29326 38276
rect 30454 38220 30492 38276
rect 30548 38220 30558 38276
rect 43474 38220 43484 38276
rect 43540 38220 43820 38276
rect 43876 38220 43886 38276
rect 26786 38108 26796 38164
rect 26852 38108 27244 38164
rect 27300 38108 27310 38164
rect 27794 38108 27804 38164
rect 27860 38108 29372 38164
rect 29428 38108 29708 38164
rect 29764 38108 29774 38164
rect 35858 38108 35868 38164
rect 35924 38108 37996 38164
rect 38052 38108 38062 38164
rect 1810 37996 1820 38052
rect 1876 37996 2492 38052
rect 2548 37996 2558 38052
rect 2818 37996 2828 38052
rect 2884 37996 3500 38052
rect 3556 37996 3566 38052
rect 4386 37996 4396 38052
rect 4452 37996 4956 38052
rect 5012 37996 5022 38052
rect 7186 37996 7196 38052
rect 7252 37996 7644 38052
rect 7700 37996 7710 38052
rect 7868 37996 8428 38052
rect 8484 37996 9436 38052
rect 9492 37996 9502 38052
rect 10322 37996 10332 38052
rect 10388 37996 11116 38052
rect 11172 37996 12908 38052
rect 12964 37996 13580 38052
rect 13636 37996 13646 38052
rect 14690 37996 14700 38052
rect 14756 37996 15372 38052
rect 15428 37996 15438 38052
rect 28914 37996 28924 38052
rect 28980 37996 29036 38052
rect 29092 37996 29102 38052
rect 32050 37996 32060 38052
rect 32116 37996 33292 38052
rect 33348 37996 33358 38052
rect 35634 37996 35644 38052
rect 35700 37996 36092 38052
rect 36148 37996 36764 38052
rect 36820 37996 36830 38052
rect 7868 37940 7924 37996
rect 2146 37884 2156 37940
rect 2212 37884 4620 37940
rect 4676 37884 4686 37940
rect 7522 37884 7532 37940
rect 7588 37884 7924 37940
rect 26562 37884 26572 37940
rect 26628 37884 27244 37940
rect 27300 37884 28252 37940
rect 28308 37884 28318 37940
rect 31266 37884 31276 37940
rect 31332 37884 31948 37940
rect 32004 37884 33740 37940
rect 33796 37884 33806 37940
rect 34262 37884 34300 37940
rect 34356 37884 34366 37940
rect 36418 37884 36428 37940
rect 36484 37884 37212 37940
rect 37268 37884 37278 37940
rect 43652 37884 44044 37940
rect 44100 37884 44110 37940
rect 11554 37772 11564 37828
rect 11620 37772 12460 37828
rect 12516 37772 12526 37828
rect 22530 37772 22540 37828
rect 22596 37772 27356 37828
rect 27412 37772 27422 37828
rect 30678 37772 30716 37828
rect 30772 37772 30782 37828
rect 42690 37772 42700 37828
rect 42756 37772 43372 37828
rect 43428 37772 43438 37828
rect 43652 37716 43708 37884
rect 23492 37660 27244 37716
rect 27300 37660 27310 37716
rect 43138 37660 43148 37716
rect 43204 37660 43708 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 3238 37548 3276 37604
rect 3332 37548 3342 37604
rect 7298 37548 7308 37604
rect 7364 37548 9548 37604
rect 9604 37548 9614 37604
rect 0 37492 400 37520
rect 23492 37492 23548 37660
rect 0 37436 1932 37492
rect 1988 37436 1998 37492
rect 4274 37436 4284 37492
rect 4340 37436 5180 37492
rect 5236 37436 9884 37492
rect 9940 37436 11004 37492
rect 11060 37436 11070 37492
rect 21186 37436 21196 37492
rect 21252 37436 21532 37492
rect 21588 37436 23548 37492
rect 26852 37548 28812 37604
rect 28868 37548 28878 37604
rect 0 37408 400 37436
rect 26852 37380 26908 37548
rect 27010 37436 27020 37492
rect 27076 37436 28476 37492
rect 28532 37436 28542 37492
rect 29474 37436 29484 37492
rect 29540 37436 30604 37492
rect 30660 37436 32732 37492
rect 32788 37436 32798 37492
rect 33954 37436 33964 37492
rect 34020 37436 41580 37492
rect 41636 37436 41646 37492
rect 2258 37324 2268 37380
rect 2324 37324 2940 37380
rect 2996 37324 3724 37380
rect 3780 37324 4396 37380
rect 4452 37324 4462 37380
rect 8530 37324 8540 37380
rect 8596 37324 9772 37380
rect 9828 37324 9838 37380
rect 16818 37324 16828 37380
rect 16884 37324 19180 37380
rect 19236 37324 19246 37380
rect 25554 37324 25564 37380
rect 25620 37324 26908 37380
rect 27346 37324 27356 37380
rect 27412 37324 28588 37380
rect 28644 37324 31836 37380
rect 31892 37324 33628 37380
rect 33684 37324 33694 37380
rect 8194 37212 8204 37268
rect 8260 37212 10556 37268
rect 10612 37212 10622 37268
rect 24434 37212 24444 37268
rect 24500 37212 25844 37268
rect 27570 37212 27580 37268
rect 27636 37212 29820 37268
rect 29876 37212 29886 37268
rect 31378 37212 31388 37268
rect 31444 37212 31948 37268
rect 32004 37212 32014 37268
rect 33730 37212 33740 37268
rect 33796 37212 34524 37268
rect 34580 37212 34590 37268
rect 34962 37212 34972 37268
rect 35028 37212 36204 37268
rect 36260 37212 37660 37268
rect 37716 37212 37726 37268
rect 25788 37156 25844 37212
rect 6178 37100 6188 37156
rect 6244 37100 7532 37156
rect 7588 37100 7598 37156
rect 14354 37100 14364 37156
rect 14420 37100 15036 37156
rect 15092 37100 15102 37156
rect 16706 37100 16716 37156
rect 16772 37100 21756 37156
rect 21812 37100 25564 37156
rect 25620 37100 25630 37156
rect 25788 37100 28812 37156
rect 28868 37100 28878 37156
rect 30930 37100 30940 37156
rect 30996 37100 31612 37156
rect 31668 37100 31678 37156
rect 34738 37100 34748 37156
rect 34804 37100 37212 37156
rect 37268 37100 37278 37156
rect 38098 37100 38108 37156
rect 38164 37100 40908 37156
rect 40964 37100 45276 37156
rect 45332 37100 45342 37156
rect 2482 36988 2492 37044
rect 2548 36988 2558 37044
rect 3378 36988 3388 37044
rect 3444 36988 3556 37044
rect 6850 36988 6860 37044
rect 6916 36988 8204 37044
rect 8260 36988 8652 37044
rect 8708 36988 8718 37044
rect 12898 36988 12908 37044
rect 12964 36988 13412 37044
rect 16482 36988 16492 37044
rect 16548 36988 16828 37044
rect 16884 36988 16894 37044
rect 27458 36988 27468 37044
rect 27524 36988 27580 37044
rect 27636 36988 27646 37044
rect 32050 36988 32060 37044
rect 32116 36988 32956 37044
rect 33012 36988 34188 37044
rect 34244 36988 34254 37044
rect 34850 36988 34860 37044
rect 34916 36988 45612 37044
rect 45668 36988 45678 37044
rect 2492 36932 2548 36988
rect 2492 36876 3388 36932
rect 2258 36764 2268 36820
rect 2324 36764 3164 36820
rect 3220 36764 3230 36820
rect 3332 36708 3388 36876
rect 3500 36820 3556 36988
rect 13356 36932 13412 36988
rect 13356 36876 14700 36932
rect 14756 36876 14766 36932
rect 18946 36876 18956 36932
rect 19012 36876 19740 36932
rect 19796 36876 19806 36932
rect 25890 36876 25900 36932
rect 25956 36876 26348 36932
rect 26404 36876 26414 36932
rect 37202 36876 37212 36932
rect 37268 36876 44268 36932
rect 44324 36876 44334 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 3500 36764 4284 36820
rect 4340 36764 4350 36820
rect 19058 36764 19068 36820
rect 19124 36764 20748 36820
rect 20804 36764 27916 36820
rect 27972 36764 27982 36820
rect 29922 36764 29932 36820
rect 29988 36764 32620 36820
rect 32676 36764 32686 36820
rect 3332 36652 4060 36708
rect 4116 36652 4126 36708
rect 5954 36652 5964 36708
rect 6020 36652 6748 36708
rect 6804 36652 6814 36708
rect 8866 36652 8876 36708
rect 8932 36652 9996 36708
rect 10052 36652 10062 36708
rect 26450 36652 26460 36708
rect 26516 36652 27804 36708
rect 27860 36652 27870 36708
rect 28578 36652 28588 36708
rect 28644 36652 30156 36708
rect 30212 36652 30222 36708
rect 34626 36652 34636 36708
rect 34692 36652 35308 36708
rect 35364 36652 36988 36708
rect 37044 36652 37054 36708
rect 4834 36540 4844 36596
rect 4900 36540 5516 36596
rect 5572 36540 5582 36596
rect 5730 36540 5740 36596
rect 5796 36540 6188 36596
rect 6244 36540 6254 36596
rect 26114 36540 26124 36596
rect 26180 36540 26908 36596
rect 26964 36540 26974 36596
rect 31714 36540 31724 36596
rect 31780 36540 32284 36596
rect 32340 36540 32350 36596
rect 37986 36540 37996 36596
rect 38052 36540 38062 36596
rect 41346 36540 41356 36596
rect 41412 36540 42364 36596
rect 42420 36540 48076 36596
rect 48132 36540 48142 36596
rect 3332 36428 3612 36484
rect 3668 36428 3678 36484
rect 3826 36428 3836 36484
rect 3892 36428 6524 36484
rect 6580 36428 6748 36484
rect 6804 36428 6814 36484
rect 14690 36428 14700 36484
rect 14756 36428 15932 36484
rect 15988 36428 15998 36484
rect 25778 36428 25788 36484
rect 25844 36428 26460 36484
rect 26516 36428 26526 36484
rect 28242 36428 28252 36484
rect 28308 36428 29820 36484
rect 29876 36428 29886 36484
rect 30146 36428 30156 36484
rect 30212 36428 36092 36484
rect 36148 36428 36158 36484
rect 3332 36372 3388 36428
rect 1922 36316 1932 36372
rect 1988 36316 2604 36372
rect 2660 36316 3388 36372
rect 6188 36260 6244 36428
rect 37996 36372 38052 36540
rect 38294 36428 38332 36484
rect 38388 36428 38398 36484
rect 7186 36316 7196 36372
rect 7252 36316 7532 36372
rect 7588 36316 7598 36372
rect 25106 36316 25116 36372
rect 25172 36316 25900 36372
rect 25956 36316 25966 36372
rect 26114 36316 26124 36372
rect 26180 36316 26572 36372
rect 26628 36316 26638 36372
rect 30790 36316 30828 36372
rect 30884 36316 30894 36372
rect 31042 36316 31052 36372
rect 31108 36316 31612 36372
rect 31668 36316 31678 36372
rect 37986 36316 37996 36372
rect 38052 36316 38062 36372
rect 2034 36204 2044 36260
rect 2100 36204 2492 36260
rect 2548 36204 2558 36260
rect 6178 36204 6188 36260
rect 6244 36204 6254 36260
rect 20066 36204 20076 36260
rect 20132 36204 21252 36260
rect 21410 36204 21420 36260
rect 21476 36204 23548 36260
rect 23604 36204 24668 36260
rect 24724 36204 24734 36260
rect 27346 36204 27356 36260
rect 27412 36204 28364 36260
rect 28420 36204 28430 36260
rect 34738 36204 34748 36260
rect 34804 36204 35532 36260
rect 35588 36204 35598 36260
rect 37762 36204 37772 36260
rect 37828 36204 38108 36260
rect 38164 36204 38174 36260
rect 21196 36148 21252 36204
rect 21196 36092 25788 36148
rect 25844 36092 25854 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 26226 35980 26236 36036
rect 26292 35980 26460 36036
rect 26516 35980 26526 36036
rect 27906 35980 27916 36036
rect 27972 35980 28140 36036
rect 28196 35980 33404 36036
rect 33460 35980 33470 36036
rect 2482 35868 2492 35924
rect 2548 35868 3500 35924
rect 3556 35868 3566 35924
rect 6962 35868 6972 35924
rect 7028 35868 7420 35924
rect 7476 35868 7486 35924
rect 10210 35868 10220 35924
rect 10276 35868 11004 35924
rect 11060 35868 12684 35924
rect 12740 35868 12750 35924
rect 30034 35868 30044 35924
rect 30100 35868 30940 35924
rect 30996 35868 31388 35924
rect 31444 35868 31454 35924
rect 11442 35756 11452 35812
rect 11508 35756 12908 35812
rect 12964 35756 18172 35812
rect 18228 35756 27020 35812
rect 27076 35756 29596 35812
rect 29652 35756 30716 35812
rect 30772 35756 30782 35812
rect 32722 35756 32732 35812
rect 32788 35756 34188 35812
rect 34244 35756 35252 35812
rect 12674 35644 12684 35700
rect 12740 35644 18060 35700
rect 18116 35644 18126 35700
rect 15250 35532 15260 35588
rect 15316 35532 16380 35588
rect 16436 35532 17836 35588
rect 17892 35532 17902 35588
rect 18386 35532 18396 35588
rect 18452 35532 19964 35588
rect 20020 35532 20412 35588
rect 20468 35532 21644 35588
rect 21700 35532 25900 35588
rect 25956 35532 25966 35588
rect 30716 35476 30772 35756
rect 35196 35700 35252 35756
rect 30930 35644 30940 35700
rect 30996 35644 33068 35700
rect 33124 35644 33134 35700
rect 35186 35644 35196 35700
rect 35252 35644 42028 35700
rect 42084 35644 43484 35700
rect 43540 35644 43550 35700
rect 31724 35532 32508 35588
rect 32564 35532 32574 35588
rect 35634 35532 35644 35588
rect 35700 35532 36652 35588
rect 36708 35532 37212 35588
rect 37268 35532 37278 35588
rect 31724 35476 31780 35532
rect 30716 35420 30940 35476
rect 30996 35420 31006 35476
rect 31154 35420 31164 35476
rect 31220 35420 31724 35476
rect 31780 35420 31790 35476
rect 32834 35420 32844 35476
rect 32900 35420 33404 35476
rect 33460 35420 33470 35476
rect 33628 35420 34300 35476
rect 34356 35420 35084 35476
rect 35140 35420 36204 35476
rect 36260 35420 36270 35476
rect 33628 35364 33684 35420
rect 25778 35308 25788 35364
rect 25844 35308 26460 35364
rect 26516 35308 26526 35364
rect 30146 35308 30156 35364
rect 30212 35308 32508 35364
rect 32564 35308 32574 35364
rect 32844 35308 33684 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 32844 35252 32900 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 13570 35196 13580 35252
rect 13636 35196 16660 35252
rect 27234 35196 27244 35252
rect 27300 35196 32900 35252
rect 16604 35028 16660 35196
rect 17378 35084 17388 35140
rect 17444 35084 18508 35140
rect 18564 35084 18574 35140
rect 28914 35084 28924 35140
rect 28980 35084 29484 35140
rect 29540 35084 29550 35140
rect 34962 35084 34972 35140
rect 35028 35084 35196 35140
rect 35252 35084 35262 35140
rect 4946 34972 4956 35028
rect 5012 34972 5022 35028
rect 10882 34972 10892 35028
rect 10948 34972 12796 35028
rect 12852 34972 15932 35028
rect 15988 34972 15998 35028
rect 16604 34972 17948 35028
rect 18004 34972 19628 35028
rect 19684 34972 19694 35028
rect 34290 34972 34300 35028
rect 34356 34972 34366 35028
rect 4956 34804 5012 34972
rect 6598 34860 6636 34916
rect 6692 34860 6702 34916
rect 8194 34860 8204 34916
rect 8260 34860 8652 34916
rect 8708 34860 8718 34916
rect 9314 34860 9324 34916
rect 9380 34860 10780 34916
rect 10836 34860 10846 34916
rect 4162 34748 4172 34804
rect 4228 34748 5012 34804
rect 5618 34748 5628 34804
rect 5684 34748 6972 34804
rect 7028 34748 7038 34804
rect 10098 34748 10108 34804
rect 10164 34748 12068 34804
rect 12012 34692 12068 34748
rect 34300 34692 34356 34972
rect 36530 34860 36540 34916
rect 36596 34860 37212 34916
rect 37268 34860 37278 34916
rect 7186 34636 7196 34692
rect 7252 34636 7756 34692
rect 7812 34636 7822 34692
rect 8194 34636 8204 34692
rect 8260 34636 10556 34692
rect 10612 34636 10622 34692
rect 10770 34636 10780 34692
rect 10836 34636 11788 34692
rect 11844 34636 11854 34692
rect 12002 34636 12012 34692
rect 12068 34636 13580 34692
rect 13636 34636 13646 34692
rect 27906 34636 27916 34692
rect 27972 34636 29148 34692
rect 29204 34636 29214 34692
rect 29362 34636 29372 34692
rect 29428 34636 29932 34692
rect 29988 34636 31836 34692
rect 31892 34636 32060 34692
rect 32116 34636 32620 34692
rect 32676 34636 32686 34692
rect 34300 34636 34972 34692
rect 35028 34636 35038 34692
rect 29036 34524 29820 34580
rect 29876 34524 29886 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 29036 34468 29092 34524
rect 15922 34412 15932 34468
rect 15988 34412 15998 34468
rect 27010 34412 27020 34468
rect 27076 34412 29036 34468
rect 29092 34412 29102 34468
rect 33170 34412 33180 34468
rect 33236 34412 33246 34468
rect 3938 34300 3948 34356
rect 4004 34300 4014 34356
rect 3948 34244 4004 34300
rect 3602 34188 3612 34244
rect 3668 34188 4844 34244
rect 4900 34188 5628 34244
rect 5684 34188 5694 34244
rect 6290 34188 6300 34244
rect 6356 34188 6636 34244
rect 6692 34188 6702 34244
rect 15474 34188 15484 34244
rect 15540 34188 15708 34244
rect 15764 34188 15774 34244
rect 5628 34020 5684 34188
rect 8278 34076 8316 34132
rect 8372 34076 8382 34132
rect 15932 34020 15988 34412
rect 33180 34356 33236 34412
rect 27468 34300 29260 34356
rect 29316 34300 29326 34356
rect 33068 34300 33236 34356
rect 33618 34300 33628 34356
rect 33684 34300 34412 34356
rect 34468 34300 34478 34356
rect 39442 34300 39452 34356
rect 39508 34300 42700 34356
rect 42756 34300 43036 34356
rect 43092 34300 44268 34356
rect 44324 34300 44334 34356
rect 27468 34244 27524 34300
rect 19618 34188 19628 34244
rect 19684 34188 27468 34244
rect 27524 34188 27534 34244
rect 29138 34188 29148 34244
rect 29204 34188 30156 34244
rect 30212 34188 31052 34244
rect 31108 34188 31118 34244
rect 26852 34020 26908 34188
rect 29026 34076 29036 34132
rect 29092 34076 29708 34132
rect 29764 34076 29774 34132
rect 5628 33964 6076 34020
rect 6132 33964 7196 34020
rect 7252 33964 7980 34020
rect 8036 33964 8046 34020
rect 15932 33964 16380 34020
rect 16436 33964 16446 34020
rect 18498 33964 18508 34020
rect 18564 33964 21756 34020
rect 21812 33964 26012 34020
rect 26068 33964 26078 34020
rect 26852 33964 27020 34020
rect 27076 33964 27086 34020
rect 15810 33852 15820 33908
rect 15876 33852 17052 33908
rect 17108 33852 17118 33908
rect 19282 33852 19292 33908
rect 19348 33852 20636 33908
rect 20692 33852 21420 33908
rect 21476 33852 24556 33908
rect 24612 33852 24622 33908
rect 26674 33852 26684 33908
rect 26740 33852 27132 33908
rect 27188 33852 27198 33908
rect 33068 33796 33124 34300
rect 34738 34188 34748 34244
rect 34804 34188 35420 34244
rect 35476 34188 35486 34244
rect 33954 33964 33964 34020
rect 34020 33964 34300 34020
rect 34356 33964 34748 34020
rect 34804 33964 36540 34020
rect 36596 33964 36606 34020
rect 6962 33740 6972 33796
rect 7028 33740 7532 33796
rect 7588 33740 7598 33796
rect 18386 33740 18396 33796
rect 18452 33740 20748 33796
rect 20804 33740 21644 33796
rect 21700 33740 21710 33796
rect 29362 33740 29372 33796
rect 29428 33740 30380 33796
rect 30436 33740 33068 33796
rect 33124 33740 33134 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 6262 33628 6300 33684
rect 6356 33628 6366 33684
rect 16370 33628 16380 33684
rect 16436 33628 17612 33684
rect 17668 33628 19068 33684
rect 19124 33628 34636 33684
rect 34692 33628 34972 33684
rect 35028 33628 35038 33684
rect 44258 33628 44268 33684
rect 44324 33628 44828 33684
rect 44884 33628 44894 33684
rect 3938 33516 3948 33572
rect 4004 33516 4508 33572
rect 4564 33516 7084 33572
rect 7140 33516 7532 33572
rect 7588 33516 7598 33572
rect 27580 33516 30604 33572
rect 30660 33516 30670 33572
rect 32498 33516 32508 33572
rect 32564 33516 33292 33572
rect 33348 33516 33358 33572
rect 6300 33460 6356 33516
rect 6290 33404 6300 33460
rect 6356 33404 6366 33460
rect 6962 33404 6972 33460
rect 7028 33404 8092 33460
rect 8148 33404 8764 33460
rect 8820 33404 8830 33460
rect 26562 33404 26572 33460
rect 26628 33404 27412 33460
rect 1922 33292 1932 33348
rect 1988 33292 2492 33348
rect 2548 33292 4172 33348
rect 4228 33292 4238 33348
rect 19506 33292 19516 33348
rect 19572 33292 22764 33348
rect 22820 33292 24220 33348
rect 24276 33292 24286 33348
rect 24994 33292 25004 33348
rect 25060 33292 25564 33348
rect 25620 33292 25630 33348
rect 24220 33236 24276 33292
rect 27356 33236 27412 33404
rect 12002 33180 12012 33236
rect 12068 33180 13804 33236
rect 13860 33180 13870 33236
rect 24220 33180 26908 33236
rect 27346 33180 27356 33236
rect 27412 33180 27422 33236
rect 26852 33124 26908 33180
rect 27580 33124 27636 33516
rect 29474 33404 29484 33460
rect 29540 33404 30268 33460
rect 30324 33404 31836 33460
rect 31892 33404 31902 33460
rect 30594 33292 30604 33348
rect 30660 33292 33964 33348
rect 34020 33292 34030 33348
rect 36054 33180 36092 33236
rect 36148 33180 36158 33236
rect 26852 33068 27636 33124
rect 34290 33068 34300 33124
rect 34356 33068 38892 33124
rect 38948 33068 39228 33124
rect 39284 33068 42028 33124
rect 42084 33068 43036 33124
rect 43092 33068 43102 33124
rect 32610 32956 32620 33012
rect 32676 32956 33180 33012
rect 33236 32956 33246 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 26114 32844 26124 32900
rect 26180 32844 28252 32900
rect 28308 32844 28588 32900
rect 28644 32844 34636 32900
rect 34692 32844 34702 32900
rect 6738 32732 6748 32788
rect 6804 32732 7084 32788
rect 7140 32732 7150 32788
rect 32610 32732 32620 32788
rect 32676 32732 34412 32788
rect 34468 32732 34478 32788
rect 42466 32732 42476 32788
rect 42532 32732 43148 32788
rect 43204 32732 43214 32788
rect 8978 32620 8988 32676
rect 9044 32620 9772 32676
rect 9828 32620 9838 32676
rect 11106 32620 11116 32676
rect 11172 32620 12236 32676
rect 12292 32620 12302 32676
rect 28242 32620 28252 32676
rect 28308 32620 28588 32676
rect 28644 32620 28654 32676
rect 0 32564 400 32592
rect 0 32508 1708 32564
rect 1764 32508 1774 32564
rect 6514 32508 6524 32564
rect 6580 32508 7084 32564
rect 7140 32508 7150 32564
rect 9538 32508 9548 32564
rect 9604 32508 10444 32564
rect 10500 32508 10780 32564
rect 10836 32508 10846 32564
rect 15474 32508 15484 32564
rect 15540 32508 15820 32564
rect 15876 32508 15886 32564
rect 25890 32508 25900 32564
rect 25956 32508 26796 32564
rect 26852 32508 26862 32564
rect 29698 32508 29708 32564
rect 29764 32508 35532 32564
rect 35588 32508 35598 32564
rect 43026 32508 43036 32564
rect 43092 32508 44268 32564
rect 44324 32508 44334 32564
rect 0 32480 400 32508
rect 8194 32396 8204 32452
rect 8260 32396 11452 32452
rect 11508 32396 11518 32452
rect 14690 32396 14700 32452
rect 14756 32396 23548 32452
rect 23604 32396 24668 32452
rect 24724 32396 25228 32452
rect 25284 32396 31276 32452
rect 31332 32396 33404 32452
rect 33460 32396 34076 32452
rect 34132 32396 34300 32452
rect 34356 32396 34366 32452
rect 36418 32396 36428 32452
rect 36484 32396 39340 32452
rect 39396 32396 40908 32452
rect 40964 32396 40974 32452
rect 3938 32284 3948 32340
rect 4004 32284 4900 32340
rect 4844 32228 4900 32284
rect 4834 32172 4844 32228
rect 4900 32172 6972 32228
rect 7028 32172 7038 32228
rect 17490 32172 17500 32228
rect 17556 32172 17948 32228
rect 18004 32172 18732 32228
rect 18788 32172 19292 32228
rect 19348 32172 19358 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 6626 32060 6636 32116
rect 6692 32060 6702 32116
rect 27346 32060 27356 32116
rect 27412 32060 28812 32116
rect 28868 32060 28878 32116
rect 43586 32060 43596 32116
rect 43652 32060 45052 32116
rect 45108 32060 46284 32116
rect 46340 32060 46350 32116
rect 4610 31948 4620 32004
rect 4676 31948 5740 32004
rect 5796 31948 5806 32004
rect 6636 31892 6692 32060
rect 16818 31948 16828 32004
rect 16884 31948 18172 32004
rect 18228 31948 25004 32004
rect 25060 31948 25070 32004
rect 33590 31948 33628 32004
rect 33684 31948 33694 32004
rect 44258 31948 44268 32004
rect 44324 31948 44828 32004
rect 44884 31948 44894 32004
rect 3332 31836 4396 31892
rect 4452 31836 6692 31892
rect 18274 31836 18284 31892
rect 18340 31836 19516 31892
rect 19572 31836 19964 31892
rect 20020 31836 20030 31892
rect 26226 31836 26236 31892
rect 26292 31836 26684 31892
rect 26740 31836 26750 31892
rect 27682 31836 27692 31892
rect 27748 31836 29260 31892
rect 29316 31836 30156 31892
rect 30212 31836 35532 31892
rect 35588 31836 35598 31892
rect 46386 31836 46396 31892
rect 46452 31836 47740 31892
rect 47796 31836 47806 31892
rect 3266 31724 3276 31780
rect 3332 31724 3388 31836
rect 26114 31724 26124 31780
rect 26180 31724 28140 31780
rect 28196 31724 28206 31780
rect 31602 31724 31612 31780
rect 31668 31724 33740 31780
rect 33796 31724 33806 31780
rect 38070 31724 38108 31780
rect 38164 31724 38174 31780
rect 30930 31612 30940 31668
rect 30996 31612 32284 31668
rect 32340 31612 33628 31668
rect 33684 31612 37660 31668
rect 37716 31612 38892 31668
rect 38948 31612 41356 31668
rect 41412 31612 41804 31668
rect 41860 31612 41870 31668
rect 6290 31500 6300 31556
rect 6356 31500 6860 31556
rect 6916 31500 8204 31556
rect 8260 31500 8270 31556
rect 24546 31500 24556 31556
rect 24612 31500 25900 31556
rect 25956 31500 26572 31556
rect 26628 31500 29372 31556
rect 29428 31500 29438 31556
rect 32050 31500 32060 31556
rect 32116 31500 33180 31556
rect 33236 31500 34860 31556
rect 34916 31500 38052 31556
rect 38210 31500 38220 31556
rect 38276 31500 40124 31556
rect 40180 31500 40572 31556
rect 40628 31500 41916 31556
rect 41972 31500 41982 31556
rect 37996 31444 38052 31500
rect 31378 31388 31388 31444
rect 31444 31388 34188 31444
rect 34244 31388 34254 31444
rect 34934 31388 34972 31444
rect 35028 31388 35038 31444
rect 37996 31388 38108 31444
rect 38164 31388 38668 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 1922 31276 1932 31332
rect 1988 31276 3052 31332
rect 3108 31276 6188 31332
rect 6244 31276 6254 31332
rect 25554 31276 25564 31332
rect 25620 31276 26796 31332
rect 26852 31276 26862 31332
rect 28690 31276 28700 31332
rect 28756 31276 28766 31332
rect 28700 31220 28756 31276
rect 3154 31164 3164 31220
rect 3220 31164 5292 31220
rect 5348 31164 5516 31220
rect 5572 31164 5582 31220
rect 26852 31164 28756 31220
rect 30482 31164 30492 31220
rect 30548 31164 31052 31220
rect 31108 31164 31118 31220
rect 32274 31164 32284 31220
rect 32340 31164 32732 31220
rect 32788 31164 34076 31220
rect 34132 31164 34748 31220
rect 34804 31164 34814 31220
rect 38612 31164 38668 31388
rect 38724 31164 40796 31220
rect 40852 31164 41244 31220
rect 41300 31164 42028 31220
rect 42084 31164 43148 31220
rect 43204 31164 43214 31220
rect 4172 31052 5068 31108
rect 5124 31052 5134 31108
rect 4172 30996 4228 31052
rect 3378 30940 3388 30996
rect 3444 30940 4172 30996
rect 4228 30940 4238 30996
rect 4834 30940 4844 30996
rect 4900 30940 5740 30996
rect 5796 30940 7084 30996
rect 7140 30940 7150 30996
rect 14802 30940 14812 30996
rect 14868 30940 15260 30996
rect 15316 30940 15326 30996
rect 19618 30828 19628 30884
rect 19684 30828 25228 30884
rect 25284 30828 25294 30884
rect 26310 30828 26348 30884
rect 26404 30828 26414 30884
rect 7410 30716 7420 30772
rect 7476 30716 10556 30772
rect 10612 30716 12908 30772
rect 12964 30716 12974 30772
rect 26852 30660 26908 31164
rect 31826 31052 31836 31108
rect 31892 31052 33964 31108
rect 34020 31052 34300 31108
rect 34356 31052 34366 31108
rect 35858 31052 35868 31108
rect 35924 31052 37436 31108
rect 37492 31052 37502 31108
rect 28130 30940 28140 30996
rect 28196 30940 29148 30996
rect 29204 30940 29214 30996
rect 33842 30940 33852 30996
rect 33908 30940 34972 30996
rect 35028 30940 35038 30996
rect 45490 30940 45500 30996
rect 45556 30940 46284 30996
rect 46340 30940 46350 30996
rect 29372 30828 35756 30884
rect 35812 30828 36764 30884
rect 36820 30828 36830 30884
rect 40898 30828 40908 30884
rect 40964 30828 43372 30884
rect 43428 30828 45052 30884
rect 45108 30828 45118 30884
rect 29372 30772 29428 30828
rect 28774 30716 28812 30772
rect 28868 30716 29372 30772
rect 29428 30716 29438 30772
rect 32386 30716 32396 30772
rect 32452 30716 33404 30772
rect 33460 30716 33470 30772
rect 34636 30716 34860 30772
rect 34916 30716 34926 30772
rect 11442 30604 11452 30660
rect 11508 30604 26908 30660
rect 32050 30604 32060 30660
rect 32116 30604 32620 30660
rect 32676 30604 33068 30660
rect 33124 30604 33134 30660
rect 33702 30604 33740 30660
rect 33796 30604 33806 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 34636 30548 34692 30716
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 25666 30492 25676 30548
rect 25732 30492 26684 30548
rect 26740 30492 26750 30548
rect 31490 30492 31500 30548
rect 31556 30492 33964 30548
rect 34020 30492 34188 30548
rect 34244 30492 34254 30548
rect 34626 30492 34636 30548
rect 34692 30492 34702 30548
rect 26226 30380 26236 30436
rect 26292 30380 27468 30436
rect 27524 30380 27534 30436
rect 31154 30380 31164 30436
rect 31220 30380 34860 30436
rect 34916 30380 34926 30436
rect 43138 30380 43148 30436
rect 43204 30380 44380 30436
rect 44436 30380 44446 30436
rect 2818 30268 2828 30324
rect 2884 30268 2894 30324
rect 4946 30268 4956 30324
rect 5012 30268 5022 30324
rect 16258 30268 16268 30324
rect 16324 30268 16940 30324
rect 16996 30268 17006 30324
rect 33730 30268 33740 30324
rect 33796 30268 33852 30324
rect 33908 30268 33918 30324
rect 34290 30268 34300 30324
rect 34356 30268 35756 30324
rect 35812 30268 35822 30324
rect 37202 30268 37212 30324
rect 37268 30268 38220 30324
rect 38276 30268 38286 30324
rect 41682 30268 41692 30324
rect 41748 30268 42252 30324
rect 42308 30268 42318 30324
rect 2828 30212 2884 30268
rect 2828 30156 3724 30212
rect 3780 30156 3790 30212
rect 4956 30100 5012 30268
rect 5954 30156 5964 30212
rect 6020 30156 7980 30212
rect 8036 30156 8046 30212
rect 13794 30156 13804 30212
rect 13860 30156 14476 30212
rect 14532 30156 14542 30212
rect 15250 30156 15260 30212
rect 15316 30156 15596 30212
rect 15652 30156 17052 30212
rect 17108 30156 18732 30212
rect 18788 30156 20076 30212
rect 20132 30156 22316 30212
rect 22372 30156 22382 30212
rect 34178 30156 34188 30212
rect 34244 30156 36204 30212
rect 36260 30156 36270 30212
rect 36418 30156 36428 30212
rect 36484 30156 40348 30212
rect 40404 30156 41580 30212
rect 41636 30156 41646 30212
rect 4956 30044 5628 30100
rect 5684 30044 5694 30100
rect 5964 29988 6020 30156
rect 7634 30044 7644 30100
rect 7700 30044 8204 30100
rect 8260 30044 8270 30100
rect 10210 30044 10220 30100
rect 10276 30044 10668 30100
rect 10724 30044 11116 30100
rect 11172 30044 11788 30100
rect 11844 30044 11854 30100
rect 12114 30044 12124 30100
rect 12180 30044 14028 30100
rect 14084 30044 14094 30100
rect 19842 30044 19852 30100
rect 19908 30044 20636 30100
rect 20692 30044 20702 30100
rect 31490 30044 31500 30100
rect 31556 30044 32060 30100
rect 32116 30044 32126 30100
rect 34402 30044 34412 30100
rect 34468 30044 35308 30100
rect 35364 30044 36652 30100
rect 36708 30044 36718 30100
rect 4162 29932 4172 29988
rect 4228 29932 6020 29988
rect 9874 29932 9884 29988
rect 9940 29932 10556 29988
rect 10612 29932 11452 29988
rect 11508 29932 11518 29988
rect 12226 29932 12236 29988
rect 12292 29932 13244 29988
rect 13300 29932 13310 29988
rect 28578 29932 28588 29988
rect 28644 29932 31724 29988
rect 31780 29932 31790 29988
rect 33282 29932 33292 29988
rect 33348 29932 34636 29988
rect 34692 29932 34702 29988
rect 36530 29932 36540 29988
rect 36596 29932 37100 29988
rect 37156 29932 38108 29988
rect 38164 29932 38174 29988
rect 12338 29820 12348 29876
rect 12404 29820 12796 29876
rect 12852 29820 12862 29876
rect 26852 29820 30044 29876
rect 30100 29820 30110 29876
rect 30818 29820 30828 29876
rect 30884 29820 31500 29876
rect 31556 29820 31948 29876
rect 32004 29820 33180 29876
rect 33236 29820 33246 29876
rect 33702 29820 33740 29876
rect 33796 29820 33806 29876
rect 34038 29820 34076 29876
rect 34132 29820 34142 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 26852 29764 26908 29820
rect 3378 29708 3388 29764
rect 3444 29708 5740 29764
rect 5796 29708 6412 29764
rect 6468 29708 6478 29764
rect 24434 29708 24444 29764
rect 24500 29708 26908 29764
rect 28588 29708 28812 29764
rect 28868 29708 28878 29764
rect 29922 29708 29932 29764
rect 29988 29708 36204 29764
rect 36260 29708 36270 29764
rect 28588 29652 28644 29708
rect 6850 29596 6860 29652
rect 6916 29596 7532 29652
rect 7588 29596 7598 29652
rect 8530 29596 8540 29652
rect 8596 29596 10668 29652
rect 10724 29596 10734 29652
rect 26450 29596 26460 29652
rect 26516 29596 26908 29652
rect 26964 29596 26974 29652
rect 27122 29596 27132 29652
rect 27188 29596 27198 29652
rect 28578 29596 28588 29652
rect 28644 29596 28654 29652
rect 32162 29596 32172 29652
rect 32228 29596 32956 29652
rect 33012 29596 35532 29652
rect 35588 29596 35598 29652
rect 42018 29596 42028 29652
rect 42084 29596 42364 29652
rect 42420 29596 42812 29652
rect 42868 29596 42878 29652
rect 27132 29540 27188 29596
rect 16034 29484 16044 29540
rect 16100 29484 17388 29540
rect 17444 29484 17454 29540
rect 20626 29484 20636 29540
rect 20692 29484 21420 29540
rect 21476 29484 23884 29540
rect 23940 29484 23950 29540
rect 25666 29484 25676 29540
rect 25732 29484 27188 29540
rect 27906 29484 27916 29540
rect 27972 29484 29372 29540
rect 29428 29484 29438 29540
rect 32386 29484 32396 29540
rect 32452 29484 34524 29540
rect 34580 29484 34590 29540
rect 34850 29484 34860 29540
rect 34916 29484 34926 29540
rect 34860 29428 34916 29484
rect 2930 29372 2940 29428
rect 2996 29372 4172 29428
rect 4228 29372 4238 29428
rect 4722 29372 4732 29428
rect 4788 29372 7084 29428
rect 7140 29372 7150 29428
rect 9762 29372 9772 29428
rect 9828 29372 10332 29428
rect 10388 29372 13244 29428
rect 13300 29372 13310 29428
rect 16594 29372 16604 29428
rect 16660 29372 17612 29428
rect 17668 29372 17678 29428
rect 26002 29372 26012 29428
rect 26068 29372 29148 29428
rect 29204 29372 29214 29428
rect 30034 29372 30044 29428
rect 30100 29372 31948 29428
rect 32004 29372 32508 29428
rect 32564 29372 32574 29428
rect 33618 29372 33628 29428
rect 33684 29372 33694 29428
rect 34626 29372 34636 29428
rect 34692 29372 36428 29428
rect 36484 29372 36494 29428
rect 33628 29316 33684 29372
rect 27346 29260 27356 29316
rect 27412 29260 33684 29316
rect 33964 29260 41020 29316
rect 41076 29260 41086 29316
rect 33964 29204 34020 29260
rect 28802 29148 28812 29204
rect 28868 29148 32620 29204
rect 32676 29148 32686 29204
rect 33954 29148 33964 29204
rect 34020 29148 34030 29204
rect 38882 29148 38892 29204
rect 38948 29148 39452 29204
rect 39508 29148 41244 29204
rect 41300 29148 41580 29204
rect 41636 29148 41646 29204
rect 10994 29036 11004 29092
rect 11060 29036 13020 29092
rect 13076 29036 13086 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 30594 28924 30604 28980
rect 30660 28924 32284 28980
rect 32340 28924 34412 28980
rect 34468 28924 34478 28980
rect 36642 28924 36652 28980
rect 36708 28924 37604 28980
rect 6402 28812 6412 28868
rect 6468 28812 8988 28868
rect 9044 28812 10668 28868
rect 10724 28812 10734 28868
rect 14466 28812 14476 28868
rect 14532 28812 16268 28868
rect 16324 28812 17500 28868
rect 17556 28812 17566 28868
rect 32162 28812 32172 28868
rect 32228 28812 33516 28868
rect 33572 28812 33582 28868
rect 34850 28812 34860 28868
rect 34916 28812 37156 28868
rect 1922 28700 1932 28756
rect 1988 28700 6636 28756
rect 6692 28700 6702 28756
rect 10770 28700 10780 28756
rect 10836 28700 11788 28756
rect 11844 28700 12684 28756
rect 12740 28700 13356 28756
rect 13412 28700 13422 28756
rect 23426 28700 23436 28756
rect 23492 28700 24444 28756
rect 24500 28700 24510 28756
rect 26674 28700 26684 28756
rect 26740 28700 29260 28756
rect 29316 28700 29708 28756
rect 29764 28700 29774 28756
rect 29922 28700 29932 28756
rect 29988 28700 31052 28756
rect 31108 28700 31118 28756
rect 33730 28700 33740 28756
rect 33796 28700 35476 28756
rect 35420 28644 35476 28700
rect 37100 28644 37156 28812
rect 6178 28588 6188 28644
rect 6244 28588 6972 28644
rect 7028 28588 7038 28644
rect 12786 28588 12796 28644
rect 12852 28588 13580 28644
rect 13636 28588 16940 28644
rect 16996 28588 17006 28644
rect 30370 28588 30380 28644
rect 30436 28588 34412 28644
rect 34468 28588 34478 28644
rect 35410 28588 35420 28644
rect 35476 28588 35486 28644
rect 35970 28588 35980 28644
rect 36036 28588 36876 28644
rect 36932 28588 36942 28644
rect 37090 28588 37100 28644
rect 37156 28588 37166 28644
rect 37548 28532 37604 28924
rect 42242 28700 42252 28756
rect 42308 28700 42924 28756
rect 42980 28700 42990 28756
rect 41010 28588 41020 28644
rect 41076 28588 41356 28644
rect 41412 28588 44268 28644
rect 44324 28588 44940 28644
rect 44996 28588 45006 28644
rect 9874 28476 9884 28532
rect 9940 28476 11116 28532
rect 11172 28476 11182 28532
rect 23986 28476 23996 28532
rect 24052 28476 25116 28532
rect 25172 28476 25182 28532
rect 37538 28476 37548 28532
rect 37604 28476 37614 28532
rect 2146 28364 2156 28420
rect 2212 28364 2222 28420
rect 23202 28364 23212 28420
rect 23268 28364 25788 28420
rect 25844 28364 25854 28420
rect 37202 28364 37212 28420
rect 37268 28364 37772 28420
rect 37828 28364 38444 28420
rect 38500 28364 38510 28420
rect 2156 27972 2212 28364
rect 22306 28252 22316 28308
rect 22372 28252 26348 28308
rect 26404 28252 26414 28308
rect 32610 28252 32620 28308
rect 32676 28252 33628 28308
rect 33684 28252 33694 28308
rect 41906 28252 41916 28308
rect 41972 28252 43820 28308
rect 43876 28252 43886 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 3826 28140 3836 28196
rect 3892 28140 4732 28196
rect 4788 28140 4798 28196
rect 7522 28140 7532 28196
rect 7588 28140 8092 28196
rect 8148 28140 8158 28196
rect 25890 28140 25900 28196
rect 25956 28140 26908 28196
rect 26964 28140 26974 28196
rect 3154 28028 3164 28084
rect 3220 28028 4060 28084
rect 4116 28028 4396 28084
rect 4452 28028 4462 28084
rect 4620 27972 4676 28140
rect 6066 28028 6076 28084
rect 6132 28028 6636 28084
rect 6692 28028 7532 28084
rect 7588 28028 7598 28084
rect 15586 28028 15596 28084
rect 15652 28028 16268 28084
rect 16324 28028 28924 28084
rect 28980 28028 28990 28084
rect 30146 28028 30156 28084
rect 30212 28028 30492 28084
rect 30548 28028 30558 28084
rect 36866 28028 36876 28084
rect 36932 28028 37548 28084
rect 37604 28028 37614 28084
rect 2156 27916 2716 27972
rect 2772 27916 6412 27972
rect 6468 27916 6478 27972
rect 6626 27916 6636 27972
rect 6692 27916 8092 27972
rect 8148 27916 9212 27972
rect 9268 27916 9660 27972
rect 9716 27916 9726 27972
rect 11890 27916 11900 27972
rect 11956 27916 14140 27972
rect 14196 27916 14206 27972
rect 22754 27916 22764 27972
rect 22820 27916 24668 27972
rect 24724 27916 24734 27972
rect 2146 27804 2156 27860
rect 2212 27804 3164 27860
rect 3220 27804 3230 27860
rect 5282 27804 5292 27860
rect 5348 27804 6860 27860
rect 6916 27804 6926 27860
rect 7410 27804 7420 27860
rect 7476 27804 10220 27860
rect 10276 27804 10286 27860
rect 24098 27804 24108 27860
rect 24164 27804 25452 27860
rect 25508 27804 25518 27860
rect 27682 27804 27692 27860
rect 27748 27804 29932 27860
rect 29988 27804 29998 27860
rect 35074 27804 35084 27860
rect 35140 27804 35420 27860
rect 35476 27804 36204 27860
rect 36260 27804 36270 27860
rect 37548 27748 37604 28028
rect 39890 27804 39900 27860
rect 39956 27804 41020 27860
rect 41076 27804 41086 27860
rect 20514 27692 20524 27748
rect 20580 27692 21868 27748
rect 21924 27692 21934 27748
rect 25218 27692 25228 27748
rect 25284 27692 25900 27748
rect 25956 27692 25966 27748
rect 32918 27692 32956 27748
rect 33012 27692 33022 27748
rect 37548 27692 43036 27748
rect 43092 27692 43102 27748
rect 43362 27692 43372 27748
rect 43428 27692 43820 27748
rect 43876 27692 43886 27748
rect 0 27636 400 27664
rect 0 27580 2604 27636
rect 2660 27580 2670 27636
rect 4172 27580 4396 27636
rect 4452 27580 4462 27636
rect 5282 27580 5292 27636
rect 5348 27580 5740 27636
rect 5796 27580 5806 27636
rect 27682 27580 27692 27636
rect 27748 27580 28476 27636
rect 28532 27580 28542 27636
rect 30818 27580 30828 27636
rect 30884 27580 31948 27636
rect 32004 27580 34860 27636
rect 34916 27580 36428 27636
rect 36484 27580 37436 27636
rect 37492 27580 37502 27636
rect 40338 27580 40348 27636
rect 40404 27580 41692 27636
rect 41748 27580 41758 27636
rect 0 27552 400 27580
rect 2146 27468 2156 27524
rect 2212 27468 3724 27524
rect 3780 27468 3790 27524
rect 4172 27300 4228 27580
rect 25666 27468 25676 27524
rect 25732 27468 29988 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 29932 27412 29988 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 5058 27356 5068 27412
rect 5124 27356 6524 27412
rect 6580 27356 6590 27412
rect 10322 27356 10332 27412
rect 10388 27356 11788 27412
rect 11844 27356 15596 27412
rect 15652 27356 15662 27412
rect 29922 27356 29932 27412
rect 29988 27356 29998 27412
rect 30594 27356 30604 27412
rect 30660 27356 31948 27412
rect 32004 27356 32676 27412
rect 37650 27356 37660 27412
rect 37716 27356 37726 27412
rect 32620 27300 32676 27356
rect 37660 27300 37716 27356
rect 4162 27244 4172 27300
rect 4228 27244 4238 27300
rect 6066 27244 6076 27300
rect 6132 27244 6636 27300
rect 6692 27244 6702 27300
rect 10546 27244 10556 27300
rect 10612 27244 11900 27300
rect 11956 27244 11966 27300
rect 26562 27244 26572 27300
rect 26628 27244 27020 27300
rect 27076 27244 27086 27300
rect 28690 27244 28700 27300
rect 28756 27244 30268 27300
rect 30324 27244 30334 27300
rect 30706 27244 30716 27300
rect 30772 27244 32172 27300
rect 32228 27244 32238 27300
rect 32610 27244 32620 27300
rect 32676 27244 37716 27300
rect 43586 27244 43596 27300
rect 43652 27244 45388 27300
rect 45444 27244 45454 27300
rect 30716 27188 30772 27244
rect 7410 27132 7420 27188
rect 7476 27132 7756 27188
rect 7812 27132 8876 27188
rect 8932 27132 8942 27188
rect 10098 27132 10108 27188
rect 10164 27132 11340 27188
rect 11396 27132 11406 27188
rect 21970 27132 21980 27188
rect 22036 27132 23996 27188
rect 24052 27132 24062 27188
rect 24658 27132 24668 27188
rect 24724 27132 26124 27188
rect 26180 27132 26684 27188
rect 26740 27132 27244 27188
rect 27300 27132 28812 27188
rect 28868 27132 28878 27188
rect 29250 27132 29260 27188
rect 29316 27132 30772 27188
rect 31042 27132 31052 27188
rect 31108 27132 32060 27188
rect 32116 27132 36988 27188
rect 37044 27132 37054 27188
rect 42690 27132 42700 27188
rect 42756 27132 43372 27188
rect 43428 27132 43438 27188
rect 6850 27020 6860 27076
rect 6916 27020 7644 27076
rect 7700 27020 8428 27076
rect 8484 27020 8764 27076
rect 8820 27020 8830 27076
rect 19394 27020 19404 27076
rect 19460 27020 21308 27076
rect 21364 27020 22316 27076
rect 22372 27020 22382 27076
rect 29474 27020 29484 27076
rect 29540 27020 29820 27076
rect 29876 27020 30828 27076
rect 30884 27020 30894 27076
rect 43026 27020 43036 27076
rect 43092 27020 43596 27076
rect 43652 27020 44268 27076
rect 44324 27020 44334 27076
rect 3266 26908 3276 26964
rect 3332 26908 3724 26964
rect 3780 26908 3790 26964
rect 7494 26908 7532 26964
rect 7588 26908 7598 26964
rect 11666 26908 11676 26964
rect 11732 26908 12124 26964
rect 12180 26908 12190 26964
rect 22530 26908 22540 26964
rect 22596 26908 23212 26964
rect 23268 26908 23278 26964
rect 25554 26908 25564 26964
rect 25620 26908 26012 26964
rect 26068 26908 26078 26964
rect 27132 26908 28476 26964
rect 28532 26908 31276 26964
rect 31332 26908 31342 26964
rect 40450 26908 40460 26964
rect 40516 26908 41132 26964
rect 41188 26908 47180 26964
rect 47236 26908 47246 26964
rect 27122 26852 27132 26908
rect 27188 26852 27198 26908
rect 6290 26796 6300 26852
rect 6356 26796 7756 26852
rect 7812 26796 7822 26852
rect 8194 26796 8204 26852
rect 8260 26796 8316 26852
rect 8372 26796 9660 26852
rect 9716 26796 9726 26852
rect 17602 26796 17612 26852
rect 17668 26796 20972 26852
rect 21028 26796 21038 26852
rect 23874 26796 23884 26852
rect 23940 26796 24556 26852
rect 24612 26796 24622 26852
rect 28242 26796 28252 26852
rect 28308 26796 31500 26852
rect 31556 26796 35196 26852
rect 35252 26796 35644 26852
rect 35700 26796 39228 26852
rect 39284 26796 39900 26852
rect 39956 26796 39966 26852
rect 24994 26684 25004 26740
rect 25060 26684 27020 26740
rect 27076 26684 27086 26740
rect 37762 26684 37772 26740
rect 37828 26684 38108 26740
rect 38164 26684 38174 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 4834 26572 4844 26628
rect 4900 26572 7644 26628
rect 7700 26572 7710 26628
rect 8278 26572 8316 26628
rect 8372 26572 8382 26628
rect 16034 26572 16044 26628
rect 16100 26572 17276 26628
rect 17332 26572 17342 26628
rect 26898 26572 26908 26628
rect 26964 26572 28476 26628
rect 28532 26572 28542 26628
rect 29026 26572 29036 26628
rect 29092 26572 32620 26628
rect 32676 26572 32686 26628
rect 4050 26460 4060 26516
rect 4116 26460 4956 26516
rect 5012 26460 5022 26516
rect 6738 26460 6748 26516
rect 6804 26460 8876 26516
rect 8932 26460 8942 26516
rect 25442 26460 25452 26516
rect 25508 26460 27244 26516
rect 27300 26460 31388 26516
rect 31444 26460 31454 26516
rect 37650 26460 37660 26516
rect 37716 26460 39116 26516
rect 39172 26460 39182 26516
rect 27570 26348 27580 26404
rect 27636 26348 28252 26404
rect 28308 26348 28318 26404
rect 28466 26348 28476 26404
rect 28532 26348 29036 26404
rect 29092 26348 29102 26404
rect 2258 26236 2268 26292
rect 2324 26236 3052 26292
rect 3108 26236 3118 26292
rect 23202 26236 23212 26292
rect 23268 26236 23884 26292
rect 23940 26236 23950 26292
rect 32386 26236 32396 26292
rect 32452 26236 33068 26292
rect 33124 26236 33134 26292
rect 6178 26124 6188 26180
rect 6244 26124 7196 26180
rect 7252 26124 7262 26180
rect 20962 26124 20972 26180
rect 21028 26124 21420 26180
rect 21476 26124 23996 26180
rect 24052 26124 24062 26180
rect 17042 26012 17052 26068
rect 17108 26012 18060 26068
rect 18116 26012 18732 26068
rect 18788 26012 18798 26068
rect 24546 26012 24556 26068
rect 24612 26012 25452 26068
rect 25508 26012 25518 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 9090 25788 9100 25844
rect 9156 25788 10220 25844
rect 10276 25788 10286 25844
rect 27010 25788 27020 25844
rect 27076 25788 31612 25844
rect 31668 25788 31678 25844
rect 7532 25676 7868 25732
rect 7924 25676 7934 25732
rect 7532 25508 7588 25676
rect 7746 25564 7756 25620
rect 7812 25564 8988 25620
rect 9044 25564 9054 25620
rect 11666 25564 11676 25620
rect 11732 25564 12572 25620
rect 12628 25564 12638 25620
rect 17266 25564 17276 25620
rect 17332 25564 22092 25620
rect 22148 25564 22158 25620
rect 29698 25564 29708 25620
rect 29764 25564 30380 25620
rect 30436 25564 30446 25620
rect 7532 25452 7980 25508
rect 8036 25452 8046 25508
rect 10322 25452 10332 25508
rect 10388 25452 10836 25508
rect 10780 25396 10836 25452
rect 7858 25340 7868 25396
rect 7924 25340 8764 25396
rect 8820 25340 8830 25396
rect 10770 25340 10780 25396
rect 10836 25340 11228 25396
rect 11284 25340 11294 25396
rect 8082 25228 8092 25284
rect 8148 25228 10108 25284
rect 10164 25228 10174 25284
rect 29698 25228 29708 25284
rect 29764 25228 29932 25284
rect 29988 25228 29998 25284
rect 32274 25228 32284 25284
rect 32340 25228 33404 25284
rect 33460 25228 36652 25284
rect 36708 25228 36718 25284
rect 10658 25116 10668 25172
rect 10724 25116 11340 25172
rect 11396 25116 11900 25172
rect 11956 25116 11966 25172
rect 44258 25116 44268 25172
rect 44324 25116 45164 25172
rect 45220 25116 45230 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 5618 25004 5628 25060
rect 5684 25004 6300 25060
rect 6356 25004 7196 25060
rect 7252 25004 7262 25060
rect 31154 25004 31164 25060
rect 31220 25004 31276 25060
rect 31332 25004 31342 25060
rect 2370 24892 2380 24948
rect 2436 24892 2940 24948
rect 2996 24892 9212 24948
rect 9268 24892 9278 24948
rect 13234 24892 13244 24948
rect 13300 24892 14476 24948
rect 14532 24892 16492 24948
rect 16548 24892 17500 24948
rect 17556 24892 17566 24948
rect 32918 24892 32956 24948
rect 33012 24892 33022 24948
rect 36418 24892 36428 24948
rect 36484 24892 37212 24948
rect 37268 24892 38780 24948
rect 38836 24892 38846 24948
rect 41010 24892 41020 24948
rect 41076 24892 41468 24948
rect 41524 24892 42812 24948
rect 42868 24892 43260 24948
rect 43316 24892 43326 24948
rect 3378 24780 3388 24836
rect 3444 24780 4396 24836
rect 4452 24780 5964 24836
rect 6020 24780 7084 24836
rect 7140 24780 7150 24836
rect 7634 24780 7644 24836
rect 7700 24780 8876 24836
rect 8932 24780 8942 24836
rect 31938 24780 31948 24836
rect 32004 24780 33180 24836
rect 33236 24780 33246 24836
rect 6262 24668 6300 24724
rect 6356 24668 6366 24724
rect 7410 24668 7420 24724
rect 7476 24668 9548 24724
rect 9604 24668 9614 24724
rect 22306 24668 22316 24724
rect 22372 24668 24668 24724
rect 24724 24668 24734 24724
rect 3938 24556 3948 24612
rect 4004 24556 9660 24612
rect 9716 24556 9726 24612
rect 15698 24556 15708 24612
rect 15764 24556 16044 24612
rect 16100 24556 19740 24612
rect 19796 24556 19806 24612
rect 22978 24556 22988 24612
rect 23044 24556 25452 24612
rect 25508 24556 36092 24612
rect 36148 24556 36158 24612
rect 6962 24444 6972 24500
rect 7028 24444 7644 24500
rect 7700 24444 7710 24500
rect 10882 24444 10892 24500
rect 10948 24444 12796 24500
rect 12852 24444 20188 24500
rect 20244 24444 20254 24500
rect 32386 24444 32396 24500
rect 32452 24444 32844 24500
rect 32900 24444 32910 24500
rect 7186 24332 7196 24388
rect 7252 24332 7868 24388
rect 7924 24332 8428 24388
rect 8484 24332 9100 24388
rect 9156 24332 9166 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 7410 24220 7420 24276
rect 7476 24220 9884 24276
rect 9940 24220 9950 24276
rect 7746 24108 7756 24164
rect 7812 24108 8316 24164
rect 8372 24108 8382 24164
rect 8530 24108 8540 24164
rect 8596 24108 11228 24164
rect 11284 24108 13468 24164
rect 13524 24108 13534 24164
rect 13906 24108 13916 24164
rect 13972 24108 16044 24164
rect 16100 24108 16110 24164
rect 41906 24108 41916 24164
rect 41972 24108 42588 24164
rect 42644 24108 43932 24164
rect 43988 24108 43998 24164
rect 5058 23996 5068 24052
rect 5124 23996 5628 24052
rect 5684 23996 5694 24052
rect 7830 23996 7868 24052
rect 7924 23996 7934 24052
rect 8194 23996 8204 24052
rect 8260 23996 8876 24052
rect 8932 23996 8942 24052
rect 13794 23996 13804 24052
rect 13860 23996 14700 24052
rect 14756 23996 14766 24052
rect 24322 23996 24332 24052
rect 24388 23996 26012 24052
rect 26068 23996 27020 24052
rect 27076 23996 27580 24052
rect 27636 23996 27646 24052
rect 27794 23996 27804 24052
rect 27860 23996 28252 24052
rect 28308 23996 38556 24052
rect 38612 23996 38622 24052
rect 42802 23996 42812 24052
rect 42868 23996 47740 24052
rect 47796 23996 47806 24052
rect 2258 23884 2268 23940
rect 2324 23884 3388 23940
rect 6514 23884 6524 23940
rect 6580 23884 10108 23940
rect 10164 23884 10174 23940
rect 15446 23884 15484 23940
rect 15540 23884 16716 23940
rect 16772 23884 16782 23940
rect 22082 23884 22092 23940
rect 22148 23884 22764 23940
rect 22820 23884 22830 23940
rect 27906 23884 27916 23940
rect 27972 23884 29596 23940
rect 29652 23884 29662 23940
rect 32498 23884 32508 23940
rect 32564 23884 33068 23940
rect 33124 23884 33134 23940
rect 43698 23884 43708 23940
rect 43764 23884 44268 23940
rect 44324 23884 44334 23940
rect 3332 23716 3388 23884
rect 6626 23772 6636 23828
rect 6692 23772 6972 23828
rect 7028 23772 7038 23828
rect 7308 23772 9772 23828
rect 9828 23772 9838 23828
rect 15026 23772 15036 23828
rect 15092 23772 16380 23828
rect 16436 23772 16446 23828
rect 24322 23772 24332 23828
rect 24388 23772 24556 23828
rect 24612 23772 26796 23828
rect 26852 23772 32396 23828
rect 32452 23772 32462 23828
rect 7308 23716 7364 23772
rect 3332 23660 5292 23716
rect 5348 23660 5358 23716
rect 5730 23660 5740 23716
rect 5796 23660 5964 23716
rect 6020 23660 6860 23716
rect 6916 23660 6926 23716
rect 7298 23660 7308 23716
rect 7364 23660 7374 23716
rect 7746 23660 7756 23716
rect 7812 23660 8428 23716
rect 8484 23660 8494 23716
rect 12562 23660 12572 23716
rect 12628 23660 12908 23716
rect 12964 23660 13580 23716
rect 13636 23660 13646 23716
rect 24658 23660 24668 23716
rect 24724 23660 31164 23716
rect 31220 23660 31230 23716
rect 31602 23660 31612 23716
rect 31668 23660 32060 23716
rect 32116 23660 32126 23716
rect 32498 23660 32508 23716
rect 32564 23660 32844 23716
rect 32900 23660 32910 23716
rect 5292 23604 5348 23660
rect 5068 23548 5348 23604
rect 6486 23548 6524 23604
rect 6580 23548 6590 23604
rect 8082 23548 8092 23604
rect 8148 23548 11676 23604
rect 11732 23548 16940 23604
rect 16996 23548 17006 23604
rect 40338 23548 40348 23604
rect 40404 23548 43708 23604
rect 5068 23492 5124 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 40348 23492 40404 23548
rect 5058 23436 5068 23492
rect 5124 23436 5134 23492
rect 5516 23436 5628 23492
rect 5684 23436 5694 23492
rect 5842 23436 5852 23492
rect 5908 23436 6412 23492
rect 6468 23436 6478 23492
rect 6738 23436 6748 23492
rect 6804 23436 7644 23492
rect 7700 23436 7868 23492
rect 7924 23436 9100 23492
rect 9156 23436 9166 23492
rect 38210 23436 38220 23492
rect 38276 23436 40404 23492
rect 4274 23324 4284 23380
rect 4340 23324 4956 23380
rect 5012 23324 5022 23380
rect 5516 23268 5572 23436
rect 14690 23324 14700 23380
rect 14756 23324 15484 23380
rect 15540 23324 15550 23380
rect 30594 23324 30604 23380
rect 30660 23324 33180 23380
rect 33236 23324 33246 23380
rect 4834 23212 4844 23268
rect 4900 23212 4910 23268
rect 5516 23212 7308 23268
rect 7364 23212 7374 23268
rect 9202 23212 9212 23268
rect 9268 23212 12124 23268
rect 12180 23212 12190 23268
rect 18946 23212 18956 23268
rect 19012 23212 19628 23268
rect 19684 23212 19694 23268
rect 4844 23156 4900 23212
rect 4844 23100 7420 23156
rect 7476 23100 7486 23156
rect 7858 23100 7868 23156
rect 7924 23100 8316 23156
rect 8372 23100 8382 23156
rect 8866 23100 8876 23156
rect 8932 23100 9100 23156
rect 9156 23100 10444 23156
rect 10500 23100 10510 23156
rect 17938 23100 17948 23156
rect 18004 23100 18508 23156
rect 18564 23100 18574 23156
rect 26852 23100 27020 23156
rect 27076 23100 27086 23156
rect 29922 23100 29932 23156
rect 29988 23100 30380 23156
rect 30436 23100 30446 23156
rect 31602 23100 31612 23156
rect 31668 23100 32172 23156
rect 32228 23100 33404 23156
rect 33460 23100 34300 23156
rect 34356 23100 34366 23156
rect 43652 23100 43708 23548
rect 43764 23100 43774 23156
rect 26852 23044 26908 23100
rect 5394 22988 5404 23044
rect 5460 22988 6748 23044
rect 6804 22988 6814 23044
rect 26674 22988 26684 23044
rect 26740 22988 26908 23044
rect 40898 22988 40908 23044
rect 40964 22988 42028 23044
rect 42084 22988 42094 23044
rect 6262 22876 6300 22932
rect 6356 22876 6366 22932
rect 17826 22876 17836 22932
rect 17892 22876 18620 22932
rect 18676 22876 18686 22932
rect 24546 22876 24556 22932
rect 24612 22876 25340 22932
rect 25396 22876 25406 22932
rect 25666 22876 25676 22932
rect 25732 22876 26012 22932
rect 26068 22876 26078 22932
rect 12114 22764 12124 22820
rect 12180 22764 18508 22820
rect 18564 22764 18574 22820
rect 0 22708 400 22736
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 0 22652 1708 22708
rect 1764 22652 1774 22708
rect 19170 22652 19180 22708
rect 19236 22652 27020 22708
rect 27076 22652 27356 22708
rect 27412 22652 27422 22708
rect 0 22624 400 22652
rect 4498 22540 4508 22596
rect 4564 22540 8316 22596
rect 8372 22540 9772 22596
rect 9828 22540 10668 22596
rect 10724 22540 10734 22596
rect 10882 22540 10892 22596
rect 10948 22540 11676 22596
rect 11732 22540 22204 22596
rect 22260 22540 22270 22596
rect 26114 22540 26124 22596
rect 26180 22540 26908 22596
rect 26964 22540 26974 22596
rect 10668 22484 10724 22540
rect 1810 22428 1820 22484
rect 1876 22428 5740 22484
rect 5796 22428 7196 22484
rect 7252 22428 7262 22484
rect 10668 22428 11228 22484
rect 11284 22428 11900 22484
rect 11956 22428 12572 22484
rect 12628 22428 12638 22484
rect 20514 22428 20524 22484
rect 20580 22428 21420 22484
rect 21476 22428 33964 22484
rect 34020 22428 34030 22484
rect 36642 22428 36652 22484
rect 36708 22428 37772 22484
rect 37828 22428 37838 22484
rect 16818 22316 16828 22372
rect 16884 22316 17612 22372
rect 17668 22316 19516 22372
rect 19572 22316 20972 22372
rect 21028 22316 23100 22372
rect 23156 22316 24332 22372
rect 24388 22316 24398 22372
rect 35074 22316 35084 22372
rect 35140 22316 37100 22372
rect 37156 22316 38220 22372
rect 38276 22316 38286 22372
rect 26898 22204 26908 22260
rect 26964 22204 27244 22260
rect 27300 22204 34076 22260
rect 34132 22204 34142 22260
rect 28018 22092 28028 22148
rect 28084 22092 28700 22148
rect 28756 22092 29260 22148
rect 29316 22092 29326 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 7970 21756 7980 21812
rect 8036 21756 9548 21812
rect 9604 21756 9614 21812
rect 23986 21756 23996 21812
rect 24052 21756 24668 21812
rect 24724 21756 25228 21812
rect 25284 21756 26684 21812
rect 26740 21756 26750 21812
rect 31938 21756 31948 21812
rect 32004 21756 33516 21812
rect 33572 21756 33582 21812
rect 33954 21756 33964 21812
rect 34020 21756 35196 21812
rect 35252 21756 39228 21812
rect 39284 21756 39294 21812
rect 31948 21700 32004 21756
rect 10322 21644 10332 21700
rect 10388 21644 10892 21700
rect 10948 21644 11564 21700
rect 11620 21644 11630 21700
rect 16370 21644 16380 21700
rect 16436 21644 17388 21700
rect 17444 21644 17454 21700
rect 30818 21644 30828 21700
rect 30884 21644 32004 21700
rect 35858 21644 35868 21700
rect 35924 21644 38892 21700
rect 38948 21644 38958 21700
rect 2482 21532 2492 21588
rect 2548 21532 3052 21588
rect 3108 21532 3388 21588
rect 7970 21532 7980 21588
rect 8036 21532 9772 21588
rect 9828 21532 9838 21588
rect 14252 21532 14700 21588
rect 14756 21532 14766 21588
rect 20850 21532 20860 21588
rect 20916 21532 23884 21588
rect 23940 21532 23950 21588
rect 30482 21532 30492 21588
rect 30548 21532 31164 21588
rect 31220 21532 31500 21588
rect 31556 21532 31566 21588
rect 36054 21532 36092 21588
rect 36148 21532 36158 21588
rect 41906 21532 41916 21588
rect 41972 21532 42476 21588
rect 42532 21532 42542 21588
rect 3332 21476 3388 21532
rect 14252 21476 14308 21532
rect 3332 21420 13692 21476
rect 13748 21420 14252 21476
rect 14308 21420 14318 21476
rect 14466 21420 14476 21476
rect 14532 21420 15820 21476
rect 15876 21420 18620 21476
rect 18676 21420 18686 21476
rect 22418 21420 22428 21476
rect 22484 21420 23436 21476
rect 23492 21420 23502 21476
rect 25890 21420 25900 21476
rect 25956 21420 28140 21476
rect 28196 21420 28206 21476
rect 35970 21420 35980 21476
rect 36036 21420 36204 21476
rect 36260 21420 36270 21476
rect 38322 21420 38332 21476
rect 38388 21420 38780 21476
rect 38836 21420 40012 21476
rect 40068 21420 40078 21476
rect 34402 21308 34412 21364
rect 34468 21308 35084 21364
rect 35140 21308 36876 21364
rect 36932 21308 36942 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 3798 21084 3836 21140
rect 3892 21084 3902 21140
rect 13458 21084 13468 21140
rect 13524 21084 17500 21140
rect 17556 21084 17566 21140
rect 22754 20972 22764 21028
rect 22820 20972 23772 21028
rect 23828 20972 23838 21028
rect 36530 20972 36540 21028
rect 36596 20972 39228 21028
rect 39284 20972 39294 21028
rect 9314 20860 9324 20916
rect 9380 20860 11004 20916
rect 11060 20860 11070 20916
rect 23874 20860 23884 20916
rect 23940 20860 24108 20916
rect 24164 20860 24174 20916
rect 31378 20860 31388 20916
rect 31444 20860 32284 20916
rect 32340 20860 32350 20916
rect 32946 20860 32956 20916
rect 33012 20860 38220 20916
rect 38276 20860 38286 20916
rect 23538 20748 23548 20804
rect 23604 20748 26012 20804
rect 26068 20748 26078 20804
rect 18946 20636 18956 20692
rect 19012 20636 29484 20692
rect 29540 20636 29550 20692
rect 9650 20524 9660 20580
rect 9716 20524 13468 20580
rect 13524 20524 13534 20580
rect 22530 20524 22540 20580
rect 22596 20524 22876 20580
rect 22932 20524 23548 20580
rect 23986 20524 23996 20580
rect 24052 20524 30380 20580
rect 30436 20524 30446 20580
rect 30828 20524 37660 20580
rect 37716 20524 37726 20580
rect 23492 20468 23548 20524
rect 23492 20412 30604 20468
rect 30660 20412 30670 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 30828 20356 30884 20524
rect 23426 20300 23436 20356
rect 23492 20300 30884 20356
rect 38210 20300 38220 20356
rect 38276 20300 40124 20356
rect 40180 20300 40348 20356
rect 40404 20300 40414 20356
rect 19506 20188 19516 20244
rect 19572 20188 21644 20244
rect 21700 20188 21710 20244
rect 22754 20132 22764 20188
rect 22820 20132 22830 20188
rect 3042 20076 3052 20132
rect 3108 20076 4284 20132
rect 4340 20076 4350 20132
rect 4834 20076 4844 20132
rect 4900 20076 5740 20132
rect 5796 20076 5806 20132
rect 22764 20020 22820 20132
rect 25330 20076 25340 20132
rect 25396 20076 26572 20132
rect 26628 20076 26638 20132
rect 32050 20076 32060 20132
rect 32116 20076 33180 20132
rect 33236 20076 34860 20132
rect 34916 20076 35532 20132
rect 35588 20076 36204 20132
rect 36260 20076 37548 20132
rect 37604 20076 37614 20132
rect 3378 19964 3388 20020
rect 3444 19964 6860 20020
rect 6916 19964 6926 20020
rect 12562 19964 12572 20020
rect 12628 19964 13020 20020
rect 13076 19964 15596 20020
rect 15652 19964 16380 20020
rect 16436 19964 19068 20020
rect 19124 19964 19134 20020
rect 22530 19964 22540 20020
rect 22596 19964 23996 20020
rect 24052 19964 26348 20020
rect 26404 19964 26414 20020
rect 34066 19964 34076 20020
rect 34132 19964 35196 20020
rect 35252 19964 38892 20020
rect 38948 19964 38958 20020
rect 33730 19852 33740 19908
rect 33796 19852 44604 19908
rect 44660 19852 44670 19908
rect 5954 19628 5964 19684
rect 6020 19628 6636 19684
rect 6692 19628 6702 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 43922 19292 43932 19348
rect 43988 19292 44940 19348
rect 44996 19292 45006 19348
rect 3490 19180 3500 19236
rect 3556 19180 3948 19236
rect 4004 19180 4014 19236
rect 23202 19180 23212 19236
rect 23268 19180 23884 19236
rect 23940 19180 24668 19236
rect 24724 19180 24734 19236
rect 1922 18956 1932 19012
rect 1988 18956 4844 19012
rect 4900 18956 4910 19012
rect 6066 18956 6076 19012
rect 6132 18956 6860 19012
rect 6916 18956 6926 19012
rect 38322 18956 38332 19012
rect 38388 18956 38668 19012
rect 38724 18956 38734 19012
rect 44482 18956 44492 19012
rect 44548 18956 45388 19012
rect 45444 18956 45454 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 6290 18732 6300 18788
rect 6356 18732 6636 18788
rect 6692 18732 6702 18788
rect 7868 18732 8204 18788
rect 8260 18732 8652 18788
rect 8708 18732 8718 18788
rect 7868 18676 7924 18732
rect 2034 18620 2044 18676
rect 2100 18620 2828 18676
rect 2884 18620 3948 18676
rect 4004 18620 4014 18676
rect 5842 18620 5852 18676
rect 5908 18620 6524 18676
rect 6580 18620 7924 18676
rect 8082 18620 8092 18676
rect 8148 18620 9436 18676
rect 9492 18620 9502 18676
rect 14802 18620 14812 18676
rect 14868 18620 17724 18676
rect 17780 18620 17790 18676
rect 23202 18620 23212 18676
rect 23268 18620 25452 18676
rect 25508 18620 25518 18676
rect 2706 18508 2716 18564
rect 2772 18508 3724 18564
rect 3780 18508 3790 18564
rect 5366 18508 5404 18564
rect 5460 18508 5470 18564
rect 6066 18508 6076 18564
rect 6132 18508 7196 18564
rect 7252 18508 7262 18564
rect 7970 18508 7980 18564
rect 8036 18508 9660 18564
rect 9716 18508 9726 18564
rect 23090 18508 23100 18564
rect 23156 18508 23166 18564
rect 31602 18508 31612 18564
rect 31668 18508 31678 18564
rect 37314 18508 37324 18564
rect 37380 18508 37884 18564
rect 37940 18508 37950 18564
rect 6524 18452 6580 18508
rect 23100 18452 23156 18508
rect 2930 18396 2940 18452
rect 2996 18396 4956 18452
rect 5012 18396 5022 18452
rect 5170 18396 5180 18452
rect 5236 18396 6300 18452
rect 6356 18396 6366 18452
rect 6514 18396 6524 18452
rect 6580 18396 6590 18452
rect 6962 18396 6972 18452
rect 7028 18396 7308 18452
rect 7364 18396 7374 18452
rect 8082 18396 8092 18452
rect 8148 18396 8540 18452
rect 8596 18396 8606 18452
rect 10994 18396 11004 18452
rect 11060 18396 11788 18452
rect 11844 18396 12460 18452
rect 12516 18396 14588 18452
rect 14644 18396 14654 18452
rect 18050 18396 18060 18452
rect 18116 18396 18732 18452
rect 18788 18396 23156 18452
rect 23538 18396 23548 18452
rect 23604 18396 24220 18452
rect 24276 18396 24286 18452
rect 24994 18396 25004 18452
rect 25060 18396 26012 18452
rect 26068 18396 26078 18452
rect 6300 18340 6356 18396
rect 31612 18340 31668 18508
rect 6300 18284 7756 18340
rect 7812 18284 8316 18340
rect 8372 18284 8382 18340
rect 18274 18284 18284 18340
rect 18340 18284 18956 18340
rect 19012 18284 19022 18340
rect 31612 18284 32396 18340
rect 32452 18284 33068 18340
rect 33124 18284 33134 18340
rect 36642 18284 36652 18340
rect 36708 18284 38332 18340
rect 38388 18284 39788 18340
rect 39844 18284 39854 18340
rect 3490 18172 3500 18228
rect 3556 18172 4060 18228
rect 4116 18172 4508 18228
rect 4564 18172 4574 18228
rect 17938 18172 17948 18228
rect 18004 18172 20412 18228
rect 20468 18172 20478 18228
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 5842 17948 5852 18004
rect 5908 17948 6188 18004
rect 6244 17948 6254 18004
rect 7186 17948 7196 18004
rect 7252 17948 7980 18004
rect 8036 17948 9436 18004
rect 9492 17948 9502 18004
rect 2034 17836 2044 17892
rect 2100 17836 10780 17892
rect 10836 17836 10846 17892
rect 18834 17836 18844 17892
rect 18900 17836 19628 17892
rect 19684 17836 19694 17892
rect 24770 17836 24780 17892
rect 24836 17836 26236 17892
rect 26292 17836 26908 17892
rect 41906 17836 41916 17892
rect 41972 17836 45276 17892
rect 45332 17836 45342 17892
rect 0 17780 400 17808
rect 0 17724 1708 17780
rect 1764 17724 1774 17780
rect 5366 17724 5404 17780
rect 5460 17724 5740 17780
rect 5796 17724 5806 17780
rect 6962 17724 6972 17780
rect 7028 17724 7868 17780
rect 7924 17724 7934 17780
rect 0 17696 400 17724
rect 6038 17612 6076 17668
rect 6132 17612 6142 17668
rect 6748 17612 7532 17668
rect 7588 17612 7598 17668
rect 8530 17612 8540 17668
rect 8596 17612 9324 17668
rect 9380 17612 9390 17668
rect 17938 17612 17948 17668
rect 18004 17612 19180 17668
rect 19236 17612 19246 17668
rect 6748 17556 6804 17612
rect 3378 17500 3388 17556
rect 3444 17500 3724 17556
rect 3780 17500 3790 17556
rect 4834 17500 4844 17556
rect 4900 17500 6300 17556
rect 6356 17500 6748 17556
rect 6804 17500 6814 17556
rect 8082 17500 8092 17556
rect 8148 17500 8158 17556
rect 8418 17500 8428 17556
rect 8484 17500 9212 17556
rect 9268 17500 9278 17556
rect 17490 17500 17500 17556
rect 17556 17500 18732 17556
rect 18788 17500 18798 17556
rect 20132 17500 21308 17556
rect 21364 17500 21374 17556
rect 4946 17388 4956 17444
rect 5012 17388 6636 17444
rect 6692 17388 7308 17444
rect 7364 17388 7374 17444
rect 8092 17332 8148 17500
rect 20132 17444 20188 17500
rect 13570 17388 13580 17444
rect 13636 17388 14700 17444
rect 14756 17388 15148 17444
rect 15204 17388 16604 17444
rect 16660 17388 20188 17444
rect 26852 17388 26908 17836
rect 31042 17724 31052 17780
rect 31108 17724 31948 17780
rect 32004 17724 33180 17780
rect 33236 17724 33516 17780
rect 33572 17724 36652 17780
rect 36708 17724 36718 17780
rect 39890 17612 39900 17668
rect 39956 17612 40908 17668
rect 40964 17612 40974 17668
rect 29138 17500 29148 17556
rect 29204 17500 32620 17556
rect 32676 17500 32686 17556
rect 26964 17388 27356 17444
rect 27412 17388 29932 17444
rect 29988 17388 29998 17444
rect 2930 17276 2940 17332
rect 2996 17276 3276 17332
rect 3332 17276 3342 17332
rect 5394 17276 5404 17332
rect 5460 17276 8148 17332
rect 20402 17276 20412 17332
rect 20468 17276 22092 17332
rect 22148 17276 22158 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 38612 17220 38668 17332
rect 38724 17276 39340 17332
rect 39396 17276 41468 17332
rect 41524 17276 41534 17332
rect 7746 17164 7756 17220
rect 7812 17164 8204 17220
rect 8260 17164 8270 17220
rect 33618 17164 33628 17220
rect 33684 17164 33964 17220
rect 34020 17164 35644 17220
rect 35700 17164 36204 17220
rect 36260 17164 36764 17220
rect 36820 17164 36830 17220
rect 38322 17164 38332 17220
rect 38388 17164 38668 17220
rect 5058 17052 5068 17108
rect 5124 17052 5740 17108
rect 5796 17052 5806 17108
rect 8082 17052 8092 17108
rect 8148 17052 9772 17108
rect 9828 17052 9838 17108
rect 19282 17052 19292 17108
rect 19348 17052 19516 17108
rect 19572 17052 20188 17108
rect 20244 17052 22316 17108
rect 22372 17052 22382 17108
rect 23650 17052 23660 17108
rect 23716 17052 30268 17108
rect 30324 17052 30334 17108
rect 33842 17052 33852 17108
rect 33908 17052 35196 17108
rect 35252 17052 35756 17108
rect 35812 17052 35822 17108
rect 38434 17052 38444 17108
rect 38500 17052 39788 17108
rect 39844 17052 39854 17108
rect 40226 17052 40236 17108
rect 40292 17052 41916 17108
rect 41972 17052 41982 17108
rect 6066 16940 6076 16996
rect 6132 16940 8540 16996
rect 8596 16940 8606 16996
rect 28802 16940 28812 16996
rect 28868 16940 29708 16996
rect 29764 16940 29774 16996
rect 33506 16940 33516 16996
rect 33572 16940 34412 16996
rect 34468 16940 34478 16996
rect 37650 16940 37660 16996
rect 37716 16940 38948 16996
rect 38892 16884 38948 16940
rect 6076 16828 6636 16884
rect 6692 16828 6702 16884
rect 7522 16828 7532 16884
rect 7588 16828 8428 16884
rect 8484 16828 8494 16884
rect 14130 16828 14140 16884
rect 14196 16828 15036 16884
rect 15092 16828 15102 16884
rect 17826 16828 17836 16884
rect 17892 16828 18620 16884
rect 18676 16828 18686 16884
rect 21298 16828 21308 16884
rect 21364 16828 24668 16884
rect 24724 16828 25116 16884
rect 25172 16828 25564 16884
rect 25620 16828 26684 16884
rect 26740 16828 28028 16884
rect 28084 16828 28094 16884
rect 36530 16828 36540 16884
rect 36596 16828 38108 16884
rect 38164 16828 38174 16884
rect 38882 16828 38892 16884
rect 38948 16828 39564 16884
rect 39620 16828 39630 16884
rect 39778 16828 39788 16884
rect 39844 16828 40460 16884
rect 40516 16828 40526 16884
rect 6076 16772 6132 16828
rect 6066 16716 6076 16772
rect 6132 16716 6142 16772
rect 10546 16716 10556 16772
rect 10612 16716 12796 16772
rect 12852 16716 12862 16772
rect 16258 16716 16268 16772
rect 16324 16716 17052 16772
rect 17108 16716 17118 16772
rect 19170 16716 19180 16772
rect 19236 16716 21084 16772
rect 21140 16716 21150 16772
rect 27346 16716 27356 16772
rect 27412 16716 33740 16772
rect 33796 16716 33806 16772
rect 34962 16716 34972 16772
rect 35028 16716 37996 16772
rect 38052 16716 38062 16772
rect 42018 16716 42028 16772
rect 42084 16716 43036 16772
rect 43092 16716 43484 16772
rect 43540 16716 43550 16772
rect 6598 16604 6636 16660
rect 6692 16604 6702 16660
rect 29474 16604 29484 16660
rect 29540 16604 29932 16660
rect 29988 16604 30268 16660
rect 30324 16604 30334 16660
rect 31378 16604 31388 16660
rect 31444 16604 32060 16660
rect 32116 16604 32126 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 34514 16268 34524 16324
rect 34580 16268 36204 16324
rect 36260 16268 38332 16324
rect 38388 16268 38398 16324
rect 41122 16268 41132 16324
rect 41188 16268 43708 16324
rect 43764 16268 43774 16324
rect 10994 16156 11004 16212
rect 11060 16156 11564 16212
rect 11620 16156 11630 16212
rect 20402 16156 20412 16212
rect 20468 16156 22764 16212
rect 22820 16156 22830 16212
rect 25778 16156 25788 16212
rect 25844 16156 33516 16212
rect 33572 16156 34076 16212
rect 34132 16156 39788 16212
rect 39844 16156 39854 16212
rect 10658 16044 10668 16100
rect 10724 16044 11116 16100
rect 11172 16044 11182 16100
rect 16370 16044 16380 16100
rect 16436 16044 18172 16100
rect 18228 16044 18238 16100
rect 20178 16044 20188 16100
rect 20244 16044 20636 16100
rect 20692 16044 20702 16100
rect 33954 16044 33964 16100
rect 34020 16044 35196 16100
rect 35252 16044 41468 16100
rect 41524 16044 41534 16100
rect 35970 15932 35980 15988
rect 36036 15932 36652 15988
rect 36708 15932 36718 15988
rect 38612 15932 39676 15988
rect 39732 15932 39742 15988
rect 38612 15876 38668 15932
rect 19730 15820 19740 15876
rect 19796 15820 22540 15876
rect 22596 15820 22606 15876
rect 30818 15820 30828 15876
rect 30884 15820 31612 15876
rect 31668 15820 31678 15876
rect 36418 15820 36428 15876
rect 36484 15820 38668 15876
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 20188 15540 20244 15820
rect 35942 15708 35980 15764
rect 36036 15708 36046 15764
rect 11330 15484 11340 15540
rect 11396 15484 12572 15540
rect 12628 15484 12638 15540
rect 20178 15484 20188 15540
rect 20244 15484 20254 15540
rect 34066 15484 34076 15540
rect 34132 15484 34748 15540
rect 34804 15484 34814 15540
rect 19394 15372 19404 15428
rect 19460 15372 21868 15428
rect 21924 15372 21934 15428
rect 39778 15372 39788 15428
rect 39844 15372 40012 15428
rect 40068 15372 41020 15428
rect 41076 15372 41086 15428
rect 10546 15260 10556 15316
rect 10612 15260 11116 15316
rect 11172 15260 11182 15316
rect 11732 15260 12796 15316
rect 12852 15260 12862 15316
rect 28578 15260 28588 15316
rect 28644 15260 29148 15316
rect 29204 15260 29214 15316
rect 35298 15260 35308 15316
rect 35364 15260 35868 15316
rect 35924 15260 35934 15316
rect 41570 15260 41580 15316
rect 41636 15260 42028 15316
rect 42084 15260 42094 15316
rect 11732 15204 11788 15260
rect 9762 15148 9772 15204
rect 9828 15148 11452 15204
rect 11508 15148 11788 15204
rect 31154 15148 31164 15204
rect 31220 15148 33068 15204
rect 33124 15148 34300 15204
rect 34356 15148 34366 15204
rect 10444 15036 11900 15092
rect 11956 15036 13020 15092
rect 13076 15036 13086 15092
rect 23314 15036 23324 15092
rect 23380 15036 23996 15092
rect 24052 15036 24062 15092
rect 10444 14980 10500 15036
rect 10434 14924 10444 14980
rect 10500 14924 10510 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 35746 14812 35756 14868
rect 35812 14812 37212 14868
rect 37268 14812 38444 14868
rect 38500 14812 38510 14868
rect 35756 14756 35812 14812
rect 29810 14700 29820 14756
rect 29876 14700 30156 14756
rect 30212 14700 30222 14756
rect 35410 14700 35420 14756
rect 35476 14700 35812 14756
rect 2034 14588 2044 14644
rect 2100 14588 2828 14644
rect 2884 14588 2894 14644
rect 14018 14588 14028 14644
rect 14084 14588 14924 14644
rect 14980 14588 14990 14644
rect 18060 14588 19740 14644
rect 19796 14588 19806 14644
rect 18060 14532 18116 14588
rect 20132 14532 20188 14644
rect 20244 14588 20254 14644
rect 22530 14588 22540 14644
rect 22596 14588 23212 14644
rect 23268 14588 24892 14644
rect 24948 14588 24958 14644
rect 28690 14588 28700 14644
rect 28756 14588 29260 14644
rect 29316 14588 30828 14644
rect 30884 14588 31724 14644
rect 31780 14588 31790 14644
rect 34962 14588 34972 14644
rect 35028 14588 36540 14644
rect 36596 14588 36606 14644
rect 9874 14476 9884 14532
rect 9940 14476 10444 14532
rect 10500 14476 10510 14532
rect 12002 14476 12012 14532
rect 12068 14476 12796 14532
rect 12852 14476 13468 14532
rect 13524 14476 13534 14532
rect 17378 14476 17388 14532
rect 17444 14476 18060 14532
rect 18116 14476 18126 14532
rect 19058 14476 19068 14532
rect 19124 14476 20188 14532
rect 6850 14364 6860 14420
rect 6916 14364 7420 14420
rect 7476 14364 7486 14420
rect 18834 14364 18844 14420
rect 18900 14364 20412 14420
rect 20468 14364 20478 14420
rect 24220 14308 24276 14588
rect 29362 14476 29372 14532
rect 29428 14476 29932 14532
rect 29988 14476 30380 14532
rect 30436 14476 30446 14532
rect 34402 14476 34412 14532
rect 34468 14476 39004 14532
rect 39060 14476 39452 14532
rect 39508 14476 40908 14532
rect 40964 14476 41580 14532
rect 41636 14476 41646 14532
rect 30146 14364 30156 14420
rect 30212 14364 30828 14420
rect 30884 14364 32060 14420
rect 32116 14364 32126 14420
rect 42914 14364 42924 14420
rect 42980 14364 43820 14420
rect 43876 14364 43886 14420
rect 1810 14252 1820 14308
rect 1876 14252 4844 14308
rect 4900 14252 4910 14308
rect 6598 14252 6636 14308
rect 6692 14252 6702 14308
rect 12450 14252 12460 14308
rect 12516 14252 14588 14308
rect 14644 14252 14654 14308
rect 16594 14252 16604 14308
rect 16660 14252 17388 14308
rect 17444 14252 17454 14308
rect 24210 14252 24220 14308
rect 24276 14252 24286 14308
rect 29586 14252 29596 14308
rect 29652 14252 30492 14308
rect 30548 14252 30558 14308
rect 40226 14252 40236 14308
rect 40292 14252 42812 14308
rect 42868 14252 42878 14308
rect 2258 14140 2268 14196
rect 2324 14140 3164 14196
rect 3220 14140 3724 14196
rect 3780 14140 3836 14196
rect 3892 14140 3902 14196
rect 10546 14140 10556 14196
rect 10612 14140 11228 14196
rect 11284 14140 11294 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 27122 14028 27132 14084
rect 27188 14028 28364 14084
rect 28420 14028 28430 14084
rect 18386 13916 18396 13972
rect 18452 13916 19852 13972
rect 19908 13916 19918 13972
rect 20066 13916 20076 13972
rect 20132 13916 22652 13972
rect 22708 13916 22718 13972
rect 23426 13916 23436 13972
rect 23492 13916 24668 13972
rect 24724 13916 24734 13972
rect 5954 13804 5964 13860
rect 6020 13804 6524 13860
rect 6580 13804 6972 13860
rect 7028 13804 7038 13860
rect 12226 13804 12236 13860
rect 12292 13804 13580 13860
rect 13636 13804 14140 13860
rect 14196 13804 14206 13860
rect 19506 13804 19516 13860
rect 19572 13804 20188 13860
rect 20244 13804 20254 13860
rect 22978 13804 22988 13860
rect 23044 13804 23324 13860
rect 23380 13804 23390 13860
rect 32050 13692 32060 13748
rect 32116 13692 33292 13748
rect 33348 13692 34076 13748
rect 34132 13692 34142 13748
rect 37986 13692 37996 13748
rect 38052 13692 39900 13748
rect 39956 13692 39966 13748
rect 6178 13580 6188 13636
rect 6244 13580 6748 13636
rect 6804 13580 6814 13636
rect 9622 13580 9660 13636
rect 9716 13580 11116 13636
rect 11172 13580 11182 13636
rect 25106 13580 25116 13636
rect 25172 13580 26684 13636
rect 26740 13580 27132 13636
rect 27188 13580 28028 13636
rect 28084 13580 28094 13636
rect 1698 13468 1708 13524
rect 1764 13468 3052 13524
rect 3108 13468 3118 13524
rect 6934 13468 6972 13524
rect 7028 13468 7038 13524
rect 11666 13468 11676 13524
rect 11732 13468 11900 13524
rect 11956 13468 12908 13524
rect 12964 13468 12974 13524
rect 13906 13468 13916 13524
rect 13972 13468 14756 13524
rect 15362 13468 15372 13524
rect 15428 13468 17388 13524
rect 17444 13468 17454 13524
rect 22530 13468 22540 13524
rect 22596 13468 24108 13524
rect 24164 13468 24174 13524
rect 14700 13412 14756 13468
rect 14690 13356 14700 13412
rect 14756 13356 14766 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 6374 13244 6412 13300
rect 6468 13244 6478 13300
rect 16930 13132 16940 13188
rect 16996 13132 17724 13188
rect 17780 13132 17790 13188
rect 21746 13132 21756 13188
rect 21812 13132 23996 13188
rect 24052 13132 24062 13188
rect 29922 13132 29932 13188
rect 29988 13132 31948 13188
rect 32004 13132 35644 13188
rect 35700 13132 36764 13188
rect 36820 13132 36830 13188
rect 2482 13020 2492 13076
rect 2548 13020 3388 13076
rect 3444 13020 3454 13076
rect 6822 13020 6860 13076
rect 6916 13020 6926 13076
rect 8428 13020 14028 13076
rect 14084 13020 14094 13076
rect 32274 13020 32284 13076
rect 32340 13020 33068 13076
rect 33124 13020 33404 13076
rect 33460 13020 34076 13076
rect 34132 13020 34142 13076
rect 35756 13020 35868 13076
rect 35924 13020 35934 13076
rect 2370 12908 2380 12964
rect 2436 12908 2828 12964
rect 2884 12908 3724 12964
rect 3780 12908 4284 12964
rect 4340 12908 4350 12964
rect 4946 12908 4956 12964
rect 5012 12908 5852 12964
rect 5908 12908 6076 12964
rect 6132 12908 6142 12964
rect 0 12852 400 12880
rect 8428 12852 8484 13020
rect 8642 12908 8652 12964
rect 8708 12908 9548 12964
rect 9604 12908 10444 12964
rect 10500 12908 10510 12964
rect 0 12796 1708 12852
rect 1764 12796 1932 12852
rect 1988 12796 1998 12852
rect 2482 12796 2492 12852
rect 2548 12796 8484 12852
rect 9426 12796 9436 12852
rect 9492 12796 9996 12852
rect 10052 12796 10062 12852
rect 31602 12796 31612 12852
rect 31668 12796 32508 12852
rect 32564 12796 32574 12852
rect 0 12768 400 12796
rect 5170 12684 5180 12740
rect 5236 12684 6076 12740
rect 6132 12684 6244 12740
rect 26002 12684 26012 12740
rect 26068 12684 27356 12740
rect 27412 12684 27422 12740
rect 29586 12684 29596 12740
rect 29652 12684 30380 12740
rect 30436 12684 30446 12740
rect 6188 12516 6244 12684
rect 35756 12628 35812 13020
rect 11778 12572 11788 12628
rect 11844 12572 12236 12628
rect 12292 12572 12302 12628
rect 35746 12572 35756 12628
rect 35812 12572 35822 12628
rect 36054 12572 36092 12628
rect 36148 12572 36158 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 6178 12460 6188 12516
rect 6244 12460 6254 12516
rect 6374 12460 6412 12516
rect 6468 12460 6478 12516
rect 12114 12460 12124 12516
rect 12180 12460 13132 12516
rect 13188 12460 13198 12516
rect 21858 12460 21868 12516
rect 21924 12460 22652 12516
rect 22708 12460 22718 12516
rect 35830 12460 35868 12516
rect 35924 12460 35934 12516
rect 10658 12348 10668 12404
rect 10724 12348 11340 12404
rect 11396 12348 11406 12404
rect 14242 12348 14252 12404
rect 14308 12348 15260 12404
rect 15316 12348 15932 12404
rect 15988 12348 17612 12404
rect 17668 12348 28588 12404
rect 28644 12348 29932 12404
rect 29988 12348 29998 12404
rect 4274 12236 4284 12292
rect 4340 12236 5180 12292
rect 5236 12236 6748 12292
rect 6804 12236 7308 12292
rect 7364 12236 7374 12292
rect 11554 12236 11564 12292
rect 11620 12236 12572 12292
rect 12628 12236 12638 12292
rect 29698 12236 29708 12292
rect 29764 12236 30940 12292
rect 30996 12236 33236 12292
rect 33180 12180 33236 12236
rect 4722 12124 4732 12180
rect 4788 12124 5740 12180
rect 5796 12124 5806 12180
rect 6066 12124 6076 12180
rect 6132 12124 6524 12180
rect 6580 12124 6590 12180
rect 18610 12124 18620 12180
rect 18676 12124 19180 12180
rect 19236 12124 19246 12180
rect 20132 12124 21420 12180
rect 21476 12124 21486 12180
rect 21858 12124 21868 12180
rect 21924 12124 23100 12180
rect 23156 12124 25228 12180
rect 25284 12124 25294 12180
rect 33170 12124 33180 12180
rect 33236 12124 33404 12180
rect 33460 12124 33740 12180
rect 33796 12124 33806 12180
rect 20132 12068 20188 12124
rect 4610 12012 4620 12068
rect 4676 12012 5068 12068
rect 5124 12012 5134 12068
rect 19058 12012 19068 12068
rect 19124 12012 20188 12068
rect 5394 11900 5404 11956
rect 5460 11900 5852 11956
rect 5908 11900 7196 11956
rect 7252 11900 7262 11956
rect 8530 11900 8540 11956
rect 8596 11900 9660 11956
rect 9716 11900 11564 11956
rect 11620 11900 11630 11956
rect 6850 11788 6860 11844
rect 6916 11788 6926 11844
rect 12002 11788 12012 11844
rect 12068 11788 12628 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 6860 11732 6916 11788
rect 4844 11676 6636 11732
rect 6692 11676 6702 11732
rect 6860 11676 7756 11732
rect 7812 11676 8092 11732
rect 8148 11676 9324 11732
rect 9380 11676 9390 11732
rect 11890 11676 11900 11732
rect 11956 11676 12348 11732
rect 12404 11676 12414 11732
rect 4844 11620 4900 11676
rect 12572 11620 12628 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 14466 11676 14476 11732
rect 14532 11676 15596 11732
rect 15652 11676 17836 11732
rect 17892 11676 18732 11732
rect 18788 11676 19068 11732
rect 19124 11676 19134 11732
rect 23314 11676 23324 11732
rect 23380 11676 25116 11732
rect 25172 11676 25182 11732
rect 3938 11564 3948 11620
rect 4004 11564 4900 11620
rect 5618 11564 5628 11620
rect 5684 11564 6524 11620
rect 6580 11564 6590 11620
rect 12572 11564 14364 11620
rect 14420 11564 14430 11620
rect 29922 11564 29932 11620
rect 29988 11564 30268 11620
rect 30324 11564 30334 11620
rect 5058 11452 5068 11508
rect 5124 11452 5516 11508
rect 5572 11452 6860 11508
rect 6916 11452 6926 11508
rect 7858 11452 7868 11508
rect 7924 11452 8652 11508
rect 8708 11452 8718 11508
rect 11330 11452 11340 11508
rect 11396 11452 12572 11508
rect 12628 11452 12638 11508
rect 12898 11452 12908 11508
rect 12964 11452 14140 11508
rect 14196 11452 14206 11508
rect 22642 11452 22652 11508
rect 22708 11452 24164 11508
rect 24434 11452 24444 11508
rect 24500 11452 25452 11508
rect 25508 11452 25518 11508
rect 34514 11452 34524 11508
rect 34580 11452 35084 11508
rect 35140 11452 35150 11508
rect 24108 11396 24164 11452
rect 6178 11340 6188 11396
rect 6244 11340 6972 11396
rect 7028 11340 7038 11396
rect 7410 11340 7420 11396
rect 7476 11340 8316 11396
rect 8372 11340 8382 11396
rect 23314 11340 23324 11396
rect 23380 11340 23390 11396
rect 24098 11340 24108 11396
rect 24164 11340 25900 11396
rect 25956 11340 28252 11396
rect 28308 11340 28318 11396
rect 35298 11340 35308 11396
rect 35364 11340 35756 11396
rect 35812 11340 39452 11396
rect 39508 11340 39518 11396
rect 4834 11228 4844 11284
rect 4900 11228 5852 11284
rect 5908 11228 6636 11284
rect 6692 11228 6702 11284
rect 8754 11228 8764 11284
rect 8820 11228 10220 11284
rect 10276 11228 10892 11284
rect 10948 11228 10958 11284
rect 23324 11172 23380 11340
rect 21634 11116 21644 11172
rect 21700 11116 22764 11172
rect 22820 11116 23380 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 23324 10948 23380 11116
rect 23314 10892 23324 10948
rect 23380 10892 23390 10948
rect 2706 10780 2716 10836
rect 2772 10780 3388 10836
rect 3444 10780 3948 10836
rect 4004 10780 4014 10836
rect 39106 10780 39116 10836
rect 39172 10780 40908 10836
rect 40964 10780 40974 10836
rect 6962 10668 6972 10724
rect 7028 10668 10668 10724
rect 10724 10668 10734 10724
rect 14578 10668 14588 10724
rect 14644 10668 16604 10724
rect 16660 10668 34636 10724
rect 34692 10668 34972 10724
rect 35028 10668 38556 10724
rect 38612 10668 38622 10724
rect 38882 10668 38892 10724
rect 38948 10668 39788 10724
rect 39844 10668 39854 10724
rect 5282 10556 5292 10612
rect 5348 10556 6076 10612
rect 6132 10556 6860 10612
rect 6916 10556 7420 10612
rect 7476 10556 7486 10612
rect 12562 10556 12572 10612
rect 12628 10556 13468 10612
rect 13524 10556 13534 10612
rect 14242 10556 14252 10612
rect 14308 10556 15820 10612
rect 15876 10556 15886 10612
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 6738 10108 6748 10164
rect 6804 10108 7756 10164
rect 7812 10108 7822 10164
rect 39554 9996 39564 10052
rect 39620 9996 40572 10052
rect 40628 9996 40638 10052
rect 9538 9884 9548 9940
rect 9604 9884 11900 9940
rect 11956 9884 12908 9940
rect 12964 9884 12974 9940
rect 15092 9884 15260 9940
rect 15316 9884 15326 9940
rect 23538 9884 23548 9940
rect 23604 9884 24220 9940
rect 24276 9884 24286 9940
rect 27906 9884 27916 9940
rect 27972 9884 28924 9940
rect 28980 9884 31388 9940
rect 31444 9884 31454 9940
rect 40114 9884 40124 9940
rect 40180 9884 43036 9940
rect 43092 9884 43102 9940
rect 15092 9828 15148 9884
rect 11554 9772 11564 9828
rect 11620 9772 15148 9828
rect 29362 9772 29372 9828
rect 29428 9772 30492 9828
rect 30548 9772 31724 9828
rect 31780 9772 31790 9828
rect 12114 9660 12124 9716
rect 12180 9660 12796 9716
rect 12852 9660 14028 9716
rect 14084 9660 14094 9716
rect 26562 9660 26572 9716
rect 26628 9660 26908 9716
rect 26852 9604 26908 9660
rect 10098 9548 10108 9604
rect 10164 9548 10780 9604
rect 10836 9548 15372 9604
rect 15428 9548 15438 9604
rect 26852 9548 27356 9604
rect 27412 9548 28588 9604
rect 28644 9548 28924 9604
rect 28980 9548 30044 9604
rect 30100 9548 30940 9604
rect 30996 9548 31006 9604
rect 3490 9436 3500 9492
rect 3556 9436 3566 9492
rect 3500 9268 3556 9436
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 2706 9212 2716 9268
rect 2772 9212 3556 9268
rect 3332 9044 3388 9212
rect 43652 9156 43708 9268
rect 43764 9212 43774 9268
rect 5842 9100 5852 9156
rect 5908 9100 7084 9156
rect 7140 9100 7150 9156
rect 10098 9100 10108 9156
rect 10164 9100 11060 9156
rect 37314 9100 37324 9156
rect 37380 9100 41020 9156
rect 41076 9100 43708 9156
rect 11004 9044 11060 9100
rect 3332 8988 3612 9044
rect 3668 8988 3678 9044
rect 5954 8988 5964 9044
rect 6020 8988 6524 9044
rect 6580 8988 6590 9044
rect 7410 8988 7420 9044
rect 7476 8988 8204 9044
rect 8260 8988 8270 9044
rect 10994 8988 11004 9044
rect 11060 8988 14924 9044
rect 14980 8988 14990 9044
rect 16594 8988 16604 9044
rect 16660 8988 17948 9044
rect 18004 8988 18014 9044
rect 26898 8988 26908 9044
rect 26964 8988 27804 9044
rect 27860 8988 27870 9044
rect 31490 8988 31500 9044
rect 31556 8988 32060 9044
rect 32116 8988 32126 9044
rect 33394 8988 33404 9044
rect 33460 8988 33628 9044
rect 33684 8988 33694 9044
rect 10546 8876 10556 8932
rect 10612 8876 11676 8932
rect 11732 8876 13356 8932
rect 13412 8876 15148 8932
rect 15204 8876 15214 8932
rect 27122 8876 27132 8932
rect 27188 8876 27468 8932
rect 27524 8876 27534 8932
rect 36306 8876 36316 8932
rect 36372 8876 37100 8932
rect 37156 8876 37548 8932
rect 37604 8876 37614 8932
rect 2706 8652 2716 8708
rect 2772 8652 3276 8708
rect 3332 8652 3342 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 20178 8540 20188 8596
rect 20244 8540 20748 8596
rect 20804 8540 21868 8596
rect 21924 8540 21934 8596
rect 12002 8428 12012 8484
rect 12068 8428 12908 8484
rect 12964 8428 12974 8484
rect 35970 8428 35980 8484
rect 36036 8428 37324 8484
rect 37380 8428 37390 8484
rect 4498 8316 4508 8372
rect 4564 8316 13916 8372
rect 13972 8316 14588 8372
rect 14644 8316 14654 8372
rect 17938 8316 17948 8372
rect 18004 8316 18844 8372
rect 18900 8316 20076 8372
rect 20132 8316 20142 8372
rect 33506 8316 33516 8372
rect 33572 8316 34412 8372
rect 34468 8316 34478 8372
rect 4162 8204 4172 8260
rect 4228 8204 4956 8260
rect 5012 8204 5852 8260
rect 5908 8204 6748 8260
rect 6804 8204 7196 8260
rect 7252 8204 7262 8260
rect 32050 8204 32060 8260
rect 32116 8204 35756 8260
rect 35812 8204 36316 8260
rect 36372 8204 37324 8260
rect 37380 8204 37390 8260
rect 29586 8092 29596 8148
rect 29652 8092 31164 8148
rect 31220 8092 31612 8148
rect 31668 8092 32732 8148
rect 32788 8092 33404 8148
rect 33460 8092 35644 8148
rect 35700 8092 35980 8148
rect 36036 8092 36046 8148
rect 36194 8092 36204 8148
rect 36260 8092 36988 8148
rect 37044 8092 37054 8148
rect 1922 7980 1932 8036
rect 1988 7980 2604 8036
rect 2660 7980 2670 8036
rect 0 7924 400 7952
rect 0 7868 1820 7924
rect 1876 7868 1886 7924
rect 0 7840 400 7868
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 7858 7756 7868 7812
rect 7924 7756 9100 7812
rect 9156 7756 9772 7812
rect 9828 7756 9838 7812
rect 15138 7756 15148 7812
rect 15204 7756 15372 7812
rect 15428 7756 15438 7812
rect 7186 7644 7196 7700
rect 7252 7644 8428 7700
rect 8484 7644 8494 7700
rect 9314 7644 9324 7700
rect 9380 7644 10444 7700
rect 10500 7644 10510 7700
rect 6514 7532 6524 7588
rect 6580 7532 7756 7588
rect 7812 7532 7822 7588
rect 9874 7532 9884 7588
rect 9940 7532 11340 7588
rect 11396 7532 11406 7588
rect 4498 7420 4508 7476
rect 4564 7420 6412 7476
rect 6468 7420 6478 7476
rect 6626 7420 6636 7476
rect 6692 7420 8428 7476
rect 8484 7420 8494 7476
rect 12674 7420 12684 7476
rect 12740 7420 14364 7476
rect 14420 7420 16044 7476
rect 16100 7420 16110 7476
rect 8306 7308 8316 7364
rect 8372 7308 10220 7364
rect 10276 7308 10286 7364
rect 3042 7196 3052 7252
rect 3108 7196 5404 7252
rect 5460 7196 5470 7252
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 37202 6972 37212 7028
rect 37268 6972 38108 7028
rect 38164 6972 38892 7028
rect 38948 6972 38958 7028
rect 2258 6860 2268 6916
rect 2324 6860 2334 6916
rect 26898 6860 26908 6916
rect 26964 6860 27580 6916
rect 27636 6860 27646 6916
rect 2268 6692 2324 6860
rect 9548 6748 10108 6804
rect 10164 6748 10174 6804
rect 12226 6748 12236 6804
rect 12292 6748 12684 6804
rect 12740 6748 12750 6804
rect 1698 6636 1708 6692
rect 1764 6636 2044 6692
rect 2100 6636 2110 6692
rect 2268 6636 3836 6692
rect 3892 6636 3902 6692
rect 9548 6580 9604 6748
rect 9986 6636 9996 6692
rect 10052 6636 10892 6692
rect 10948 6636 13356 6692
rect 13412 6636 13422 6692
rect 13794 6636 13804 6692
rect 13860 6636 14252 6692
rect 14308 6636 14318 6692
rect 19058 6636 19068 6692
rect 19124 6636 20300 6692
rect 20356 6636 21420 6692
rect 21476 6636 21486 6692
rect 27234 6636 27244 6692
rect 27300 6636 27916 6692
rect 27972 6636 27982 6692
rect 2930 6524 2940 6580
rect 2996 6524 3388 6580
rect 3444 6524 4508 6580
rect 4564 6524 4574 6580
rect 5058 6524 5068 6580
rect 5124 6524 5964 6580
rect 6020 6524 6030 6580
rect 7746 6524 7756 6580
rect 7812 6524 8540 6580
rect 8596 6524 8606 6580
rect 9538 6524 9548 6580
rect 9604 6524 9614 6580
rect 13010 6524 13020 6580
rect 13076 6524 13692 6580
rect 13748 6524 13758 6580
rect 13916 6468 13972 6636
rect 17490 6524 17500 6580
rect 17556 6524 19404 6580
rect 19460 6524 20748 6580
rect 20804 6524 20814 6580
rect 1810 6412 1820 6468
rect 1876 6412 2268 6468
rect 2324 6412 3948 6468
rect 4004 6412 4284 6468
rect 4340 6412 4350 6468
rect 7298 6412 7308 6468
rect 7364 6412 9100 6468
rect 9156 6412 9166 6468
rect 12562 6412 12572 6468
rect 12628 6412 13972 6468
rect 18274 6412 18284 6468
rect 18340 6412 18620 6468
rect 18676 6412 19516 6468
rect 19572 6412 19582 6468
rect 11778 6300 11788 6356
rect 11844 6300 13804 6356
rect 13860 6300 13870 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 14578 6188 14588 6244
rect 14644 6188 15484 6244
rect 15540 6188 15550 6244
rect 7522 6076 7532 6132
rect 7588 6076 8092 6132
rect 8148 6076 11228 6132
rect 11284 6076 11294 6132
rect 26852 6076 27244 6132
rect 27300 6076 27692 6132
rect 27748 6076 27758 6132
rect 28802 6076 28812 6132
rect 28868 6076 30380 6132
rect 30436 6076 30940 6132
rect 30996 6076 31006 6132
rect 8866 5964 8876 6020
rect 8932 5964 10220 6020
rect 10276 5964 10948 6020
rect 12450 5964 12460 6020
rect 12516 5964 13132 6020
rect 13188 5964 14476 6020
rect 14532 5964 14542 6020
rect 23090 5964 23100 6020
rect 23156 5964 25788 6020
rect 25844 5964 26684 6020
rect 26740 5964 26750 6020
rect 10892 5908 10948 5964
rect 26852 5908 26908 6076
rect 29586 5964 29596 6020
rect 29652 5964 30716 6020
rect 30772 5964 30782 6020
rect 6626 5852 6636 5908
rect 6692 5852 7644 5908
rect 7700 5852 7980 5908
rect 8036 5852 8046 5908
rect 9314 5852 9324 5908
rect 9380 5852 9884 5908
rect 9940 5852 9950 5908
rect 10882 5852 10892 5908
rect 10948 5852 10958 5908
rect 13682 5852 13692 5908
rect 13748 5852 14700 5908
rect 14756 5852 14766 5908
rect 18610 5852 18620 5908
rect 18676 5852 19964 5908
rect 20020 5852 20030 5908
rect 23874 5852 23884 5908
rect 23940 5852 26908 5908
rect 11106 5740 11116 5796
rect 11172 5740 14924 5796
rect 14980 5740 14990 5796
rect 25218 5740 25228 5796
rect 25284 5740 26012 5796
rect 26068 5740 26078 5796
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 20132 5404 28140 5460
rect 28196 5404 28206 5460
rect 20132 5348 20188 5404
rect 10322 5292 10332 5348
rect 10388 5292 12460 5348
rect 12516 5292 12526 5348
rect 14802 5292 14812 5348
rect 14868 5292 15708 5348
rect 15764 5292 18732 5348
rect 18788 5292 20188 5348
rect 21522 5292 21532 5348
rect 21588 5292 23324 5348
rect 23380 5292 23390 5348
rect 33058 5292 33068 5348
rect 33124 5292 33516 5348
rect 33572 5292 34076 5348
rect 34132 5292 34972 5348
rect 35028 5292 35644 5348
rect 35700 5292 35710 5348
rect 7410 5180 7420 5236
rect 7476 5180 8876 5236
rect 8932 5180 8942 5236
rect 12338 5180 12348 5236
rect 12404 5180 13804 5236
rect 13860 5180 13870 5236
rect 15474 5180 15484 5236
rect 15540 5180 15820 5236
rect 15876 5180 17724 5236
rect 17780 5180 17790 5236
rect 20402 5180 20412 5236
rect 20468 5180 22652 5236
rect 22708 5180 22718 5236
rect 34290 5180 34300 5236
rect 34356 5180 34748 5236
rect 34804 5180 36092 5236
rect 36148 5180 36158 5236
rect 6402 5068 6412 5124
rect 6468 5068 8316 5124
rect 8372 5068 8382 5124
rect 12226 5068 12236 5124
rect 12292 5068 13468 5124
rect 13524 5068 13534 5124
rect 19618 5068 19628 5124
rect 19684 5068 21868 5124
rect 21924 5068 23100 5124
rect 23156 5068 23166 5124
rect 24434 5068 24444 5124
rect 24500 5068 25452 5124
rect 25508 5068 25518 5124
rect 25778 5068 25788 5124
rect 25844 5068 26460 5124
rect 26516 5068 27132 5124
rect 27188 5068 28532 5124
rect 28476 5012 28532 5068
rect 6066 4956 6076 5012
rect 6132 4956 10332 5012
rect 10388 4956 10398 5012
rect 23426 4956 23436 5012
rect 23492 4956 24220 5012
rect 24276 4956 24286 5012
rect 28476 4956 30156 5012
rect 30212 4956 30940 5012
rect 30996 4956 33628 5012
rect 33684 4956 33694 5012
rect 35858 4956 35868 5012
rect 35924 4956 36988 5012
rect 37044 4956 37054 5012
rect 7522 4844 7532 4900
rect 7588 4844 8764 4900
rect 8820 4844 8830 4900
rect 15138 4844 15148 4900
rect 15204 4844 16492 4900
rect 16548 4844 17052 4900
rect 17108 4844 17500 4900
rect 17556 4844 17566 4900
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 7186 4620 7196 4676
rect 7252 4620 8204 4676
rect 8260 4620 9660 4676
rect 9716 4620 9726 4676
rect 7746 4508 7756 4564
rect 7812 4508 8876 4564
rect 8932 4508 8942 4564
rect 10322 4508 10332 4564
rect 10388 4508 10668 4564
rect 10724 4508 11788 4564
rect 11844 4508 11854 4564
rect 18386 4508 18396 4564
rect 18452 4508 33740 4564
rect 33796 4508 33806 4564
rect 10434 4396 10444 4452
rect 10500 4396 12124 4452
rect 12180 4396 12190 4452
rect 24658 4396 24668 4452
rect 24724 4396 26012 4452
rect 26068 4396 26078 4452
rect 32498 4396 32508 4452
rect 32564 4396 33852 4452
rect 33908 4396 33918 4452
rect 35970 4396 35980 4452
rect 36036 4396 36204 4452
rect 36260 4396 36764 4452
rect 36820 4396 38668 4452
rect 38612 4340 38668 4396
rect 13234 4284 13244 4340
rect 13300 4284 15148 4340
rect 15204 4284 15214 4340
rect 17490 4284 17500 4340
rect 17556 4284 18284 4340
rect 18340 4284 18350 4340
rect 38612 4284 39116 4340
rect 39172 4284 39788 4340
rect 39844 4284 39854 4340
rect 14690 4172 14700 4228
rect 14756 4172 19068 4228
rect 19124 4172 20300 4228
rect 20356 4172 20366 4228
rect 27458 4172 27468 4228
rect 27524 4172 28140 4228
rect 28196 4172 28206 4228
rect 35746 4172 35756 4228
rect 35812 4172 38444 4228
rect 38500 4172 38510 4228
rect 8866 4060 8876 4116
rect 8932 4060 10444 4116
rect 10500 4060 10510 4116
rect 33954 4060 33964 4116
rect 34020 4060 36316 4116
rect 36372 4060 36382 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 7382 3724 7420 3780
rect 7476 3724 7486 3780
rect 8418 3724 8428 3780
rect 8484 3724 11340 3780
rect 11396 3724 11406 3780
rect 33730 3724 33740 3780
rect 33796 3724 34412 3780
rect 34468 3724 34478 3780
rect 3602 3612 3612 3668
rect 3668 3612 4620 3668
rect 4676 3612 4686 3668
rect 18050 3612 18060 3668
rect 18116 3612 18956 3668
rect 19012 3612 19022 3668
rect 1698 3276 1708 3332
rect 1764 3276 3388 3332
rect 3444 3276 4956 3332
rect 5012 3276 6748 3332
rect 6804 3276 6814 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 0 2996 400 3024
rect 0 2940 5852 2996
rect 5908 2940 5918 2996
rect 18274 2940 18284 2996
rect 18340 2940 19180 2996
rect 19236 2940 19628 2996
rect 19684 2940 19694 2996
rect 0 2912 400 2940
rect 24220 2828 25788 2884
rect 25844 2828 25854 2884
rect 24220 2772 24276 2828
rect 23426 2716 23436 2772
rect 23492 2716 24220 2772
rect 24276 2716 24286 2772
rect 25330 2716 25340 2772
rect 25396 2716 26796 2772
rect 26852 2716 26862 2772
rect 7298 2492 7308 2548
rect 7364 2492 10108 2548
rect 10164 2492 10174 2548
rect 4466 2324 4476 2380
rect 4532 2324 4580 2380
rect 4636 2324 4684 2380
rect 4740 2324 4750 2380
rect 35186 2324 35196 2380
rect 35252 2324 35300 2380
rect 35356 2324 35404 2380
rect 35460 2324 35470 2380
rect 19826 1540 19836 1596
rect 19892 1540 19940 1596
rect 19996 1540 20044 1596
rect 20100 1540 20110 1596
<< via3 >>
rect 19836 78372 19892 78428
rect 19940 78372 19996 78428
rect 20044 78372 20100 78428
rect 4476 77588 4532 77644
rect 4580 77588 4636 77644
rect 4684 77588 4740 77644
rect 35196 77588 35252 77644
rect 35300 77588 35356 77644
rect 35404 77588 35460 77644
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 22652 67564 22708 67620
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 28700 63868 28756 63924
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 34860 62860 34916 62916
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 22652 59052 22708 59108
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 25564 58268 25620 58324
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 25564 57596 25620 57652
rect 23100 57260 23156 57316
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 25676 56924 25732 56980
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 23100 55020 23156 55076
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 25676 53116 25732 53172
rect 39900 53116 39956 53172
rect 4284 52892 4340 52948
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 39900 51996 39956 52052
rect 4284 51884 4340 51940
rect 31052 51884 31108 51940
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 29484 50652 29540 50708
rect 30156 50540 30212 50596
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 31276 50092 31332 50148
rect 30156 49756 30212 49812
rect 31052 49532 31108 49588
rect 31276 49532 31332 49588
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 3388 48860 3444 48916
rect 23100 48748 23156 48804
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 28924 48300 28980 48356
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 5180 46732 5236 46788
rect 3276 46396 3332 46452
rect 30716 46396 30772 46452
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 28812 45500 28868 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 2268 44492 2324 44548
rect 35980 44380 36036 44436
rect 29372 44268 29428 44324
rect 29036 44044 29092 44100
rect 29596 44044 29652 44100
rect 3388 43932 3444 43988
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 22428 43708 22484 43764
rect 29820 43708 29876 43764
rect 38332 43484 38388 43540
rect 4956 43372 5012 43428
rect 4060 43148 4116 43204
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 33964 43260 34020 43316
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 4060 42364 4116 42420
rect 29260 42364 29316 42420
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 2492 42140 2548 42196
rect 28812 42140 28868 42196
rect 29708 42140 29764 42196
rect 4956 42028 5012 42084
rect 34300 41916 34356 41972
rect 22428 41580 22484 41636
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 35980 41468 36036 41524
rect 30828 40908 30884 40964
rect 28924 40796 28980 40852
rect 29260 40796 29316 40852
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 2604 40572 2660 40628
rect 2492 40348 2548 40404
rect 28924 40012 28980 40068
rect 29596 40012 29652 40068
rect 29820 40012 29876 40068
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 5180 39788 5236 39844
rect 27580 39452 27636 39508
rect 29596 39340 29652 39396
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 26460 39116 26516 39172
rect 2604 38556 2660 38612
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 2268 38220 2324 38276
rect 30492 38220 30548 38276
rect 29372 38108 29428 38164
rect 29036 37996 29092 38052
rect 34300 37884 34356 37940
rect 30716 37772 30772 37828
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 3276 37548 3332 37604
rect 28812 37548 28868 37604
rect 34972 37212 35028 37268
rect 27580 36988 27636 37044
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 38332 36428 38388 36484
rect 30828 36316 30884 36372
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 26460 35980 26516 36036
rect 34300 35420 34356 35476
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 34972 35084 35028 35140
rect 6636 34860 6692 34916
rect 8204 34636 8260 34692
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 15484 34188 15540 34244
rect 8316 34076 8372 34132
rect 6972 33740 7028 33796
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 6300 33628 6356 33684
rect 29484 33404 29540 33460
rect 36092 33180 36148 33236
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 31276 32396 31332 32452
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 33628 31948 33684 32004
rect 38108 31724 38164 31780
rect 8204 31500 8260 31556
rect 34860 31500 34916 31556
rect 34972 31388 35028 31444
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 34076 31164 34132 31220
rect 7084 30940 7140 30996
rect 26348 30828 26404 30884
rect 33852 30940 33908 30996
rect 28812 30716 28868 30772
rect 33740 30604 33796 30660
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 34188 30492 34244 30548
rect 33852 30268 33908 30324
rect 34188 30156 34244 30212
rect 33740 29820 33796 29876
rect 34076 29820 34132 29876
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 7084 29372 7140 29428
rect 33628 29372 33684 29428
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 29932 28700 29988 28756
rect 26348 28252 26404 28308
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 7532 28140 7588 28196
rect 6636 28028 6692 28084
rect 30492 28028 30548 28084
rect 32956 27692 33012 27748
rect 34860 27580 34916 27636
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 6524 27356 6580 27412
rect 29932 27356 29988 27412
rect 28700 27244 28756 27300
rect 7532 26908 7588 26964
rect 6300 26796 6356 26852
rect 8204 26796 8260 26852
rect 27020 26684 27076 26740
rect 38108 26684 38164 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 8316 26572 8372 26628
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 27020 25788 27076 25844
rect 29932 25228 29988 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 31276 25004 31332 25060
rect 32956 24892 33012 24948
rect 6300 24668 6356 24724
rect 36092 24556 36148 24612
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 7868 23996 7924 24052
rect 15484 23884 15540 23940
rect 29596 23884 29652 23940
rect 6972 23772 7028 23828
rect 6524 23548 6580 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 7868 23100 7924 23156
rect 6300 22876 6356 22932
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 33964 22428 34020 22484
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 36092 21532 36148 21588
rect 35980 21420 36036 21476
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 3836 21084 3892 21140
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 6860 19964 6916 20020
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 6636 18732 6692 18788
rect 5404 18508 5460 18564
rect 6076 18508 6132 18564
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 5404 17724 5460 17780
rect 6972 17724 7028 17780
rect 6076 17612 6132 17668
rect 31948 17724 32004 17780
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 29708 16940 29764 16996
rect 6636 16604 6692 16660
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 35980 15708 36036 15764
rect 35868 15260 35924 15316
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 6636 14252 6692 14308
rect 3836 14140 3892 14196
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 6972 13804 7028 13860
rect 9660 13580 9716 13636
rect 6972 13468 7028 13524
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 6412 13244 6468 13300
rect 31948 13132 32004 13188
rect 6860 13020 6916 13076
rect 6076 12684 6132 12740
rect 36092 12572 36148 12628
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 6412 12460 6468 12516
rect 35868 12460 35924 12516
rect 9660 11900 9716 11956
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 6636 11676 6692 11732
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 7420 11340 7476 11396
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 7420 3724 7476 3780
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 4476 2324 4532 2380
rect 4580 2324 4636 2380
rect 4684 2324 4740 2380
rect 35196 2324 35252 2380
rect 35300 2324 35356 2380
rect 35404 2324 35460 2380
rect 19836 1540 19892 1596
rect 19940 1540 19996 1596
rect 20044 1540 20100 1596
<< metal4 >>
rect 4448 77644 4768 78460
rect 4448 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4768 77644
rect 4448 76076 4768 77588
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4284 52948 4340 52958
rect 4284 51940 4340 52892
rect 4284 51874 4340 51884
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 3388 48916 3444 48926
rect 3276 46452 3332 46462
rect 2268 44548 2324 44558
rect 2268 38276 2324 44492
rect 2492 42196 2548 42206
rect 2492 40404 2548 42140
rect 2492 40338 2548 40348
rect 2604 40628 2660 40638
rect 2604 38612 2660 40572
rect 2604 38546 2660 38556
rect 2268 38210 2324 38220
rect 3276 37604 3332 46396
rect 3388 43988 3444 48860
rect 3388 43922 3444 43932
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 19808 78428 20128 78460
rect 19808 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20128 78428
rect 19808 76860 20128 78372
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 35168 77644 35488 78460
rect 35168 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35488 77644
rect 35168 76076 35488 77588
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 22652 67620 22708 67630
rect 22652 59108 22708 67564
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 22652 59042 22708 59052
rect 28700 63924 28756 63934
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 25564 58324 25620 58334
rect 25564 57652 25620 58268
rect 25564 57586 25620 57596
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 23100 57316 23156 57326
rect 23100 55076 23156 57260
rect 23100 48804 23156 55020
rect 25676 56980 25732 56990
rect 25676 53172 25732 56924
rect 25676 53106 25732 53116
rect 23100 48738 23156 48748
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4060 43204 4116 43214
rect 4060 42420 4116 43148
rect 4060 42354 4116 42364
rect 4448 43148 4768 44660
rect 5180 46788 5236 46798
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 3276 37538 3332 37548
rect 4448 41580 4768 43092
rect 4956 43428 5012 43438
rect 4956 42084 5012 43372
rect 4956 42018 5012 42028
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 5180 39844 5236 46732
rect 5180 39778 5236 39788
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 22428 43764 22484 43774
rect 22428 41636 22484 43708
rect 22428 41570 22484 41580
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 27580 39508 27636 39518
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 6636 34916 6692 34926
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 6300 33684 6356 33694
rect 6300 26852 6356 33628
rect 6636 28084 6692 34860
rect 8204 34692 8260 34702
rect 6636 28018 6692 28028
rect 6972 33796 7028 33806
rect 6300 26786 6356 26796
rect 6524 27412 6580 27422
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 6300 24724 6356 24734
rect 6300 22932 6356 24668
rect 6524 23604 6580 27356
rect 6972 23828 7028 33740
rect 8204 31556 8260 34636
rect 19808 34524 20128 36036
rect 26460 39172 26516 39182
rect 26460 36036 26516 39116
rect 27580 37044 27636 39452
rect 27580 36978 27636 36988
rect 26460 35970 26516 35980
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 15484 34244 15540 34254
rect 7084 30996 7140 31006
rect 7084 29428 7140 30940
rect 7084 29362 7140 29372
rect 7532 28196 7588 28206
rect 7532 26964 7588 28140
rect 7532 26898 7588 26908
rect 8204 26852 8260 31500
rect 8204 26786 8260 26796
rect 8316 34132 8372 34142
rect 8316 26628 8372 34076
rect 8316 26562 8372 26572
rect 6972 23762 7028 23772
rect 7868 24052 7924 24062
rect 6524 23538 6580 23548
rect 7868 23156 7924 23996
rect 15484 23940 15540 34188
rect 15484 23874 15540 23884
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 26348 30884 26404 30894
rect 26348 28308 26404 30828
rect 26348 28242 26404 28252
rect 19808 26684 20128 28196
rect 28700 27300 28756 63868
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 34860 62916 34916 62926
rect 34860 62188 34916 62860
rect 34860 62132 35028 62188
rect 31052 51940 31108 51950
rect 29484 50708 29540 50718
rect 28924 48356 28980 48366
rect 28812 45556 28868 45566
rect 28812 42196 28868 45500
rect 28812 42130 28868 42140
rect 28924 40852 28980 48300
rect 29372 44324 29428 44334
rect 28924 40068 28980 40796
rect 28924 40002 28980 40012
rect 29036 44100 29092 44110
rect 29036 38052 29092 44044
rect 29260 42420 29316 42430
rect 29260 40852 29316 42364
rect 29260 40786 29316 40796
rect 29372 38164 29428 44268
rect 29372 38098 29428 38108
rect 29036 37986 29092 37996
rect 28812 37604 28868 37614
rect 28812 30772 28868 37548
rect 29484 33460 29540 50652
rect 30156 50596 30212 50606
rect 30156 49812 30212 50540
rect 30156 49746 30212 49756
rect 31052 49588 31108 51884
rect 31052 49522 31108 49532
rect 31276 50148 31332 50158
rect 31276 49588 31332 50092
rect 31276 49522 31332 49532
rect 30716 46452 30772 46462
rect 29596 44100 29652 44110
rect 29596 40068 29652 44044
rect 29820 43764 29876 43774
rect 29596 40002 29652 40012
rect 29708 42196 29764 42206
rect 29484 33394 29540 33404
rect 29596 39396 29652 39406
rect 28812 30706 28868 30716
rect 28700 27234 28756 27244
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 27020 26740 27076 26750
rect 27020 25844 27076 26684
rect 27020 25778 27076 25788
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 7868 23090 7924 23100
rect 19808 23548 20128 25060
rect 29596 23940 29652 39340
rect 29596 23874 29652 23884
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 6300 22866 6356 22876
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 3836 21140 3892 21150
rect 3836 14196 3892 21084
rect 3836 14130 3892 14140
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 6860 20020 6916 20030
rect 6636 18788 6692 18798
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 5404 18564 5460 18574
rect 5404 17780 5460 18508
rect 5404 17714 5460 17724
rect 6076 18564 6132 18574
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 6076 17668 6132 18508
rect 6076 12740 6132 17612
rect 6636 16660 6692 18732
rect 6636 16594 6692 16604
rect 6636 14308 6692 14318
rect 6076 12674 6132 12684
rect 6412 13300 6468 13310
rect 6412 12516 6468 13244
rect 6412 12450 6468 12460
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 6636 11732 6692 14252
rect 6860 13076 6916 19964
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 6972 17780 7028 17790
rect 6972 13860 7028 17724
rect 6972 13524 7028 13804
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 29708 16996 29764 42140
rect 29820 40068 29876 43708
rect 29820 40002 29876 40012
rect 30492 38276 30548 38286
rect 29932 28756 29988 28766
rect 29932 27412 29988 28700
rect 30492 28084 30548 38220
rect 30716 37828 30772 46396
rect 33964 43316 34020 43326
rect 30716 37762 30772 37772
rect 30828 40964 30884 40974
rect 30828 36372 30884 40908
rect 30828 36306 30884 36316
rect 30492 28018 30548 28028
rect 31276 32452 31332 32462
rect 29932 25284 29988 27356
rect 29932 25218 29988 25228
rect 31276 25060 31332 32396
rect 33628 32004 33684 32014
rect 33628 29428 33684 31948
rect 33852 30996 33908 31006
rect 33740 30660 33796 30670
rect 33740 29876 33796 30604
rect 33852 30324 33908 30940
rect 33852 30258 33908 30268
rect 33740 29810 33796 29820
rect 33628 29362 33684 29372
rect 31276 24994 31332 25004
rect 32956 27748 33012 27758
rect 32956 24948 33012 27692
rect 32956 24882 33012 24892
rect 33964 22484 34020 43260
rect 34300 41972 34356 41982
rect 34300 37940 34356 41916
rect 34300 35476 34356 37884
rect 34972 37268 35028 62132
rect 34972 37202 35028 37212
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 39900 53172 39956 53182
rect 39900 52052 39956 53116
rect 39900 51986 39956 51996
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35980 44436 36036 44446
rect 35980 41524 36036 44380
rect 35980 41458 36036 41468
rect 38332 43540 38388 43550
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 34300 35410 34356 35420
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 38332 36484 38388 43484
rect 38332 36418 38388 36428
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 34972 35140 35028 35150
rect 34860 31556 34916 31566
rect 34076 31220 34132 31230
rect 34076 29876 34132 31164
rect 34188 30548 34244 30558
rect 34188 30212 34244 30492
rect 34188 30146 34244 30156
rect 34076 29810 34132 29820
rect 34860 27636 34916 31500
rect 34972 31444 35028 35084
rect 34972 31378 35028 31388
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 34860 27570 34916 27580
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 33964 22418 34020 22428
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 36092 33236 36148 33246
rect 36092 24612 36148 33180
rect 38108 31780 38164 31790
rect 38108 26740 38164 31724
rect 38108 26674 38164 26684
rect 36092 24546 36148 24556
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 36092 21588 36148 21598
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 29708 16930 29764 16940
rect 31948 17780 32004 17790
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 6972 13458 7028 13468
rect 9660 13636 9716 13646
rect 6860 13010 6916 13020
rect 9660 11956 9716 13580
rect 9660 11890 9716 11900
rect 19808 12572 20128 14084
rect 31948 13188 32004 17724
rect 31948 13122 32004 13132
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35980 21476 36036 21486
rect 35980 15764 36036 21420
rect 35980 15698 36036 15708
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 6636 11666 6692 11676
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 2380 4768 3892
rect 7420 11396 7476 11406
rect 7420 3780 7476 11340
rect 7420 3714 7476 3724
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 4448 2324 4476 2380
rect 4532 2324 4580 2380
rect 4636 2324 4684 2380
rect 4740 2324 4768 2380
rect 4448 1508 4768 2324
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 1596 20128 3108
rect 19808 1540 19836 1596
rect 19892 1540 19940 1596
rect 19996 1540 20044 1596
rect 20100 1540 20128 1596
rect 19808 1508 20128 1540
rect 35168 11788 35488 13300
rect 35868 15316 35924 15326
rect 35868 12516 35924 15260
rect 36092 12628 36148 21532
rect 36092 12562 36148 12572
rect 35868 12450 35924 12460
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 2380 35488 3892
rect 35168 2324 35196 2380
rect 35252 2324 35300 2380
rect 35356 2324 35404 2380
rect 35460 2324 35488 2380
rect 35168 1508 35488 2324
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _0812_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6608 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0813_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0814_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7952 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0815_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12656 0 -1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0816_
timestamp 1698431365
transform -1 0 14896 0 1 53312
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0817_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4032 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0818_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7056 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0819_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7840 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0820_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0821_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9296 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0822_
timestamp 1698431365
transform 1 0 2800 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0823_
timestamp 1698431365
transform -1 0 3584 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0824_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4704 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _0825_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4704 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _0826_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13664 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_8  _0827_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _0828_
timestamp 1698431365
transform 1 0 2016 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0829_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8288 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _0830_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15232 0 1 37632
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_12  _0831_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20160 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _0832_
timestamp 1698431365
transform 1 0 30912 0 1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0833_
timestamp 1698431365
transform 1 0 30016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _0834_
timestamp 1698431365
transform 1 0 14112 0 1 34496
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_12  _0835_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12768 0 -1 45472
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_8  _0836_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 31024 0 1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_12  _0837_
timestamp 1698431365
transform 1 0 11088 0 -1 36064
box -86 -86 4342 870
use gf180mcu_fd_sc_mcu7t5v0__inv_4  _0838_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 26096 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0839_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34160 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _0840_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20160 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0841_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32256 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0842_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 30128 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0843_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 29568 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _0844_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0845_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31024 0 -1 29792
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0846_
timestamp 1698431365
transform -1 0 19264 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0847_
timestamp 1698431365
transform -1 0 20048 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _0848_
timestamp 1698431365
transform 1 0 41552 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0849_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0850_
timestamp 1698431365
transform -1 0 31248 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0851_
timestamp 1698431365
transform -1 0 24416 0 -1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0852_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22960 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0853_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 32480 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0854_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0855_
timestamp 1698431365
transform -1 0 33264 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0856_
timestamp 1698431365
transform 1 0 19824 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0857_
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _0858_
timestamp 1698431365
transform 1 0 25312 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0859_
timestamp 1698431365
transform -1 0 19712 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0860_
timestamp 1698431365
transform -1 0 22176 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0861_
timestamp 1698431365
transform 1 0 33264 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_8  _0862_
timestamp 1698431365
transform 1 0 19600 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0863_
timestamp 1698431365
transform 1 0 30688 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and4_4  _0864_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32256 0 1 36064
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0865_
timestamp 1698431365
transform -1 0 40544 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _0866_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18256 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0867_
timestamp 1698431365
transform -1 0 28784 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0868_
timestamp 1698431365
transform 1 0 30688 0 -1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0869_
timestamp 1698431365
transform 1 0 31248 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0870_
timestamp 1698431365
transform -1 0 45584 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _0871_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40768 0 1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0872_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34048 0 -1 21952
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0873_
timestamp 1698431365
transform -1 0 35840 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0874_
timestamp 1698431365
transform 1 0 30800 0 1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__and3_4  _0875_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29232 0 -1 40768
box -86 -86 2326 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0876_
timestamp 1698431365
transform 1 0 33376 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0877_
timestamp 1698431365
transform 1 0 29456 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _0878_
timestamp 1698431365
transform 1 0 31136 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0879_
timestamp 1698431365
transform 1 0 32032 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0880_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0881_
timestamp 1698431365
transform -1 0 35840 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _0882_
timestamp 1698431365
transform -1 0 36512 0 1 68992
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0883_
timestamp 1698431365
transform 1 0 34048 0 -1 65856
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0884_
timestamp 1698431365
transform 1 0 16800 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  _0885_
timestamp 1698431365
transform -1 0 32704 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0886_
timestamp 1698431365
transform 1 0 23968 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0887_
timestamp 1698431365
transform 1 0 18144 0 -1 58016
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0888_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18928 0 -1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0889_
timestamp 1698431365
transform -1 0 23072 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0890_
timestamp 1698431365
transform 1 0 24640 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0891_
timestamp 1698431365
transform -1 0 22960 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0892_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21504 0 -1 56448
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0893_
timestamp 1698431365
transform -1 0 20608 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0894_
timestamp 1698431365
transform 1 0 20608 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0895_
timestamp 1698431365
transform -1 0 28672 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0896_
timestamp 1698431365
transform 1 0 19488 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0897_
timestamp 1698431365
transform -1 0 22624 0 -1 68992
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0898_
timestamp 1698431365
transform 1 0 16352 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0899_
timestamp 1698431365
transform -1 0 24864 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0900_
timestamp 1698431365
transform -1 0 22960 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0901_
timestamp 1698431365
transform -1 0 20832 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0902_
timestamp 1698431365
transform 1 0 21168 0 1 56448
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0903_
timestamp 1698431365
transform 1 0 37856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0904_
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0905_
timestamp 1698431365
transform 1 0 22176 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0906_
timestamp 1698431365
transform -1 0 39760 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0907_
timestamp 1698431365
transform -1 0 40432 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0908_
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0909_
timestamp 1698431365
transform -1 0 40320 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0910_
timestamp 1698431365
transform 1 0 38640 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0911_
timestamp 1698431365
transform 1 0 38416 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0912_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0913_
timestamp 1698431365
transform 1 0 30352 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0914_
timestamp 1698431365
transform 1 0 38304 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0915_
timestamp 1698431365
transform -1 0 40432 0 1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0916_
timestamp 1698431365
transform -1 0 39200 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0917_
timestamp 1698431365
transform -1 0 35056 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0918_
timestamp 1698431365
transform 1 0 37408 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0919_
timestamp 1698431365
transform -1 0 38976 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0920_
timestamp 1698431365
transform 1 0 37968 0 1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0921_
timestamp 1698431365
transform 1 0 33712 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _0922_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20944 0 1 21952
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0923_
timestamp 1698431365
transform -1 0 10528 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0924_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12096 0 1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0925_
timestamp 1698431365
transform 1 0 30128 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0926_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29120 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0927_
timestamp 1698431365
transform 1 0 29232 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0928_
timestamp 1698431365
transform 1 0 30128 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0929_
timestamp 1698431365
transform -1 0 18928 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0930_
timestamp 1698431365
transform -1 0 18816 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0931_
timestamp 1698431365
transform 1 0 22176 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0932_
timestamp 1698431365
transform -1 0 18928 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0933_
timestamp 1698431365
transform -1 0 20944 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0934_
timestamp 1698431365
transform -1 0 41216 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0935_
timestamp 1698431365
transform -1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _0936_
timestamp 1698431365
transform -1 0 41216 0 1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0937_
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0938_
timestamp 1698431365
transform -1 0 36624 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0939_
timestamp 1698431365
transform -1 0 38640 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _0940_
timestamp 1698431365
transform -1 0 36624 0 1 70560
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0941_
timestamp 1698431365
transform 1 0 34944 0 -1 67424
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0942_
timestamp 1698431365
transform 1 0 18368 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0943_
timestamp 1698431365
transform 1 0 18704 0 1 58016
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0944_
timestamp 1698431365
transform 1 0 18928 0 1 56448
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0945_
timestamp 1698431365
transform 1 0 21616 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0946_
timestamp 1698431365
transform 1 0 21504 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0947_
timestamp 1698431365
transform 1 0 21392 0 -1 59584
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0948_
timestamp 1698431365
transform 1 0 21168 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0949_
timestamp 1698431365
transform 1 0 20720 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0950_
timestamp 1698431365
transform -1 0 23744 0 1 68992
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0951_
timestamp 1698431365
transform 1 0 18592 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0952_
timestamp 1698431365
transform 1 0 18704 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0953_
timestamp 1698431365
transform 1 0 19264 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0954_
timestamp 1698431365
transform 1 0 20608 0 -1 58016
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0955_
timestamp 1698431365
transform -1 0 40544 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0956_
timestamp 1698431365
transform -1 0 42672 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0957_
timestamp 1698431365
transform 1 0 42224 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0958_
timestamp 1698431365
transform 1 0 41664 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0959_
timestamp 1698431365
transform 1 0 42336 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0960_
timestamp 1698431365
transform -1 0 42560 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0961_
timestamp 1698431365
transform -1 0 41328 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0962_
timestamp 1698431365
transform -1 0 42896 0 1 53312
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0963_
timestamp 1698431365
transform 1 0 41440 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0964_
timestamp 1698431365
transform -1 0 42672 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0965_
timestamp 1698431365
transform 1 0 40768 0 1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0966_
timestamp 1698431365
transform 1 0 40880 0 -1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0967_
timestamp 1698431365
transform 1 0 35168 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _0968_
timestamp 1698431365
transform -1 0 22848 0 -1 21952
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0969_
timestamp 1698431365
transform -1 0 14448 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _0970_
timestamp 1698431365
transform -1 0 13776 0 -1 23520
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0971_
timestamp 1698431365
transform -1 0 31920 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0972_
timestamp 1698431365
transform 1 0 30352 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0973_
timestamp 1698431365
transform 1 0 31136 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0974_
timestamp 1698431365
transform -1 0 20944 0 1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0975_
timestamp 1698431365
transform -1 0 20272 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0976_
timestamp 1698431365
transform 1 0 22176 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0977_
timestamp 1698431365
transform -1 0 19936 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0978_
timestamp 1698431365
transform -1 0 22736 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0979_
timestamp 1698431365
transform -1 0 41216 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0980_
timestamp 1698431365
transform -1 0 43120 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _0981_
timestamp 1698431365
transform -1 0 40544 0 -1 14112
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0982_
timestamp 1698431365
transform 1 0 36064 0 -1 17248
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0983_
timestamp 1698431365
transform -1 0 37296 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0984_
timestamp 1698431365
transform -1 0 39088 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _0985_
timestamp 1698431365
transform -1 0 36736 0 -1 72128
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0986_
timestamp 1698431365
transform 1 0 34944 0 -1 64288
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0987_
timestamp 1698431365
transform 1 0 19488 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0988_
timestamp 1698431365
transform -1 0 20272 0 -1 54880
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0989_
timestamp 1698431365
transform 1 0 19264 0 1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0990_
timestamp 1698431365
transform 1 0 24304 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0991_
timestamp 1698431365
transform -1 0 24080 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0992_
timestamp 1698431365
transform -1 0 25424 0 1 58016
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0993_
timestamp 1698431365
transform -1 0 23744 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0994_
timestamp 1698431365
transform -1 0 24752 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0995_
timestamp 1698431365
transform 1 0 22288 0 -1 70560
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0996_
timestamp 1698431365
transform 1 0 18928 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0997_
timestamp 1698431365
transform 1 0 19152 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0998_
timestamp 1698431365
transform -1 0 20608 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0999_
timestamp 1698431365
transform 1 0 22624 0 1 54880
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1000_
timestamp 1698431365
transform 1 0 44016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1001_
timestamp 1698431365
transform 1 0 42672 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1002_
timestamp 1698431365
transform -1 0 46592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1003_
timestamp 1698431365
transform -1 0 44576 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1004_
timestamp 1698431365
transform 1 0 42672 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1005_
timestamp 1698431365
transform -1 0 44240 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1006_
timestamp 1698431365
transform -1 0 42560 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1007_
timestamp 1698431365
transform -1 0 43456 0 -1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1008_
timestamp 1698431365
transform -1 0 45136 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1009_
timestamp 1698431365
transform -1 0 43344 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1010_
timestamp 1698431365
transform 1 0 41440 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1011_
timestamp 1698431365
transform 1 0 41552 0 -1 43904
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1012_
timestamp 1698431365
transform 1 0 35392 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _1013_
timestamp 1698431365
transform -1 0 24304 0 -1 25088
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1014_
timestamp 1698431365
transform -1 0 12208 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1015_
timestamp 1698431365
transform -1 0 12992 0 -1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1016_
timestamp 1698431365
transform -1 0 31136 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1017_
timestamp 1698431365
transform -1 0 31920 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1018_
timestamp 1698431365
transform -1 0 30800 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1019_
timestamp 1698431365
transform -1 0 23184 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1020_
timestamp 1698431365
transform -1 0 23520 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1021_
timestamp 1698431365
transform 1 0 22848 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1022_
timestamp 1698431365
transform -1 0 22960 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1023_
timestamp 1698431365
transform 1 0 21280 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1024_
timestamp 1698431365
transform -1 0 39760 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1025_
timestamp 1698431365
transform -1 0 41776 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1026_
timestamp 1698431365
transform 1 0 34496 0 1 15680
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1027_
timestamp 1698431365
transform 1 0 34832 0 -1 15680
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1028_
timestamp 1698431365
transform -1 0 33712 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1029_
timestamp 1698431365
transform -1 0 33376 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1030_
timestamp 1698431365
transform 1 0 32256 0 1 70560
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1031_
timestamp 1698431365
transform 1 0 32144 0 1 62720
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1032_
timestamp 1698431365
transform 1 0 23856 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1033_
timestamp 1698431365
transform 1 0 23408 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1034_
timestamp 1698431365
transform -1 0 24192 0 1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1035_
timestamp 1698431365
transform 1 0 25200 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1036_
timestamp 1698431365
transform 1 0 26096 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1037_
timestamp 1698431365
transform 1 0 25088 0 -1 58016
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1038_
timestamp 1698431365
transform 1 0 23968 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1039_
timestamp 1698431365
transform 1 0 25424 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1040_
timestamp 1698431365
transform 1 0 25088 0 -1 70560
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1041_
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1042_
timestamp 1698431365
transform 1 0 19152 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1043_
timestamp 1698431365
transform 1 0 20944 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1044_
timestamp 1698431365
transform 1 0 24192 0 1 53312
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1045_
timestamp 1698431365
transform -1 0 46704 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1046_
timestamp 1698431365
transform 1 0 41440 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1047_
timestamp 1698431365
transform -1 0 46592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1048_
timestamp 1698431365
transform 1 0 41440 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1049_
timestamp 1698431365
transform 1 0 44352 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1050_
timestamp 1698431365
transform -1 0 45360 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1051_
timestamp 1698431365
transform -1 0 43008 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1052_
timestamp 1698431365
transform -1 0 43232 0 1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1053_
timestamp 1698431365
transform -1 0 46144 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1054_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41776 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1055_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42784 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1056_
timestamp 1698431365
transform 1 0 41328 0 -1 37632
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1057_
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _1058_
timestamp 1698431365
transform -1 0 26544 0 1 21952
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1059_
timestamp 1698431365
transform -1 0 12544 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1060_
timestamp 1698431365
transform -1 0 13104 0 1 21952
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1061_
timestamp 1698431365
transform -1 0 10864 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1062_
timestamp 1698431365
transform -1 0 30912 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1063_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27552 0 -1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1064_
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1065_
timestamp 1698431365
transform -1 0 28112 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1066_
timestamp 1698431365
transform -1 0 26656 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1067_
timestamp 1698431365
transform 1 0 20720 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1068_
timestamp 1698431365
transform -1 0 28000 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1069_
timestamp 1698431365
transform 1 0 26880 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1070_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28000 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1071_
timestamp 1698431365
transform -1 0 26880 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1072_
timestamp 1698431365
transform -1 0 27328 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1073_
timestamp 1698431365
transform 1 0 25760 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1074_
timestamp 1698431365
transform 1 0 26208 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1075_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30688 0 -1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1076_
timestamp 1698431365
transform -1 0 30800 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1077_
timestamp 1698431365
transform -1 0 31696 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1078_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30800 0 -1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1079_
timestamp 1698431365
transform 1 0 26544 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1080_
timestamp 1698431365
transform -1 0 29232 0 -1 40768
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1081_
timestamp 1698431365
transform 1 0 29456 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1082_
timestamp 1698431365
transform 1 0 31696 0 -1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1083_
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1084_
timestamp 1698431365
transform -1 0 33600 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1085_
timestamp 1698431365
transform 1 0 31696 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1086_
timestamp 1698431365
transform -1 0 37296 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1087_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 34384 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1088_
timestamp 1698431365
transform -1 0 27328 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1089_
timestamp 1698431365
transform -1 0 45920 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1090_
timestamp 1698431365
transform 1 0 31360 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1091_
timestamp 1698431365
transform -1 0 36288 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1092_
timestamp 1698431365
transform -1 0 37856 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1093_
timestamp 1698431365
transform 1 0 35168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1094_
timestamp 1698431365
transform -1 0 47488 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1095_
timestamp 1698431365
transform -1 0 42672 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1096_
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1097_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33152 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1098_
timestamp 1698431365
transform -1 0 26096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1099_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25536 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1100_
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1101_
timestamp 1698431365
transform -1 0 37968 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1102_
timestamp 1698431365
transform 1 0 31584 0 1 37632
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1103_
timestamp 1698431365
transform 1 0 34160 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1104_
timestamp 1698431365
transform -1 0 27776 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1105_
timestamp 1698431365
transform 1 0 27552 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1106_
timestamp 1698431365
transform -1 0 27440 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1107_
timestamp 1698431365
transform -1 0 28784 0 1 26656
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1108_
timestamp 1698431365
transform -1 0 33824 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1109_
timestamp 1698431365
transform -1 0 33152 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1110_
timestamp 1698431365
transform 1 0 27776 0 -1 28224
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1111_
timestamp 1698431365
transform -1 0 31472 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1112_
timestamp 1698431365
transform -1 0 12544 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1113_
timestamp 1698431365
transform -1 0 13552 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1114_
timestamp 1698431365
transform 1 0 9632 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1115_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14000 0 -1 28224
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1116_
timestamp 1698431365
transform -1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1117_
timestamp 1698431365
transform 1 0 28224 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1118_
timestamp 1698431365
transform -1 0 30352 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1119_
timestamp 1698431365
transform -1 0 31360 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1120_
timestamp 1698431365
transform 1 0 30688 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1121_
timestamp 1698431365
transform 1 0 28896 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1122_
timestamp 1698431365
transform -1 0 30800 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1123_
timestamp 1698431365
transform 1 0 30464 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1124_
timestamp 1698431365
transform -1 0 30352 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1125_
timestamp 1698431365
transform 1 0 27216 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1126_
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1127_
timestamp 1698431365
transform 1 0 25984 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1128_
timestamp 1698431365
transform 1 0 25536 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1129_
timestamp 1698431365
transform 1 0 25536 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1130_
timestamp 1698431365
transform 1 0 28672 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1131_
timestamp 1698431365
transform -1 0 30128 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1132_
timestamp 1698431365
transform 1 0 26544 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1133_
timestamp 1698431365
transform 1 0 28336 0 -1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1134_
timestamp 1698431365
transform -1 0 31808 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1135_
timestamp 1698431365
transform -1 0 36064 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1136_
timestamp 1698431365
transform 1 0 34496 0 1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1137_
timestamp 1698431365
transform 1 0 34832 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1138_
timestamp 1698431365
transform -1 0 35952 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1139_
timestamp 1698431365
transform 1 0 35056 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1140_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27776 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1141_
timestamp 1698431365
transform -1 0 31360 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1142_
timestamp 1698431365
transform 1 0 27104 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1143_
timestamp 1698431365
transform 1 0 26768 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1144_
timestamp 1698431365
transform 1 0 25424 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1145_
timestamp 1698431365
transform 1 0 26880 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1146_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29120 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _1147_
timestamp 1698431365
transform -1 0 30464 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1148_
timestamp 1698431365
transform 1 0 11424 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1149_
timestamp 1698431365
transform -1 0 16016 0 -1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__inv_4  _1150_
timestamp 1698431365
transform 1 0 3808 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1151_
timestamp 1698431365
transform -1 0 4592 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1152_
timestamp 1698431365
transform -1 0 4256 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1153_
timestamp 1698431365
transform -1 0 4704 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1154_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3920 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1155_
timestamp 1698431365
transform -1 0 3584 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _1156_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2912 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1157_
timestamp 1698431365
transform -1 0 6384 0 -1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1158_
timestamp 1698431365
transform -1 0 7056 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1159_
timestamp 1698431365
transform -1 0 7168 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1160_
timestamp 1698431365
transform -1 0 8176 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1161_
timestamp 1698431365
transform -1 0 7728 0 -1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1162_
timestamp 1698431365
transform -1 0 9072 0 -1 50176
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1163_
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1164_
timestamp 1698431365
transform 1 0 3360 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1165_
timestamp 1698431365
transform -1 0 3920 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1166_
timestamp 1698431365
transform 1 0 2016 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_3  _1167_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2464 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1168_
timestamp 1698431365
transform 1 0 1792 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1169_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3360 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1170_
timestamp 1698431365
transform -1 0 3136 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _1171_
timestamp 1698431365
transform -1 0 2800 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1172_
timestamp 1698431365
transform 1 0 2464 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1173_
timestamp 1698431365
transform 1 0 2352 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1174_
timestamp 1698431365
transform 1 0 4816 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1175_
timestamp 1698431365
transform 1 0 2352 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1176_
timestamp 1698431365
transform 1 0 2016 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1177_
timestamp 1698431365
transform -1 0 6720 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1178_
timestamp 1698431365
transform 1 0 2352 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1179_
timestamp 1698431365
transform 1 0 3360 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1180_
timestamp 1698431365
transform 1 0 4592 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1181_
timestamp 1698431365
transform -1 0 7728 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1182_
timestamp 1698431365
transform -1 0 5264 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1183_
timestamp 1698431365
transform -1 0 5040 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1184_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4928 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1185_
timestamp 1698431365
transform -1 0 5152 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1186_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2352 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1187_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3584 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1188_
timestamp 1698431365
transform -1 0 3136 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1189_
timestamp 1698431365
transform -1 0 4816 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1190_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4368 0 -1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1191_
timestamp 1698431365
transform 1 0 4368 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1192_
timestamp 1698431365
transform -1 0 5264 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1193_
timestamp 1698431365
transform 1 0 2352 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1194_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2464 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _1195_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 2800 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1196_
timestamp 1698431365
transform 1 0 2912 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1197_
timestamp 1698431365
transform -1 0 8288 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1198_
timestamp 1698431365
transform -1 0 9072 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1199_
timestamp 1698431365
transform -1 0 7952 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1200_
timestamp 1698431365
transform 1 0 8624 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1201_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1202_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4592 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1203_
timestamp 1698431365
transform 1 0 3808 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1204_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5376 0 -1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1205_
timestamp 1698431365
transform -1 0 4592 0 1 37632
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1206_
timestamp 1698431365
transform -1 0 3360 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1207_
timestamp 1698431365
transform -1 0 9408 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1208_
timestamp 1698431365
transform -1 0 6944 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1209_
timestamp 1698431365
transform -1 0 6048 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1210_
timestamp 1698431365
transform 1 0 7504 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1211_
timestamp 1698431365
transform 1 0 7168 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1212_
timestamp 1698431365
transform -1 0 5264 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1213_
timestamp 1698431365
transform 1 0 5376 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1214_
timestamp 1698431365
transform -1 0 6384 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1215_
timestamp 1698431365
transform 1 0 5600 0 -1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1216_
timestamp 1698431365
transform -1 0 5264 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1217_
timestamp 1698431365
transform 1 0 4256 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1218_
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1219_
timestamp 1698431365
transform -1 0 6048 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1220__1
timestamp 1698431365
transform -1 0 8736 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1221_
timestamp 1698431365
transform -1 0 3696 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1222_
timestamp 1698431365
transform -1 0 11088 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1223_
timestamp 1698431365
transform 1 0 7728 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1224_
timestamp 1698431365
transform -1 0 9184 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1225_
timestamp 1698431365
transform 1 0 8064 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1226_
timestamp 1698431365
transform 1 0 7728 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1227_
timestamp 1698431365
transform -1 0 8512 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1228_
timestamp 1698431365
transform 1 0 6832 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1229_
timestamp 1698431365
transform -1 0 8512 0 -1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1230_
timestamp 1698431365
transform -1 0 8848 0 -1 40768
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1231_
timestamp 1698431365
transform -1 0 6384 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1232_
timestamp 1698431365
transform -1 0 7392 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1233_
timestamp 1698431365
transform -1 0 9856 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1234_
timestamp 1698431365
transform -1 0 11088 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1235_
timestamp 1698431365
transform 1 0 5264 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1236_
timestamp 1698431365
transform 1 0 5824 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1237_
timestamp 1698431365
transform 1 0 6048 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1238_
timestamp 1698431365
transform -1 0 6944 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1239_
timestamp 1698431365
transform 1 0 5936 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1240_
timestamp 1698431365
transform -1 0 7728 0 1 32928
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1241_
timestamp 1698431365
transform 1 0 5600 0 1 39200
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1242_
timestamp 1698431365
transform 1 0 7392 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1243_
timestamp 1698431365
transform 1 0 3472 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1244_
timestamp 1698431365
transform -1 0 9072 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1245_
timestamp 1698431365
transform -1 0 11312 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1246_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10192 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1247_
timestamp 1698431365
transform -1 0 9184 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1248_
timestamp 1698431365
transform -1 0 7280 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1249_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4592 0 1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1250_
timestamp 1698431365
transform 1 0 7280 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1251_
timestamp 1698431365
transform -1 0 6832 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1252_
timestamp 1698431365
transform 1 0 6832 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1253_
timestamp 1698431365
transform -1 0 3136 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1254_
timestamp 1698431365
transform 1 0 4256 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1255_
timestamp 1698431365
transform 1 0 3360 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1256_
timestamp 1698431365
transform -1 0 10976 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1257_
timestamp 1698431365
transform 1 0 5712 0 -1 28224
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1258_
timestamp 1698431365
transform -1 0 5936 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1259_
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1260_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6048 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1261_
timestamp 1698431365
transform 1 0 5824 0 1 37632
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1262_
timestamp 1698431365
transform 1 0 3920 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1263_
timestamp 1698431365
transform -1 0 3360 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1264_
timestamp 1698431365
transform -1 0 2352 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1265_
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1266_
timestamp 1698431365
transform -1 0 4480 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1267_
timestamp 1698431365
transform -1 0 5152 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1268_
timestamp 1698431365
transform -1 0 2688 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1269_
timestamp 1698431365
transform -1 0 2688 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1270_
timestamp 1698431365
transform 1 0 2800 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1271_
timestamp 1698431365
transform 1 0 1904 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1272_
timestamp 1698431365
transform 1 0 2016 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1273_
timestamp 1698431365
transform 1 0 14112 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1274_
timestamp 1698431365
transform 1 0 10640 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1275_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11088 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_4  _1276_
timestamp 1698431365
transform 1 0 15680 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1277_
timestamp 1698431365
transform 1 0 14000 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1278_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1279_
timestamp 1698431365
transform -1 0 14896 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1280_
timestamp 1698431365
transform 1 0 14336 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1281_
timestamp 1698431365
transform -1 0 16576 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1282_
timestamp 1698431365
transform -1 0 15904 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1283_
timestamp 1698431365
transform -1 0 15680 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1284_
timestamp 1698431365
transform 1 0 15904 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1285_
timestamp 1698431365
transform -1 0 17920 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1286_
timestamp 1698431365
transform -1 0 14224 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1287_
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1288_
timestamp 1698431365
transform 1 0 13664 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1289_
timestamp 1698431365
transform -1 0 15568 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1290_
timestamp 1698431365
transform -1 0 19712 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1291_
timestamp 1698431365
transform -1 0 19376 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1292_
timestamp 1698431365
transform 1 0 17584 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1293_
timestamp 1698431365
transform -1 0 21840 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1294_
timestamp 1698431365
transform 1 0 13888 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1295_
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1296_
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1297_
timestamp 1698431365
transform 1 0 30016 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1298_
timestamp 1698431365
transform 1 0 33488 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1299_
timestamp 1698431365
transform 1 0 34720 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1300_
timestamp 1698431365
transform -1 0 38976 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1301_
timestamp 1698431365
transform 1 0 39872 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1302_
timestamp 1698431365
transform 1 0 40768 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1303_
timestamp 1698431365
transform 1 0 41664 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1304_
timestamp 1698431365
transform 1 0 27888 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1305_
timestamp 1698431365
transform 1 0 28784 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1306_
timestamp 1698431365
transform 1 0 31696 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1307_
timestamp 1698431365
transform 1 0 32928 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1308_
timestamp 1698431365
transform 1 0 34272 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1309_
timestamp 1698431365
transform 1 0 37072 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1310_
timestamp 1698431365
transform 1 0 32928 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1311_
timestamp 1698431365
transform -1 0 30576 0 1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1312_
timestamp 1698431365
transform -1 0 28000 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1313_
timestamp 1698431365
transform -1 0 27104 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1314_
timestamp 1698431365
transform -1 0 28448 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1315_
timestamp 1698431365
transform -1 0 27104 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1316_
timestamp 1698431365
transform -1 0 14672 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1317_
timestamp 1698431365
transform 1 0 14224 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1318_
timestamp 1698431365
transform -1 0 15120 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1319_
timestamp 1698431365
transform -1 0 14672 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1320_
timestamp 1698431365
transform -1 0 16800 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1321_
timestamp 1698431365
transform -1 0 15680 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1322_
timestamp 1698431365
transform 1 0 17360 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1323_
timestamp 1698431365
transform -1 0 19488 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1324_
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1325_
timestamp 1698431365
transform -1 0 20384 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1326_
timestamp 1698431365
transform -1 0 19600 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1327_
timestamp 1698431365
transform -1 0 19264 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1328_
timestamp 1698431365
transform -1 0 17584 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1329_
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1330_
timestamp 1698431365
transform -1 0 17024 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1331_
timestamp 1698431365
transform -1 0 15792 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1332_
timestamp 1698431365
transform 1 0 17584 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1333_
timestamp 1698431365
transform -1 0 18480 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1334_
timestamp 1698431365
transform -1 0 20832 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1335_
timestamp 1698431365
transform 1 0 19824 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1336_
timestamp 1698431365
transform -1 0 22512 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1337_
timestamp 1698431365
transform 1 0 21840 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1338_
timestamp 1698431365
transform -1 0 24304 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1339_
timestamp 1698431365
transform -1 0 23856 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1340_
timestamp 1698431365
transform -1 0 19824 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1341_
timestamp 1698431365
transform -1 0 19712 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1342_
timestamp 1698431365
transform 1 0 19152 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1343_
timestamp 1698431365
transform -1 0 21840 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1344_
timestamp 1698431365
transform 1 0 22624 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1345_
timestamp 1698431365
transform 1 0 25088 0 -1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1346_
timestamp 1698431365
transform -1 0 28560 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1347_
timestamp 1698431365
transform 1 0 27664 0 1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1348_
timestamp 1698431365
transform 1 0 29792 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1349_
timestamp 1698431365
transform 1 0 30464 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1350_
timestamp 1698431365
transform 1 0 34384 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1351_
timestamp 1698431365
transform -1 0 36176 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1352_
timestamp 1698431365
transform 1 0 33264 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1353_
timestamp 1698431365
transform 1 0 30128 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1354_
timestamp 1698431365
transform -1 0 29456 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1355_
timestamp 1698431365
transform -1 0 28784 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1356_
timestamp 1698431365
transform 1 0 29568 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1357_
timestamp 1698431365
transform -1 0 31024 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1358_
timestamp 1698431365
transform 1 0 32928 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1359_
timestamp 1698431365
transform -1 0 33600 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1360_
timestamp 1698431365
transform -1 0 33936 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1361_
timestamp 1698431365
transform 1 0 33376 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1362_
timestamp 1698431365
transform -1 0 31696 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1363_
timestamp 1698431365
transform -1 0 31024 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1364_
timestamp 1698431365
transform -1 0 30800 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1365_
timestamp 1698431365
transform -1 0 30240 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1366_
timestamp 1698431365
transform -1 0 30800 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1367_
timestamp 1698431365
transform 1 0 29680 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1368_
timestamp 1698431365
transform -1 0 29904 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1369_
timestamp 1698431365
transform -1 0 29008 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1370_
timestamp 1698431365
transform -1 0 24640 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1371_
timestamp 1698431365
transform 1 0 23856 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1372_
timestamp 1698431365
transform -1 0 22848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1373_
timestamp 1698431365
transform -1 0 22512 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1374_
timestamp 1698431365
transform 1 0 22960 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1375_
timestamp 1698431365
transform -1 0 24640 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1376_
timestamp 1698431365
transform 1 0 24416 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1377_
timestamp 1698431365
transform 1 0 24528 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1378_
timestamp 1698431365
transform -1 0 25760 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1379_
timestamp 1698431365
transform -1 0 26656 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1380_
timestamp 1698431365
transform 1 0 25536 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1381_
timestamp 1698431365
transform -1 0 22064 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1382_
timestamp 1698431365
transform -1 0 20720 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1383_
timestamp 1698431365
transform -1 0 22064 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1384_
timestamp 1698431365
transform -1 0 21392 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1385_
timestamp 1698431365
transform -1 0 22288 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1386_
timestamp 1698431365
transform 1 0 21168 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1387_
timestamp 1698431365
transform -1 0 23632 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1388_
timestamp 1698431365
transform 1 0 23072 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1389_
timestamp 1698431365
transform -1 0 25648 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1390_
timestamp 1698431365
transform -1 0 19376 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1391_
timestamp 1698431365
transform -1 0 17920 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1392_
timestamp 1698431365
transform -1 0 18144 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1393_
timestamp 1698431365
transform -1 0 15568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1394_
timestamp 1698431365
transform -1 0 17248 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1395_
timestamp 1698431365
transform -1 0 16240 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1396_
timestamp 1698431365
transform 1 0 17584 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1397_
timestamp 1698431365
transform 1 0 18032 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1398_
timestamp 1698431365
transform 1 0 20272 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1399_
timestamp 1698431365
transform -1 0 21840 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1400_
timestamp 1698431365
transform 1 0 22400 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1401_
timestamp 1698431365
transform 1 0 23296 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1402_
timestamp 1698431365
transform -1 0 18704 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1403_
timestamp 1698431365
transform -1 0 17472 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1404_
timestamp 1698431365
transform -1 0 18480 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1405_
timestamp 1698431365
transform -1 0 15008 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1406_
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1407_
timestamp 1698431365
transform -1 0 16688 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1408_
timestamp 1698431365
transform -1 0 16464 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1409_
timestamp 1698431365
transform -1 0 18480 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1410_
timestamp 1698431365
transform 1 0 17920 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1411_
timestamp 1698431365
transform -1 0 22064 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1412_
timestamp 1698431365
transform 1 0 21280 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1413_
timestamp 1698431365
transform -1 0 24416 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1414_
timestamp 1698431365
transform 1 0 22848 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1415_
timestamp 1698431365
transform -1 0 23408 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1416_
timestamp 1698431365
transform -1 0 22624 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1417_
timestamp 1698431365
transform 1 0 19600 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1418_
timestamp 1698431365
transform 1 0 21504 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1419_
timestamp 1698431365
transform 1 0 23520 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1420_
timestamp 1698431365
transform 1 0 24192 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1421_
timestamp 1698431365
transform -1 0 27216 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1422_
timestamp 1698431365
transform -1 0 26992 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1423_
timestamp 1698431365
transform -1 0 28224 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1424_
timestamp 1698431365
transform -1 0 18480 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1425_
timestamp 1698431365
transform -1 0 19264 0 1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1426_
timestamp 1698431365
transform -1 0 21840 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1427_
timestamp 1698431365
transform -1 0 24304 0 -1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1428_
timestamp 1698431365
transform -1 0 26544 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1429_
timestamp 1698431365
transform -1 0 28224 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1430_
timestamp 1698431365
transform -1 0 27888 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1431_
timestamp 1698431365
transform -1 0 29904 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1432_
timestamp 1698431365
transform -1 0 18592 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1433_
timestamp 1698431365
transform -1 0 18144 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1434_
timestamp 1698431365
transform -1 0 17920 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1435_
timestamp 1698431365
transform -1 0 18256 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1436_
timestamp 1698431365
transform -1 0 17920 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1437_
timestamp 1698431365
transform 1 0 19264 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1438_
timestamp 1698431365
transform 1 0 20160 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1439_
timestamp 1698431365
transform -1 0 23856 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1440_
timestamp 1698431365
transform 1 0 23184 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1441_
timestamp 1698431365
transform -1 0 25984 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1442_
timestamp 1698431365
transform 1 0 25088 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1443_
timestamp 1698431365
transform 1 0 34720 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1444_
timestamp 1698431365
transform 1 0 29008 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1445_
timestamp 1698431365
transform 1 0 35392 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1446_
timestamp 1698431365
transform 1 0 39088 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1447_
timestamp 1698431365
transform 1 0 39872 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1448_
timestamp 1698431365
transform 1 0 43232 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1449_
timestamp 1698431365
transform -1 0 44352 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1450_
timestamp 1698431365
transform -1 0 45584 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1451_
timestamp 1698431365
transform 1 0 44688 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1452_
timestamp 1698431365
transform -1 0 43008 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1453_
timestamp 1698431365
transform 1 0 41776 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1454_
timestamp 1698431365
transform 1 0 42112 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1455_
timestamp 1698431365
transform -1 0 43008 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1456_
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1457_
timestamp 1698431365
transform -1 0 44688 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1458_
timestamp 1698431365
transform 1 0 41664 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1459_
timestamp 1698431365
transform 1 0 40880 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1460_
timestamp 1698431365
transform 1 0 39872 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1461_
timestamp 1698431365
transform -1 0 34272 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1462_
timestamp 1698431365
transform -1 0 25312 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1463_
timestamp 1698431365
transform -1 0 24304 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1464_
timestamp 1698431365
transform -1 0 16912 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1465_
timestamp 1698431365
transform -1 0 15904 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1466_
timestamp 1698431365
transform -1 0 16912 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1467_
timestamp 1698431365
transform -1 0 18032 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1468_
timestamp 1698431365
transform -1 0 19376 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1469_
timestamp 1698431365
transform -1 0 23632 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1470_
timestamp 1698431365
transform -1 0 25984 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1471_
timestamp 1698431365
transform 1 0 24416 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1472_
timestamp 1698431365
transform 1 0 31808 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1473_
timestamp 1698431365
transform 1 0 35840 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1474_
timestamp 1698431365
transform 1 0 38976 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1475_
timestamp 1698431365
transform 1 0 39424 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1476_
timestamp 1698431365
transform 1 0 42560 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1477_
timestamp 1698431365
transform 1 0 43680 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1478_
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1479_
timestamp 1698431365
transform 1 0 45584 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1480_
timestamp 1698431365
transform -1 0 41552 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1481_
timestamp 1698431365
transform -1 0 41104 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1482_
timestamp 1698431365
transform -1 0 37968 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1483_
timestamp 1698431365
transform 1 0 37184 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1484_
timestamp 1698431365
transform 1 0 31808 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1485_
timestamp 1698431365
transform -1 0 33376 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1486_
timestamp 1698431365
transform -1 0 34496 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1487_
timestamp 1698431365
transform 1 0 33824 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1488_
timestamp 1698431365
transform -1 0 37744 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1489_
timestamp 1698431365
transform 1 0 35952 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1490_
timestamp 1698431365
transform 1 0 37072 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1491_
timestamp 1698431365
transform 1 0 37968 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1492_
timestamp 1698431365
transform -1 0 36064 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1493_
timestamp 1698431365
transform 1 0 35280 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1494_
timestamp 1698431365
transform -1 0 34160 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1495_
timestamp 1698431365
transform 1 0 32032 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1496_
timestamp 1698431365
transform -1 0 34496 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1497_
timestamp 1698431365
transform -1 0 18592 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1498_
timestamp 1698431365
transform -1 0 14896 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1499_
timestamp 1698431365
transform -1 0 15008 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1500_
timestamp 1698431365
transform 1 0 15344 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1501_
timestamp 1698431365
transform -1 0 16912 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1502_
timestamp 1698431365
transform 1 0 18816 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1503_
timestamp 1698431365
transform 1 0 19712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1504_
timestamp 1698431365
transform 1 0 23072 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1505_
timestamp 1698431365
transform -1 0 24080 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1506_
timestamp 1698431365
transform -1 0 26208 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1507_
timestamp 1698431365
transform 1 0 24192 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1508_
timestamp 1698431365
transform -1 0 27664 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1509_
timestamp 1698431365
transform -1 0 27664 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1510_
timestamp 1698431365
transform -1 0 29232 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1511_
timestamp 1698431365
transform -1 0 28672 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1512_
timestamp 1698431365
transform 1 0 29792 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1513_
timestamp 1698431365
transform 1 0 30240 0 -1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1514_
timestamp 1698431365
transform 1 0 30576 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1515_
timestamp 1698431365
transform -1 0 31024 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1516_
timestamp 1698431365
transform 1 0 31696 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1517_
timestamp 1698431365
transform -1 0 32816 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _1518_
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1519_
timestamp 1698431365
transform 1 0 31024 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1520_
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1521_
timestamp 1698431365
transform 1 0 34272 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1522_
timestamp 1698431365
transform 1 0 35952 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1523_
timestamp 1698431365
transform 1 0 39984 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1524_
timestamp 1698431365
transform -1 0 45360 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1525_
timestamp 1698431365
transform 1 0 39536 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1526_
timestamp 1698431365
transform 1 0 35728 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1527_
timestamp 1698431365
transform -1 0 37520 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1528_
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1529_
timestamp 1698431365
transform 1 0 37408 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1530_
timestamp 1698431365
transform 1 0 39312 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1531_
timestamp 1698431365
transform 1 0 42896 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1532_
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1533_
timestamp 1698431365
transform 1 0 45024 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1534_
timestamp 1698431365
transform 1 0 40096 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1535_
timestamp 1698431365
transform -1 0 28448 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1536_
timestamp 1698431365
transform -1 0 28224 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1537_
timestamp 1698431365
transform 1 0 36512 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1538_
timestamp 1698431365
transform -1 0 29904 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1539_
timestamp 1698431365
transform -1 0 28784 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1540_
timestamp 1698431365
transform -1 0 30576 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1541_
timestamp 1698431365
transform 1 0 29120 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1542_
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1543_
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1544_
timestamp 1698431365
transform -1 0 31808 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1545_
timestamp 1698431365
transform 1 0 30912 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1546_
timestamp 1698431365
transform 1 0 30128 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1547_
timestamp 1698431365
transform 1 0 31024 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1548_
timestamp 1698431365
transform -1 0 31024 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1549_
timestamp 1698431365
transform -1 0 28448 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1550_
timestamp 1698431365
transform -1 0 21952 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1551_
timestamp 1698431365
transform -1 0 22624 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1552_
timestamp 1698431365
transform 1 0 23184 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1553_
timestamp 1698431365
transform 1 0 25312 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1554_
timestamp 1698431365
transform 1 0 27440 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1555_
timestamp 1698431365
transform 1 0 30240 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1556_
timestamp 1698431365
transform 1 0 30912 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1557_
timestamp 1698431365
transform -1 0 35280 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1558_
timestamp 1698431365
transform -1 0 35280 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1559_
timestamp 1698431365
transform 1 0 36736 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1560_
timestamp 1698431365
transform 1 0 37072 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1561_
timestamp 1698431365
transform 1 0 37520 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1562_
timestamp 1698431365
transform 1 0 38416 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1563_
timestamp 1698431365
transform -1 0 36624 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1564_
timestamp 1698431365
transform -1 0 36288 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1565_
timestamp 1698431365
transform -1 0 35056 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1566_
timestamp 1698431365
transform 1 0 35280 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1567_
timestamp 1698431365
transform 1 0 35840 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1568_
timestamp 1698431365
transform 1 0 38528 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1569_
timestamp 1698431365
transform 1 0 41440 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1570_
timestamp 1698431365
transform 1 0 43456 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1571_
timestamp 1698431365
transform 1 0 37184 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1572_
timestamp 1698431365
transform -1 0 34832 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1573_
timestamp 1698431365
transform -1 0 34384 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1574_
timestamp 1698431365
transform 1 0 35728 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1575_
timestamp 1698431365
transform 1 0 36288 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1576_
timestamp 1698431365
transform 1 0 38416 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1577_
timestamp 1698431365
transform -1 0 42224 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1578_
timestamp 1698431365
transform 1 0 43568 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1579_
timestamp 1698431365
transform 1 0 43680 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1580_
timestamp 1698431365
transform -1 0 34384 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1581_
timestamp 1698431365
transform 1 0 34944 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1582_
timestamp 1698431365
transform 1 0 35392 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1583_
timestamp 1698431365
transform -1 0 37744 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1584_
timestamp 1698431365
transform 1 0 35952 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1585_
timestamp 1698431365
transform -1 0 39424 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1586_
timestamp 1698431365
transform 1 0 38304 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1587_
timestamp 1698431365
transform -1 0 37744 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1588_
timestamp 1698431365
transform 1 0 36960 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1589_
timestamp 1698431365
transform -1 0 33376 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1590_
timestamp 1698431365
transform -1 0 32704 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1591_
timestamp 1698431365
transform -1 0 34720 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1592_
timestamp 1698431365
transform -1 0 33936 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1593_
timestamp 1698431365
transform 1 0 38976 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1594_
timestamp 1698431365
transform 1 0 36176 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1595_
timestamp 1698431365
transform 1 0 39088 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1596_
timestamp 1698431365
transform 1 0 39648 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1597_
timestamp 1698431365
transform 1 0 38752 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1598_
timestamp 1698431365
transform 1 0 34832 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1599_
timestamp 1698431365
transform 1 0 34608 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1600_
timestamp 1698431365
transform 1 0 3136 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1601_
timestamp 1698431365
transform -1 0 4032 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1602_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7728 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1603_
timestamp 1698431365
transform 1 0 12096 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1604_
timestamp 1698431365
transform 1 0 11200 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1605_
timestamp 1698431365
transform 1 0 9520 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1606_
timestamp 1698431365
transform -1 0 9184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1607_
timestamp 1698431365
transform -1 0 10864 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1608_
timestamp 1698431365
transform -1 0 11760 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1609_
timestamp 1698431365
transform 1 0 11648 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1610_
timestamp 1698431365
transform 1 0 10752 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1611_
timestamp 1698431365
transform -1 0 11760 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1612_
timestamp 1698431365
transform -1 0 12656 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1613_
timestamp 1698431365
transform 1 0 10304 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1614_
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1615_
timestamp 1698431365
transform 1 0 1792 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1616_
timestamp 1698431365
transform 1 0 2352 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1617_
timestamp 1698431365
transform -1 0 12880 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1618_
timestamp 1698431365
transform -1 0 2912 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1619_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5600 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1620_
timestamp 1698431365
transform 1 0 8400 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1621_
timestamp 1698431365
transform -1 0 6608 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1622_
timestamp 1698431365
transform 1 0 8176 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1623_
timestamp 1698431365
transform -1 0 7840 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1624_
timestamp 1698431365
transform 1 0 8736 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1625_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1626_
timestamp 1698431365
transform 1 0 11088 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1627_
timestamp 1698431365
transform 1 0 9520 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1628_
timestamp 1698431365
transform 1 0 10080 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1629_
timestamp 1698431365
transform 1 0 11424 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1630_
timestamp 1698431365
transform -1 0 10752 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1631_
timestamp 1698431365
transform -1 0 9968 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1632_
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1633_
timestamp 1698431365
transform -1 0 2800 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1634_
timestamp 1698431365
transform 1 0 2688 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1635_
timestamp 1698431365
transform 1 0 3248 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1636_
timestamp 1698431365
transform -1 0 2800 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1637_
timestamp 1698431365
transform 1 0 2128 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1638_
timestamp 1698431365
transform -1 0 2464 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1639_
timestamp 1698431365
transform 1 0 3136 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1640_
timestamp 1698431365
transform -1 0 3248 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1641_
timestamp 1698431365
transform 1 0 2240 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1642_
timestamp 1698431365
transform 1 0 2464 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1643_
timestamp 1698431365
transform -1 0 3472 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1644_
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1645_
timestamp 1698431365
transform 1 0 3024 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1646_
timestamp 1698431365
transform -1 0 2912 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1647_
timestamp 1698431365
transform 1 0 3696 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1648_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12768 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1649_
timestamp 1698431365
transform 1 0 12768 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1650_
timestamp 1698431365
transform 1 0 12992 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1651_
timestamp 1698431365
transform 1 0 14224 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1652_
timestamp 1698431365
transform -1 0 17024 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1653_
timestamp 1698431365
transform -1 0 15120 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1654_
timestamp 1698431365
transform 1 0 13552 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1655_
timestamp 1698431365
transform 1 0 15456 0 1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1656_
timestamp 1698431365
transform 1 0 17248 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1657_
timestamp 1698431365
transform 1 0 20384 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1658_
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1659_
timestamp 1698431365
transform 1 0 30016 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1660_
timestamp 1698431365
transform 1 0 35168 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1661_
timestamp 1698431365
transform 1 0 37632 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1662_
timestamp 1698431365
transform 1 0 39760 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1663_
timestamp 1698431365
transform 1 0 40768 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1664_
timestamp 1698431365
transform -1 0 44464 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1665_
timestamp 1698431365
transform 1 0 28336 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1666_
timestamp 1698431365
transform 1 0 32928 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1667_
timestamp 1698431365
transform 1 0 34944 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1668_
timestamp 1698431365
transform 1 0 36848 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1669_
timestamp 1698431365
transform 1 0 30576 0 1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1670_
timestamp 1698431365
transform 1 0 25760 0 -1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1671_
timestamp 1698431365
transform 1 0 25536 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1672_
timestamp 1698431365
transform -1 0 18928 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1673_
timestamp 1698431365
transform -1 0 15904 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1674_
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1675_
timestamp 1698431365
transform 1 0 13776 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1676_
timestamp 1698431365
transform 1 0 17024 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1677_
timestamp 1698431365
transform 1 0 17696 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1678_
timestamp 1698431365
transform 1 0 14896 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1679_
timestamp 1698431365
transform 1 0 14112 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1680_
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1681_
timestamp 1698431365
transform 1 0 19152 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1682_
timestamp 1698431365
transform 1 0 21168 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1683_
timestamp 1698431365
transform 1 0 22176 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1684_
timestamp 1698431365
transform 1 0 17696 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1685_
timestamp 1698431365
transform 1 0 17696 0 1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1686_
timestamp 1698431365
transform 1 0 18368 0 -1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1687_
timestamp 1698431365
transform 1 0 21616 0 -1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1688_
timestamp 1698431365
transform 1 0 24416 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1689_
timestamp 1698431365
transform 1 0 26992 0 -1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1690_
timestamp 1698431365
transform 1 0 30240 0 1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1691_
timestamp 1698431365
transform 1 0 33824 0 -1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1692_
timestamp 1698431365
transform 1 0 34832 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1693_
timestamp 1698431365
transform 1 0 31136 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1694_
timestamp 1698431365
transform -1 0 32256 0 -1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1695_
timestamp 1698431365
transform 1 0 27104 0 -1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1696_
timestamp 1698431365
transform 1 0 29456 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1697_
timestamp 1698431365
transform 1 0 31696 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1698_
timestamp 1698431365
transform 1 0 32704 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1699_
timestamp 1698431365
transform 1 0 29232 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1700_
timestamp 1698431365
transform 1 0 28224 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1701_
timestamp 1698431365
transform -1 0 31696 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1702_
timestamp 1698431365
transform -1 0 28560 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1703_
timestamp 1698431365
transform -1 0 26096 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1704_
timestamp 1698431365
transform 1 0 20608 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1705_
timestamp 1698431365
transform 1 0 21616 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1706_
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1707_
timestamp 1698431365
transform 1 0 23632 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1708_
timestamp 1698431365
transform -1 0 28336 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1709_
timestamp 1698431365
transform 1 0 18928 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1710_
timestamp 1698431365
transform 1 0 19600 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1711_
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1712_
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1713_
timestamp 1698431365
transform 1 0 23968 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1714_
timestamp 1698431365
transform 1 0 15456 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1715_
timestamp 1698431365
transform 1 0 13776 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1716_
timestamp 1698431365
transform 1 0 14336 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1717_
timestamp 1698431365
transform 1 0 17584 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1718_
timestamp 1698431365
transform 1 0 19824 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1719_
timestamp 1698431365
transform -1 0 24864 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1720_
timestamp 1698431365
transform 1 0 15344 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1721_
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1722_
timestamp 1698431365
transform 1 0 14896 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1723_
timestamp 1698431365
transform 1 0 17472 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1724_
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1725_
timestamp 1698431365
transform 1 0 22624 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1726_
timestamp 1698431365
transform 1 0 20496 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1727_
timestamp 1698431365
transform 1 0 17696 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1728_
timestamp 1698431365
transform 1 0 20832 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1729_
timestamp 1698431365
transform 1 0 22848 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1730_
timestamp 1698431365
transform 1 0 25088 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1731_
timestamp 1698431365
transform 1 0 25424 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1732_
timestamp 1698431365
transform 1 0 16576 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1733_
timestamp 1698431365
transform 1 0 17472 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1734_
timestamp 1698431365
transform 1 0 20496 0 -1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1735_
timestamp 1698431365
transform 1 0 22624 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1736_
timestamp 1698431365
transform 1 0 24752 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1737_
timestamp 1698431365
transform 1 0 26208 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1738_
timestamp 1698431365
transform 1 0 14784 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1739_
timestamp 1698431365
transform 1 0 15344 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1740_
timestamp 1698431365
transform 1 0 16128 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1741_
timestamp 1698431365
transform 1 0 19712 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1742_
timestamp 1698431365
transform 1 0 22736 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1743_
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1744_
timestamp 1698431365
transform 1 0 36512 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1745_
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1746_
timestamp 1698431365
transform 1 0 43008 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1747_
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1748_
timestamp 1698431365
transform -1 0 44016 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1749_
timestamp 1698431365
transform 1 0 41552 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1750_
timestamp 1698431365
transform 1 0 43232 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1751_
timestamp 1698431365
transform 1 0 41440 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1752_
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1753_
timestamp 1698431365
transform 1 0 39200 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1754_
timestamp 1698431365
transform -1 0 28336 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1755_
timestamp 1698431365
transform -1 0 24864 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1756_
timestamp 1698431365
transform 1 0 13776 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1757_
timestamp 1698431365
transform 1 0 15344 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1758_
timestamp 1698431365
transform 1 0 15904 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1759_
timestamp 1698431365
transform 1 0 18032 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1760_
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1761_
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1762_
timestamp 1698431365
transform 1 0 37296 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1763_
timestamp 1698431365
transform 1 0 39200 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1764_
timestamp 1698431365
transform 1 0 45024 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1765_
timestamp 1698431365
transform 1 0 45024 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1766_
timestamp 1698431365
transform -1 0 41552 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1767_
timestamp 1698431365
transform -1 0 40096 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1768_
timestamp 1698431365
transform 1 0 31584 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1769_
timestamp 1698431365
transform 1 0 33264 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1770_
timestamp 1698431365
transform 1 0 35840 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1771_
timestamp 1698431365
transform -1 0 40096 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1772_
timestamp 1698431365
transform -1 0 39424 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1773_
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1774_
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1775_
timestamp 1698431365
transform 1 0 12992 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1776_
timestamp 1698431365
transform 1 0 15008 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1777_
timestamp 1698431365
transform 1 0 19376 0 -1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1778_
timestamp 1698431365
transform 1 0 22848 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1779_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1780_
timestamp 1698431365
transform 1 0 26208 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1781_
timestamp 1698431365
transform 1 0 26992 0 -1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1782_
timestamp 1698431365
transform -1 0 32816 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1783_
timestamp 1698431365
transform 1 0 29456 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1784_
timestamp 1698431365
transform 1 0 31360 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1785_
timestamp 1698431365
transform 1 0 30464 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1786_
timestamp 1698431365
transform 1 0 34496 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1787_
timestamp 1698431365
transform 1 0 37408 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1788_
timestamp 1698431365
transform 1 0 40768 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1789_
timestamp 1698431365
transform 1 0 43456 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1790_
timestamp 1698431365
transform -1 0 41104 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1791_
timestamp 1698431365
transform -1 0 37744 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1792_
timestamp 1698431365
transform 1 0 36960 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1793_
timestamp 1698431365
transform 1 0 39088 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1794_
timestamp 1698431365
transform 1 0 42896 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1795_
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1796_
timestamp 1698431365
transform 1 0 44800 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1797_
timestamp 1698431365
transform -1 0 41664 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1798_
timestamp 1698431365
transform 1 0 26768 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1799_
timestamp 1698431365
transform 1 0 26880 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1800_
timestamp 1698431365
transform 1 0 29456 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1801_
timestamp 1698431365
transform -1 0 34608 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1802_
timestamp 1698431365
transform -1 0 32704 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1803_
timestamp 1698431365
transform -1 0 32592 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1804_
timestamp 1698431365
transform -1 0 28784 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1805_
timestamp 1698431365
transform 1 0 17808 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1806_
timestamp 1698431365
transform 1 0 21056 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1807_
timestamp 1698431365
transform 1 0 22176 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1808_
timestamp 1698431365
transform 1 0 25088 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1809_
timestamp 1698431365
transform 1 0 26880 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1810_
timestamp 1698431365
transform 1 0 31360 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1811_
timestamp 1698431365
transform 1 0 33376 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1812_
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1813_
timestamp 1698431365
transform -1 0 40096 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1814_
timestamp 1698431365
transform 1 0 34496 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1815_
timestamp 1698431365
transform 1 0 33264 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1816_
timestamp 1698431365
transform 1 0 35392 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1817_
timestamp 1698431365
transform 1 0 38192 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1818_
timestamp 1698431365
transform 1 0 41216 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1819_
timestamp 1698431365
transform 1 0 43008 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1820_
timestamp 1698431365
transform -1 0 39648 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1821_
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1822_
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1823_
timestamp 1698431365
transform 1 0 38080 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1824_
timestamp 1698431365
transform 1 0 42224 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1825_
timestamp 1698431365
transform 1 0 43344 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1826_
timestamp 1698431365
transform 1 0 43120 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1827_
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1828_
timestamp 1698431365
transform 1 0 34832 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1829_
timestamp 1698431365
transform 1 0 36848 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1830_
timestamp 1698431365
transform -1 0 41104 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1831_
timestamp 1698431365
transform -1 0 39424 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1832_
timestamp 1698431365
transform 1 0 30688 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1833_
timestamp 1698431365
transform 1 0 32592 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1834_
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1835_
timestamp 1698431365
transform 1 0 38528 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1836_
timestamp 1698431365
transform -1 0 44016 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1837_
timestamp 1698431365
transform 1 0 37520 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1838_
timestamp 1698431365
transform 1 0 33600 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1839_
timestamp 1698431365
transform 1 0 33376 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1840_
timestamp 1698431365
transform 1 0 10864 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1841_
timestamp 1698431365
transform 1 0 8288 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1842_
timestamp 1698431365
transform 1 0 9856 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1843_
timestamp 1698431365
transform 1 0 11312 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1844_
timestamp 1698431365
transform 1 0 11648 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1845_
timestamp 1698431365
transform 1 0 8400 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1846_
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1847_
timestamp 1698431365
transform 1 0 10976 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1848_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1849_
timestamp 1698431365
transform -1 0 9856 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1850_
timestamp 1698431365
transform -1 0 10080 0 1 45472
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1851_
timestamp 1698431365
transform 1 0 7728 0 1 50176
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1852_
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1853_
timestamp 1698431365
transform -1 0 13552 0 -1 48608
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1854_
timestamp 1698431365
transform -1 0 10864 0 1 42336
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1855_
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1856_
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1857_
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1858_
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1859_
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1860_
timestamp 1698431365
transform 1 0 3248 0 -1 3136
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0814__I open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0817__A1
timestamp 1698431365
transform 1 0 5040 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0818__A2
timestamp 1698431365
transform -1 0 6160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0819__A1
timestamp 1698431365
transform 1 0 10304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0820__A1
timestamp 1698431365
transform 1 0 11088 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0822__A3
timestamp 1698431365
transform -1 0 4704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__I
timestamp 1698431365
transform 1 0 15344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0829__A1
timestamp 1698431365
transform -1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0829__A2
timestamp 1698431365
transform 1 0 6608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0831__I
timestamp 1698431365
transform 1 0 19936 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0832__I
timestamp 1698431365
transform 1 0 30688 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0836__I
timestamp 1698431365
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0838__I
timestamp 1698431365
transform 1 0 25872 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0839__A1
timestamp 1698431365
transform 1 0 29792 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0839__A4
timestamp 1698431365
transform 1 0 30352 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0840__I
timestamp 1698431365
transform 1 0 20384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0841__A1
timestamp 1698431365
transform 1 0 30016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0841__A2
timestamp 1698431365
transform 1 0 30912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__A1
timestamp 1698431365
transform 1 0 29904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0843__A1
timestamp 1698431365
transform 1 0 28560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0843__A3
timestamp 1698431365
transform -1 0 30688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0844__A1
timestamp 1698431365
transform 1 0 31136 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0844__A3
timestamp 1698431365
transform -1 0 32256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0845__A1
timestamp 1698431365
transform 1 0 26432 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0845__A3
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0845__A4
timestamp 1698431365
transform 1 0 26656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0846__A1
timestamp 1698431365
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0846__A2
timestamp 1698431365
transform 1 0 19712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0846__A3
timestamp 1698431365
transform 1 0 20160 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0847__A1
timestamp 1698431365
transform 1 0 17696 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0847__A3
timestamp 1698431365
transform -1 0 21616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0848__I
timestamp 1698431365
transform 1 0 41328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0849__A1
timestamp 1698431365
transform 1 0 32592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0849__A2
timestamp 1698431365
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0850__A1
timestamp 1698431365
transform 1 0 27440 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0850__A3
timestamp 1698431365
transform 1 0 26992 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0850__A4
timestamp 1698431365
transform 1 0 27888 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0851__A1
timestamp 1698431365
transform 1 0 24416 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0851__A2
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0852__A2
timestamp 1698431365
transform -1 0 24752 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0852__B1
timestamp 1698431365
transform -1 0 25200 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0853__A1
timestamp 1698431365
transform 1 0 31248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0854__A1
timestamp 1698431365
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0854__A2
timestamp 1698431365
transform 1 0 34944 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0855__A1
timestamp 1698431365
transform 1 0 30128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0856__A1
timestamp 1698431365
transform 1 0 19936 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0856__A2
timestamp 1698431365
transform 1 0 18144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0856__A3
timestamp 1698431365
transform -1 0 18816 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0857__A1
timestamp 1698431365
transform 1 0 35504 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0857__A2
timestamp 1698431365
transform 1 0 35056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0858__A1
timestamp 1698431365
transform 1 0 24640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0859__A2
timestamp 1698431365
transform -1 0 17920 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0859__B1
timestamp 1698431365
transform 1 0 19264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0861__A1
timestamp 1698431365
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__I
timestamp 1698431365
transform 1 0 18704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0863__A1
timestamp 1698431365
transform 1 0 30240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0863__A2
timestamp 1698431365
transform 1 0 30688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0864__A1
timestamp 1698431365
transform 1 0 35168 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0864__A2
timestamp 1698431365
transform 1 0 31808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0864__A3
timestamp 1698431365
transform 1 0 32032 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0864__A4
timestamp 1698431365
transform 1 0 31584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__A1
timestamp 1698431365
transform 1 0 18480 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__A2
timestamp 1698431365
transform 1 0 17584 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__A3
timestamp 1698431365
transform 1 0 17136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__A4
timestamp 1698431365
transform 1 0 18032 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0867__A1
timestamp 1698431365
transform 1 0 26096 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0867__A2
timestamp 1698431365
transform 1 0 26544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0868__A1
timestamp 1698431365
transform -1 0 33376 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0868__A2
timestamp 1698431365
transform 1 0 28112 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0869__A1
timestamp 1698431365
transform -1 0 31248 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0869__A3
timestamp 1698431365
transform 1 0 32032 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0871__A2
timestamp 1698431365
transform 1 0 38416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0871__B1
timestamp 1698431365
transform 1 0 38192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0872__A2
timestamp 1698431365
transform 1 0 38752 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0872__B1
timestamp 1698431365
transform 1 0 39200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0873__A1
timestamp 1698431365
transform 1 0 36064 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0873__A2
timestamp 1698431365
transform 1 0 34608 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0874__A1
timestamp 1698431365
transform 1 0 29792 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0874__A3
timestamp 1698431365
transform 1 0 35728 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__A1
timestamp 1698431365
transform 1 0 28112 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__A3
timestamp 1698431365
transform 1 0 28560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0877__A1
timestamp 1698431365
transform 1 0 29232 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0877__A2
timestamp 1698431365
transform 1 0 28560 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0879__A1
timestamp 1698431365
transform 1 0 31808 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0879__A2
timestamp 1698431365
transform -1 0 31920 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0879__A3
timestamp 1698431365
transform -1 0 32368 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0879__A4
timestamp 1698431365
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0880__A1
timestamp 1698431365
transform 1 0 32704 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0880__A3
timestamp 1698431365
transform 1 0 36512 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0882__A2
timestamp 1698431365
transform 1 0 34160 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0882__B1
timestamp 1698431365
transform 1 0 37072 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__A2
timestamp 1698431365
transform 1 0 34048 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__B1
timestamp 1698431365
transform 1 0 33600 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0886__A1
timestamp 1698431365
transform 1 0 24080 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0886__A3
timestamp 1698431365
transform 1 0 23296 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0886__A4
timestamp 1698431365
transform 1 0 28896 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0887__A1
timestamp 1698431365
transform 1 0 18704 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0887__A3
timestamp 1698431365
transform -1 0 19936 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0890__A1
timestamp 1698431365
transform 1 0 23968 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0890__A3
timestamp 1698431365
transform 1 0 24416 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0892__A1
timestamp 1698431365
transform 1 0 22400 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0892__A3
timestamp 1698431365
transform 1 0 24528 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0893__I
timestamp 1698431365
transform 1 0 21392 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__A1
timestamp 1698431365
transform -1 0 18928 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__A2
timestamp 1698431365
transform 1 0 19936 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__A3
timestamp 1698431365
transform 1 0 19488 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__A4
timestamp 1698431365
transform 1 0 20384 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0895__A1
timestamp 1698431365
transform 1 0 24192 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0895__A2
timestamp 1698431365
transform -1 0 23968 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0895__A3
timestamp 1698431365
transform 1 0 24640 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0897__A1
timestamp 1698431365
transform 1 0 23296 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0897__A3
timestamp 1698431365
transform 1 0 22848 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0897__B1
timestamp 1698431365
transform 1 0 23072 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__A1
timestamp 1698431365
transform -1 0 22064 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__A2
timestamp 1698431365
transform 1 0 20608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__A3
timestamp 1698431365
transform 1 0 21392 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__A4
timestamp 1698431365
transform 1 0 25312 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0900__A1
timestamp 1698431365
transform 1 0 21504 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0900__A2
timestamp 1698431365
transform 1 0 21056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0900__A4
timestamp 1698431365
transform -1 0 23184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0904__A1
timestamp 1698431365
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0904__A2
timestamp 1698431365
transform 1 0 33600 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0904__A3
timestamp 1698431365
transform 1 0 34048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0904__A4
timestamp 1698431365
transform 1 0 39424 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0905__A1
timestamp 1698431365
transform 1 0 21952 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0905__A2
timestamp 1698431365
transform 1 0 24192 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0906__B
timestamp 1698431365
transform 1 0 39312 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__A1
timestamp 1698431365
transform -1 0 34720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__A2
timestamp 1698431365
transform 1 0 34048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__A4
timestamp 1698431365
transform 1 0 33600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0909__A1
timestamp 1698431365
transform 1 0 40544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0909__A3
timestamp 1698431365
transform 1 0 37632 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0909__A4
timestamp 1698431365
transform 1 0 38080 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__A1
timestamp 1698431365
transform 1 0 42784 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__A2
timestamp 1698431365
transform 1 0 40992 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0913__A1
timestamp 1698431365
transform 1 0 31024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0913__A2
timestamp 1698431365
transform 1 0 29568 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0913__A3
timestamp 1698431365
transform 1 0 31472 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0913__A4
timestamp 1698431365
transform 1 0 35056 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0915__A2
timestamp 1698431365
transform 1 0 37632 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0915__A3
timestamp 1698431365
transform 1 0 40992 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0917__A1
timestamp 1698431365
transform 1 0 31808 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0917__A3
timestamp 1698431365
transform 1 0 32256 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0918__A1
timestamp 1698431365
transform 1 0 40768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0918__A3
timestamp 1698431365
transform 1 0 38192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0918__A4
timestamp 1698431365
transform 1 0 40320 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__A2
timestamp 1698431365
transform 1 0 38640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__A1
timestamp 1698431365
transform 1 0 37296 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__A2
timestamp 1698431365
transform 1 0 37744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__A3
timestamp 1698431365
transform 1 0 34608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0922__A3
timestamp 1698431365
transform 1 0 21392 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0922__B1
timestamp 1698431365
transform 1 0 20944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__A1
timestamp 1698431365
transform -1 0 11424 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__A2
timestamp 1698431365
transform 1 0 9184 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__A1
timestamp 1698431365
transform 1 0 8400 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0925__A1
timestamp 1698431365
transform 1 0 31472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0925__A2
timestamp 1698431365
transform 1 0 31920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0926__A2
timestamp 1698431365
transform -1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0927__A1
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0927__A3
timestamp 1698431365
transform -1 0 30240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0929__A1
timestamp 1698431365
transform -1 0 19824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0929__A3
timestamp 1698431365
transform 1 0 19152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0930__A1
timestamp 1698431365
transform 1 0 19488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0930__A3
timestamp 1698431365
transform 1 0 19040 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0931__A2
timestamp 1698431365
transform 1 0 24640 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0931__B1
timestamp 1698431365
transform 1 0 24192 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0932__A2
timestamp 1698431365
transform -1 0 18704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0932__B1
timestamp 1698431365
transform -1 0 19152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0936__A2
timestamp 1698431365
transform 1 0 41440 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0936__B1
timestamp 1698431365
transform 1 0 40320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0937__A2
timestamp 1698431365
transform -1 0 37296 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0937__B1
timestamp 1698431365
transform -1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0940__A2
timestamp 1698431365
transform 1 0 34272 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0940__B1
timestamp 1698431365
transform 1 0 37072 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__A2
timestamp 1698431365
transform -1 0 34272 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__B1
timestamp 1698431365
transform 1 0 34496 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0943__A1
timestamp 1698431365
transform -1 0 19712 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0943__A3
timestamp 1698431365
transform -1 0 20384 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0947__A1
timestamp 1698431365
transform -1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0947__A3
timestamp 1698431365
transform -1 0 24416 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0950__A1
timestamp 1698431365
transform 1 0 23744 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0950__A3
timestamp 1698431365
transform 1 0 24640 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0950__B1
timestamp 1698431365
transform 1 0 24192 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0952__A1
timestamp 1698431365
transform 1 0 21392 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0952__A2
timestamp 1698431365
transform 1 0 18480 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0952__A4
timestamp 1698431365
transform -1 0 18704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0956__B
timestamp 1698431365
transform -1 0 42560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0958__A1
timestamp 1698431365
transform 1 0 43680 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0958__A3
timestamp 1698431365
transform 1 0 41440 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0958__A4
timestamp 1698431365
transform 1 0 41216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0962__A2
timestamp 1698431365
transform -1 0 40320 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0962__A3
timestamp 1698431365
transform 1 0 43120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0964__A1
timestamp 1698431365
transform 1 0 43008 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0964__A3
timestamp 1698431365
transform 1 0 42112 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0964__A4
timestamp 1698431365
transform 1 0 42896 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0965__A2
timestamp 1698431365
transform -1 0 41216 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__A1
timestamp 1698431365
transform 1 0 39312 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__A2
timestamp 1698431365
transform 1 0 40320 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__A3
timestamp 1698431365
transform 1 0 35504 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0968__A1
timestamp 1698431365
transform -1 0 23968 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0968__A3
timestamp 1698431365
transform -1 0 23520 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0968__B1
timestamp 1698431365
transform 1 0 24192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0969__A1
timestamp 1698431365
transform -1 0 14896 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0969__A2
timestamp 1698431365
transform 1 0 12880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0970__A1
timestamp 1698431365
transform 1 0 9744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0971__A2
timestamp 1698431365
transform 1 0 32144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0972__A1
timestamp 1698431365
transform 1 0 30128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0972__A3
timestamp 1698431365
transform 1 0 31136 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__A1
timestamp 1698431365
transform 1 0 22960 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__A3
timestamp 1698431365
transform 1 0 22512 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0975__A1
timestamp 1698431365
transform 1 0 18592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0975__A3
timestamp 1698431365
transform 1 0 20272 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0976__A2
timestamp 1698431365
transform 1 0 23968 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0976__B1
timestamp 1698431365
transform 1 0 24864 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0977__A2
timestamp 1698431365
transform 1 0 19936 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0977__B1
timestamp 1698431365
transform 1 0 20160 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0981__A2
timestamp 1698431365
transform 1 0 38416 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0981__B1
timestamp 1698431365
transform 1 0 37968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0982__A2
timestamp 1698431365
transform 1 0 35168 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0982__B1
timestamp 1698431365
transform 1 0 35616 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__A2
timestamp 1698431365
transform -1 0 35280 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__B1
timestamp 1698431365
transform -1 0 34384 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__A2
timestamp 1698431365
transform 1 0 33152 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__B1
timestamp 1698431365
transform 1 0 34496 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A1
timestamp 1698431365
transform 1 0 20272 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A3
timestamp 1698431365
transform 1 0 18816 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0992__A1
timestamp 1698431365
transform 1 0 26096 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0992__A3
timestamp 1698431365
transform 1 0 25648 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__A1
timestamp 1698431365
transform 1 0 25760 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__A3
timestamp 1698431365
transform 1 0 25312 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__B1
timestamp 1698431365
transform 1 0 24528 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0997__A1
timestamp 1698431365
transform 1 0 21392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0997__A2
timestamp 1698431365
transform 1 0 19600 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0997__A4
timestamp 1698431365
transform 1 0 21840 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1001__B
timestamp 1698431365
transform -1 0 43008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A1
timestamp 1698431365
transform 1 0 44800 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A3
timestamp 1698431365
transform 1 0 43344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A4
timestamp 1698431365
transform 1 0 42336 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1007__A2
timestamp 1698431365
transform 1 0 40320 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1007__A3
timestamp 1698431365
transform 1 0 43680 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__A1
timestamp 1698431365
transform 1 0 44016 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__A3
timestamp 1698431365
transform 1 0 42672 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__A4
timestamp 1698431365
transform 1 0 43120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1010__A2
timestamp 1698431365
transform 1 0 41216 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__A1
timestamp 1698431365
transform 1 0 39872 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__A2
timestamp 1698431365
transform 1 0 39872 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__A3
timestamp 1698431365
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1013__A1
timestamp 1698431365
transform -1 0 24752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1013__A3
timestamp 1698431365
transform -1 0 25536 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1013__B1
timestamp 1698431365
transform 1 0 24304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1014__A1
timestamp 1698431365
transform -1 0 12656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1014__A2
timestamp 1698431365
transform 1 0 10864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1015__A1
timestamp 1698431365
transform 1 0 9296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__A2
timestamp 1698431365
transform 1 0 31360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__A1
timestamp 1698431365
transform 1 0 30912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__A3
timestamp 1698431365
transform 1 0 31920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1019__A1
timestamp 1698431365
transform 1 0 22848 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1019__A3
timestamp 1698431365
transform 1 0 23968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1020__A1
timestamp 1698431365
transform 1 0 21840 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1020__A3
timestamp 1698431365
transform -1 0 23968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__A2
timestamp 1698431365
transform 1 0 24304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__B1
timestamp 1698431365
transform 1 0 25424 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1022__A2
timestamp 1698431365
transform 1 0 22176 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1022__B1
timestamp 1698431365
transform 1 0 23184 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__A2
timestamp 1698431365
transform 1 0 24864 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1026__A2
timestamp 1698431365
transform 1 0 34496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1026__B1
timestamp 1698431365
transform 1 0 34048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A2
timestamp 1698431365
transform -1 0 35504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__B1
timestamp 1698431365
transform -1 0 35056 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1030__A2
timestamp 1698431365
transform 1 0 33824 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1030__B1
timestamp 1698431365
transform -1 0 34832 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1031__A2
timestamp 1698431365
transform 1 0 37968 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1031__B1
timestamp 1698431365
transform 1 0 31920 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1033__A1
timestamp 1698431365
transform 1 0 23184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1033__A3
timestamp 1698431365
transform 1 0 22736 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1037__A1
timestamp 1698431365
transform -1 0 25536 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1037__A3
timestamp 1698431365
transform 1 0 27888 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A1
timestamp 1698431365
transform -1 0 28112 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A3
timestamp 1698431365
transform -1 0 26992 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__B1
timestamp 1698431365
transform 1 0 28336 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__A1
timestamp 1698431365
transform 1 0 21840 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__A2
timestamp 1698431365
transform 1 0 18928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__A4
timestamp 1698431365
transform 1 0 22288 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__B
timestamp 1698431365
transform 1 0 41888 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__A1
timestamp 1698431365
transform 1 0 40320 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__A3
timestamp 1698431365
transform 1 0 41216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__A4
timestamp 1698431365
transform 1 0 40768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__A2
timestamp 1698431365
transform 1 0 41440 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__A3
timestamp 1698431365
transform 1 0 44128 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1054__A1
timestamp 1698431365
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1054__A3
timestamp 1698431365
transform 1 0 41328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1054__A4
timestamp 1698431365
transform 1 0 42336 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__A2
timestamp 1698431365
transform 1 0 42784 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__A1
timestamp 1698431365
transform 1 0 37184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__A2
timestamp 1698431365
transform 1 0 37632 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__A3
timestamp 1698431365
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1058__A3
timestamp 1698431365
transform 1 0 27216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1058__B1
timestamp 1698431365
transform 1 0 26768 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1059__A1
timestamp 1698431365
transform 1 0 12768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1059__A2
timestamp 1698431365
transform 1 0 11200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1060__A1
timestamp 1698431365
transform 1 0 10192 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1062__A1
timestamp 1698431365
transform -1 0 30464 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1062__A2
timestamp 1698431365
transform 1 0 29792 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__A1
timestamp 1698431365
transform 1 0 29008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__A3
timestamp 1698431365
transform 1 0 27328 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__A4
timestamp 1698431365
transform 1 0 29232 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1064__A1
timestamp 1698431365
transform 1 0 28000 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1065__I
timestamp 1698431365
transform 1 0 28112 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1066__A1
timestamp 1698431365
transform 1 0 25872 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__A1
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__A2
timestamp 1698431365
transform 1 0 20496 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__A4
timestamp 1698431365
transform 1 0 21952 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1068__A2
timestamp 1698431365
transform 1 0 28224 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__A1
timestamp 1698431365
transform 1 0 28224 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__A2
timestamp 1698431365
transform 1 0 29232 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__A2
timestamp 1698431365
transform 1 0 28224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__B2
timestamp 1698431365
transform 1 0 29680 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1071__A1
timestamp 1698431365
transform 1 0 27104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1071__A2
timestamp 1698431365
transform 1 0 25760 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1072__A1
timestamp 1698431365
transform 1 0 25984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1072__A2
timestamp 1698431365
transform 1 0 29232 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__A1
timestamp 1698431365
transform 1 0 30688 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__A3
timestamp 1698431365
transform 1 0 31136 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__A1
timestamp 1698431365
transform 1 0 31920 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__A2
timestamp 1698431365
transform -1 0 31472 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__A3
timestamp 1698431365
transform 1 0 32368 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__A1
timestamp 1698431365
transform 1 0 30240 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__B2
timestamp 1698431365
transform 1 0 30688 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__A1
timestamp 1698431365
transform 1 0 28112 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__A2
timestamp 1698431365
transform 1 0 28560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__A3
timestamp 1698431365
transform 1 0 28560 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__A4
timestamp 1698431365
transform -1 0 34384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__B1
timestamp 1698431365
transform -1 0 26544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__A1
timestamp 1698431365
transform 1 0 29232 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__A2
timestamp 1698431365
transform 1 0 24640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__A1
timestamp 1698431365
transform -1 0 30128 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__A2
timestamp 1698431365
transform -1 0 31584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__B2
timestamp 1698431365
transform -1 0 29456 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__A2
timestamp 1698431365
transform 1 0 34048 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__B1
timestamp 1698431365
transform 1 0 33152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__A1
timestamp 1698431365
transform 1 0 34496 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__A2
timestamp 1698431365
transform 1 0 32704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__A4
timestamp 1698431365
transform 1 0 35280 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__A1
timestamp 1698431365
transform 1 0 34944 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__A2
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__A3
timestamp 1698431365
transform 1 0 35728 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__A1
timestamp 1698431365
transform 1 0 33600 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__A3
timestamp 1698431365
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__B1
timestamp 1698431365
transform -1 0 35616 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__B2
timestamp 1698431365
transform -1 0 34944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__A1
timestamp 1698431365
transform 1 0 38080 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__A3
timestamp 1698431365
transform 1 0 36400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__A4
timestamp 1698431365
transform 1 0 36624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__A2
timestamp 1698431365
transform 1 0 35504 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__A1
timestamp 1698431365
transform 1 0 43792 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__A3
timestamp 1698431365
transform 1 0 42896 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__A4
timestamp 1698431365
transform 1 0 41888 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__A1
timestamp 1698431365
transform 1 0 25312 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__A3
timestamp 1698431365
transform 1 0 26656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__A1
timestamp 1698431365
transform 1 0 25872 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__A3
timestamp 1698431365
transform 1 0 26096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__A1
timestamp 1698431365
transform 1 0 39424 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__A2
timestamp 1698431365
transform -1 0 36848 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__A1
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__A2
timestamp 1698431365
transform 1 0 31360 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1104__A3
timestamp 1698431365
transform 1 0 27328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1105__I
timestamp 1698431365
transform 1 0 28224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__A1
timestamp 1698431365
transform 1 0 25760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__A3
timestamp 1698431365
transform 1 0 27664 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__A1
timestamp 1698431365
transform 1 0 28448 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__A3
timestamp 1698431365
transform 1 0 29232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__B
timestamp 1698431365
transform 1 0 31248 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__A2
timestamp 1698431365
transform 1 0 34048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1109__A1
timestamp 1698431365
transform 1 0 32368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1112__A2
timestamp 1698431365
transform 1 0 12768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1112__B
timestamp 1698431365
transform 1 0 10640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1114__A1
timestamp 1698431365
transform -1 0 9968 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1115__A2
timestamp 1698431365
transform 1 0 10752 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__A1
timestamp 1698431365
transform 1 0 28784 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1118__A2
timestamp 1698431365
transform 1 0 29232 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__A1
timestamp 1698431365
transform 1 0 29568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__A3
timestamp 1698431365
transform 1 0 32480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A1
timestamp 1698431365
transform 1 0 30464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A2
timestamp 1698431365
transform -1 0 33824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A3
timestamp 1698431365
transform 1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A4
timestamp 1698431365
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__A1
timestamp 1698431365
transform -1 0 28896 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__A2
timestamp 1698431365
transform 1 0 31136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__B2
timestamp 1698431365
transform 1 0 30912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1123__A4
timestamp 1698431365
transform 1 0 30240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1124__A2
timestamp 1698431365
transform -1 0 30800 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__B1
timestamp 1698431365
transform 1 0 26992 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__A2
timestamp 1698431365
transform 1 0 26768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1128__A1
timestamp 1698431365
transform 1 0 26544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1128__A3
timestamp 1698431365
transform -1 0 27216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__B1
timestamp 1698431365
transform 1 0 26544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1130__A1
timestamp 1698431365
transform 1 0 29680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1130__A2
timestamp 1698431365
transform 1 0 29568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1131__A2
timestamp 1698431365
transform 1 0 32144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1134__A1
timestamp 1698431365
transform 1 0 32480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1135__I
timestamp 1698431365
transform -1 0 36288 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__B1
timestamp 1698431365
transform 1 0 36176 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__B1
timestamp 1698431365
transform -1 0 37296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__B2
timestamp 1698431365
transform 1 0 37072 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1138__B1
timestamp 1698431365
transform 1 0 34720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1138__B2
timestamp 1698431365
transform 1 0 35952 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1140__B
timestamp 1698431365
transform -1 0 27104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1140__C
timestamp 1698431365
transform 1 0 27328 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1141__A1
timestamp 1698431365
transform 1 0 29904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1141__A3
timestamp 1698431365
transform -1 0 31920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1141__A4
timestamp 1698431365
transform -1 0 32368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1143__A1
timestamp 1698431365
transform 1 0 26544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1143__A3
timestamp 1698431365
transform 1 0 27776 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1144__A2
timestamp 1698431365
transform 1 0 26656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1145__A2
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1146__A1
timestamp 1698431365
transform -1 0 30688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1148__A2
timestamp 1698431365
transform 1 0 13552 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1148__B
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__A1
timestamp 1698431365
transform 1 0 16240 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1151__A1
timestamp 1698431365
transform 1 0 4816 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__A1
timestamp 1698431365
transform 1 0 3808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__A3
timestamp 1698431365
transform 1 0 4256 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1156__I
timestamp 1698431365
transform 1 0 6160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1157__A2
timestamp 1698431365
transform 1 0 4144 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1159__A1
timestamp 1698431365
transform -1 0 7392 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1160__A1
timestamp 1698431365
transform -1 0 8624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1161__A1
timestamp 1698431365
transform -1 0 8176 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1163__A1
timestamp 1698431365
transform -1 0 9072 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1164__A1
timestamp 1698431365
transform 1 0 3136 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__A1
timestamp 1698431365
transform 1 0 2576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__B
timestamp 1698431365
transform -1 0 2352 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__A2
timestamp 1698431365
transform -1 0 2576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1177__A1
timestamp 1698431365
transform -1 0 6832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1177__A2
timestamp 1698431365
transform 1 0 5600 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1187__A1
timestamp 1698431365
transform 1 0 2800 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1190__A1
timestamp 1698431365
transform 1 0 7168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1191__A1
timestamp 1698431365
transform -1 0 3920 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__B
timestamp 1698431365
transform 1 0 3808 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__A1
timestamp 1698431365
transform 1 0 3248 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1194__A1
timestamp 1698431365
transform 1 0 2240 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1194__A2
timestamp 1698431365
transform 1 0 4592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1196__A2
timestamp 1698431365
transform 1 0 1904 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1196__B
timestamp 1698431365
transform 1 0 2352 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1197__A1
timestamp 1698431365
transform 1 0 7168 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1200__A1
timestamp 1698431365
transform -1 0 7504 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1205__A1
timestamp 1698431365
transform 1 0 5152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1206__A1
timestamp 1698431365
transform 1 0 2800 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1207__A1
timestamp 1698431365
transform 1 0 8288 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__A1
timestamp 1698431365
transform -1 0 9072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1215__A1
timestamp 1698431365
transform 1 0 8064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__A2
timestamp 1698431365
transform 1 0 3696 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__B
timestamp 1698431365
transform 1 0 4144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1217__A1
timestamp 1698431365
transform 1 0 3696 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1217__A2
timestamp 1698431365
transform 1 0 2688 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1219__B2
timestamp 1698431365
transform 1 0 6048 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1220__1_I
timestamp 1698431365
transform 1 0 8960 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1222__A1
timestamp 1698431365
transform 1 0 9744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1225__A1
timestamp 1698431365
transform 1 0 9632 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1227__I0
timestamp 1698431365
transform 1 0 6160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1228__A1
timestamp 1698431365
transform 1 0 7728 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1230__A1
timestamp 1698431365
transform 1 0 10080 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1231__A1
timestamp 1698431365
transform -1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1231__A2
timestamp 1698431365
transform -1 0 4368 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1231__B
timestamp 1698431365
transform -1 0 4816 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1234__A1
timestamp 1698431365
transform 1 0 9744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1238__I0
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1239__A1
timestamp 1698431365
transform 1 0 6608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1241__A1
timestamp 1698431365
transform -1 0 4368 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1242__A1
timestamp 1698431365
transform 1 0 8400 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1242__A2
timestamp 1698431365
transform 1 0 8848 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1242__B
timestamp 1698431365
transform 1 0 9408 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1245__I
timestamp 1698431365
transform 1 0 10192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1246__B1
timestamp 1698431365
transform 1 0 11424 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1248__A1
timestamp 1698431365
transform -1 0 7728 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1249__A1
timestamp 1698431365
transform -1 0 4144 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1251__A1
timestamp 1698431365
transform 1 0 6832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1254__A1
timestamp 1698431365
transform -1 0 4256 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1254__A2
timestamp 1698431365
transform 1 0 4144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1254__B
timestamp 1698431365
transform 1 0 3584 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__A1
timestamp 1698431365
transform 1 0 4928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1256__A1
timestamp 1698431365
transform -1 0 11872 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1258__A1
timestamp 1698431365
transform -1 0 5040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1261__A1
timestamp 1698431365
transform 1 0 10528 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__A2
timestamp 1698431365
transform 1 0 2240 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__B
timestamp 1698431365
transform 1 0 3248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1263__A1
timestamp 1698431365
transform 1 0 3248 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1263__A2
timestamp 1698431365
transform 1 0 2352 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1263__B1
timestamp 1698431365
transform -1 0 3024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1264__A1
timestamp 1698431365
transform -1 0 2016 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1265__B2
timestamp 1698431365
transform 1 0 4368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1266__A1
timestamp 1698431365
transform 1 0 4704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1268__C
timestamp 1698431365
transform -1 0 2576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1269__A1
timestamp 1698431365
transform -1 0 2016 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1269__A2
timestamp 1698431365
transform -1 0 3584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__A2
timestamp 1698431365
transform 1 0 2352 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__A1
timestamp 1698431365
transform 1 0 2800 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1273__I
timestamp 1698431365
transform 1 0 13888 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1274__A2
timestamp 1698431365
transform 1 0 11760 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1276__I
timestamp 1698431365
transform 1 0 15456 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1277__I
timestamp 1698431365
transform 1 0 15904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1278__A2
timestamp 1698431365
transform 1 0 14224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__A2
timestamp 1698431365
transform 1 0 15456 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1282__A2
timestamp 1698431365
transform 1 0 16800 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1284__A2
timestamp 1698431365
transform 1 0 17472 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1286__A2
timestamp 1698431365
transform 1 0 14448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1288__A2
timestamp 1698431365
transform 1 0 14560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1289__I
timestamp 1698431365
transform 1 0 14896 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1290__I
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1291__A2
timestamp 1698431365
transform 1 0 18928 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1292__A2
timestamp 1698431365
transform 1 0 18480 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1293__A2
timestamp 1698431365
transform 1 0 20944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1294__I
timestamp 1698431365
transform 1 0 17472 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1295__A2
timestamp 1698431365
transform 1 0 25872 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A2
timestamp 1698431365
transform 1 0 28560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1298__A1
timestamp 1698431365
transform -1 0 33376 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1298__A2
timestamp 1698431365
transform -1 0 33824 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1300__A2
timestamp 1698431365
transform 1 0 38080 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1301__A2
timestamp 1698431365
transform 1 0 39648 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1302__A2
timestamp 1698431365
transform 1 0 40544 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1303__A2
timestamp 1698431365
transform 1 0 42448 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1304__A1
timestamp 1698431365
transform 1 0 29680 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1304__A2
timestamp 1698431365
transform -1 0 27888 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1306__A2
timestamp 1698431365
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1308__A2
timestamp 1698431365
transform 1 0 34048 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1309__A2
timestamp 1698431365
transform 1 0 37520 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1310__A2
timestamp 1698431365
transform 1 0 32480 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1311__A2
timestamp 1698431365
transform 1 0 29792 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1312__A1
timestamp 1698431365
transform 1 0 28224 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1312__A2
timestamp 1698431365
transform 1 0 26208 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1314__A2
timestamp 1698431365
transform 1 0 29232 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1316__A2
timestamp 1698431365
transform 1 0 14896 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1318__A2
timestamp 1698431365
transform 1 0 15120 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1320__A2
timestamp 1698431365
transform 1 0 17472 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1322__A2
timestamp 1698431365
transform 1 0 16128 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1324__I
timestamp 1698431365
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1325__A2
timestamp 1698431365
transform 1 0 21392 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1327__A2
timestamp 1698431365
transform 1 0 19488 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1329__I
timestamp 1698431365
transform 1 0 19040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1330__A1
timestamp 1698431365
transform 1 0 17248 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1330__A2
timestamp 1698431365
transform 1 0 16800 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1332__A2
timestamp 1698431365
transform -1 0 18928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1334__A2
timestamp 1698431365
transform 1 0 20384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1336__A2
timestamp 1698431365
transform 1 0 22736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1338__A2
timestamp 1698431365
transform 1 0 24528 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1340__A2
timestamp 1698431365
transform 1 0 19824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1342__A2
timestamp 1698431365
transform 1 0 18928 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1343__A2
timestamp 1698431365
transform 1 0 20720 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1344__A2
timestamp 1698431365
transform 1 0 22400 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__A2
timestamp 1698431365
transform 1 0 25872 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1346__A1
timestamp 1698431365
transform -1 0 27664 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1346__A2
timestamp 1698431365
transform 1 0 29232 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1348__A1
timestamp 1698431365
transform 1 0 30912 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1348__A2
timestamp 1698431365
transform 1 0 30912 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1350__A2
timestamp 1698431365
transform 1 0 34160 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__A2
timestamp 1698431365
transform 1 0 35280 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1352__A2
timestamp 1698431365
transform 1 0 32480 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1353__A2
timestamp 1698431365
transform 1 0 29904 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1354__A1
timestamp 1698431365
transform 1 0 30688 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1354__A2
timestamp 1698431365
transform 1 0 29456 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1356__A1
timestamp 1698431365
transform 1 0 31584 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1356__A2
timestamp 1698431365
transform 1 0 31136 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__A2
timestamp 1698431365
transform -1 0 32704 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1360__A2
timestamp 1698431365
transform 1 0 32032 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__A2
timestamp 1698431365
transform 1 0 30576 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1364__A2
timestamp 1698431365
transform 1 0 31024 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1366__A2
timestamp 1698431365
transform 1 0 31024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1368__A1
timestamp 1698431365
transform 1 0 28784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1368__A2
timestamp 1698431365
transform -1 0 30352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1370__A2
timestamp 1698431365
transform 1 0 23520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__A2
timestamp 1698431365
transform -1 0 21952 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1374__A2
timestamp 1698431365
transform 1 0 22736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__A2
timestamp 1698431365
transform 1 0 27328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1378__A2
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1379__A2
timestamp 1698431365
transform 1 0 26880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1381__A2
timestamp 1698431365
transform 1 0 20944 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1383__A2
timestamp 1698431365
transform 1 0 20720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1385__A2
timestamp 1698431365
transform 1 0 22064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1387__A2
timestamp 1698431365
transform 1 0 23856 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1389__A2
timestamp 1698431365
transform 1 0 25312 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1390__A2
timestamp 1698431365
transform 1 0 19600 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__A2
timestamp 1698431365
transform 1 0 18368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1394__A2
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1396__A2
timestamp 1698431365
transform 1 0 18480 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1398__A2
timestamp 1698431365
transform 1 0 21392 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__A2
timestamp 1698431365
transform 1 0 24192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__A2
timestamp 1698431365
transform 1 0 19936 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1404__A2
timestamp 1698431365
transform 1 0 18704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1406__I
timestamp 1698431365
transform 1 0 17920 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1407__A2
timestamp 1698431365
transform 1 0 16800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A2
timestamp 1698431365
transform 1 0 18704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1411__A2
timestamp 1698431365
transform 1 0 20720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1413__A2
timestamp 1698431365
transform 1 0 23632 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1415__A2
timestamp 1698431365
transform 1 0 22288 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1417__A2
timestamp 1698431365
transform 1 0 19376 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1418__A2
timestamp 1698431365
transform 1 0 22288 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1419__A2
timestamp 1698431365
transform 1 0 23296 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1420__A2
timestamp 1698431365
transform 1 0 24304 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1421__A2
timestamp 1698431365
transform 1 0 26096 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1423__A1
timestamp 1698431365
transform -1 0 28672 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1423__A2
timestamp 1698431365
transform -1 0 27328 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1425__A2
timestamp 1698431365
transform 1 0 18480 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1426__A2
timestamp 1698431365
transform 1 0 20720 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1427__A2
timestamp 1698431365
transform 1 0 23520 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1428__A2
timestamp 1698431365
transform 1 0 26096 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1429__A1
timestamp 1698431365
transform 1 0 28448 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1429__A2
timestamp 1698431365
transform 1 0 27104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__A2
timestamp 1698431365
transform 1 0 30128 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1433__A2
timestamp 1698431365
transform 1 0 18144 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1435__A2
timestamp 1698431365
transform 1 0 18480 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1437__A2
timestamp 1698431365
transform 1 0 19040 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1439__A2
timestamp 1698431365
transform 1 0 23184 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__A2
timestamp 1698431365
transform 1 0 24864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1443__I
timestamp 1698431365
transform 1 0 34496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1444__A2
timestamp 1698431365
transform 1 0 28784 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1446__A2
timestamp 1698431365
transform 1 0 38864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1448__A2
timestamp 1698431365
transform 1 0 43008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1450__A2
timestamp 1698431365
transform 1 0 44240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1452__A2
timestamp 1698431365
transform 1 0 41888 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__A2
timestamp 1698431365
transform 1 0 41888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__A1
timestamp 1698431365
transform -1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__A2
timestamp 1698431365
transform 1 0 43792 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1458__A2
timestamp 1698431365
transform 1 0 41440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1459__A2
timestamp 1698431365
transform 1 0 40992 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1460__A2
timestamp 1698431365
transform -1 0 39872 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1461__A2
timestamp 1698431365
transform 1 0 33488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__A1
timestamp 1698431365
transform 1 0 25536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__A2
timestamp 1698431365
transform 1 0 25312 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1464__A2
timestamp 1698431365
transform 1 0 16800 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__A2
timestamp 1698431365
transform 1 0 16128 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1467__A2
timestamp 1698431365
transform 1 0 18256 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1468__A2
timestamp 1698431365
transform 1 0 18592 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__A2
timestamp 1698431365
transform 1 0 23856 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1470__A2
timestamp 1698431365
transform -1 0 26656 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1472__A2
timestamp 1698431365
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1474__A2
timestamp 1698431365
transform 1 0 40096 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1476__A2
timestamp 1698431365
transform 1 0 43344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__A2
timestamp 1698431365
transform 1 0 44240 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1480__A2
timestamp 1698431365
transform 1 0 40432 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1482__A2
timestamp 1698431365
transform 1 0 36848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__A2
timestamp 1698431365
transform 1 0 31584 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1486__A2
timestamp 1698431365
transform 1 0 33376 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A2
timestamp 1698431365
transform 1 0 35728 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__A2
timestamp 1698431365
transform 1 0 36400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1492__A2
timestamp 1698431365
transform 1 0 34944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__A2
timestamp 1698431365
transform 1 0 34384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1496__A1
timestamp 1698431365
transform 1 0 34720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1496__A2
timestamp 1698431365
transform -1 0 33600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1498__A2
timestamp 1698431365
transform -1 0 14000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__A2
timestamp 1698431365
transform 1 0 15456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1502__A2
timestamp 1698431365
transform -1 0 18816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1504__A2
timestamp 1698431365
transform 1 0 24192 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1506__A2
timestamp 1698431365
transform 1 0 26432 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A2
timestamp 1698431365
transform 1 0 27888 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1510__A2
timestamp 1698431365
transform 1 0 28112 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__A2
timestamp 1698431365
transform 1 0 30912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__A2
timestamp 1698431365
transform 1 0 30352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__A2
timestamp 1698431365
transform 1 0 31472 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1518__I
timestamp 1698431365
transform 1 0 32368 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__A1
timestamp 1698431365
transform 1 0 32144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__A2
timestamp 1698431365
transform 1 0 31696 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__A2
timestamp 1698431365
transform 1 0 32480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__A2
timestamp 1698431365
transform 1 0 35952 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1523__A2
timestamp 1698431365
transform 1 0 40992 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__A2
timestamp 1698431365
transform 1 0 44576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__A2
timestamp 1698431365
transform 1 0 41440 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__A2
timestamp 1698431365
transform 1 0 36736 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1528__A2
timestamp 1698431365
transform 1 0 36624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1530__A2
timestamp 1698431365
transform 1 0 39088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__A2
timestamp 1698431365
transform 1 0 42672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1532__A2
timestamp 1698431365
transform 1 0 44240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1533__A2
timestamp 1698431365
transform 1 0 44912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1534__A2
timestamp 1698431365
transform 1 0 39872 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1535__A2
timestamp 1698431365
transform 1 0 29232 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1537__I
timestamp 1698431365
transform 1 0 38416 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1538__A2
timestamp 1698431365
transform 1 0 29904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1540__A2
timestamp 1698431365
transform 1 0 30800 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1542__A2
timestamp 1698431365
transform 1 0 34048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1544__A2
timestamp 1698431365
transform 1 0 32032 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__A1
timestamp 1698431365
transform 1 0 30016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__A2
timestamp 1698431365
transform 1 0 31920 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1548__A2
timestamp 1698431365
transform 1 0 32592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1549__I
timestamp 1698431365
transform 1 0 28672 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1550__A2
timestamp 1698431365
transform 1 0 21952 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A2
timestamp 1698431365
transform 1 0 22848 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__A2
timestamp 1698431365
transform 1 0 24080 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1553__A2
timestamp 1698431365
transform 1 0 26208 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1554__A2
timestamp 1698431365
transform -1 0 28336 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__A2
timestamp 1698431365
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1557__A2
timestamp 1698431365
transform 1 0 35504 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1559__A2
timestamp 1698431365
transform 1 0 37856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1561__A2
timestamp 1698431365
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1563__A2
timestamp 1698431365
transform 1 0 37520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1565__A2
timestamp 1698431365
transform 1 0 35840 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__A1
timestamp 1698431365
transform 1 0 35056 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__A2
timestamp 1698431365
transform 1 0 36400 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1568__A2
timestamp 1698431365
transform 1 0 38304 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1569__A2
timestamp 1698431365
transform 1 0 41216 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1570__A2
timestamp 1698431365
transform 1 0 42784 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__A2
timestamp 1698431365
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1572__A2
timestamp 1698431365
transform 1 0 36288 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__A2
timestamp 1698431365
transform 1 0 37184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A2
timestamp 1698431365
transform 1 0 38192 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__A2
timestamp 1698431365
transform 1 0 41328 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1578__A2
timestamp 1698431365
transform 1 0 43344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__A2
timestamp 1698431365
transform 1 0 43456 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A1
timestamp 1698431365
transform -1 0 34608 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A2
timestamp 1698431365
transform 1 0 33488 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1581__A2
timestamp 1698431365
transform 1 0 36064 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1583__A2
timestamp 1698431365
transform 1 0 39648 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1585__A2
timestamp 1698431365
transform 1 0 39648 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1587__A2
timestamp 1698431365
transform 1 0 39200 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1589__A2
timestamp 1698431365
transform 1 0 33600 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1591__A2
timestamp 1698431365
transform 1 0 34944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1593__A2
timestamp 1698431365
transform 1 0 38864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1594__I
timestamp 1698431365
transform -1 0 37296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1595__A2
timestamp 1698431365
transform 1 0 38864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1596__A2
timestamp 1698431365
transform 1 0 39984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A2
timestamp 1698431365
transform 1 0 38528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__A2
timestamp 1698431365
transform 1 0 34608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__A2
timestamp 1698431365
transform 1 0 34384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1600__A3
timestamp 1698431365
transform -1 0 3584 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__A1
timestamp 1698431365
transform -1 0 12656 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__B
timestamp 1698431365
transform 1 0 13552 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__A1
timestamp 1698431365
transform 1 0 10976 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__B
timestamp 1698431365
transform 1 0 10640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A1
timestamp 1698431365
transform 1 0 8064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__A1
timestamp 1698431365
transform 1 0 10864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__B
timestamp 1698431365
transform -1 0 12208 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1608__A1
timestamp 1698431365
transform 1 0 11760 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1609__A1
timestamp 1698431365
transform 1 0 13552 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1609__B
timestamp 1698431365
transform 1 0 12768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A1
timestamp 1698431365
transform 1 0 10528 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__A1
timestamp 1698431365
transform 1 0 10640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__B
timestamp 1698431365
transform 1 0 12880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__B
timestamp 1698431365
transform -1 0 11424 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1614__A1
timestamp 1698431365
transform 1 0 8960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A1
timestamp 1698431365
transform 1 0 2240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1617__A1
timestamp 1698431365
transform 1 0 12096 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1617__A2
timestamp 1698431365
transform 1 0 13104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1618__B
timestamp 1698431365
transform -1 0 2016 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__A1
timestamp 1698431365
transform 1 0 10304 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__B
timestamp 1698431365
transform 1 0 6384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__B
timestamp 1698431365
transform 1 0 8848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1623__A1
timestamp 1698431365
transform 1 0 9632 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__B
timestamp 1698431365
transform 1 0 9856 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__A1
timestamp 1698431365
transform 1 0 11088 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__A1
timestamp 1698431365
transform -1 0 12096 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A1
timestamp 1698431365
transform 1 0 9296 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1629__A1
timestamp 1698431365
transform 1 0 12208 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__A1
timestamp 1698431365
transform 1 0 10976 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__A1
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A2
timestamp 1698431365
transform 1 0 2912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1633__A1
timestamp 1698431365
transform 1 0 3024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__A2
timestamp 1698431365
transform -1 0 2128 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1637__A1
timestamp 1698431365
transform 1 0 2128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__B
timestamp 1698431365
transform 1 0 4256 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1640__A1
timestamp 1698431365
transform 1 0 3920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__A1
timestamp 1698431365
transform 1 0 3024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A1
timestamp 1698431365
transform -1 0 2352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A1
timestamp 1698431365
transform 1 0 4592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__B
timestamp 1698431365
transform 1 0 4144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__A1
timestamp 1698431365
transform -1 0 3136 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__A1
timestamp 1698431365
transform -1 0 4480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__CLK
timestamp 1698431365
transform 1 0 12768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__CLK
timestamp 1698431365
transform -1 0 16464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__CLK
timestamp 1698431365
transform 1 0 16464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__CLK
timestamp 1698431365
transform 1 0 14000 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__CLK
timestamp 1698431365
transform 1 0 17024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__CLK
timestamp 1698431365
transform 1 0 15344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__CLK
timestamp 1698431365
transform 1 0 18144 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__CLK
timestamp 1698431365
transform 1 0 19600 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__CLK
timestamp 1698431365
transform 1 0 19264 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__CLK
timestamp 1698431365
transform 1 0 34608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__CLK
timestamp 1698431365
transform 1 0 38640 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__CLK
timestamp 1698431365
transform -1 0 37632 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__CLK
timestamp 1698431365
transform 1 0 39536 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__CLK
timestamp 1698431365
transform 1 0 40096 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__CLK
timestamp 1698431365
transform 1 0 40992 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__CLK
timestamp 1698431365
transform 1 0 33600 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__CLK
timestamp 1698431365
transform 1 0 32704 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__CLK
timestamp 1698431365
transform 1 0 33600 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__CLK
timestamp 1698431365
transform 1 0 37968 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__CLK
timestamp 1698431365
transform 1 0 33824 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__CLK
timestamp 1698431365
transform 1 0 25536 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1671__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__CLK
timestamp 1698431365
transform 1 0 15456 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__CLK
timestamp 1698431365
transform 1 0 16128 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__CLK
timestamp 1698431365
transform 1 0 16800 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__CLK
timestamp 1698431365
transform 1 0 17024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__CLK
timestamp 1698431365
transform 1 0 16352 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__CLK
timestamp 1698431365
transform 1 0 14784 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__CLK
timestamp 1698431365
transform 1 0 17920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__CLK
timestamp 1698431365
transform -1 0 19152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__CLK
timestamp 1698431365
transform 1 0 20944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__CLK
timestamp 1698431365
transform 1 0 21952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__CLK
timestamp 1698431365
transform 1 0 17472 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__CLK
timestamp 1698431365
transform 1 0 18144 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__CLK
timestamp 1698431365
transform -1 0 21616 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__CLK
timestamp 1698431365
transform 1 0 24192 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__CLK
timestamp 1698431365
transform 1 0 26768 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__CLK
timestamp 1698431365
transform 1 0 33712 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__CLK
timestamp 1698431365
transform 1 0 34608 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__CLK
timestamp 1698431365
transform 1 0 35280 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__CLK
timestamp 1698431365
transform 1 0 29232 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__CLK
timestamp 1698431365
transform 1 0 26880 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__CLK
timestamp 1698431365
transform 1 0 32928 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__CLK
timestamp 1698431365
transform 1 0 31472 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__CLK
timestamp 1698431365
transform 1 0 31696 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__CLK
timestamp 1698431365
transform -1 0 33824 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__CLK
timestamp 1698431365
transform 1 0 24080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__CLK
timestamp 1698431365
transform 1 0 22624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__CLK
timestamp 1698431365
transform 1 0 20384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1705__CLK
timestamp 1698431365
transform 1 0 21392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__CLK
timestamp 1698431365
transform 1 0 25536 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__CLK
timestamp 1698431365
transform 1 0 23408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__CLK
timestamp 1698431365
transform 1 0 25088 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__CLK
timestamp 1698431365
transform 1 0 18704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__CLK
timestamp 1698431365
transform 1 0 19376 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__CLK
timestamp 1698431365
transform 1 0 20944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__CLK
timestamp 1698431365
transform -1 0 23968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1714__CLK
timestamp 1698431365
transform 1 0 15232 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__CLK
timestamp 1698431365
transform 1 0 17360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__CLK
timestamp 1698431365
transform 1 0 17808 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1717__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__CLK
timestamp 1698431365
transform 1 0 18704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__CLK
timestamp 1698431365
transform 1 0 21392 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__CLK
timestamp 1698431365
transform 1 0 15120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__CLK
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__CLK
timestamp 1698431365
transform 1 0 14672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__CLK
timestamp 1698431365
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__CLK
timestamp 1698431365
transform 1 0 22400 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__CLK
timestamp 1698431365
transform 1 0 18032 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__CLK
timestamp 1698431365
transform 1 0 17472 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__CLK
timestamp 1698431365
transform 1 0 20608 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1729__CLK
timestamp 1698431365
transform 1 0 22624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__CLK
timestamp 1698431365
transform 1 0 24864 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__CLK
timestamp 1698431365
transform 1 0 16352 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__CLK
timestamp 1698431365
transform 1 0 20272 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__CLK
timestamp 1698431365
transform 1 0 22400 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__CLK
timestamp 1698431365
transform 1 0 24080 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__CLK
timestamp 1698431365
transform 1 0 25984 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__CLK
timestamp 1698431365
transform 1 0 18256 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__CLK
timestamp 1698431365
transform 1 0 18816 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__CLK
timestamp 1698431365
transform 1 0 15904 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__CLK
timestamp 1698431365
transform 1 0 19488 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__CLK
timestamp 1698431365
transform 1 0 22512 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1744__CLK
timestamp 1698431365
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__CLK
timestamp 1698431365
transform 1 0 39648 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__CLK
timestamp 1698431365
transform 1 0 42784 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__CLK
timestamp 1698431365
transform 1 0 44240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__CLK
timestamp 1698431365
transform 1 0 41328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__CLK
timestamp 1698431365
transform 1 0 43008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__CLK
timestamp 1698431365
transform 1 0 42000 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__CLK
timestamp 1698431365
transform 1 0 40544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__CLK
timestamp 1698431365
transform 1 0 38976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__CLK
timestamp 1698431365
transform 1 0 21392 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__CLK
timestamp 1698431365
transform -1 0 16352 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1757__CLK
timestamp 1698431365
transform 1 0 14000 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__CLK
timestamp 1698431365
transform 1 0 15680 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__CLK
timestamp 1698431365
transform 1 0 17808 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__CLK
timestamp 1698431365
transform 1 0 20720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__CLK
timestamp 1698431365
transform 1 0 41216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__CLK
timestamp 1698431365
transform 1 0 44912 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__CLK
timestamp 1698431365
transform 1 0 44912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__CLK
timestamp 1698431365
transform 1 0 38080 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__CLK
timestamp 1698431365
transform 1 0 36624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__CLK
timestamp 1698431365
transform 1 0 35056 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__CLK
timestamp 1698431365
transform 1 0 33824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__CLK
timestamp 1698431365
transform 1 0 35616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__CLK
timestamp 1698431365
transform -1 0 36848 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__CLK
timestamp 1698431365
transform 1 0 36176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1773__CLK
timestamp 1698431365
transform 1 0 32704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__CLK
timestamp 1698431365
transform 1 0 17024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__CLK
timestamp 1698431365
transform 1 0 16464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__CLK
timestamp 1698431365
transform 1 0 18256 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1777__CLK
timestamp 1698431365
transform 1 0 19152 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__CLK
timestamp 1698431365
transform 1 0 22624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__CLK
timestamp 1698431365
transform 1 0 24864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__CLK
timestamp 1698431365
transform 1 0 25984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__CLK
timestamp 1698431365
transform 1 0 26768 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__CLK
timestamp 1698431365
transform 1 0 33040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1784__CLK
timestamp 1698431365
transform 1 0 31136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__CLK
timestamp 1698431365
transform 1 0 33936 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1786__CLK
timestamp 1698431365
transform 1 0 34272 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__CLK
timestamp 1698431365
transform -1 0 41440 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__CLK
timestamp 1698431365
transform -1 0 40992 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__CLK
timestamp 1698431365
transform 1 0 43232 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__CLK
timestamp 1698431365
transform 1 0 38080 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__CLK
timestamp 1698431365
transform -1 0 38192 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__CLK
timestamp 1698431365
transform 1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__CLK
timestamp 1698431365
transform 1 0 38864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__CLK
timestamp 1698431365
transform 1 0 42000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__CLK
timestamp 1698431365
transform 1 0 44240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__CLK
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__CLK
timestamp 1698431365
transform 1 0 38192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__CLK
timestamp 1698431365
transform 1 0 26544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__CLK
timestamp 1698431365
transform 1 0 26656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__CLK
timestamp 1698431365
transform 1 0 31136 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__CLK
timestamp 1698431365
transform 1 0 33376 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__CLK
timestamp 1698431365
transform 1 0 25312 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__CLK
timestamp 1698431365
transform 1 0 17584 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__CLK
timestamp 1698431365
transform 1 0 20720 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__CLK
timestamp 1698431365
transform 1 0 21392 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__CLK
timestamp 1698431365
transform -1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__CLK
timestamp 1698431365
transform 1 0 26656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__CLK
timestamp 1698431365
transform 1 0 31584 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__CLK
timestamp 1698431365
transform 1 0 33152 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__CLK
timestamp 1698431365
transform 1 0 35616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__CLK
timestamp 1698431365
transform 1 0 36624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__CLK
timestamp 1698431365
transform 1 0 34272 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__CLK
timestamp 1698431365
transform 1 0 34048 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__CLK
timestamp 1698431365
transform 1 0 38864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__CLK
timestamp 1698431365
transform 1 0 42784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__CLK
timestamp 1698431365
transform 1 0 42336 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__CLK
timestamp 1698431365
transform 1 0 39872 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__CLK
timestamp 1698431365
transform 1 0 37632 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__CLK
timestamp 1698431365
transform 1 0 40096 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__CLK
timestamp 1698431365
transform 1 0 42560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__CLK
timestamp 1698431365
transform 1 0 42000 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__CLK
timestamp 1698431365
transform 1 0 43568 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__CLK
timestamp 1698431365
transform 1 0 42896 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__CLK
timestamp 1698431365
transform 1 0 32256 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__CLK
timestamp 1698431365
transform 1 0 34608 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__CLK
timestamp 1698431365
transform 1 0 35728 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__CLK
timestamp 1698431365
transform 1 0 36400 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__CLK
timestamp 1698431365
transform 1 0 35952 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1832__CLK
timestamp 1698431365
transform -1 0 34384 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__CLK
timestamp 1698431365
transform 1 0 32368 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__CLK
timestamp 1698431365
transform -1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1835__CLK
timestamp 1698431365
transform 1 0 38304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__CLK
timestamp 1698431365
transform 1 0 37296 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__CLK
timestamp 1698431365
transform 1 0 33376 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__CLK
timestamp 1698431365
transform 1 0 33152 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__CLK
timestamp 1698431365
transform 1 0 13664 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__CLK
timestamp 1698431365
transform 1 0 8512 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__CLK
timestamp 1698431365
transform 1 0 13552 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__CLK
timestamp 1698431365
transform 1 0 11648 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__CLK
timestamp 1698431365
transform 1 0 11424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__CLK
timestamp 1698431365
transform 1 0 8176 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__CLK
timestamp 1698431365
transform 1 0 5040 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__CLK
timestamp 1698431365
transform 1 0 14448 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__CLK
timestamp 1698431365
transform 1 0 5264 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1849__CLK
timestamp 1698431365
transform 1 0 9856 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1850__CLK
timestamp 1698431365
transform 1 0 10304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__CLK
timestamp 1698431365
transform 1 0 11424 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__CLK
timestamp 1698431365
transform 1 0 12656 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__CLK
timestamp 1698431365
transform 1 0 13776 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__CLK
timestamp 1698431365
transform 1 0 11312 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__CLK
timestamp 1698431365
transform 1 0 5712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__CLK
timestamp 1698431365
transform 1 0 4816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1857__CLK
timestamp 1698431365
transform 1 0 4816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__CLK
timestamp 1698431365
transform 1 0 5040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__CLK
timestamp 1698431365
transform 1 0 5040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__CLK
timestamp 1698431365
transform -1 0 6944 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_io_in[0]_I
timestamp 1698431365
transform 1 0 6160 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_0__f_io_in[0]_I
timestamp 1698431365
transform 1 0 9296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_1__f_io_in[0]_I
timestamp 1698431365
transform 1 0 13552 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._060__I
timestamp 1698431365
transform -1 0 5712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._061__I
timestamp 1698431365
transform -1 0 5488 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._063__B
timestamp 1698431365
transform 1 0 15232 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._066__A1
timestamp 1698431365
transform 1 0 13552 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._070__A1
timestamp 1698431365
transform 1 0 14112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._071__I
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._072__A1
timestamp 1698431365
transform -1 0 9632 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._074__A1
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._078__A1
timestamp 1698431365
transform 1 0 10752 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._080__B
timestamp 1698431365
transform 1 0 12768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._084__A1
timestamp 1698431365
transform 1 0 10640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._085__A1
timestamp 1698431365
transform 1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._086__B
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._087__I
timestamp 1698431365
transform -1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._090__A1
timestamp 1698431365
transform -1 0 15232 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._093__A1
timestamp 1698431365
transform 1 0 9632 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._094__C
timestamp 1698431365
transform 1 0 16016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._101__A1
timestamp 1698431365
transform 1 0 6720 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._108__I
timestamp 1698431365
transform -1 0 8064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._114__A1
timestamp 1698431365
transform 1 0 6832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._118__A1
timestamp 1698431365
transform 1 0 9296 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_dec1._123__B2
timestamp 1698431365
transform 1 0 7728 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout8_I
timestamp 1698431365
transform -1 0 17696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout9_I
timestamp 1698431365
transform 1 0 13776 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout10_I
timestamp 1698431365
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout11_I
timestamp 1698431365
transform 1 0 14784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout12_I
timestamp 1698431365
transform 1 0 30912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout13_I
timestamp 1698431365
transform 1 0 14000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout14_I
timestamp 1698431365
transform 1 0 40320 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout15_I
timestamp 1698431365
transform 1 0 12880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout16_I
timestamp 1698431365
transform -1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout17_I
timestamp 1698431365
transform 1 0 30688 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout18_I
timestamp 1698431365
transform -1 0 15232 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 1792 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 1792 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 1792 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 1792 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 2464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 1792 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 2128 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac._4__I
timestamp 1698431365
transform 1 0 4704 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac._5__A2
timestamp 1698431365
transform 1 0 4032 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._3__I
timestamp 1698431365
transform -1 0 5488 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._4__A1
timestamp 1698431365
transform -1 0 2016 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._4__A2
timestamp 1698431365
transform 1 0 4144 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._5__A1
timestamp 1698431365
transform 1 0 2576 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 2128 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 4592 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._4__A2
timestamp 1698431365
transform 1 0 5040 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._5__A1
timestamp 1698431365
transform 1 0 4032 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 4928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 5264 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref_I
timestamp 1698431365
transform 1 0 4480 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._4__A2
timestamp 1698431365
transform 1 0 7168 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._5__A1
timestamp 1698431365
transform 1 0 5824 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 5040 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 7952 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref_I
timestamp 1698431365
transform 1 0 9632 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref_I
timestamp 1698431365
transform 1 0 4592 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref_I
timestamp 1698431365
transform 1 0 6384 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._3__I
timestamp 1698431365
transform -1 0 6160 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._4__A1
timestamp 1698431365
transform 1 0 7616 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._4__A2
timestamp 1698431365
transform 1 0 7168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._5__A1
timestamp 1698431365
transform 1 0 4592 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 6160 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 6608 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref_I
timestamp 1698431365
transform 1 0 5712 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref_I
timestamp 1698431365
transform 1 0 5824 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref_I
timestamp 1698431365
transform 1 0 5040 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref_I
timestamp 1698431365
transform 1 0 5488 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref_I
timestamp 1698431365
transform 1 0 6160 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref_I
timestamp 1698431365
transform 1 0 6608 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref_I
timestamp 1698431365
transform 1 0 5040 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._3__I
timestamp 1698431365
transform 1 0 8960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._4__A1
timestamp 1698431365
transform 1 0 8176 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._4__A2
timestamp 1698431365
transform 1 0 7728 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._5__A1
timestamp 1698431365
transform 1 0 7280 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch._7__I
timestamp 1698431365
transform 1 0 6496 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 10304 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref_I
timestamp 1698431365
transform 1 0 8960 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref_I
timestamp 1698431365
transform 1 0 8960 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref_I
timestamp 1698431365
transform 1 0 12656 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref_I
timestamp 1698431365
transform 1 0 10080 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref_I
timestamp 1698431365
transform 1 0 11984 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref_I
timestamp 1698431365
transform 1 0 9520 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref_I
timestamp 1698431365
transform 1 0 10304 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref_I
timestamp 1698431365
transform 1 0 8960 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref_I
timestamp 1698431365
transform 1 0 8288 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref_I
timestamp 1698431365
transform 1 0 7280 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref_I
timestamp 1698431365
transform 1 0 10192 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref_I
timestamp 1698431365
transform 1 0 10304 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref_I
timestamp 1698431365
transform 1 0 11760 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref_I
timestamp 1698431365
transform 1 0 9408 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref_I
timestamp 1698431365
transform 1 0 8736 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dac.vdac_single.einvp_batch\[0\].vref_I
timestamp 1698431365
transform 1 0 6048 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_temp1.dcdc_EN
timestamp 1698431365
transform 1 0 1904 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0__0316_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3136 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0__0318_
timestamp 1698431365
transform 1 0 10416 0 -1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_io_in[0]
timestamp 1698431365
transform 1 0 6832 0 1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_net23
timestamp 1698431365
transform 1 0 3360 0 -1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_temp1.i_precharge_n
timestamp 1698431365
transform 1 0 3472 0 -1 54880
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f__0316_
timestamp 1698431365
transform -1 0 9184 0 -1 39200
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f__0318_
timestamp 1698431365
transform -1 0 15680 0 -1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_io_in[0]
timestamp 1698431365
transform -1 0 9184 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_net23
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_temp1.i_precharge_n
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f__0316_
timestamp 1698431365
transform -1 0 7280 0 -1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f__0318_
timestamp 1698431365
transform -1 0 17024 0 -1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_io_in[0]
timestamp 1698431365
transform -1 0 13104 0 1 39200
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_net23
timestamp 1698431365
transform -1 0 8624 0 -1 48608
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_temp1.i_precharge_n
timestamp 1698431365
transform -1 0 7728 0 -1 56448
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._060_
timestamp 1698431365
transform 1 0 5712 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  dec1._061_
timestamp 1698431365
transform 1 0 4816 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  dec1._062_
timestamp 1698431365
transform 1 0 5824 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  dec1._063_
timestamp 1698431365
transform 1 0 11312 0 -1 17248
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  dec1._064_
timestamp 1698431365
transform -1 0 12544 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  dec1._065_
timestamp 1698431365
transform 1 0 12432 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  dec1._066_
timestamp 1698431365
transform -1 0 12768 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  dec1._067_
timestamp 1698431365
transform 1 0 12768 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  dec1._068_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11088 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._069_
timestamp 1698431365
transform 1 0 13328 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  dec1._070_
timestamp 1698431365
transform 1 0 12208 0 -1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_3  dec1._071_
timestamp 1698431365
transform 1 0 10528 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  dec1._072_
timestamp 1698431365
transform 1 0 11088 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  dec1._073_
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  dec1._074_
timestamp 1698431365
transform 1 0 12096 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  dec1._075_
timestamp 1698431365
transform -1 0 14336 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  dec1._076_
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  dec1._077_
timestamp 1698431365
transform -1 0 14112 0 -1 10976
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  dec1._078_
timestamp 1698431365
transform -1 0 10752 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  dec1._079_
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  dec1._080_
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  dec1._081_
timestamp 1698431365
transform 1 0 9408 0 1 14112
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  dec1._082_
timestamp 1698431365
transform 1 0 10640 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  dec1._083_
timestamp 1698431365
transform -1 0 12432 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  dec1._084_
timestamp 1698431365
transform 1 0 10976 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  dec1._085_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  dec1._086_
timestamp 1698431365
transform 1 0 9744 0 1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._087_
timestamp 1698431365
transform -1 0 12880 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  dec1._088_
timestamp 1698431365
transform -1 0 12992 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  dec1._089_
timestamp 1698431365
transform 1 0 10864 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  dec1._090_
timestamp 1698431365
transform 1 0 14224 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  dec1._091_
timestamp 1698431365
transform -1 0 14336 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  dec1._092_
timestamp 1698431365
transform 1 0 11088 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  dec1._093_
timestamp 1698431365
transform -1 0 9184 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  dec1._094_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11088 0 -1 7840
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  dec1._095_
timestamp 1698431365
transform -1 0 15232 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  dec1._096_
timestamp 1698431365
transform -1 0 11088 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  dec1._097_
timestamp 1698431365
transform 1 0 9744 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  dec1._098_
timestamp 1698431365
transform 1 0 10640 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  dec1._099_
timestamp 1698431365
transform -1 0 13328 0 -1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  dec1._100_
timestamp 1698431365
transform -1 0 11088 0 1 3136
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  dec1._101_
timestamp 1698431365
transform 1 0 6944 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  dec1._102_
timestamp 1698431365
transform 1 0 6160 0 -1 9408
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  dec1._103_
timestamp 1698431365
transform 1 0 10080 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  dec1._104_
timestamp 1698431365
transform -1 0 10080 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  dec1._105_
timestamp 1698431365
transform -1 0 9856 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  dec1._106_
timestamp 1698431365
transform 1 0 9744 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  dec1._107_
timestamp 1698431365
transform 1 0 8064 0 1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  dec1._108_
timestamp 1698431365
transform 1 0 8064 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  dec1._109_
timestamp 1698431365
transform -1 0 9744 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  dec1._110_
timestamp 1698431365
transform -1 0 10640 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  dec1._111_
timestamp 1698431365
transform -1 0 11088 0 -1 3136
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  dec1._112_
timestamp 1698431365
transform 1 0 5824 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  dec1._113_
timestamp 1698431365
transform -1 0 11424 0 1 4704
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  dec1._114_
timestamp 1698431365
transform 1 0 6496 0 -1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  dec1._115_
timestamp 1698431365
transform -1 0 9072 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  dec1._116_
timestamp 1698431365
transform 1 0 6272 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  dec1._117_
timestamp 1698431365
transform -1 0 8848 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  dec1._118_
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  dec1._119_
timestamp 1698431365
transform 1 0 7616 0 1 7840
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  dec1._120_
timestamp 1698431365
transform -1 0 8176 0 -1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  dec1._121_
timestamp 1698431365
transform -1 0 7952 0 -1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  dec1._122_
timestamp 1698431365
transform 1 0 6496 0 1 3136
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  dec1._123_
timestamp 1698431365
transform 1 0 7952 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout8
timestamp 1698431365
transform 1 0 14896 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  fanout9 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 14000 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout10
timestamp 1698431365
transform 1 0 29792 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout11
timestamp 1698431365
transform -1 0 14784 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout12
timestamp 1698431365
transform 1 0 31136 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  fanout13
timestamp 1698431365
transform 1 0 14224 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout14
timestamp 1698431365
transform 1 0 37632 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout15
timestamp 1698431365
transform 1 0 14112 0 -1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout16
timestamp 1698431365
transform -1 0 16576 0 -1 59584
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  fanout17
timestamp 1698431365
transform 1 0 30912 0 1 59584
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  fanout18
timestamp 1698431365
transform 1 0 15232 0 -1 61152
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 1568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_36 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 1568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_44 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6272 0 1 1568
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_50 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6944 0 1 1568
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_66 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8736 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 1568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 1568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 1568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 1568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 1568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 1568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 1568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 1568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 1568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 1568
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 1568
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_418
timestamp 1698431365
transform 1 0 48160 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_10
timestamp 1698431365
transform 1 0 2464 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_14
timestamp 1698431365
transform 1 0 2912 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_16 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3136 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_48
timestamp 1698431365
transform 1 0 6720 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_59
timestamp 1698431365
transform 1 0 7952 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_67
timestamp 1698431365
transform 1 0 8848 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_69
timestamp 1698431365
transform 1 0 9072 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_87
timestamp 1698431365
transform 1 0 11088 0 -1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_119
timestamp 1698431365
transform 1 0 14672 0 -1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_135
timestamp 1698431365
transform 1 0 16464 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_150
timestamp 1698431365
transform 1 0 18144 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_153
timestamp 1698431365
transform 1 0 18480 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_157
timestamp 1698431365
transform 1 0 18928 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_190
timestamp 1698431365
transform 1 0 22624 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_202
timestamp 1698431365
transform 1 0 23968 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_224
timestamp 1698431365
transform 1 0 26432 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_226
timestamp 1698431365
transform 1 0 26656 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_264
timestamp 1698431365
transform 1 0 30912 0 -1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_314
timestamp 1698431365
transform 1 0 36512 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_317
timestamp 1698431365
transform 1 0 36848 0 -1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_352 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 3136
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698431365
transform 1 0 47936 0 -1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_31
timestamp 1698431365
transform 1 0 4816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_45
timestamp 1698431365
transform 1 0 6384 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_56
timestamp 1698431365
transform 1 0 7616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_121
timestamp 1698431365
transform 1 0 14896 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_151
timestamp 1698431365
transform 1 0 18256 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_153
timestamp 1698431365
transform 1 0 18480 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_170
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_174
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_185
timestamp 1698431365
transform 1 0 22064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_189
timestamp 1698431365
transform 1 0 22512 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_221
timestamp 1698431365
transform 1 0 26096 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_244
timestamp 1698431365
transform 1 0 28672 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_251
timestamp 1698431365
transform 1 0 29456 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_281
timestamp 1698431365
transform 1 0 32816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_293
timestamp 1698431365
transform 1 0 34160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_297
timestamp 1698431365
transform 1 0 34608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_301
timestamp 1698431365
transform 1 0 35056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_309
timestamp 1698431365
transform 1 0 35952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_313
timestamp 1698431365
transform 1 0 36400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_346
timestamp 1698431365
transform 1 0 40096 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_378
timestamp 1698431365
transform 1 0 43680 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_382
timestamp 1698431365
transform 1 0 44128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_384
timestamp 1698431365
transform 1 0 44352 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_419
timestamp 1698431365
transform 1 0 48272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_34
timestamp 1698431365
transform 1 0 5152 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_42
timestamp 1698431365
transform 1 0 6048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_76
timestamp 1698431365
transform 1 0 9856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_103
timestamp 1698431365
transform 1 0 12880 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_171
timestamp 1698431365
transform 1 0 20496 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_187
timestamp 1698431365
transform 1 0 22288 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_195
timestamp 1698431365
transform 1 0 23184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_203
timestamp 1698431365
transform 1 0 24080 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_249
timestamp 1698431365
transform 1 0 29232 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_253
timestamp 1698431365
transform 1 0 29680 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_262
timestamp 1698431365
transform 1 0 30688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_266
timestamp 1698431365
transform 1 0 31136 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_340
timestamp 1698431365
transform 1 0 39424 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_348
timestamp 1698431365
transform 1 0 40320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698431365
transform 1 0 47936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_31
timestamp 1698431365
transform 1 0 4816 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_39
timestamp 1698431365
transform 1 0 5712 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_90
timestamp 1698431365
transform 1 0 11424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_92
timestamp 1698431365
transform 1 0 11648 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_104
timestamp 1698431365
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_122
timestamp 1698431365
transform 1 0 15008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_124
timestamp 1698431365
transform 1 0 15232 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_133
timestamp 1698431365
transform 1 0 16240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_137
timestamp 1698431365
transform 1 0 16688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_139
timestamp 1698431365
transform 1 0 16912 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_142
timestamp 1698431365
transform 1 0 17248 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_167
timestamp 1698431365
transform 1 0 20048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_169
timestamp 1698431365
transform 1 0 20272 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_174
timestamp 1698431365
transform 1 0 20832 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_181
timestamp 1698431365
transform 1 0 21616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_198
timestamp 1698431365
transform 1 0 23520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_202
timestamp 1698431365
transform 1 0 23968 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_212
timestamp 1698431365
transform 1 0 25088 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_222
timestamp 1698431365
transform 1 0 26208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_226
timestamp 1698431365
transform 1 0 26656 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_234
timestamp 1698431365
transform 1 0 27552 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_238
timestamp 1698431365
transform 1 0 28000 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_279
timestamp 1698431365
transform 1 0 32592 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_282
timestamp 1698431365
transform 1 0 32928 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_296
timestamp 1698431365
transform 1 0 34496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_300
timestamp 1698431365
transform 1 0 34944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_310
timestamp 1698431365
transform 1 0 36064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_312
timestamp 1698431365
transform 1 0 36288 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_333
timestamp 1698431365
transform 1 0 38640 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_365
timestamp 1698431365
transform 1 0 42224 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_419
timestamp 1698431365
transform 1 0 48272 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_6
timestamp 1698431365
transform 1 0 2016 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_9
timestamp 1698431365
transform 1 0 2352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_13
timestamp 1698431365
transform 1 0 2800 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_16
timestamp 1698431365
transform 1 0 3136 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_24
timestamp 1698431365
transform 1 0 4032 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_28
timestamp 1698431365
transform 1 0 4480 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_32
timestamp 1698431365
transform 1 0 4928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_34
timestamp 1698431365
transform 1 0 5152 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_37
timestamp 1698431365
transform 1 0 5488 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_53
timestamp 1698431365
transform 1 0 7280 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 9072 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_74
timestamp 1698431365
transform 1 0 9632 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_124
timestamp 1698431365
transform 1 0 15232 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_128
timestamp 1698431365
transform 1 0 15680 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_169
timestamp 1698431365
transform 1 0 20272 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_171
timestamp 1698431365
transform 1 0 20496 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_201
timestamp 1698431365
transform 1 0 23856 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_233
timestamp 1698431365
transform 1 0 27440 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_237
timestamp 1698431365
transform 1 0 27888 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_253
timestamp 1698431365
transform 1 0 29680 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_257
timestamp 1698431365
transform 1 0 30128 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_269
timestamp 1698431365
transform 1 0 31472 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_277
timestamp 1698431365
transform 1 0 32368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_298
timestamp 1698431365
transform 1 0 34720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_302
timestamp 1698431365
transform 1 0 35168 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_334
timestamp 1698431365
transform 1 0 38752 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1698431365
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_19
timestamp 1698431365
transform 1 0 3472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_30
timestamp 1698431365
transform 1 0 4704 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_39
timestamp 1698431365
transform 1 0 5712 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_56
timestamp 1698431365
transform 1 0 7616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_66
timestamp 1698431365
transform 1 0 8736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_68
timestamp 1698431365
transform 1 0 8960 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_99
timestamp 1698431365
transform 1 0 12432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_103
timestamp 1698431365
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_120
timestamp 1698431365
transform 1 0 14784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_124
timestamp 1698431365
transform 1 0 15232 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_140
timestamp 1698431365
transform 1 0 17024 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_148
timestamp 1698431365
transform 1 0 17920 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_152
timestamp 1698431365
transform 1 0 18368 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_156
timestamp 1698431365
transform 1 0 18816 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_160
timestamp 1698431365
transform 1 0 19264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_164
timestamp 1698431365
transform 1 0 19712 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_168
timestamp 1698431365
transform 1 0 20160 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_181
timestamp 1698431365
transform 1 0 21616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_189
timestamp 1698431365
transform 1 0 22512 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_221
timestamp 1698431365
transform 1 0 26096 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_225
timestamp 1698431365
transform 1 0 26544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_235
timestamp 1698431365
transform 1 0 27664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_239
timestamp 1698431365
transform 1 0 28112 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_243
timestamp 1698431365
transform 1 0 28560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_265
timestamp 1698431365
transform 1 0 31024 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_297
timestamp 1698431365
transform 1 0 34608 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_313
timestamp 1698431365
transform 1 0 36400 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_419
timestamp 1698431365
transform 1 0 48272 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_8
timestamp 1698431365
transform 1 0 2240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_67
timestamp 1698431365
transform 1 0 8848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_78
timestamp 1698431365
transform 1 0 10080 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_129
timestamp 1698431365
transform 1 0 15792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_133
timestamp 1698431365
transform 1 0 16240 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_137
timestamp 1698431365
transform 1 0 16688 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_146
timestamp 1698431365
transform 1 0 17696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_150
timestamp 1698431365
transform 1 0 18144 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_158
timestamp 1698431365
transform 1 0 19040 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_160
timestamp 1698431365
transform 1 0 19264 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_192
timestamp 1698431365
transform 1 0 22848 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_208
timestamp 1698431365
transform 1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_286
timestamp 1698431365
transform 1 0 33376 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_302
timestamp 1698431365
transform 1 0 35168 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_337
timestamp 1698431365
transform 1 0 39088 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_345
timestamp 1698431365
transform 1 0 39984 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_349
timestamp 1698431365
transform 1 0 40432 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698431365
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_47
timestamp 1698431365
transform 1 0 6608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_49
timestamp 1698431365
transform 1 0 6832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_55
timestamp 1698431365
transform 1 0 7504 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_99
timestamp 1698431365
transform 1 0 12432 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_111
timestamp 1698431365
transform 1 0 13776 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_143
timestamp 1698431365
transform 1 0 17360 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_153
timestamp 1698431365
transform 1 0 18480 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_157
timestamp 1698431365
transform 1 0 18928 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_173
timestamp 1698431365
transform 1 0 20720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_181
timestamp 1698431365
transform 1 0 21616 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_221
timestamp 1698431365
transform 1 0 26096 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_235
timestamp 1698431365
transform 1 0 27664 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_243
timestamp 1698431365
transform 1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_263
timestamp 1698431365
transform 1 0 30800 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_265
timestamp 1698431365
transform 1 0 31024 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_297
timestamp 1698431365
transform 1 0 34608 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_305
timestamp 1698431365
transform 1 0 35504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_357
timestamp 1698431365
transform 1 0 41328 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_373
timestamp 1698431365
transform 1 0 43120 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_381
timestamp 1698431365
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_419
timestamp 1698431365
transform 1 0 48272 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_23
timestamp 1698431365
transform 1 0 3920 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_27
timestamp 1698431365
transform 1 0 4368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_31
timestamp 1698431365
transform 1 0 4816 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_35
timestamp 1698431365
transform 1 0 5264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_130
timestamp 1698431365
transform 1 0 15904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_171
timestamp 1698431365
transform 1 0 20496 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_179
timestamp 1698431365
transform 1 0 21392 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_187
timestamp 1698431365
transform 1 0 22288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_189
timestamp 1698431365
transform 1 0 22512 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_192
timestamp 1698431365
transform 1 0 22848 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_200
timestamp 1698431365
transform 1 0 23744 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_207
timestamp 1698431365
transform 1 0 24528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_220
timestamp 1698431365
transform 1 0 25984 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_224
timestamp 1698431365
transform 1 0 26432 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_234
timestamp 1698431365
transform 1 0 27552 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_238
timestamp 1698431365
transform 1 0 28000 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_242
timestamp 1698431365
transform 1 0 28448 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_252
timestamp 1698431365
transform 1 0 29568 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_258
timestamp 1698431365
transform 1 0 30240 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_262
timestamp 1698431365
transform 1 0 30688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_266
timestamp 1698431365
transform 1 0 31136 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_268
timestamp 1698431365
transform 1 0 31360 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_284
timestamp 1698431365
transform 1 0 33152 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_314
timestamp 1698431365
transform 1 0 36512 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_356
timestamp 1698431365
transform 1 0 41216 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_6
timestamp 1698431365
transform 1 0 2016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_13
timestamp 1698431365
transform 1 0 2800 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_17
timestamp 1698431365
transform 1 0 3248 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_33
timestamp 1698431365
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_47
timestamp 1698431365
transform 1 0 6608 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_50
timestamp 1698431365
transform 1 0 6944 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_66
timestamp 1698431365
transform 1 0 8736 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_70
timestamp 1698431365
transform 1 0 9184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_84
timestamp 1698431365
transform 1 0 10752 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_86
timestamp 1698431365
transform 1 0 10976 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_102
timestamp 1698431365
transform 1 0 12768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_133
timestamp 1698431365
transform 1 0 16240 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_137
timestamp 1698431365
transform 1 0 16688 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_140
timestamp 1698431365
transform 1 0 17024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_144
timestamp 1698431365
transform 1 0 17472 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_146
timestamp 1698431365
transform 1 0 17696 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_153
timestamp 1698431365
transform 1 0 18480 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_169
timestamp 1698431365
transform 1 0 20272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_185
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_193
timestamp 1698431365
transform 1 0 22960 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_197
timestamp 1698431365
transform 1 0 23408 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_208
timestamp 1698431365
transform 1 0 24640 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_240
timestamp 1698431365
transform 1 0 28224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_242
timestamp 1698431365
transform 1 0 28448 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_256
timestamp 1698431365
transform 1 0 30016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_258
timestamp 1698431365
transform 1 0 30240 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_273
timestamp 1698431365
transform 1 0 31920 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_281
timestamp 1698431365
transform 1 0 32816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_283
timestamp 1698431365
transform 1 0 33040 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_288
timestamp 1698431365
transform 1 0 33600 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_292
timestamp 1698431365
transform 1 0 34048 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_308
timestamp 1698431365
transform 1 0 35840 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_312
timestamp 1698431365
transform 1 0 36288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_314
timestamp 1698431365
transform 1 0 36512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_419
timestamp 1698431365
transform 1 0 48272 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_4
timestamp 1698431365
transform 1 0 1792 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_21
timestamp 1698431365
transform 1 0 3696 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_25
timestamp 1698431365
transform 1 0 4144 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_33
timestamp 1698431365
transform 1 0 5040 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_37
timestamp 1698431365
transform 1 0 5488 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_39
timestamp 1698431365
transform 1 0 5712 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_44
timestamp 1698431365
transform 1 0 6272 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_60
timestamp 1698431365
transform 1 0 8064 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_68
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_162
timestamp 1698431365
transform 1 0 19488 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_170
timestamp 1698431365
transform 1 0 20384 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_174
timestamp 1698431365
transform 1 0 20832 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_177
timestamp 1698431365
transform 1 0 21168 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_244
timestamp 1698431365
transform 1 0 28672 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_252
timestamp 1698431365
transform 1 0 29568 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_256
timestamp 1698431365
transform 1 0 30016 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_259
timestamp 1698431365
transform 1 0 30352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_263
timestamp 1698431365
transform 1 0 30800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_265
timestamp 1698431365
transform 1 0 31024 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_268
timestamp 1698431365
transform 1 0 31360 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_272
timestamp 1698431365
transform 1 0 31808 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_275
timestamp 1698431365
transform 1 0 32144 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_290
timestamp 1698431365
transform 1 0 33824 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_294
timestamp 1698431365
transform 1 0 34272 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_296
timestamp 1698431365
transform 1 0 34496 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_299
timestamp 1698431365
transform 1 0 34832 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_331
timestamp 1698431365
transform 1 0 38416 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_340
timestamp 1698431365
transform 1 0 39424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_348
timestamp 1698431365
transform 1 0 40320 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_356
timestamp 1698431365
transform 1 0 41216 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_18
timestamp 1698431365
transform 1 0 3360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_26
timestamp 1698431365
transform 1 0 4256 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_28
timestamp 1698431365
transform 1 0 4480 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_53
timestamp 1698431365
transform 1 0 7280 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_69
timestamp 1698431365
transform 1 0 9072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_73
timestamp 1698431365
transform 1 0 9520 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_81
timestamp 1698431365
transform 1 0 10416 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_83
timestamp 1698431365
transform 1 0 10640 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_99
timestamp 1698431365
transform 1 0 12432 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_112
timestamp 1698431365
transform 1 0 13888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_145
timestamp 1698431365
transform 1 0 17584 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_149
timestamp 1698431365
transform 1 0 18032 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_153
timestamp 1698431365
transform 1 0 18480 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_157
timestamp 1698431365
transform 1 0 18928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_161
timestamp 1698431365
transform 1 0 19376 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_165
timestamp 1698431365
transform 1 0 19824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_173
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_189
timestamp 1698431365
transform 1 0 22512 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_201
timestamp 1698431365
transform 1 0 23856 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_205
timestamp 1698431365
transform 1 0 24304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_209
timestamp 1698431365
transform 1 0 24752 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_213
timestamp 1698431365
transform 1 0 25200 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698431365
transform 1 0 28560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_279
timestamp 1698431365
transform 1 0 32592 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_283
timestamp 1698431365
transform 1 0 33040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_285
timestamp 1698431365
transform 1 0 33264 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_288
timestamp 1698431365
transform 1 0 33600 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_296
timestamp 1698431365
transform 1 0 34496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_298
timestamp 1698431365
transform 1 0 34720 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_305
timestamp 1698431365
transform 1 0 35504 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_313
timestamp 1698431365
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_333
timestamp 1698431365
transform 1 0 38640 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_337
timestamp 1698431365
transform 1 0 39088 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_343
timestamp 1698431365
transform 1 0 39760 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_347
timestamp 1698431365
transform 1 0 40208 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_379
timestamp 1698431365
transform 1 0 43792 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_383
timestamp 1698431365
transform 1 0 44240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_419
timestamp 1698431365
transform 1 0 48272 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_6
timestamp 1698431365
transform 1 0 2016 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_22
timestamp 1698431365
transform 1 0 3808 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_43
timestamp 1698431365
transform 1 0 6160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_45
timestamp 1698431365
transform 1 0 6384 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_81
timestamp 1698431365
transform 1 0 10416 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_135
timestamp 1698431365
transform 1 0 16464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_137
timestamp 1698431365
transform 1 0 16688 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_186
timestamp 1698431365
transform 1 0 22176 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_190
timestamp 1698431365
transform 1 0 22624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_192
timestamp 1698431365
transform 1 0 22848 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_247
timestamp 1698431365
transform 1 0 29008 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_286
timestamp 1698431365
transform 1 0 33376 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_317
timestamp 1698431365
transform 1 0 36848 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_325
timestamp 1698431365
transform 1 0 37744 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_341
timestamp 1698431365
transform 1 0 39536 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698431365
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_24
timestamp 1698431365
transform 1 0 4032 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_28
timestamp 1698431365
transform 1 0 4480 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_47
timestamp 1698431365
transform 1 0 6608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_51
timestamp 1698431365
transform 1 0 7056 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_83
timestamp 1698431365
transform 1 0 10640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_85
timestamp 1698431365
transform 1 0 10864 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_133
timestamp 1698431365
transform 1 0 16240 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_142
timestamp 1698431365
transform 1 0 17248 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_210
timestamp 1698431365
transform 1 0 24864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_214
timestamp 1698431365
transform 1 0 25312 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_222
timestamp 1698431365
transform 1 0 26208 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_238
timestamp 1698431365
transform 1 0 28000 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_242
timestamp 1698431365
transform 1 0 28448 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_273
timestamp 1698431365
transform 1 0 31920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_277
timestamp 1698431365
transform 1 0 32368 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_285
timestamp 1698431365
transform 1 0 33264 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_296
timestamp 1698431365
transform 1 0 34496 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_304
timestamp 1698431365
transform 1 0 35392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_312
timestamp 1698431365
transform 1 0 36288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_346
timestamp 1698431365
transform 1 0 40096 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_352
timestamp 1698431365
transform 1 0 40768 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_384
timestamp 1698431365
transform 1 0 44352 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_419
timestamp 1698431365
transform 1 0 48272 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_31
timestamp 1698431365
transform 1 0 4816 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_46
timestamp 1698431365
transform 1 0 6496 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_52
timestamp 1698431365
transform 1 0 7168 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1698431365
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_76
timestamp 1698431365
transform 1 0 9856 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_84
timestamp 1698431365
transform 1 0 10752 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_86
timestamp 1698431365
transform 1 0 10976 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_150
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_202
timestamp 1698431365
transform 1 0 23968 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_224
timestamp 1698431365
transform 1 0 26432 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_275
timestamp 1698431365
transform 1 0 32144 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_290
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_294
timestamp 1698431365
transform 1 0 34272 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_310
timestamp 1698431365
transform 1 0 36064 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_314
timestamp 1698431365
transform 1 0 36512 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_324
timestamp 1698431365
transform 1 0 37632 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_328
timestamp 1698431365
transform 1 0 38080 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_330
timestamp 1698431365
transform 1 0 38304 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_381
timestamp 1698431365
transform 1 0 44016 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_413
timestamp 1698431365
transform 1 0 47600 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_417
timestamp 1698431365
transform 1 0 48048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_419
timestamp 1698431365
transform 1 0 48272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_24
timestamp 1698431365
transform 1 0 4032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_28
timestamp 1698431365
transform 1 0 4480 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_30
timestamp 1698431365
transform 1 0 4704 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_33
timestamp 1698431365
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_69
timestamp 1698431365
transform 1 0 9072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_71
timestamp 1698431365
transform 1 0 9296 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_111
timestamp 1698431365
transform 1 0 13776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_141
timestamp 1698431365
transform 1 0 17136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_145
timestamp 1698431365
transform 1 0 17584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_160
timestamp 1698431365
transform 1 0 19264 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_166
timestamp 1698431365
transform 1 0 19936 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_170
timestamp 1698431365
transform 1 0 20384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_185
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_208
timestamp 1698431365
transform 1 0 24640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_212
timestamp 1698431365
transform 1 0 25088 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_228
timestamp 1698431365
transform 1 0 26880 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_236
timestamp 1698431365
transform 1 0 27776 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_240
timestamp 1698431365
transform 1 0 28224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_242
timestamp 1698431365
transform 1 0 28448 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_261
timestamp 1698431365
transform 1 0 30576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_265
timestamp 1698431365
transform 1 0 31024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_267
timestamp 1698431365
transform 1 0 31248 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_297
timestamp 1698431365
transform 1 0 34608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_301
timestamp 1698431365
transform 1 0 35056 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_305
timestamp 1698431365
transform 1 0 35504 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_321
timestamp 1698431365
transform 1 0 37296 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_325
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_329
timestamp 1698431365
transform 1 0 38192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_333
timestamp 1698431365
transform 1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_335
timestamp 1698431365
transform 1 0 38864 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_367
timestamp 1698431365
transform 1 0 42448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_373
timestamp 1698431365
transform 1 0 43120 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_419
timestamp 1698431365
transform 1 0 48272 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_10
timestamp 1698431365
transform 1 0 2464 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_14
timestamp 1698431365
transform 1 0 2912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_23
timestamp 1698431365
transform 1 0 3920 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_55
timestamp 1698431365
transform 1 0 7504 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_63
timestamp 1698431365
transform 1 0 8400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_67
timestamp 1698431365
transform 1 0 8848 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_100
timestamp 1698431365
transform 1 0 12544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_104
timestamp 1698431365
transform 1 0 12992 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698431365
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_150
timestamp 1698431365
transform 1 0 18144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_152
timestamp 1698431365
transform 1 0 18368 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_155
timestamp 1698431365
transform 1 0 18704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_191
timestamp 1698431365
transform 1 0 22736 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_199
timestamp 1698431365
transform 1 0 23632 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_201
timestamp 1698431365
transform 1 0 23856 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_204
timestamp 1698431365
transform 1 0 24192 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698431365
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_228
timestamp 1698431365
transform 1 0 26880 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_236
timestamp 1698431365
transform 1 0 27776 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_238
timestamp 1698431365
transform 1 0 28000 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_245
timestamp 1698431365
transform 1 0 28784 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_253
timestamp 1698431365
transform 1 0 29680 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_257
timestamp 1698431365
transform 1 0 30128 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_265
timestamp 1698431365
transform 1 0 31024 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_268
timestamp 1698431365
transform 1 0 31360 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_288
timestamp 1698431365
transform 1 0 33600 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_294
timestamp 1698431365
transform 1 0 34272 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_298
timestamp 1698431365
transform 1 0 34720 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_339
timestamp 1698431365
transform 1 0 39312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_341
timestamp 1698431365
transform 1 0 39536 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_387
timestamp 1698431365
transform 1 0 44688 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_419
timestamp 1698431365
transform 1 0 48272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_45
timestamp 1698431365
transform 1 0 6384 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_77
timestamp 1698431365
transform 1 0 9968 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_81
timestamp 1698431365
transform 1 0 10416 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_95
timestamp 1698431365
transform 1 0 11984 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_103
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_136
timestamp 1698431365
transform 1 0 16576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_140
timestamp 1698431365
transform 1 0 17024 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_157
timestamp 1698431365
transform 1 0 18928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_159
timestamp 1698431365
transform 1 0 19152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_187
timestamp 1698431365
transform 1 0 22288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_191
timestamp 1698431365
transform 1 0 22736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_195
timestamp 1698431365
transform 1 0 23184 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_227
timestamp 1698431365
transform 1 0 26768 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_243
timestamp 1698431365
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_255
timestamp 1698431365
transform 1 0 29904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_259
timestamp 1698431365
transform 1 0 30352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_266
timestamp 1698431365
transform 1 0 31136 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_270
timestamp 1698431365
transform 1 0 31584 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_286
timestamp 1698431365
transform 1 0 33376 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_294
timestamp 1698431365
transform 1 0 34272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_361
timestamp 1698431365
transform 1 0 41776 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_365
timestamp 1698431365
transform 1 0 42224 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_373
timestamp 1698431365
transform 1 0 43120 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_419
timestamp 1698431365
transform 1 0 48272 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_6
timestamp 1698431365
transform 1 0 2016 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_22
timestamp 1698431365
transform 1 0 3808 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_30
timestamp 1698431365
transform 1 0 4704 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_61
timestamp 1698431365
transform 1 0 8176 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_88
timestamp 1698431365
transform 1 0 11200 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_122
timestamp 1698431365
transform 1 0 15008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_126
timestamp 1698431365
transform 1 0 15456 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_128
timestamp 1698431365
transform 1 0 15680 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698431365
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_164
timestamp 1698431365
transform 1 0 19712 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_170
timestamp 1698431365
transform 1 0 20384 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_174
timestamp 1698431365
transform 1 0 20832 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_183
timestamp 1698431365
transform 1 0 21840 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_187
timestamp 1698431365
transform 1 0 22288 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_203
timestamp 1698431365
transform 1 0 24080 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_241
timestamp 1698431365
transform 1 0 28336 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_255
timestamp 1698431365
transform 1 0 29904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_257
timestamp 1698431365
transform 1 0 30128 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_263
timestamp 1698431365
transform 1 0 30800 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_272
timestamp 1698431365
transform 1 0 31808 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_284
timestamp 1698431365
transform 1 0 33152 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_290
timestamp 1698431365
transform 1 0 33824 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_294
timestamp 1698431365
transform 1 0 34272 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_304
timestamp 1698431365
transform 1 0 35392 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_308
timestamp 1698431365
transform 1 0 35840 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_356
timestamp 1698431365
transform 1 0 41216 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_365
timestamp 1698431365
transform 1 0 42224 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_369
timestamp 1698431365
transform 1 0 42672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_371
timestamp 1698431365
transform 1 0 42896 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_403
timestamp 1698431365
transform 1 0 46480 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_419
timestamp 1698431365
transform 1 0 48272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_26
timestamp 1698431365
transform 1 0 4256 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_74
timestamp 1698431365
transform 1 0 9632 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_90
timestamp 1698431365
transform 1 0 11424 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_98
timestamp 1698431365
transform 1 0 12320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_102
timestamp 1698431365
transform 1 0 12768 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_104
timestamp 1698431365
transform 1 0 12992 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_115
timestamp 1698431365
transform 1 0 14224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_214
timestamp 1698431365
transform 1 0 25312 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_226
timestamp 1698431365
transform 1 0 26656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_230
timestamp 1698431365
transform 1 0 27104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_234
timestamp 1698431365
transform 1 0 27552 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_242
timestamp 1698431365
transform 1 0 28448 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_261
timestamp 1698431365
transform 1 0 30576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_263
timestamp 1698431365
transform 1 0 30800 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_270
timestamp 1698431365
transform 1 0 31584 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_278
timestamp 1698431365
transform 1 0 32480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_282
timestamp 1698431365
transform 1 0 32928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_356
timestamp 1698431365
transform 1 0 41216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_360
timestamp 1698431365
transform 1 0 41664 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_376
timestamp 1698431365
transform 1 0 43456 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_384
timestamp 1698431365
transform 1 0 44352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_395
timestamp 1698431365
transform 1 0 45584 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_411
timestamp 1698431365
transform 1 0 47376 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_419
timestamp 1698431365
transform 1 0 48272 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_31
timestamp 1698431365
transform 1 0 4816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_33
timestamp 1698431365
transform 1 0 5040 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_42
timestamp 1698431365
transform 1 0 6048 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_77
timestamp 1698431365
transform 1 0 9968 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_81
timestamp 1698431365
transform 1 0 10416 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_91
timestamp 1698431365
transform 1 0 11536 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_95
timestamp 1698431365
transform 1 0 11984 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_127
timestamp 1698431365
transform 1 0 15568 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_135
timestamp 1698431365
transform 1 0 16464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_153
timestamp 1698431365
transform 1 0 18480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_157
timestamp 1698431365
transform 1 0 18928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_165
timestamp 1698431365
transform 1 0 19824 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_168
timestamp 1698431365
transform 1 0 20160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_172
timestamp 1698431365
transform 1 0 20608 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_188
timestamp 1698431365
transform 1 0 22400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_208
timestamp 1698431365
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_241
timestamp 1698431365
transform 1 0 28336 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_249
timestamp 1698431365
transform 1 0 29232 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_286
timestamp 1698431365
transform 1 0 33376 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_302
timestamp 1698431365
transform 1 0 35168 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_310
timestamp 1698431365
transform 1 0 36064 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_314
timestamp 1698431365
transform 1 0 36512 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_356
timestamp 1698431365
transform 1 0 41216 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_372
timestamp 1698431365
transform 1 0 43008 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_380
timestamp 1698431365
transform 1 0 43904 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_387
timestamp 1698431365
transform 1 0 44688 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_419
timestamp 1698431365
transform 1 0 48272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_4
timestamp 1698431365
transform 1 0 1792 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_26
timestamp 1698431365
transform 1 0 4256 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_30
timestamp 1698431365
transform 1 0 4704 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_33
timestamp 1698431365
transform 1 0 5040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_39
timestamp 1698431365
transform 1 0 5712 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_50
timestamp 1698431365
transform 1 0 6944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_52
timestamp 1698431365
transform 1 0 7168 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_61
timestamp 1698431365
transform 1 0 8176 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_70
timestamp 1698431365
transform 1 0 9184 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_86
timestamp 1698431365
transform 1 0 10976 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_93
timestamp 1698431365
transform 1 0 11760 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_139
timestamp 1698431365
transform 1 0 16912 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_155
timestamp 1698431365
transform 1 0 18704 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_163
timestamp 1698431365
transform 1 0 19600 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_185
timestamp 1698431365
transform 1 0 22064 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_189
timestamp 1698431365
transform 1 0 22512 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_199
timestamp 1698431365
transform 1 0 23632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_203
timestamp 1698431365
transform 1 0 24080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_213
timestamp 1698431365
transform 1 0 25200 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_217
timestamp 1698431365
transform 1 0 25648 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_225
timestamp 1698431365
transform 1 0 26544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_227
timestamp 1698431365
transform 1 0 26768 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_232
timestamp 1698431365
transform 1 0 27328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_240
timestamp 1698431365
transform 1 0 28224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_279
timestamp 1698431365
transform 1 0 32592 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_295
timestamp 1698431365
transform 1 0 34384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_303
timestamp 1698431365
transform 1 0 35280 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_325
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_329
timestamp 1698431365
transform 1 0 38192 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_361
timestamp 1698431365
transform 1 0 41776 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_377
timestamp 1698431365
transform 1 0 43568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_381
timestamp 1698431365
transform 1 0 44016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_395
timestamp 1698431365
transform 1 0 45584 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_411
timestamp 1698431365
transform 1 0 47376 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_419
timestamp 1698431365
transform 1 0 48272 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_6
timestamp 1698431365
transform 1 0 2016 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_131
timestamp 1698431365
transform 1 0 16016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_135
timestamp 1698431365
transform 1 0 16464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698431365
transform 1 0 16912 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_154
timestamp 1698431365
transform 1 0 18592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_156
timestamp 1698431365
transform 1 0 18816 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_188
timestamp 1698431365
transform 1 0 22400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_200
timestamp 1698431365
transform 1 0 23744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_204
timestamp 1698431365
transform 1 0 24192 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698431365
transform 1 0 24640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_220
timestamp 1698431365
transform 1 0 25984 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_224
timestamp 1698431365
transform 1 0 26432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_260
timestamp 1698431365
transform 1 0 30464 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_264
timestamp 1698431365
transform 1 0 30912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_268
timestamp 1698431365
transform 1 0 31360 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_272
timestamp 1698431365
transform 1 0 31808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_290
timestamp 1698431365
transform 1 0 33824 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_294
timestamp 1698431365
transform 1 0 34272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_303
timestamp 1698431365
transform 1 0 35280 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_307
timestamp 1698431365
transform 1 0 35728 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_323
timestamp 1698431365
transform 1 0 37520 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_333
timestamp 1698431365
transform 1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_343
timestamp 1698431365
transform 1 0 39760 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_347
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_356
timestamp 1698431365
transform 1 0 41216 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_388
timestamp 1698431365
transform 1 0 44800 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_6
timestamp 1698431365
transform 1 0 2016 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_24
timestamp 1698431365
transform 1 0 4032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698431365
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698431365
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_53
timestamp 1698431365
transform 1 0 7280 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_57
timestamp 1698431365
transform 1 0 7728 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_64
timestamp 1698431365
transform 1 0 8512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_69
timestamp 1698431365
transform 1 0 9072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_73
timestamp 1698431365
transform 1 0 9520 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_121
timestamp 1698431365
transform 1 0 14896 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_123
timestamp 1698431365
transform 1 0 15120 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_155
timestamp 1698431365
transform 1 0 18704 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_181
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_195
timestamp 1698431365
transform 1 0 23184 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_199
timestamp 1698431365
transform 1 0 23632 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_231
timestamp 1698431365
transform 1 0 27216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_233
timestamp 1698431365
transform 1 0 27440 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_240
timestamp 1698431365
transform 1 0 28224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_266
timestamp 1698431365
transform 1 0 31136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_297
timestamp 1698431365
transform 1 0 34608 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_305
timestamp 1698431365
transform 1 0 35504 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698431365
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_325
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_331
timestamp 1698431365
transform 1 0 38416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_352
timestamp 1698431365
transform 1 0 40768 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_360
timestamp 1698431365
transform 1 0 41664 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_364
timestamp 1698431365
transform 1 0 42112 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_372
timestamp 1698431365
transform 1 0 43008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_380
timestamp 1698431365
transform 1 0 43904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_384
timestamp 1698431365
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_419
timestamp 1698431365
transform 1 0 48272 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_13
timestamp 1698431365
transform 1 0 2800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_17
timestamp 1698431365
transform 1 0 3248 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_49
timestamp 1698431365
transform 1 0 6832 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_65
timestamp 1698431365
transform 1 0 8624 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_78
timestamp 1698431365
transform 1 0 10080 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_86
timestamp 1698431365
transform 1 0 10976 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_100
timestamp 1698431365
transform 1 0 12544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_104
timestamp 1698431365
transform 1 0 12992 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_112
timestamp 1698431365
transform 1 0 13888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_114
timestamp 1698431365
transform 1 0 14112 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_117
timestamp 1698431365
transform 1 0 14448 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_133
timestamp 1698431365
transform 1 0 16240 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698431365
transform 1 0 16688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_148
timestamp 1698431365
transform 1 0 17920 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_192
timestamp 1698431365
transform 1 0 22848 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_198
timestamp 1698431365
transform 1 0 23520 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_202
timestamp 1698431365
transform 1 0 23968 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_206
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_241
timestamp 1698431365
transform 1 0 28336 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_267
timestamp 1698431365
transform 1 0 31248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_271
timestamp 1698431365
transform 1 0 31696 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_275
timestamp 1698431365
transform 1 0 32144 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_290
timestamp 1698431365
transform 1 0 33824 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_332
timestamp 1698431365
transform 1 0 38528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_336
timestamp 1698431365
transform 1 0 38976 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_340
timestamp 1698431365
transform 1 0 39424 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_348
timestamp 1698431365
transform 1 0 40320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_360
timestamp 1698431365
transform 1 0 41664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_372
timestamp 1698431365
transform 1 0 43008 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_404
timestamp 1698431365
transform 1 0 46592 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_41
timestamp 1698431365
transform 1 0 5936 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_62
timestamp 1698431365
transform 1 0 8288 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_70
timestamp 1698431365
transform 1 0 9184 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_74
timestamp 1698431365
transform 1 0 9632 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_77
timestamp 1698431365
transform 1 0 9968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_123
timestamp 1698431365
transform 1 0 15120 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_131
timestamp 1698431365
transform 1 0 16016 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_181
timestamp 1698431365
transform 1 0 21616 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_225
timestamp 1698431365
transform 1 0 26544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_229
timestamp 1698431365
transform 1 0 26992 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_233
timestamp 1698431365
transform 1 0 27440 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698431365
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_251
timestamp 1698431365
transform 1 0 29456 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_259
timestamp 1698431365
transform 1 0 30352 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_263
timestamp 1698431365
transform 1 0 30800 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_299
timestamp 1698431365
transform 1 0 34832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_303
timestamp 1698431365
transform 1 0 35280 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_305
timestamp 1698431365
transform 1 0 35504 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698431365
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_350
timestamp 1698431365
transform 1 0 40544 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_382
timestamp 1698431365
transform 1 0 44128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_419
timestamp 1698431365
transform 1 0 48272 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_50
timestamp 1698431365
transform 1 0 6944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_60
timestamp 1698431365
transform 1 0 8064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_74
timestamp 1698431365
transform 1 0 9632 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_111
timestamp 1698431365
transform 1 0 13776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_115
timestamp 1698431365
transform 1 0 14224 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_124
timestamp 1698431365
transform 1 0 15232 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_128
timestamp 1698431365
transform 1 0 15680 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_144
timestamp 1698431365
transform 1 0 17472 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_161
timestamp 1698431365
transform 1 0 19376 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_165
timestamp 1698431365
transform 1 0 19824 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_173
timestamp 1698431365
transform 1 0 20720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_177
timestamp 1698431365
transform 1 0 21168 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_221
timestamp 1698431365
transform 1 0 26096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_225
timestamp 1698431365
transform 1 0 26544 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_257
timestamp 1698431365
transform 1 0 30128 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_286
timestamp 1698431365
transform 1 0 33376 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_325
timestamp 1698431365
transform 1 0 37744 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_341
timestamp 1698431365
transform 1 0 39536 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_345
timestamp 1698431365
transform 1 0 39984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_347
timestamp 1698431365
transform 1 0 40208 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_381
timestamp 1698431365
transform 1 0 44016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_385
timestamp 1698431365
transform 1 0 44464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_393
timestamp 1698431365
transform 1 0 45360 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_409
timestamp 1698431365
transform 1 0 47152 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_417
timestamp 1698431365
transform 1 0 48048 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_419
timestamp 1698431365
transform 1 0 48272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_29
timestamp 1698431365
transform 1 0 4592 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_96
timestamp 1698431365
transform 1 0 12096 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_100
timestamp 1698431365
transform 1 0 12544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_102
timestamp 1698431365
transform 1 0 12768 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_117
timestamp 1698431365
transform 1 0 14448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_121
timestamp 1698431365
transform 1 0 14896 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_136
timestamp 1698431365
transform 1 0 16576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_140
timestamp 1698431365
transform 1 0 17024 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_148
timestamp 1698431365
transform 1 0 17920 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_152
timestamp 1698431365
transform 1 0 18368 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_155
timestamp 1698431365
transform 1 0 18704 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_189
timestamp 1698431365
transform 1 0 22512 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_193
timestamp 1698431365
transform 1 0 22960 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_201
timestamp 1698431365
transform 1 0 23856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_207
timestamp 1698431365
transform 1 0 24528 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_209
timestamp 1698431365
transform 1 0 24752 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_212
timestamp 1698431365
transform 1 0 25088 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_216
timestamp 1698431365
transform 1 0 25536 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_224
timestamp 1698431365
transform 1 0 26432 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_228
timestamp 1698431365
transform 1 0 26880 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_240
timestamp 1698431365
transform 1 0 28224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_263
timestamp 1698431365
transform 1 0 30800 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_266
timestamp 1698431365
transform 1 0 31136 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_286
timestamp 1698431365
transform 1 0 33376 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_302
timestamp 1698431365
transform 1 0 35168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_310
timestamp 1698431365
transform 1 0 36064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_321
timestamp 1698431365
transform 1 0 37296 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_360
timestamp 1698431365
transform 1 0 41664 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_372
timestamp 1698431365
transform 1 0 43008 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_380
timestamp 1698431365
transform 1 0 43904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_382
timestamp 1698431365
transform 1 0 44128 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_416
timestamp 1698431365
transform 1 0 47936 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_10
timestamp 1698431365
transform 1 0 2464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_16
timestamp 1698431365
transform 1 0 3136 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_50
timestamp 1698431365
transform 1 0 6944 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_59
timestamp 1698431365
transform 1 0 7952 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_133
timestamp 1698431365
transform 1 0 16240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_137
timestamp 1698431365
transform 1 0 16688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_146
timestamp 1698431365
transform 1 0 17696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_148
timestamp 1698431365
transform 1 0 17920 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_155
timestamp 1698431365
transform 1 0 18704 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_159
timestamp 1698431365
transform 1 0 19152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_161
timestamp 1698431365
transform 1 0 19376 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_205
timestamp 1698431365
transform 1 0 24304 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_216
timestamp 1698431365
transform 1 0 25536 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_248
timestamp 1698431365
transform 1 0 29120 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_254
timestamp 1698431365
transform 1 0 29792 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_258
timestamp 1698431365
transform 1 0 30240 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_274
timestamp 1698431365
transform 1 0 32032 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_298
timestamp 1698431365
transform 1 0 34720 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_306
timestamp 1698431365
transform 1 0 35616 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_310
timestamp 1698431365
transform 1 0 36064 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_317
timestamp 1698431365
transform 1 0 36848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_321
timestamp 1698431365
transform 1 0 37296 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_337
timestamp 1698431365
transform 1 0 39088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_345
timestamp 1698431365
transform 1 0 39984 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_360
timestamp 1698431365
transform 1 0 41664 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_367
timestamp 1698431365
transform 1 0 42448 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_369
timestamp 1698431365
transform 1 0 42672 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_401
timestamp 1698431365
transform 1 0 46256 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_417
timestamp 1698431365
transform 1 0 48048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_419
timestamp 1698431365
transform 1 0 48272 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_6
timestamp 1698431365
transform 1 0 2016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_10
timestamp 1698431365
transform 1 0 2464 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_26
timestamp 1698431365
transform 1 0 4256 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_53
timestamp 1698431365
transform 1 0 7280 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_65
timestamp 1698431365
transform 1 0 8624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_69
timestamp 1698431365
transform 1 0 9072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_73
timestamp 1698431365
transform 1 0 9520 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_97
timestamp 1698431365
transform 1 0 12208 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698431365
transform 1 0 13776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_144
timestamp 1698431365
transform 1 0 17472 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698431365
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_181
timestamp 1698431365
transform 1 0 21616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_189
timestamp 1698431365
transform 1 0 22512 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_228
timestamp 1698431365
transform 1 0 26880 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_236
timestamp 1698431365
transform 1 0 27776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_238
timestamp 1698431365
transform 1 0 28000 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_251
timestamp 1698431365
transform 1 0 29456 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_255
timestamp 1698431365
transform 1 0 29904 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_271
timestamp 1698431365
transform 1 0 31696 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_275
timestamp 1698431365
transform 1 0 32144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_284
timestamp 1698431365
transform 1 0 33152 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_288
timestamp 1698431365
transform 1 0 33600 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_304
timestamp 1698431365
transform 1 0 35392 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_381
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_395
timestamp 1698431365
transform 1 0 45584 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_411
timestamp 1698431365
transform 1 0 47376 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_419
timestamp 1698431365
transform 1 0 48272 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_26
timestamp 1698431365
transform 1 0 4256 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_34
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_40
timestamp 1698431365
transform 1 0 5824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_42
timestamp 1698431365
transform 1 0 6048 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_45
timestamp 1698431365
transform 1 0 6384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_64
timestamp 1698431365
transform 1 0 8512 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_80
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_84
timestamp 1698431365
transform 1 0 10752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_87
timestamp 1698431365
transform 1 0 11088 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_103
timestamp 1698431365
transform 1 0 12880 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_105
timestamp 1698431365
transform 1 0 13104 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_120
timestamp 1698431365
transform 1 0 14784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_128
timestamp 1698431365
transform 1 0 15680 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_144
timestamp 1698431365
transform 1 0 17472 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_153
timestamp 1698431365
transform 1 0 18480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_157
timestamp 1698431365
transform 1 0 18928 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_173
timestamp 1698431365
transform 1 0 20720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_218
timestamp 1698431365
transform 1 0 25760 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_222
timestamp 1698431365
transform 1 0 26208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_228
timestamp 1698431365
transform 1 0 26880 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_232
timestamp 1698431365
transform 1 0 27328 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_239
timestamp 1698431365
transform 1 0 28112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_241
timestamp 1698431365
transform 1 0 28336 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_308
timestamp 1698431365
transform 1 0 35840 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_312
timestamp 1698431365
transform 1 0 36288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_314
timestamp 1698431365
transform 1 0 36512 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_317
timestamp 1698431365
transform 1 0 36848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_319
timestamp 1698431365
transform 1 0 37072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_326
timestamp 1698431365
transform 1 0 37856 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_342
timestamp 1698431365
transform 1 0 39648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_346
timestamp 1698431365
transform 1 0 40096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_368
timestamp 1698431365
transform 1 0 42560 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_376
timestamp 1698431365
transform 1 0 43456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_384
timestamp 1698431365
transform 1 0 44352 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_416
timestamp 1698431365
transform 1 0 47936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_6
timestamp 1698431365
transform 1 0 2016 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_8
timestamp 1698431365
transform 1 0 2240 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_39
timestamp 1698431365
transform 1 0 5712 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_48
timestamp 1698431365
transform 1 0 6720 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_52
timestamp 1698431365
transform 1 0 7168 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_65
timestamp 1698431365
transform 1 0 8624 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_69
timestamp 1698431365
transform 1 0 9072 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_72
timestamp 1698431365
transform 1 0 9408 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_76
timestamp 1698431365
transform 1 0 9856 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_86
timestamp 1698431365
transform 1 0 10976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_90
timestamp 1698431365
transform 1 0 11424 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_94
timestamp 1698431365
transform 1 0 11872 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_102
timestamp 1698431365
transform 1 0 12768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_115
timestamp 1698431365
transform 1 0 14224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_119
timestamp 1698431365
transform 1 0 14672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_122
timestamp 1698431365
transform 1 0 15008 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_138
timestamp 1698431365
transform 1 0 16800 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_146
timestamp 1698431365
transform 1 0 17696 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_154
timestamp 1698431365
transform 1 0 18592 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_170
timestamp 1698431365
transform 1 0 20384 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_193
timestamp 1698431365
transform 1 0 22960 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_205
timestamp 1698431365
transform 1 0 24304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_209
timestamp 1698431365
transform 1 0 24752 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_213
timestamp 1698431365
transform 1 0 25200 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_265
timestamp 1698431365
transform 1 0 31024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_269
timestamp 1698431365
transform 1 0 31472 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_273
timestamp 1698431365
transform 1 0 31920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_277
timestamp 1698431365
transform 1 0 32368 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_281
timestamp 1698431365
transform 1 0 32816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_283
timestamp 1698431365
transform 1 0 33040 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_352
timestamp 1698431365
transform 1 0 40768 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_368
timestamp 1698431365
transform 1 0 42560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_382
timestamp 1698431365
transform 1 0 44128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_384
timestamp 1698431365
transform 1 0 44352 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_419
timestamp 1698431365
transform 1 0 48272 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_25
timestamp 1698431365
transform 1 0 4144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_62
timestamp 1698431365
transform 1 0 8288 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_64
timestamp 1698431365
transform 1 0 8512 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_82
timestamp 1698431365
transform 1 0 10528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_131
timestamp 1698431365
transform 1 0 16016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_135
timestamp 1698431365
transform 1 0 16464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_137
timestamp 1698431365
transform 1 0 16688 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_173
timestamp 1698431365
transform 1 0 20720 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_181
timestamp 1698431365
transform 1 0 21616 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_185
timestamp 1698431365
transform 1 0 22064 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_219
timestamp 1698431365
transform 1 0 25872 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_273
timestamp 1698431365
transform 1 0 31920 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_277
timestamp 1698431365
transform 1 0 32368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_286
timestamp 1698431365
transform 1 0 33376 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_290
timestamp 1698431365
transform 1 0 33824 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_294
timestamp 1698431365
transform 1 0 34272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_303
timestamp 1698431365
transform 1 0 35280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_307
timestamp 1698431365
transform 1 0 35728 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_311
timestamp 1698431365
transform 1 0 36176 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_315
timestamp 1698431365
transform 1 0 36624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_327
timestamp 1698431365
transform 1 0 37968 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_335
timestamp 1698431365
transform 1 0 38864 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_339
timestamp 1698431365
transform 1 0 39312 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_341
timestamp 1698431365
transform 1 0 39536 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_381
timestamp 1698431365
transform 1 0 44016 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_397
timestamp 1698431365
transform 1 0 45808 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_405
timestamp 1698431365
transform 1 0 46704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_407
timestamp 1698431365
transform 1 0 46928 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_412
timestamp 1698431365
transform 1 0 47488 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_41
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_45
timestamp 1698431365
transform 1 0 6384 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_99
timestamp 1698431365
transform 1 0 12432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_103
timestamp 1698431365
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_111
timestamp 1698431365
transform 1 0 13776 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_127
timestamp 1698431365
transform 1 0 15568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_129
timestamp 1698431365
transform 1 0 15792 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_138
timestamp 1698431365
transform 1 0 16800 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_142
timestamp 1698431365
transform 1 0 17248 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_146
timestamp 1698431365
transform 1 0 17696 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_162
timestamp 1698431365
transform 1 0 19488 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_170
timestamp 1698431365
transform 1 0 20384 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_193
timestamp 1698431365
transform 1 0 22960 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_201
timestamp 1698431365
transform 1 0 23856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_205
timestamp 1698431365
transform 1 0 24304 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_208
timestamp 1698431365
transform 1 0 24640 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_216
timestamp 1698431365
transform 1 0 25536 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_218
timestamp 1698431365
transform 1 0 25760 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_221
timestamp 1698431365
transform 1 0 26096 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_225
timestamp 1698431365
transform 1 0 26544 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_228
timestamp 1698431365
transform 1 0 26880 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_238
timestamp 1698431365
transform 1 0 28000 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_242
timestamp 1698431365
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_268
timestamp 1698431365
transform 1 0 31360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_270
timestamp 1698431365
transform 1 0 31584 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_273
timestamp 1698431365
transform 1 0 31920 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_277
timestamp 1698431365
transform 1 0 32368 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_281
timestamp 1698431365
transform 1 0 32816 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_283
timestamp 1698431365
transform 1 0 33040 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_296
timestamp 1698431365
transform 1 0 34496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_300
timestamp 1698431365
transform 1 0 34944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_326
timestamp 1698431365
transform 1 0 37856 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_359
timestamp 1698431365
transform 1 0 41552 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_369
timestamp 1698431365
transform 1 0 42672 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_373
timestamp 1698431365
transform 1 0 43120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_377
timestamp 1698431365
transform 1 0 43568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_381
timestamp 1698431365
transform 1 0 44016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_417
timestamp 1698431365
transform 1 0 48048 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_419
timestamp 1698431365
transform 1 0 48272 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_42
timestamp 1698431365
transform 1 0 6048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_44
timestamp 1698431365
transform 1 0 6272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_53
timestamp 1698431365
transform 1 0 7280 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_57
timestamp 1698431365
transform 1 0 7728 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_59
timestamp 1698431365
transform 1 0 7952 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_109
timestamp 1698431365
transform 1 0 13552 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_148
timestamp 1698431365
transform 1 0 17920 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_164
timestamp 1698431365
transform 1 0 19712 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_168
timestamp 1698431365
transform 1 0 20160 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_177
timestamp 1698431365
transform 1 0 21168 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_181
timestamp 1698431365
transform 1 0 21616 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_183
timestamp 1698431365
transform 1 0 21840 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_186
timestamp 1698431365
transform 1 0 22176 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_202
timestamp 1698431365
transform 1 0 23968 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_222
timestamp 1698431365
transform 1 0 26208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_226
timestamp 1698431365
transform 1 0 26656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_265
timestamp 1698431365
transform 1 0 31024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_267
timestamp 1698431365
transform 1 0 31248 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_286
timestamp 1698431365
transform 1 0 33376 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_290
timestamp 1698431365
transform 1 0 33824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_294
timestamp 1698431365
transform 1 0 34272 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_298
timestamp 1698431365
transform 1 0 34720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_302
timestamp 1698431365
transform 1 0 35168 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_306
timestamp 1698431365
transform 1 0 35616 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_310
timestamp 1698431365
transform 1 0 36064 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_314
timestamp 1698431365
transform 1 0 36512 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_317
timestamp 1698431365
transform 1 0 36848 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_325
timestamp 1698431365
transform 1 0 37744 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_327
timestamp 1698431365
transform 1 0 37968 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_330
timestamp 1698431365
transform 1 0 38304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_334
timestamp 1698431365
transform 1 0 38752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_345
timestamp 1698431365
transform 1 0 39984 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_360
timestamp 1698431365
transform 1 0 41664 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_364
timestamp 1698431365
transform 1 0 42112 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_368
timestamp 1698431365
transform 1 0 42560 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_386
timestamp 1698431365
transform 1 0 44576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_396
timestamp 1698431365
transform 1 0 45696 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_412
timestamp 1698431365
transform 1 0 47488 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_10
timestamp 1698431365
transform 1 0 2464 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_29
timestamp 1698431365
transform 1 0 4592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_33
timestamp 1698431365
transform 1 0 5040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_52
timestamp 1698431365
transform 1 0 7168 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_61
timestamp 1698431365
transform 1 0 8176 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_69
timestamp 1698431365
transform 1 0 9072 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_73
timestamp 1698431365
transform 1 0 9520 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_77
timestamp 1698431365
transform 1 0 9968 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_81
timestamp 1698431365
transform 1 0 10416 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_89
timestamp 1698431365
transform 1 0 11312 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_91
timestamp 1698431365
transform 1 0 11536 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_100
timestamp 1698431365
transform 1 0 12544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_115
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_119
timestamp 1698431365
transform 1 0 14672 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_154
timestamp 1698431365
transform 1 0 18592 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_162
timestamp 1698431365
transform 1 0 19488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_164
timestamp 1698431365
transform 1 0 19712 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_167
timestamp 1698431365
transform 1 0 20048 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_183
timestamp 1698431365
transform 1 0 21840 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_185
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_215
timestamp 1698431365
transform 1 0 25424 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_223
timestamp 1698431365
transform 1 0 26320 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_227
timestamp 1698431365
transform 1 0 26768 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_231
timestamp 1698431365
transform 1 0 27216 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_239
timestamp 1698431365
transform 1 0 28112 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_301
timestamp 1698431365
transform 1 0 35056 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_305
timestamp 1698431365
transform 1 0 35504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_309
timestamp 1698431365
transform 1 0 35952 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_313
timestamp 1698431365
transform 1 0 36400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_321
timestamp 1698431365
transform 1 0 37296 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_337
timestamp 1698431365
transform 1 0 39088 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_345
timestamp 1698431365
transform 1 0 39984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_347
timestamp 1698431365
transform 1 0 40208 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_350
timestamp 1698431365
transform 1 0 40544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_354
timestamp 1698431365
transform 1 0 40992 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_374
timestamp 1698431365
transform 1 0 43232 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_382
timestamp 1698431365
transform 1 0 44128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_384
timestamp 1698431365
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_391
timestamp 1698431365
transform 1 0 45136 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_407
timestamp 1698431365
transform 1 0 46928 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_415
timestamp 1698431365
transform 1 0 47824 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_419
timestamp 1698431365
transform 1 0 48272 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_13
timestamp 1698431365
transform 1 0 2800 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_20
timestamp 1698431365
transform 1 0 3584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_22
timestamp 1698431365
transform 1 0 3808 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_41
timestamp 1698431365
transform 1 0 5936 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_45
timestamp 1698431365
transform 1 0 6384 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_61
timestamp 1698431365
transform 1 0 8176 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_80
timestamp 1698431365
transform 1 0 10304 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_85
timestamp 1698431365
transform 1 0 10864 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_89
timestamp 1698431365
transform 1 0 11312 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_92
timestamp 1698431365
transform 1 0 11648 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_123
timestamp 1698431365
transform 1 0 15120 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_127
timestamp 1698431365
transform 1 0 15568 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_135
timestamp 1698431365
transform 1 0 16464 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_150
timestamp 1698431365
transform 1 0 18144 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_154
timestamp 1698431365
transform 1 0 18592 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_194
timestamp 1698431365
transform 1 0 23072 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_224
timestamp 1698431365
transform 1 0 26432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_227
timestamp 1698431365
transform 1 0 26768 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_243
timestamp 1698431365
transform 1 0 28560 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_255
timestamp 1698431365
transform 1 0 29904 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_259
timestamp 1698431365
transform 1 0 30352 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_262
timestamp 1698431365
transform 1 0 30688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_264
timestamp 1698431365
transform 1 0 30912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_343
timestamp 1698431365
transform 1 0 39760 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_347
timestamp 1698431365
transform 1 0 40208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_356
timestamp 1698431365
transform 1 0 41216 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_360
timestamp 1698431365
transform 1 0 41664 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_368
timestamp 1698431365
transform 1 0 42560 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_399
timestamp 1698431365
transform 1 0 46032 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_404
timestamp 1698431365
transform 1 0 46592 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_6
timestamp 1698431365
transform 1 0 2016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_8
timestamp 1698431365
transform 1 0 2240 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_28
timestamp 1698431365
transform 1 0 4480 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_32
timestamp 1698431365
transform 1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_45
timestamp 1698431365
transform 1 0 6384 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_51
timestamp 1698431365
transform 1 0 7056 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_83
timestamp 1698431365
transform 1 0 10640 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_87
timestamp 1698431365
transform 1 0 11088 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_90
timestamp 1698431365
transform 1 0 11424 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_94
timestamp 1698431365
transform 1 0 11872 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_102
timestamp 1698431365
transform 1 0 12768 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_113
timestamp 1698431365
transform 1 0 14000 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_117
timestamp 1698431365
transform 1 0 14448 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_120
timestamp 1698431365
transform 1 0 14784 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_136
timestamp 1698431365
transform 1 0 16576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_144
timestamp 1698431365
transform 1 0 17472 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_146
timestamp 1698431365
transform 1 0 17696 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_155
timestamp 1698431365
transform 1 0 18704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_157
timestamp 1698431365
transform 1 0 18928 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_164
timestamp 1698431365
transform 1 0 19712 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_168
timestamp 1698431365
transform 1 0 20160 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_172
timestamp 1698431365
transform 1 0 20608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_174
timestamp 1698431365
transform 1 0 20832 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_209
timestamp 1698431365
transform 1 0 24752 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_213
timestamp 1698431365
transform 1 0 25200 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_215
timestamp 1698431365
transform 1 0 25424 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_259
timestamp 1698431365
transform 1 0 30352 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_261
timestamp 1698431365
transform 1 0 30576 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_278
timestamp 1698431365
transform 1 0 32480 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_282
timestamp 1698431365
transform 1 0 32928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_284
timestamp 1698431365
transform 1 0 33152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698431365
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_321
timestamp 1698431365
transform 1 0 37296 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_323
timestamp 1698431365
transform 1 0 37520 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_326
timestamp 1698431365
transform 1 0 37856 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_330
timestamp 1698431365
transform 1 0 38304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_348
timestamp 1698431365
transform 1 0 40320 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_352
timestamp 1698431365
transform 1 0 40768 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_358
timestamp 1698431365
transform 1 0 41440 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_376
timestamp 1698431365
transform 1 0 43456 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_380
timestamp 1698431365
transform 1 0 43904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_382
timestamp 1698431365
transform 1 0 44128 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_416
timestamp 1698431365
transform 1 0 47936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_36
timestamp 1698431365
transform 1 0 5376 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_40
timestamp 1698431365
transform 1 0 5824 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_58
timestamp 1698431365
transform 1 0 7840 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_60
timestamp 1698431365
transform 1 0 8064 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_63
timestamp 1698431365
transform 1 0 8400 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_67
timestamp 1698431365
transform 1 0 8848 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_88
timestamp 1698431365
transform 1 0 11200 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_118
timestamp 1698431365
transform 1 0 14560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_122
timestamp 1698431365
transform 1 0 15008 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_128
timestamp 1698431365
transform 1 0 15680 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_175
timestamp 1698431365
transform 1 0 20944 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_207
timestamp 1698431365
transform 1 0 24528 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_259
timestamp 1698431365
transform 1 0 30352 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_286
timestamp 1698431365
transform 1 0 33376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_290
timestamp 1698431365
transform 1 0 33824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_294
timestamp 1698431365
transform 1 0 34272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_298
timestamp 1698431365
transform 1 0 34720 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_302
timestamp 1698431365
transform 1 0 35168 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_310
timestamp 1698431365
transform 1 0 36064 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_326
timestamp 1698431365
transform 1 0 37856 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_330
timestamp 1698431365
transform 1 0 38304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_332
timestamp 1698431365
transform 1 0 38528 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_348
timestamp 1698431365
transform 1 0 40320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_360
timestamp 1698431365
transform 1 0 41664 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_362
timestamp 1698431365
transform 1 0 41888 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_369
timestamp 1698431365
transform 1 0 42672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_404
timestamp 1698431365
transform 1 0 46592 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_6
timestamp 1698431365
transform 1 0 2016 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_8
timestamp 1698431365
transform 1 0 2240 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_39
timestamp 1698431365
transform 1 0 5712 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_57
timestamp 1698431365
transform 1 0 7728 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_92
timestamp 1698431365
transform 1 0 11648 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_100
timestamp 1698431365
transform 1 0 12544 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_109
timestamp 1698431365
transform 1 0 13552 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_118
timestamp 1698431365
transform 1 0 14560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_120
timestamp 1698431365
transform 1 0 14784 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_150
timestamp 1698431365
transform 1 0 18144 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_166
timestamp 1698431365
transform 1 0 19936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_170
timestamp 1698431365
transform 1 0 20384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_172
timestamp 1698431365
transform 1 0 20608 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_185
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_187
timestamp 1698431365
transform 1 0 22288 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_202
timestamp 1698431365
transform 1 0 23968 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_206
timestamp 1698431365
transform 1 0 24416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_218
timestamp 1698431365
transform 1 0 25760 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_220
timestamp 1698431365
transform 1 0 25984 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_223
timestamp 1698431365
transform 1 0 26320 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_227
timestamp 1698431365
transform 1 0 26768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_255
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_257
timestamp 1698431365
transform 1 0 30128 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_289
timestamp 1698431365
transform 1 0 33712 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_293
timestamp 1698431365
transform 1 0 34160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_295
timestamp 1698431365
transform 1 0 34384 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_312
timestamp 1698431365
transform 1 0 36288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_314
timestamp 1698431365
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_333
timestamp 1698431365
transform 1 0 38640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_381
timestamp 1698431365
transform 1 0 44016 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_393
timestamp 1698431365
transform 1 0 45360 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_409
timestamp 1698431365
transform 1 0 47152 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_417
timestamp 1698431365
transform 1 0 48048 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_419
timestamp 1698431365
transform 1 0 48272 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_14
timestamp 1698431365
transform 1 0 2912 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_18
timestamp 1698431365
transform 1 0 3360 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_64
timestamp 1698431365
transform 1 0 8512 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_68
timestamp 1698431365
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_76
timestamp 1698431365
transform 1 0 9856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_138
timestamp 1698431365
transform 1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_156
timestamp 1698431365
transform 1 0 18816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_160
timestamp 1698431365
transform 1 0 19264 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_176
timestamp 1698431365
transform 1 0 21056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_178
timestamp 1698431365
transform 1 0 21280 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_228
timestamp 1698431365
transform 1 0 26880 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_232
timestamp 1698431365
transform 1 0 27328 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_234
timestamp 1698431365
transform 1 0 27552 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_267
timestamp 1698431365
transform 1 0 31248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_275
timestamp 1698431365
transform 1 0 32144 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_277
timestamp 1698431365
transform 1 0 32368 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_290
timestamp 1698431365
transform 1 0 33824 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_325
timestamp 1698431365
transform 1 0 37744 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_333
timestamp 1698431365
transform 1 0 38640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_349
timestamp 1698431365
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_368
timestamp 1698431365
transform 1 0 42560 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_377
timestamp 1698431365
transform 1 0 43568 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_409
timestamp 1698431365
transform 1 0 47152 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_417
timestamp 1698431365
transform 1 0 48048 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_419
timestamp 1698431365
transform 1 0 48272 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_6
timestamp 1698431365
transform 1 0 2016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_18
timestamp 1698431365
transform 1 0 3360 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_28
timestamp 1698431365
transform 1 0 4480 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_45
timestamp 1698431365
transform 1 0 6384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_55
timestamp 1698431365
transform 1 0 7504 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_59
timestamp 1698431365
transform 1 0 7952 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_71
timestamp 1698431365
transform 1 0 9296 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_79
timestamp 1698431365
transform 1 0 10192 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_81
timestamp 1698431365
transform 1 0 10416 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_100
timestamp 1698431365
transform 1 0 12544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_104
timestamp 1698431365
transform 1 0 12992 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_111
timestamp 1698431365
transform 1 0 13776 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_113
timestamp 1698431365
transform 1 0 14000 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_160
timestamp 1698431365
transform 1 0 19264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_164
timestamp 1698431365
transform 1 0 19712 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_172
timestamp 1698431365
transform 1 0 20608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_184
timestamp 1698431365
transform 1 0 21952 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_216
timestamp 1698431365
transform 1 0 25536 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_220
timestamp 1698431365
transform 1 0 25984 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_228
timestamp 1698431365
transform 1 0 26880 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_231
timestamp 1698431365
transform 1 0 27216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_235
timestamp 1698431365
transform 1 0 27664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_239
timestamp 1698431365
transform 1 0 28112 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_243
timestamp 1698431365
transform 1 0 28560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_283
timestamp 1698431365
transform 1 0 33040 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_291
timestamp 1698431365
transform 1 0 33936 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_293
timestamp 1698431365
transform 1 0 34160 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_300
timestamp 1698431365
transform 1 0 34944 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_308
timestamp 1698431365
transform 1 0 35840 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_312
timestamp 1698431365
transform 1 0 36288 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_347
timestamp 1698431365
transform 1 0 40208 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_355
timestamp 1698431365
transform 1 0 41104 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_371
timestamp 1698431365
transform 1 0 42896 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_379
timestamp 1698431365
transform 1 0 43792 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_383
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_391
timestamp 1698431365
transform 1 0 45136 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_407
timestamp 1698431365
transform 1 0 46928 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_415
timestamp 1698431365
transform 1 0 47824 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_419
timestamp 1698431365
transform 1 0 48272 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_6
timestamp 1698431365
transform 1 0 2016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_8
timestamp 1698431365
transform 1 0 2240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_16
timestamp 1698431365
transform 1 0 3136 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_20
timestamp 1698431365
transform 1 0 3584 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_36
timestamp 1698431365
transform 1 0 5376 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_45
timestamp 1698431365
transform 1 0 6384 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_53
timestamp 1698431365
transform 1 0 7280 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_57
timestamp 1698431365
transform 1 0 7728 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_59
timestamp 1698431365
transform 1 0 7952 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_62
timestamp 1698431365
transform 1 0 8288 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_80
timestamp 1698431365
transform 1 0 10304 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_82
timestamp 1698431365
transform 1 0 10528 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_85
timestamp 1698431365
transform 1 0 10864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_125
timestamp 1698431365
transform 1 0 15344 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_129
timestamp 1698431365
transform 1 0 15792 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_132
timestamp 1698431365
transform 1 0 16128 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_168
timestamp 1698431365
transform 1 0 20160 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_172
timestamp 1698431365
transform 1 0 20608 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_204
timestamp 1698431365
transform 1 0 24192 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_218
timestamp 1698431365
transform 1 0 25760 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_234
timestamp 1698431365
transform 1 0 27552 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_238
timestamp 1698431365
transform 1 0 28000 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_241
timestamp 1698431365
transform 1 0 28336 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_249
timestamp 1698431365
transform 1 0 29232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_251
timestamp 1698431365
transform 1 0 29456 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_254
timestamp 1698431365
transform 1 0 29792 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_258
timestamp 1698431365
transform 1 0 30240 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_260
timestamp 1698431365
transform 1 0 30464 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_268
timestamp 1698431365
transform 1 0 31360 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_272
timestamp 1698431365
transform 1 0 31808 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_300
timestamp 1698431365
transform 1 0 34944 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_304
timestamp 1698431365
transform 1 0 35392 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_308
timestamp 1698431365
transform 1 0 35840 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_311
timestamp 1698431365
transform 1 0 36176 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_317
timestamp 1698431365
transform 1 0 36848 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_321
timestamp 1698431365
transform 1 0 37296 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_328
timestamp 1698431365
transform 1 0 38080 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_344
timestamp 1698431365
transform 1 0 39872 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_348
timestamp 1698431365
transform 1 0 40320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_356
timestamp 1698431365
transform 1 0 41216 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_359
timestamp 1698431365
transform 1 0 41552 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_367
timestamp 1698431365
transform 1 0 42448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_402
timestamp 1698431365
transform 1 0 46368 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_418
timestamp 1698431365
transform 1 0 48160 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_31
timestamp 1698431365
transform 1 0 4816 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_41
timestamp 1698431365
transform 1 0 5936 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_55
timestamp 1698431365
transform 1 0 7504 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_59
timestamp 1698431365
transform 1 0 7952 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_91
timestamp 1698431365
transform 1 0 11536 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_99
timestamp 1698431365
transform 1 0 12432 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_103
timestamp 1698431365
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_111
timestamp 1698431365
transform 1 0 13776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_145
timestamp 1698431365
transform 1 0 17584 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_181
timestamp 1698431365
transform 1 0 21616 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_197
timestamp 1698431365
transform 1 0 23408 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_205
timestamp 1698431365
transform 1 0 24304 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_214
timestamp 1698431365
transform 1 0 25312 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_224
timestamp 1698431365
transform 1 0 26432 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_239
timestamp 1698431365
transform 1 0 28112 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_243
timestamp 1698431365
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_309
timestamp 1698431365
transform 1 0 35952 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_313
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_325
timestamp 1698431365
transform 1 0 37744 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_330
timestamp 1698431365
transform 1 0 38304 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698431365
transform 1 0 40096 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698431365
transform 1 0 40320 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_389
timestamp 1698431365
transform 1 0 44912 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_419
timestamp 1698431365
transform 1 0 48272 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_32
timestamp 1698431365
transform 1 0 4928 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_36
timestamp 1698431365
transform 1 0 5376 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_61
timestamp 1698431365
transform 1 0 8176 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_146
timestamp 1698431365
transform 1 0 17696 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_150
timestamp 1698431365
transform 1 0 18144 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_154
timestamp 1698431365
transform 1 0 18592 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_216
timestamp 1698431365
transform 1 0 25536 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_218
timestamp 1698431365
transform 1 0 25760 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_226
timestamp 1698431365
transform 1 0 26656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_230
timestamp 1698431365
transform 1 0 27104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_234
timestamp 1698431365
transform 1 0 27552 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_246
timestamp 1698431365
transform 1 0 28896 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_258
timestamp 1698431365
transform 1 0 30240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_262
timestamp 1698431365
transform 1 0 30688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_266
timestamp 1698431365
transform 1 0 31136 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_270
timestamp 1698431365
transform 1 0 31584 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_274
timestamp 1698431365
transform 1 0 32032 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_314
timestamp 1698431365
transform 1 0 36512 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_318
timestamp 1698431365
transform 1 0 36960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_322
timestamp 1698431365
transform 1 0 37408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_326
timestamp 1698431365
transform 1 0 37856 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_330
timestamp 1698431365
transform 1 0 38304 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_346
timestamp 1698431365
transform 1 0 40096 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_354
timestamp 1698431365
transform 1 0 40992 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_398
timestamp 1698431365
transform 1 0 45920 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_414
timestamp 1698431365
transform 1 0 47712 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_418
timestamp 1698431365
transform 1 0 48160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_39
timestamp 1698431365
transform 1 0 5712 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_80
timestamp 1698431365
transform 1 0 10304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_82
timestamp 1698431365
transform 1 0 10528 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_111
timestamp 1698431365
transform 1 0 13776 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_119
timestamp 1698431365
transform 1 0 14672 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_123
timestamp 1698431365
transform 1 0 15120 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_170
timestamp 1698431365
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_172
timestamp 1698431365
transform 1 0 20608 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_206
timestamp 1698431365
transform 1 0 24416 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_222
timestamp 1698431365
transform 1 0 26208 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_226
timestamp 1698431365
transform 1 0 26656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_228
timestamp 1698431365
transform 1 0 26880 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_238
timestamp 1698431365
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_242
timestamp 1698431365
transform 1 0 28448 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_251
timestamp 1698431365
transform 1 0 29456 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_255
timestamp 1698431365
transform 1 0 29904 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_259
timestamp 1698431365
transform 1 0 30352 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_263
timestamp 1698431365
transform 1 0 30800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_269
timestamp 1698431365
transform 1 0 31472 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_323
timestamp 1698431365
transform 1 0 37520 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_325
timestamp 1698431365
transform 1 0 37744 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_355
timestamp 1698431365
transform 1 0 41104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_359
timestamp 1698431365
transform 1 0 41552 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_419
timestamp 1698431365
transform 1 0 48272 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_76
timestamp 1698431365
transform 1 0 9856 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_80
timestamp 1698431365
transform 1 0 10304 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_84
timestamp 1698431365
transform 1 0 10752 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_88
timestamp 1698431365
transform 1 0 11200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_121
timestamp 1698431365
transform 1 0 14896 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_123
timestamp 1698431365
transform 1 0 15120 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_130
timestamp 1698431365
transform 1 0 15904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_134
timestamp 1698431365
transform 1 0 16352 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_138
timestamp 1698431365
transform 1 0 16800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_168
timestamp 1698431365
transform 1 0 20160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_170
timestamp 1698431365
transform 1 0 20384 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_182
timestamp 1698431365
transform 1 0 21728 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_186
timestamp 1698431365
transform 1 0 22176 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_202
timestamp 1698431365
transform 1 0 23968 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_220
timestamp 1698431365
transform 1 0 25984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_233
timestamp 1698431365
transform 1 0 27440 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_278
timestamp 1698431365
transform 1 0 32480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_286
timestamp 1698431365
transform 1 0 33376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_290
timestamp 1698431365
transform 1 0 33824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_294
timestamp 1698431365
transform 1 0 34272 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_325
timestamp 1698431365
transform 1 0 37744 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_329
timestamp 1698431365
transform 1 0 38192 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_333
timestamp 1698431365
transform 1 0 38640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_337
timestamp 1698431365
transform 1 0 39088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_347
timestamp 1698431365
transform 1 0 40208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_349
timestamp 1698431365
transform 1 0 40432 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_356
timestamp 1698431365
transform 1 0 41216 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_360
timestamp 1698431365
transform 1 0 41664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_364
timestamp 1698431365
transform 1 0 42112 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_368
timestamp 1698431365
transform 1 0 42560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_372
timestamp 1698431365
transform 1 0 43008 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_378
timestamp 1698431365
transform 1 0 43680 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_410
timestamp 1698431365
transform 1 0 47264 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_418
timestamp 1698431365
transform 1 0 48160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_8
timestamp 1698431365
transform 1 0 2240 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_12
timestamp 1698431365
transform 1 0 2688 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_15
timestamp 1698431365
transform 1 0 3024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_19
timestamp 1698431365
transform 1 0 3472 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_23
timestamp 1698431365
transform 1 0 3920 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_169
timestamp 1698431365
transform 1 0 20272 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_173
timestamp 1698431365
transform 1 0 20720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_181
timestamp 1698431365
transform 1 0 21616 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_183
timestamp 1698431365
transform 1 0 21840 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_202
timestamp 1698431365
transform 1 0 23968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_206
timestamp 1698431365
transform 1 0 24416 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_214
timestamp 1698431365
transform 1 0 25312 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_227
timestamp 1698431365
transform 1 0 26768 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_229
timestamp 1698431365
transform 1 0 26992 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_235
timestamp 1698431365
transform 1 0 27664 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_251
timestamp 1698431365
transform 1 0 29456 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_321
timestamp 1698431365
transform 1 0 37296 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_323
timestamp 1698431365
transform 1 0 37520 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_338
timestamp 1698431365
transform 1 0 39200 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_342
timestamp 1698431365
transform 1 0 39648 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_346
timestamp 1698431365
transform 1 0 40096 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_350
timestamp 1698431365
transform 1 0 40544 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_354
timestamp 1698431365
transform 1 0 40992 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_373
timestamp 1698431365
transform 1 0 43120 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_381
timestamp 1698431365
transform 1 0 44016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_405
timestamp 1698431365
transform 1 0 46704 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_413
timestamp 1698431365
transform 1 0 47600 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_417
timestamp 1698431365
transform 1 0 48048 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_419
timestamp 1698431365
transform 1 0 48272 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_6
timestamp 1698431365
transform 1 0 2016 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_17
timestamp 1698431365
transform 1 0 3248 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_24
timestamp 1698431365
transform 1 0 4032 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_26
timestamp 1698431365
transform 1 0 4256 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_67
timestamp 1698431365
transform 1 0 8848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_69
timestamp 1698431365
transform 1 0 9072 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_84
timestamp 1698431365
transform 1 0 10752 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_88
timestamp 1698431365
transform 1 0 11200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_146
timestamp 1698431365
transform 1 0 17696 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_152
timestamp 1698431365
transform 1 0 18368 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_162
timestamp 1698431365
transform 1 0 19488 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_164
timestamp 1698431365
transform 1 0 19712 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_191
timestamp 1698431365
transform 1 0 22736 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_207
timestamp 1698431365
transform 1 0 24528 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_269
timestamp 1698431365
transform 1 0 31472 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_271
timestamp 1698431365
transform 1 0 31696 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_343
timestamp 1698431365
transform 1 0 39760 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_345
timestamp 1698431365
transform 1 0 39984 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_368
timestamp 1698431365
transform 1 0 42560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_372
timestamp 1698431365
transform 1 0 43008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_405
timestamp 1698431365
transform 1 0 46704 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_413
timestamp 1698431365
transform 1 0 47600 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_417
timestamp 1698431365
transform 1 0 48048 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_419
timestamp 1698431365
transform 1 0 48272 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_31
timestamp 1698431365
transform 1 0 4816 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_87
timestamp 1698431365
transform 1 0 11088 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698431365
transform 1 0 12992 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_109
timestamp 1698431365
transform 1 0 13552 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_164
timestamp 1698431365
transform 1 0 19712 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_168
timestamp 1698431365
transform 1 0 20160 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_172
timestamp 1698431365
transform 1 0 20608 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_220
timestamp 1698431365
transform 1 0 25984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_238
timestamp 1698431365
transform 1 0 28000 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_242
timestamp 1698431365
transform 1 0 28448 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_244
timestamp 1698431365
transform 1 0 28672 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_260
timestamp 1698431365
transform 1 0 30464 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_321
timestamp 1698431365
transform 1 0 37296 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_351
timestamp 1698431365
transform 1 0 40656 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_393
timestamp 1698431365
transform 1 0 45360 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_409
timestamp 1698431365
transform 1 0 47152 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_417
timestamp 1698431365
transform 1 0 48048 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_419
timestamp 1698431365
transform 1 0 48272 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_6
timestamp 1698431365
transform 1 0 2016 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_66
timestamp 1698431365
transform 1 0 8736 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_128
timestamp 1698431365
transform 1 0 15680 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_138
timestamp 1698431365
transform 1 0 16800 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_164
timestamp 1698431365
transform 1 0 19712 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_199
timestamp 1698431365
transform 1 0 23632 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_203
timestamp 1698431365
transform 1 0 24080 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_207
timestamp 1698431365
transform 1 0 24528 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_241
timestamp 1698431365
transform 1 0 28336 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_243
timestamp 1698431365
transform 1 0 28560 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_298
timestamp 1698431365
transform 1 0 34720 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_302
timestamp 1698431365
transform 1 0 35168 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_344
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_384
timestamp 1698431365
transform 1 0 44352 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_388
timestamp 1698431365
transform 1 0 44800 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_50
timestamp 1698431365
transform 1 0 6944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_93
timestamp 1698431365
transform 1 0 11760 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_97
timestamp 1698431365
transform 1 0 12208 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_101
timestamp 1698431365
transform 1 0 12656 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_109
timestamp 1698431365
transform 1 0 13552 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_136
timestamp 1698431365
transform 1 0 16576 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_140
timestamp 1698431365
transform 1 0 17024 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_143
timestamp 1698431365
transform 1 0 17360 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_147
timestamp 1698431365
transform 1 0 17808 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_151
timestamp 1698431365
transform 1 0 18256 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_155
timestamp 1698431365
transform 1 0 18704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_181
timestamp 1698431365
transform 1 0 21616 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_185
timestamp 1698431365
transform 1 0 22064 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_189
timestamp 1698431365
transform 1 0 22512 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_205
timestamp 1698431365
transform 1 0 24304 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_213
timestamp 1698431365
transform 1 0 25200 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_217
timestamp 1698431365
transform 1 0 25648 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_219
timestamp 1698431365
transform 1 0 25872 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_222
timestamp 1698431365
transform 1 0 26208 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_226
timestamp 1698431365
transform 1 0 26656 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_238
timestamp 1698431365
transform 1 0 28000 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_242
timestamp 1698431365
transform 1 0 28448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_251
timestamp 1698431365
transform 1 0 29456 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_253
timestamp 1698431365
transform 1 0 29680 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_256
timestamp 1698431365
transform 1 0 30016 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_260
timestamp 1698431365
transform 1 0 30464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_264
timestamp 1698431365
transform 1 0 30912 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_268
timestamp 1698431365
transform 1 0 31360 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_312
timestamp 1698431365
transform 1 0 36288 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_364
timestamp 1698431365
transform 1 0 42112 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_368
timestamp 1698431365
transform 1 0 42560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_372
timestamp 1698431365
transform 1 0 43008 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_380
timestamp 1698431365
transform 1 0 43904 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_384
timestamp 1698431365
transform 1 0 44352 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_419
timestamp 1698431365
transform 1 0 48272 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_68
timestamp 1698431365
transform 1 0 8960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_78
timestamp 1698431365
transform 1 0 10080 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_82
timestamp 1698431365
transform 1 0 10528 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_84
timestamp 1698431365
transform 1 0 10752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_87
timestamp 1698431365
transform 1 0 11088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_91
timestamp 1698431365
transform 1 0 11536 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_95
timestamp 1698431365
transform 1 0 11984 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_146
timestamp 1698431365
transform 1 0 17696 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_216
timestamp 1698431365
transform 1 0 25536 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_232
timestamp 1698431365
transform 1 0 27328 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_240
timestamp 1698431365
transform 1 0 28224 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_244
timestamp 1698431365
transform 1 0 28672 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_247
timestamp 1698431365
transform 1 0 29008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_251
timestamp 1698431365
transform 1 0 29456 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_257
timestamp 1698431365
transform 1 0 30128 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_261
timestamp 1698431365
transform 1 0 30576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_263
timestamp 1698431365
transform 1 0 30800 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_266
timestamp 1698431365
transform 1 0 31136 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_270
timestamp 1698431365
transform 1 0 31584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_274
timestamp 1698431365
transform 1 0 32032 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_278
timestamp 1698431365
transform 1 0 32480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_286
timestamp 1698431365
transform 1 0 33376 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_288
timestamp 1698431365
transform 1 0 33600 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_356
timestamp 1698431365
transform 1 0 41216 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_358
timestamp 1698431365
transform 1 0 41440 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_400
timestamp 1698431365
transform 1 0 46144 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_416
timestamp 1698431365
transform 1 0 47936 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_6
timestamp 1698431365
transform 1 0 2016 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_8
timestamp 1698431365
transform 1 0 2240 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_16
timestamp 1698431365
transform 1 0 3136 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_20
timestamp 1698431365
transform 1 0 3584 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_33
timestamp 1698431365
transform 1 0 5040 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_111
timestamp 1698431365
transform 1 0 13776 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_119
timestamp 1698431365
transform 1 0 14672 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_121
timestamp 1698431365
transform 1 0 14896 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_128
timestamp 1698431365
transform 1 0 15680 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_138
timestamp 1698431365
transform 1 0 16800 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_142
timestamp 1698431365
transform 1 0 17248 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_146
timestamp 1698431365
transform 1 0 17696 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_161
timestamp 1698431365
transform 1 0 19376 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_169
timestamp 1698431365
transform 1 0 20272 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_171
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_174
timestamp 1698431365
transform 1 0 20832 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_181
timestamp 1698431365
transform 1 0 21616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_185
timestamp 1698431365
transform 1 0 22064 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_187
timestamp 1698431365
transform 1 0 22288 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_219
timestamp 1698431365
transform 1 0 25872 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_225
timestamp 1698431365
transform 1 0 26544 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_229
timestamp 1698431365
transform 1 0 26992 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_231
timestamp 1698431365
transform 1 0 27216 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_234
timestamp 1698431365
transform 1 0 27552 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_263
timestamp 1698431365
transform 1 0 30800 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_321
timestamp 1698431365
transform 1 0 37296 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_338
timestamp 1698431365
transform 1 0 39200 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_342
timestamp 1698431365
transform 1 0 39648 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_346
timestamp 1698431365
transform 1 0 40096 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_350
timestamp 1698431365
transform 1 0 40544 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_354
timestamp 1698431365
transform 1 0 40992 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_373
timestamp 1698431365
transform 1 0 43120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_383
timestamp 1698431365
transform 1 0 44240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_419
timestamp 1698431365
transform 1 0 48272 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_6
timestamp 1698431365
transform 1 0 2016 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_8
timestamp 1698431365
transform 1 0 2240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_11
timestamp 1698431365
transform 1 0 2576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_15
timestamp 1698431365
transform 1 0 3024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_17
timestamp 1698431365
transform 1 0 3248 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_68
timestamp 1698431365
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_88
timestamp 1698431365
transform 1 0 11200 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_96
timestamp 1698431365
transform 1 0 12096 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_100
timestamp 1698431365
transform 1 0 12544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_150
timestamp 1698431365
transform 1 0 18144 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_154
timestamp 1698431365
transform 1 0 18592 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_156
timestamp 1698431365
transform 1 0 18816 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_161
timestamp 1698431365
transform 1 0 19376 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_165
timestamp 1698431365
transform 1 0 19824 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_173
timestamp 1698431365
transform 1 0 20720 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_190
timestamp 1698431365
transform 1 0 22624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_206
timestamp 1698431365
transform 1 0 24416 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_223
timestamp 1698431365
transform 1 0 26320 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_272
timestamp 1698431365
transform 1 0 31808 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_276
timestamp 1698431365
transform 1 0 32256 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_291
timestamp 1698431365
transform 1 0 33936 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_295
timestamp 1698431365
transform 1 0 34384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_299
timestamp 1698431365
transform 1 0 34832 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_303
timestamp 1698431365
transform 1 0 35280 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_307
timestamp 1698431365
transform 1 0 35728 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_311
timestamp 1698431365
transform 1 0 36176 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_317
timestamp 1698431365
transform 1 0 36848 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_344
timestamp 1698431365
transform 1 0 39872 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_348
timestamp 1698431365
transform 1 0 40320 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_358
timestamp 1698431365
transform 1 0 41440 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_404
timestamp 1698431365
transform 1 0 46592 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_4
timestamp 1698431365
transform 1 0 1792 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_23
timestamp 1698431365
transform 1 0 3920 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_27
timestamp 1698431365
transform 1 0 4368 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_31
timestamp 1698431365
transform 1 0 4816 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_43
timestamp 1698431365
transform 1 0 6160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_78
timestamp 1698431365
transform 1 0 10080 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_82
timestamp 1698431365
transform 1 0 10528 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_98
timestamp 1698431365
transform 1 0 12320 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_102
timestamp 1698431365
transform 1 0 12768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_104
timestamp 1698431365
transform 1 0 12992 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_125
timestamp 1698431365
transform 1 0 15344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_127
timestamp 1698431365
transform 1 0 15568 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_181
timestamp 1698431365
transform 1 0 21616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_185
timestamp 1698431365
transform 1 0 22064 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_197
timestamp 1698431365
transform 1 0 23408 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_201
timestamp 1698431365
transform 1 0 23856 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_217
timestamp 1698431365
transform 1 0 25648 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_221
timestamp 1698431365
transform 1 0 26096 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_225
timestamp 1698431365
transform 1 0 26544 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_233
timestamp 1698431365
transform 1 0 27440 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_237
timestamp 1698431365
transform 1 0 27888 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_241
timestamp 1698431365
transform 1 0 28336 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_264
timestamp 1698431365
transform 1 0 30912 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_308
timestamp 1698431365
transform 1 0 35840 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_312
timestamp 1698431365
transform 1 0 36288 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_314
timestamp 1698431365
transform 1 0 36512 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_323
timestamp 1698431365
transform 1 0 37520 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_327
timestamp 1698431365
transform 1 0 37968 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_331
timestamp 1698431365
transform 1 0 38416 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_335
timestamp 1698431365
transform 1 0 38864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_337
timestamp 1698431365
transform 1 0 39088 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_367
timestamp 1698431365
transform 1 0 42448 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_371
timestamp 1698431365
transform 1 0 42896 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_375
timestamp 1698431365
transform 1 0 43344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_379
timestamp 1698431365
transform 1 0 43792 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_383
timestamp 1698431365
transform 1 0 44240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_391
timestamp 1698431365
transform 1 0 45136 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_407
timestamp 1698431365
transform 1 0 46928 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_415
timestamp 1698431365
transform 1 0 47824 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_419
timestamp 1698431365
transform 1 0 48272 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_6
timestamp 1698431365
transform 1 0 2016 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_18
timestamp 1698431365
transform 1 0 3360 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_22
timestamp 1698431365
transform 1 0 3808 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_34
timestamp 1698431365
transform 1 0 5152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_69
timestamp 1698431365
transform 1 0 9072 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_85
timestamp 1698431365
transform 1 0 10864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_89
timestamp 1698431365
transform 1 0 11312 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_121
timestamp 1698431365
transform 1 0 14896 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_127
timestamp 1698431365
transform 1 0 15568 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_135
timestamp 1698431365
transform 1 0 16464 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_139
timestamp 1698431365
transform 1 0 16912 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_149
timestamp 1698431365
transform 1 0 18032 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_153
timestamp 1698431365
transform 1 0 18480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_204
timestamp 1698431365
transform 1 0 24192 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_208
timestamp 1698431365
transform 1 0 24640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_216
timestamp 1698431365
transform 1 0 25536 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_218
timestamp 1698431365
transform 1 0 25760 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_231
timestamp 1698431365
transform 1 0 27216 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_241
timestamp 1698431365
transform 1 0 28336 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_245
timestamp 1698431365
transform 1 0 28784 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_249
timestamp 1698431365
transform 1 0 29232 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_253
timestamp 1698431365
transform 1 0 29680 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_256
timestamp 1698431365
transform 1 0 30016 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_260
timestamp 1698431365
transform 1 0 30464 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_286
timestamp 1698431365
transform 1 0 33376 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_288
timestamp 1698431365
transform 1 0 33600 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_295
timestamp 1698431365
transform 1 0 34384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_299
timestamp 1698431365
transform 1 0 34832 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_301
timestamp 1698431365
transform 1 0 35056 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_338
timestamp 1698431365
transform 1 0 39200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_346
timestamp 1698431365
transform 1 0 40096 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_419
timestamp 1698431365
transform 1 0 48272 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_30
timestamp 1698431365
transform 1 0 4704 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_64
timestamp 1698431365
transform 1 0 8512 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_66
timestamp 1698431365
transform 1 0 8736 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_69
timestamp 1698431365
transform 1 0 9072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_95
timestamp 1698431365
transform 1 0 11984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_99
timestamp 1698431365
transform 1 0 12432 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_103
timestamp 1698431365
transform 1 0 12880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_136
timestamp 1698431365
transform 1 0 16576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_140
timestamp 1698431365
transform 1 0 17024 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_148
timestamp 1698431365
transform 1 0 17920 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_152
timestamp 1698431365
transform 1 0 18368 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_155
timestamp 1698431365
transform 1 0 18704 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_159
timestamp 1698431365
transform 1 0 19152 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_161
timestamp 1698431365
transform 1 0 19376 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_164
timestamp 1698431365
transform 1 0 19712 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_168
timestamp 1698431365
transform 1 0 20160 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_172
timestamp 1698431365
transform 1 0 20608 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_174
timestamp 1698431365
transform 1 0 20832 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_181
timestamp 1698431365
transform 1 0 21616 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_183
timestamp 1698431365
transform 1 0 21840 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_190
timestamp 1698431365
transform 1 0 22624 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_198
timestamp 1698431365
transform 1 0 23520 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_204
timestamp 1698431365
transform 1 0 24192 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_240
timestamp 1698431365
transform 1 0 28224 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_242
timestamp 1698431365
transform 1 0 28448 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_299
timestamp 1698431365
transform 1 0 34832 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_303
timestamp 1698431365
transform 1 0 35280 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_346
timestamp 1698431365
transform 1 0 40096 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_350
timestamp 1698431365
transform 1 0 40544 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_367
timestamp 1698431365
transform 1 0 42448 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_376
timestamp 1698431365
transform 1 0 43456 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_384
timestamp 1698431365
transform 1 0 44352 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_419
timestamp 1698431365
transform 1 0 48272 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_4
timestamp 1698431365
transform 1 0 1792 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_7
timestamp 1698431365
transform 1 0 2128 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_11
timestamp 1698431365
transform 1 0 2576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_65
timestamp 1698431365
transform 1 0 8624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_69
timestamp 1698431365
transform 1 0 9072 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_76
timestamp 1698431365
transform 1 0 9856 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_109
timestamp 1698431365
transform 1 0 13552 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_119
timestamp 1698431365
transform 1 0 14672 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_125
timestamp 1698431365
transform 1 0 15344 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_129
timestamp 1698431365
transform 1 0 15792 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_131
timestamp 1698431365
transform 1 0 16016 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_139
timestamp 1698431365
transform 1 0 16912 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_146
timestamp 1698431365
transform 1 0 17696 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_148
timestamp 1698431365
transform 1 0 17920 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_151
timestamp 1698431365
transform 1 0 18256 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_200
timestamp 1698431365
transform 1 0 23744 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_206
timestamp 1698431365
transform 1 0 24416 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_244
timestamp 1698431365
transform 1 0 28672 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_248
timestamp 1698431365
transform 1 0 29120 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_311
timestamp 1698431365
transform 1 0 36176 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_318
timestamp 1698431365
transform 1 0 36960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_322
timestamp 1698431365
transform 1 0 37408 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_326
timestamp 1698431365
transform 1 0 37856 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_328
timestamp 1698431365
transform 1 0 38080 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_337
timestamp 1698431365
transform 1 0 39088 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_341
timestamp 1698431365
transform 1 0 39536 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_345
timestamp 1698431365
transform 1 0 39984 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_348
timestamp 1698431365
transform 1 0 40320 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_369
timestamp 1698431365
transform 1 0 42672 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_373
timestamp 1698431365
transform 1 0 43120 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_377
timestamp 1698431365
transform 1 0 43568 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_409
timestamp 1698431365
transform 1 0 47152 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_417
timestamp 1698431365
transform 1 0 48048 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_419
timestamp 1698431365
transform 1 0 48272 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_32
timestamp 1698431365
transform 1 0 4928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_74
timestamp 1698431365
transform 1 0 9632 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_78
timestamp 1698431365
transform 1 0 10080 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_82
timestamp 1698431365
transform 1 0 10528 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_98
timestamp 1698431365
transform 1 0 12320 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_102
timestamp 1698431365
transform 1 0 12768 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_104
timestamp 1698431365
transform 1 0 12992 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_111
timestamp 1698431365
transform 1 0 13776 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_123
timestamp 1698431365
transform 1 0 15120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_158
timestamp 1698431365
transform 1 0 19040 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_193
timestamp 1698431365
transform 1 0 22960 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_195
timestamp 1698431365
transform 1 0 23184 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_198
timestamp 1698431365
transform 1 0 23520 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_242
timestamp 1698431365
transform 1 0 28448 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_244
timestamp 1698431365
transform 1 0 28672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_251
timestamp 1698431365
transform 1 0 29456 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_263
timestamp 1698431365
transform 1 0 30800 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_267
timestamp 1698431365
transform 1 0 31248 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_271
timestamp 1698431365
transform 1 0 31696 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_273
timestamp 1698431365
transform 1 0 31920 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_310
timestamp 1698431365
transform 1 0 36064 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_314
timestamp 1698431365
transform 1 0 36512 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_321
timestamp 1698431365
transform 1 0 37296 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_325
timestamp 1698431365
transform 1 0 37744 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_327
timestamp 1698431365
transform 1 0 37968 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_357
timestamp 1698431365
transform 1 0 41328 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_362
timestamp 1698431365
transform 1 0 41888 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_366
timestamp 1698431365
transform 1 0 42336 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_370
timestamp 1698431365
transform 1 0 42784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_374
timestamp 1698431365
transform 1 0 43232 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_382
timestamp 1698431365
transform 1 0 44128 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_384
timestamp 1698431365
transform 1 0 44352 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_391
timestamp 1698431365
transform 1 0 45136 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_407
timestamp 1698431365
transform 1 0 46928 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_415
timestamp 1698431365
transform 1 0 47824 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_419
timestamp 1698431365
transform 1 0 48272 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_33
timestamp 1698431365
transform 1 0 5040 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_37
timestamp 1698431365
transform 1 0 5488 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_41
timestamp 1698431365
transform 1 0 5936 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_69
timestamp 1698431365
transform 1 0 9072 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_85
timestamp 1698431365
transform 1 0 10864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_89
timestamp 1698431365
transform 1 0 11312 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_97
timestamp 1698431365
transform 1 0 12208 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_130
timestamp 1698431365
transform 1 0 15904 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_134
timestamp 1698431365
transform 1 0 16352 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_138
timestamp 1698431365
transform 1 0 16800 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_158
timestamp 1698431365
transform 1 0 19040 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_174
timestamp 1698431365
transform 1 0 20832 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_178
timestamp 1698431365
transform 1 0 21280 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_182
timestamp 1698431365
transform 1 0 21728 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_190
timestamp 1698431365
transform 1 0 22624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_192
timestamp 1698431365
transform 1 0 22848 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_201
timestamp 1698431365
transform 1 0 23856 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_205
timestamp 1698431365
transform 1 0 24304 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_209
timestamp 1698431365
transform 1 0 24752 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_245
timestamp 1698431365
transform 1 0 28784 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_247
timestamp 1698431365
transform 1 0 29008 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_271
timestamp 1698431365
transform 1 0 31696 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_275
timestamp 1698431365
transform 1 0 32144 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_279
timestamp 1698431365
transform 1 0 32592 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_308
timestamp 1698431365
transform 1 0 35840 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_312
timestamp 1698431365
transform 1 0 36288 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_316
timestamp 1698431365
transform 1 0 36736 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_348
timestamp 1698431365
transform 1 0 40320 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_356
timestamp 1698431365
transform 1 0 41216 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_358
timestamp 1698431365
transform 1 0 41440 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_394
timestamp 1698431365
transform 1 0 45472 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_410
timestamp 1698431365
transform 1 0 47264 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_418
timestamp 1698431365
transform 1 0 48160 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_2
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_18
timestamp 1698431365
transform 1 0 3360 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_29
timestamp 1698431365
transform 1 0 4592 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_33
timestamp 1698431365
transform 1 0 5040 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_41
timestamp 1698431365
transform 1 0 5936 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_44
timestamp 1698431365
transform 1 0 6272 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_54
timestamp 1698431365
transform 1 0 7392 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_56
timestamp 1698431365
transform 1 0 7616 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_88
timestamp 1698431365
transform 1 0 11200 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_92
timestamp 1698431365
transform 1 0 11648 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_100
timestamp 1698431365
transform 1 0 12544 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_103
timestamp 1698431365
transform 1 0 12880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_119
timestamp 1698431365
transform 1 0 14672 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_123
timestamp 1698431365
transform 1 0 15120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_125
timestamp 1698431365
transform 1 0 15344 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_157
timestamp 1698431365
transform 1 0 18928 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_173
timestamp 1698431365
transform 1 0 20720 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_185
timestamp 1698431365
transform 1 0 22064 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_220
timestamp 1698431365
transform 1 0 25984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_238
timestamp 1698431365
transform 1 0 28000 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_242
timestamp 1698431365
transform 1 0 28448 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_244
timestamp 1698431365
transform 1 0 28672 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_295
timestamp 1698431365
transform 1 0 34384 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_305
timestamp 1698431365
transform 1 0 35504 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_309
timestamp 1698431365
transform 1 0 35952 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_313
timestamp 1698431365
transform 1 0 36400 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_321
timestamp 1698431365
transform 1 0 37296 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_323
timestamp 1698431365
transform 1 0 37520 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_326
timestamp 1698431365
transform 1 0 37856 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_342
timestamp 1698431365
transform 1 0 39648 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_350
timestamp 1698431365
transform 1 0 40544 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_354
timestamp 1698431365
transform 1 0 40992 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_356
timestamp 1698431365
transform 1 0 41216 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_359
timestamp 1698431365
transform 1 0 41552 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_365
timestamp 1698431365
transform 1 0 42224 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_381
timestamp 1698431365
transform 1 0 44016 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_419
timestamp 1698431365
transform 1 0 48272 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_10
timestamp 1698431365
transform 1 0 2464 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_14
timestamp 1698431365
transform 1 0 2912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_16
timestamp 1698431365
transform 1 0 3136 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_19
timestamp 1698431365
transform 1 0 3472 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_23
timestamp 1698431365
transform 1 0 3920 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_45
timestamp 1698431365
transform 1 0 6384 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_61
timestamp 1698431365
transform 1 0 8176 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_65
timestamp 1698431365
transform 1 0 8624 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_69
timestamp 1698431365
transform 1 0 9072 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_121
timestamp 1698431365
transform 1 0 14896 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_137
timestamp 1698431365
transform 1 0 16688 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_139
timestamp 1698431365
transform 1 0 16912 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_158
timestamp 1698431365
transform 1 0 19040 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_201
timestamp 1698431365
transform 1 0 23856 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_209
timestamp 1698431365
transform 1 0 24752 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_220
timestamp 1698431365
transform 1 0 25984 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_230
timestamp 1698431365
transform 1 0 27104 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_246
timestamp 1698431365
transform 1 0 28896 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_256
timestamp 1698431365
transform 1 0 30016 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_260
timestamp 1698431365
transform 1 0 30464 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_264
timestamp 1698431365
transform 1 0 30912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_266
timestamp 1698431365
transform 1 0 31136 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_269
timestamp 1698431365
transform 1 0 31472 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_273
timestamp 1698431365
transform 1 0 31920 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_277
timestamp 1698431365
transform 1 0 32368 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_279
timestamp 1698431365
transform 1 0 32592 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_311
timestamp 1698431365
transform 1 0 36176 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_342
timestamp 1698431365
transform 1 0 39648 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_346
timestamp 1698431365
transform 1 0 40096 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_376
timestamp 1698431365
transform 1 0 43456 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_380
timestamp 1698431365
transform 1 0 43904 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_384
timestamp 1698431365
transform 1 0 44352 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_416
timestamp 1698431365
transform 1 0 47936 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_6
timestamp 1698431365
transform 1 0 2016 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_10
timestamp 1698431365
transform 1 0 2464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_14
timestamp 1698431365
transform 1 0 2912 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_32
timestamp 1698431365
transform 1 0 4928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_92
timestamp 1698431365
transform 1 0 11648 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_96
timestamp 1698431365
transform 1 0 12096 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_104
timestamp 1698431365
transform 1 0 12992 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_171
timestamp 1698431365
transform 1 0 20496 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_185
timestamp 1698431365
transform 1 0 22064 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_193
timestamp 1698431365
transform 1 0 22960 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_197
timestamp 1698431365
transform 1 0 23408 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_229
timestamp 1698431365
transform 1 0 26992 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_255
timestamp 1698431365
transform 1 0 29904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_259
timestamp 1698431365
transform 1 0 30352 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_261
timestamp 1698431365
transform 1 0 30576 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_264
timestamp 1698431365
transform 1 0 30912 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_268
timestamp 1698431365
transform 1 0 31360 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_274
timestamp 1698431365
transform 1 0 32032 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_278
timestamp 1698431365
transform 1 0 32480 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_282
timestamp 1698431365
transform 1 0 32928 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_286
timestamp 1698431365
transform 1 0 33376 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_289
timestamp 1698431365
transform 1 0 33712 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_293
timestamp 1698431365
transform 1 0 34160 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_297
timestamp 1698431365
transform 1 0 34608 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_311
timestamp 1698431365
transform 1 0 36176 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_319
timestamp 1698431365
transform 1 0 37072 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_349
timestamp 1698431365
transform 1 0 40432 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_374
timestamp 1698431365
transform 1 0 43232 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_382
timestamp 1698431365
transform 1 0 44128 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_384
timestamp 1698431365
transform 1 0 44352 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_393
timestamp 1698431365
transform 1 0 45360 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_409
timestamp 1698431365
transform 1 0 47152 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_417
timestamp 1698431365
transform 1 0 48048 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_419
timestamp 1698431365
transform 1 0 48272 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_2
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_6
timestamp 1698431365
transform 1 0 2016 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_9
timestamp 1698431365
transform 1 0 2352 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_31
timestamp 1698431365
transform 1 0 4816 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_57
timestamp 1698431365
transform 1 0 7728 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_61
timestamp 1698431365
transform 1 0 8176 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_65
timestamp 1698431365
transform 1 0 8624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_69
timestamp 1698431365
transform 1 0 9072 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_80
timestamp 1698431365
transform 1 0 10304 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_84
timestamp 1698431365
transform 1 0 10752 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_115
timestamp 1698431365
transform 1 0 14224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_119
timestamp 1698431365
transform 1 0 14672 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_123
timestamp 1698431365
transform 1 0 15120 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_139
timestamp 1698431365
transform 1 0 16912 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_174
timestamp 1698431365
transform 1 0 20832 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_190
timestamp 1698431365
transform 1 0 22624 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_193
timestamp 1698431365
transform 1 0 22960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_204
timestamp 1698431365
transform 1 0 24192 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_270
timestamp 1698431365
transform 1 0 31584 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_279
timestamp 1698431365
transform 1 0 32592 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_286
timestamp 1698431365
transform 1 0 33376 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_290
timestamp 1698431365
transform 1 0 33824 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_298
timestamp 1698431365
transform 1 0 34720 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_302
timestamp 1698431365
transform 1 0 35168 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_333
timestamp 1698431365
transform 1 0 38640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_337
timestamp 1698431365
transform 1 0 39088 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_345
timestamp 1698431365
transform 1 0 39984 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_349
timestamp 1698431365
transform 1 0 40432 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_352
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_356
timestamp 1698431365
transform 1 0 41216 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_360
timestamp 1698431365
transform 1 0 41664 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_364
timestamp 1698431365
transform 1 0 42112 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_368
timestamp 1698431365
transform 1 0 42560 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_401
timestamp 1698431365
transform 1 0 46256 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_417
timestamp 1698431365
transform 1 0 48048 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_419
timestamp 1698431365
transform 1 0 48272 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_18
timestamp 1698431365
transform 1 0 3360 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_42
timestamp 1698431365
transform 1 0 6048 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_66
timestamp 1698431365
transform 1 0 8736 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_70
timestamp 1698431365
transform 1 0 9184 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_74
timestamp 1698431365
transform 1 0 9632 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_90
timestamp 1698431365
transform 1 0 11424 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_94
timestamp 1698431365
transform 1 0 11872 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_103
timestamp 1698431365
transform 1 0 12880 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_127
timestamp 1698431365
transform 1 0 15568 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_129
timestamp 1698431365
transform 1 0 15792 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_161
timestamp 1698431365
transform 1 0 19376 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_171
timestamp 1698431365
transform 1 0 20496 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_185
timestamp 1698431365
transform 1 0 22064 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_241
timestamp 1698431365
transform 1 0 28336 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_255
timestamp 1698431365
transform 1 0 29904 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_285
timestamp 1698431365
transform 1 0 33264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_295
timestamp 1698431365
transform 1 0 34384 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_299
timestamp 1698431365
transform 1 0 34832 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_307
timestamp 1698431365
transform 1 0 35728 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_314
timestamp 1698431365
transform 1 0 36512 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_325
timestamp 1698431365
transform 1 0 37744 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_329
timestamp 1698431365
transform 1 0 38192 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_335
timestamp 1698431365
transform 1 0 38864 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_343
timestamp 1698431365
transform 1 0 39760 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_345
timestamp 1698431365
transform 1 0 39984 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_371
timestamp 1698431365
transform 1 0 42896 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_375
timestamp 1698431365
transform 1 0 43344 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_383
timestamp 1698431365
transform 1 0 44240 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_419
timestamp 1698431365
transform 1 0 48272 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_69
timestamp 1698431365
transform 1 0 9072 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_104
timestamp 1698431365
transform 1 0 12992 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_107
timestamp 1698431365
transform 1 0 13328 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_138
timestamp 1698431365
transform 1 0 16800 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_148
timestamp 1698431365
transform 1 0 17920 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_152
timestamp 1698431365
transform 1 0 18368 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_158
timestamp 1698431365
transform 1 0 19040 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_169
timestamp 1698431365
transform 1 0 20272 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_199
timestamp 1698431365
transform 1 0 23632 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_205
timestamp 1698431365
transform 1 0 24304 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_209
timestamp 1698431365
transform 1 0 24752 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_217
timestamp 1698431365
transform 1 0 25648 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_221
timestamp 1698431365
transform 1 0 26096 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_229
timestamp 1698431365
transform 1 0 26992 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_233
timestamp 1698431365
transform 1 0 27440 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_251
timestamp 1698431365
transform 1 0 29456 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_255
timestamp 1698431365
transform 1 0 29904 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_262
timestamp 1698431365
transform 1 0 30688 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_278
timestamp 1698431365
transform 1 0 32480 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_286
timestamp 1698431365
transform 1 0 33376 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_290
timestamp 1698431365
transform 1 0 33824 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_304
timestamp 1698431365
transform 1 0 35392 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_320
timestamp 1698431365
transform 1 0 37184 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_328
timestamp 1698431365
transform 1 0 38080 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_338
timestamp 1698431365
transform 1 0 39200 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_346
timestamp 1698431365
transform 1 0 40096 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_352
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_385
timestamp 1698431365
transform 1 0 44464 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_417
timestamp 1698431365
transform 1 0 48048 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_419
timestamp 1698431365
transform 1 0 48272 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_4
timestamp 1698431365
transform 1 0 1792 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_7
timestamp 1698431365
transform 1 0 2128 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_11
timestamp 1698431365
transform 1 0 2576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_15
timestamp 1698431365
transform 1 0 3024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_19
timestamp 1698431365
transform 1 0 3472 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_23
timestamp 1698431365
transform 1 0 3920 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_27
timestamp 1698431365
transform 1 0 4368 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_31
timestamp 1698431365
transform 1 0 4816 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_45
timestamp 1698431365
transform 1 0 6384 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_70
timestamp 1698431365
transform 1 0 9184 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_102
timestamp 1698431365
transform 1 0 12768 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_104
timestamp 1698431365
transform 1 0 12992 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_123
timestamp 1698431365
transform 1 0 15120 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_131
timestamp 1698431365
transform 1 0 16016 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_135
timestamp 1698431365
transform 1 0 16464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_137
timestamp 1698431365
transform 1 0 16688 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_142
timestamp 1698431365
transform 1 0 17248 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_151
timestamp 1698431365
transform 1 0 18256 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_155
timestamp 1698431365
transform 1 0 18704 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_159
timestamp 1698431365
transform 1 0 19152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_183
timestamp 1698431365
transform 1 0 21840 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_187
timestamp 1698431365
transform 1 0 22288 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_227
timestamp 1698431365
transform 1 0 26768 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_243
timestamp 1698431365
transform 1 0 28560 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_263
timestamp 1698431365
transform 1 0 30800 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_271
timestamp 1698431365
transform 1 0 31696 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_275
timestamp 1698431365
transform 1 0 32144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_308
timestamp 1698431365
transform 1 0 35840 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_312
timestamp 1698431365
transform 1 0 36288 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_314
timestamp 1698431365
transform 1 0 36512 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_325
timestamp 1698431365
transform 1 0 37744 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_368
timestamp 1698431365
transform 1 0 42560 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_372
timestamp 1698431365
transform 1 0 43008 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_380
timestamp 1698431365
transform 1 0 43904 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_384
timestamp 1698431365
transform 1 0 44352 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_419
timestamp 1698431365
transform 1 0 48272 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_6
timestamp 1698431365
transform 1 0 2016 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_57
timestamp 1698431365
transform 1 0 7728 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_61
timestamp 1698431365
transform 1 0 8176 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_69
timestamp 1698431365
transform 1 0 9072 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_76
timestamp 1698431365
transform 1 0 9856 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_142
timestamp 1698431365
transform 1 0 17248 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_174
timestamp 1698431365
transform 1 0 20832 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_177
timestamp 1698431365
transform 1 0 21168 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_179
timestamp 1698431365
transform 1 0 21392 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_203
timestamp 1698431365
transform 1 0 24080 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_207
timestamp 1698431365
transform 1 0 24528 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_241
timestamp 1698431365
transform 1 0 28336 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_273
timestamp 1698431365
transform 1 0 31920 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_277
timestamp 1698431365
transform 1 0 32368 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_279
timestamp 1698431365
transform 1 0 32592 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_282
timestamp 1698431365
transform 1 0 32928 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_284
timestamp 1698431365
transform 1 0 33152 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_291
timestamp 1698431365
transform 1 0 33936 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_299
timestamp 1698431365
transform 1 0 34832 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_301
timestamp 1698431365
transform 1 0 35056 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_331
timestamp 1698431365
transform 1 0 38416 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_335
timestamp 1698431365
transform 1 0 38864 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_343
timestamp 1698431365
transform 1 0 39760 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_347
timestamp 1698431365
transform 1 0 40208 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_349
timestamp 1698431365
transform 1 0 40432 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_352
timestamp 1698431365
transform 1 0 40768 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_358
timestamp 1698431365
transform 1 0 41440 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_365
timestamp 1698431365
transform 1 0 42224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_369
timestamp 1698431365
transform 1 0 42672 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_401
timestamp 1698431365
transform 1 0 46256 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_417
timestamp 1698431365
transform 1 0 48048 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_419
timestamp 1698431365
transform 1 0 48272 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_2
timestamp 1698431365
transform 1 0 1568 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_6
timestamp 1698431365
transform 1 0 2016 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_9
timestamp 1698431365
transform 1 0 2352 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_21
timestamp 1698431365
transform 1 0 3696 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_27
timestamp 1698431365
transform 1 0 4368 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_37
timestamp 1698431365
transform 1 0 5488 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_99
timestamp 1698431365
transform 1 0 12432 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_103
timestamp 1698431365
transform 1 0 12880 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_107
timestamp 1698431365
transform 1 0 13328 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_139
timestamp 1698431365
transform 1 0 16912 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_147
timestamp 1698431365
transform 1 0 17808 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_149
timestamp 1698431365
transform 1 0 18032 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_152
timestamp 1698431365
transform 1 0 18368 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_154
timestamp 1698431365
transform 1 0 18592 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_172
timestamp 1698431365
transform 1 0 20608 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_174
timestamp 1698431365
transform 1 0 20832 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_220
timestamp 1698431365
transform 1 0 25984 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_224
timestamp 1698431365
transform 1 0 26432 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_240
timestamp 1698431365
transform 1 0 28224 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_244
timestamp 1698431365
transform 1 0 28672 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_247
timestamp 1698431365
transform 1 0 29008 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_251
timestamp 1698431365
transform 1 0 29456 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_259
timestamp 1698431365
transform 1 0 30352 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_261
timestamp 1698431365
transform 1 0 30576 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_298
timestamp 1698431365
transform 1 0 34720 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_302
timestamp 1698431365
transform 1 0 35168 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_310
timestamp 1698431365
transform 1 0 36064 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_314
timestamp 1698431365
transform 1 0 36512 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_317
timestamp 1698431365
transform 1 0 36848 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_325
timestamp 1698431365
transform 1 0 37744 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_329
timestamp 1698431365
transform 1 0 38192 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_334
timestamp 1698431365
transform 1 0 38752 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_350
timestamp 1698431365
transform 1 0 40544 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_387
timestamp 1698431365
transform 1 0 44688 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_419
timestamp 1698431365
transform 1 0 48272 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_2
timestamp 1698431365
transform 1 0 1568 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_40
timestamp 1698431365
transform 1 0 5824 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_44
timestamp 1698431365
transform 1 0 6272 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_72
timestamp 1698431365
transform 1 0 9408 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_80
timestamp 1698431365
transform 1 0 10304 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_99
timestamp 1698431365
transform 1 0 12432 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_118
timestamp 1698431365
transform 1 0 14560 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_134
timestamp 1698431365
transform 1 0 16352 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_138
timestamp 1698431365
transform 1 0 16800 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_209
timestamp 1698431365
transform 1 0 24752 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_235
timestamp 1698431365
transform 1 0 27664 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_239
timestamp 1698431365
transform 1 0 28112 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_241
timestamp 1698431365
transform 1 0 28336 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_282
timestamp 1698431365
transform 1 0 32928 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_286
timestamp 1698431365
transform 1 0 33376 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_290
timestamp 1698431365
transform 1 0 33824 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_294
timestamp 1698431365
transform 1 0 34272 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_298
timestamp 1698431365
transform 1 0 34720 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_308
timestamp 1698431365
transform 1 0 35840 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_312
timestamp 1698431365
transform 1 0 36288 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_336
timestamp 1698431365
transform 1 0 38976 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_344
timestamp 1698431365
transform 1 0 39872 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_348
timestamp 1698431365
transform 1 0 40320 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_352
timestamp 1698431365
transform 1 0 40768 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_416
timestamp 1698431365
transform 1 0 47936 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_31
timestamp 1698431365
transform 1 0 4816 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_50
timestamp 1698431365
transform 1 0 6944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_54
timestamp 1698431365
transform 1 0 7392 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_70
timestamp 1698431365
transform 1 0 9184 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_78
timestamp 1698431365
transform 1 0 10080 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_99
timestamp 1698431365
transform 1 0 12432 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_103
timestamp 1698431365
transform 1 0 12880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_124
timestamp 1698431365
transform 1 0 15232 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_154
timestamp 1698431365
transform 1 0 18592 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_162
timestamp 1698431365
transform 1 0 19488 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_166
timestamp 1698431365
transform 1 0 19936 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_170
timestamp 1698431365
transform 1 0 20384 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_174
timestamp 1698431365
transform 1 0 20832 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_177
timestamp 1698431365
transform 1 0 21168 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_185
timestamp 1698431365
transform 1 0 22064 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_189
timestamp 1698431365
transform 1 0 22512 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_191
timestamp 1698431365
transform 1 0 22736 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_215
timestamp 1698431365
transform 1 0 25424 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_219
timestamp 1698431365
transform 1 0 25872 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_223
timestamp 1698431365
transform 1 0 26320 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_227
timestamp 1698431365
transform 1 0 26768 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_229
timestamp 1698431365
transform 1 0 26992 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_240
timestamp 1698431365
transform 1 0 28224 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_244
timestamp 1698431365
transform 1 0 28672 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_255
timestamp 1698431365
transform 1 0 29904 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_259
timestamp 1698431365
transform 1 0 30352 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_261
timestamp 1698431365
transform 1 0 30576 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_291
timestamp 1698431365
transform 1 0 33936 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_295
timestamp 1698431365
transform 1 0 34384 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_303
timestamp 1698431365
transform 1 0 35280 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_310
timestamp 1698431365
transform 1 0 36064 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_314
timestamp 1698431365
transform 1 0 36512 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_317
timestamp 1698431365
transform 1 0 36848 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_321
timestamp 1698431365
transform 1 0 37296 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_357
timestamp 1698431365
transform 1 0 41328 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_373
timestamp 1698431365
transform 1 0 43120 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_381
timestamp 1698431365
transform 1 0 44016 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_387
timestamp 1698431365
transform 1 0 44688 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_419
timestamp 1698431365
transform 1 0 48272 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_2
timestamp 1698431365
transform 1 0 1568 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_6
timestamp 1698431365
transform 1 0 2016 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_13
timestamp 1698431365
transform 1 0 2800 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_21
timestamp 1698431365
transform 1 0 3696 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_27
timestamp 1698431365
transform 1 0 4368 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_31
timestamp 1698431365
transform 1 0 4816 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_37
timestamp 1698431365
transform 1 0 5488 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_39
timestamp 1698431365
transform 1 0 5712 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_50
timestamp 1698431365
transform 1 0 6944 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_66
timestamp 1698431365
transform 1 0 8736 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_72
timestamp 1698431365
transform 1 0 9408 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_80
timestamp 1698431365
transform 1 0 10304 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_99
timestamp 1698431365
transform 1 0 12432 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_118
timestamp 1698431365
transform 1 0 14560 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_136
timestamp 1698431365
transform 1 0 16576 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_154
timestamp 1698431365
transform 1 0 18592 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_158
timestamp 1698431365
transform 1 0 19040 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_164
timestamp 1698431365
transform 1 0 19712 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_172
timestamp 1698431365
transform 1 0 20608 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_176
timestamp 1698431365
transform 1 0 21056 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_178
timestamp 1698431365
transform 1 0 21280 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_202
timestamp 1698431365
transform 1 0 23968 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_206
timestamp 1698431365
transform 1 0 24416 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_212
timestamp 1698431365
transform 1 0 25088 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_216
timestamp 1698431365
transform 1 0 25536 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_251
timestamp 1698431365
transform 1 0 29456 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_263
timestamp 1698431365
transform 1 0 30800 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_267
timestamp 1698431365
transform 1 0 31248 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_275
timestamp 1698431365
transform 1 0 32144 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_279
timestamp 1698431365
transform 1 0 32592 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_288
timestamp 1698431365
transform 1 0 33600 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_296
timestamp 1698431365
transform 1 0 34496 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_328
timestamp 1698431365
transform 1 0 38080 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_344
timestamp 1698431365
transform 1 0 39872 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_348
timestamp 1698431365
transform 1 0 40320 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_352
timestamp 1698431365
transform 1 0 40768 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_416
timestamp 1698431365
transform 1 0 47936 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_2
timestamp 1698431365
transform 1 0 1568 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_34
timestamp 1698431365
transform 1 0 5152 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_37
timestamp 1698431365
transform 1 0 5488 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_45
timestamp 1698431365
transform 1 0 6384 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_53
timestamp 1698431365
transform 1 0 7280 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_58
timestamp 1698431365
transform 1 0 7840 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_90
timestamp 1698431365
transform 1 0 11424 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_98
timestamp 1698431365
transform 1 0 12320 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_102
timestamp 1698431365
transform 1 0 12768 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_104
timestamp 1698431365
transform 1 0 12992 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_107
timestamp 1698431365
transform 1 0 13328 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_115
timestamp 1698431365
transform 1 0 14224 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_119
timestamp 1698431365
transform 1 0 14672 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_149
timestamp 1698431365
transform 1 0 18032 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_153
timestamp 1698431365
transform 1 0 18480 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_169
timestamp 1698431365
transform 1 0 20272 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_173
timestamp 1698431365
transform 1 0 20720 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_177
timestamp 1698431365
transform 1 0 21168 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_179
timestamp 1698431365
transform 1 0 21392 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_185
timestamp 1698431365
transform 1 0 22064 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_189
timestamp 1698431365
transform 1 0 22512 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_197
timestamp 1698431365
transform 1 0 23408 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_203
timestamp 1698431365
transform 1 0 24080 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_207
timestamp 1698431365
transform 1 0 24528 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_209
timestamp 1698431365
transform 1 0 24752 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_212
timestamp 1698431365
transform 1 0 25088 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_220
timestamp 1698431365
transform 1 0 25984 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_237
timestamp 1698431365
transform 1 0 27888 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_247
timestamp 1698431365
transform 1 0 29008 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_255
timestamp 1698431365
transform 1 0 29904 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_259
timestamp 1698431365
transform 1 0 30352 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_261
timestamp 1698431365
transform 1 0 30576 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_278
timestamp 1698431365
transform 1 0 32480 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_282
timestamp 1698431365
transform 1 0 32928 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_314
timestamp 1698431365
transform 1 0 36512 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_317
timestamp 1698431365
transform 1 0 36848 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_333
timestamp 1698431365
transform 1 0 38640 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_341
timestamp 1698431365
transform 1 0 39536 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_345
timestamp 1698431365
transform 1 0 39984 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_348
timestamp 1698431365
transform 1 0 40320 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_358
timestamp 1698431365
transform 1 0 41440 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_362
timestamp 1698431365
transform 1 0 41888 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_372
timestamp 1698431365
transform 1 0 43008 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_380
timestamp 1698431365
transform 1 0 43904 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_384
timestamp 1698431365
transform 1 0 44352 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_387
timestamp 1698431365
transform 1 0 44688 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_419
timestamp 1698431365
transform 1 0 48272 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_2
timestamp 1698431365
transform 1 0 1568 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_18
timestamp 1698431365
transform 1 0 3360 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_24
timestamp 1698431365
transform 1 0 4032 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_32
timestamp 1698431365
transform 1 0 4928 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_35
timestamp 1698431365
transform 1 0 5264 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_51
timestamp 1698431365
transform 1 0 7056 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_72
timestamp 1698431365
transform 1 0 9408 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_104
timestamp 1698431365
transform 1 0 12992 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_120
timestamp 1698431365
transform 1 0 14784 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_138
timestamp 1698431365
transform 1 0 16800 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_142
timestamp 1698431365
transform 1 0 17248 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_158
timestamp 1698431365
transform 1 0 19040 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_160
timestamp 1698431365
transform 1 0 19264 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_169
timestamp 1698431365
transform 1 0 20272 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_171
timestamp 1698431365
transform 1 0 20496 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_203
timestamp 1698431365
transform 1 0 24080 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_241
timestamp 1698431365
transform 1 0 28336 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_273
timestamp 1698431365
transform 1 0 31920 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_311
timestamp 1698431365
transform 1 0 36176 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_327
timestamp 1698431365
transform 1 0 37968 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_335
timestamp 1698431365
transform 1 0 38864 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_339
timestamp 1698431365
transform 1 0 39312 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_341
timestamp 1698431365
transform 1 0 39536 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_381
timestamp 1698431365
transform 1 0 44016 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_413
timestamp 1698431365
transform 1 0 47600 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_417
timestamp 1698431365
transform 1 0 48048 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_419
timestamp 1698431365
transform 1 0 48272 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_2
timestamp 1698431365
transform 1 0 1568 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_33
timestamp 1698431365
transform 1 0 5040 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_43
timestamp 1698431365
transform 1 0 6160 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_51
timestamp 1698431365
transform 1 0 7056 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_53
timestamp 1698431365
transform 1 0 7280 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_88
timestamp 1698431365
transform 1 0 11200 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_104
timestamp 1698431365
transform 1 0 12992 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_124
timestamp 1698431365
transform 1 0 15232 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_140
timestamp 1698431365
transform 1 0 17024 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_177
timestamp 1698431365
transform 1 0 21168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_179
timestamp 1698431365
transform 1 0 21392 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_184
timestamp 1698431365
transform 1 0 21952 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_188
timestamp 1698431365
transform 1 0 22400 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_225
timestamp 1698431365
transform 1 0 26544 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_241
timestamp 1698431365
transform 1 0 28336 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_247
timestamp 1698431365
transform 1 0 29008 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_251
timestamp 1698431365
transform 1 0 29456 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_258
timestamp 1698431365
transform 1 0 30240 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_274
timestamp 1698431365
transform 1 0 32032 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_286
timestamp 1698431365
transform 1 0 33376 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_290
timestamp 1698431365
transform 1 0 33824 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_306
timestamp 1698431365
transform 1 0 35616 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_314
timestamp 1698431365
transform 1 0 36512 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_317
timestamp 1698431365
transform 1 0 36848 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_324
timestamp 1698431365
transform 1 0 37632 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_340
timestamp 1698431365
transform 1 0 39424 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_372
timestamp 1698431365
transform 1 0 43008 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_380
timestamp 1698431365
transform 1 0 43904 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_384
timestamp 1698431365
transform 1 0 44352 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_387
timestamp 1698431365
transform 1 0 44688 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_419
timestamp 1698431365
transform 1 0 48272 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_2
timestamp 1698431365
transform 1 0 1568 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_55
timestamp 1698431365
transform 1 0 7504 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_63
timestamp 1698431365
transform 1 0 8400 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_67
timestamp 1698431365
transform 1 0 8848 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_69
timestamp 1698431365
transform 1 0 9072 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_72
timestamp 1698431365
transform 1 0 9408 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_76
timestamp 1698431365
transform 1 0 9856 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_95
timestamp 1698431365
transform 1 0 11984 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_120
timestamp 1698431365
transform 1 0 14784 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_136
timestamp 1698431365
transform 1 0 16576 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_142
timestamp 1698431365
transform 1 0 17248 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_144
timestamp 1698431365
transform 1 0 17472 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_151
timestamp 1698431365
transform 1 0 18256 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_155
timestamp 1698431365
transform 1 0 18704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_159
timestamp 1698431365
transform 1 0 19152 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_161
timestamp 1698431365
transform 1 0 19376 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_166
timestamp 1698431365
transform 1 0 19936 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_182
timestamp 1698431365
transform 1 0 21728 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_190
timestamp 1698431365
transform 1 0 22624 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_194
timestamp 1698431365
transform 1 0 23072 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_203
timestamp 1698431365
transform 1 0 24080 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_207
timestamp 1698431365
transform 1 0 24528 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_209
timestamp 1698431365
transform 1 0 24752 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_212
timestamp 1698431365
transform 1 0 25088 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_228
timestamp 1698431365
transform 1 0 26880 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_236
timestamp 1698431365
transform 1 0 27776 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_269
timestamp 1698431365
transform 1 0 31472 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_273
timestamp 1698431365
transform 1 0 31920 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_277
timestamp 1698431365
transform 1 0 32368 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_279
timestamp 1698431365
transform 1 0 32592 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_282
timestamp 1698431365
transform 1 0 32928 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_298
timestamp 1698431365
transform 1 0 34720 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_306
timestamp 1698431365
transform 1 0 35616 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_308
timestamp 1698431365
transform 1 0 35840 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_340
timestamp 1698431365
transform 1 0 39424 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_348
timestamp 1698431365
transform 1 0 40320 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_352
timestamp 1698431365
transform 1 0 40768 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_416
timestamp 1698431365
transform 1 0 47936 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_2
timestamp 1698431365
transform 1 0 1568 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_6
timestamp 1698431365
transform 1 0 2016 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_14
timestamp 1698431365
transform 1 0 2912 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_22
timestamp 1698431365
transform 1 0 3808 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_26
timestamp 1698431365
transform 1 0 4256 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_30
timestamp 1698431365
transform 1 0 4704 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_34
timestamp 1698431365
transform 1 0 5152 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_77
timestamp 1698431365
transform 1 0 9968 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_93
timestamp 1698431365
transform 1 0 11760 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_101
timestamp 1698431365
transform 1 0 12656 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_124
timestamp 1698431365
transform 1 0 15232 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_161
timestamp 1698431365
transform 1 0 19376 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_165
timestamp 1698431365
transform 1 0 19824 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_173
timestamp 1698431365
transform 1 0 20720 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_177
timestamp 1698431365
transform 1 0 21168 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_241
timestamp 1698431365
transform 1 0 28336 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_247
timestamp 1698431365
transform 1 0 29008 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_263
timestamp 1698431365
transform 1 0 30800 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_267
timestamp 1698431365
transform 1 0 31248 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_271
timestamp 1698431365
transform 1 0 31696 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_325
timestamp 1698431365
transform 1 0 37744 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_329
timestamp 1698431365
transform 1 0 38192 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_336
timestamp 1698431365
transform 1 0 38976 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_340
timestamp 1698431365
transform 1 0 39424 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_372
timestamp 1698431365
transform 1 0 43008 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_380
timestamp 1698431365
transform 1 0 43904 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_384
timestamp 1698431365
transform 1 0 44352 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_387
timestamp 1698431365
transform 1 0 44688 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_419
timestamp 1698431365
transform 1 0 48272 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_2
timestamp 1698431365
transform 1 0 1568 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_34
timestamp 1698431365
transform 1 0 5152 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_37
timestamp 1698431365
transform 1 0 5488 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_69
timestamp 1698431365
transform 1 0 9072 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_72
timestamp 1698431365
transform 1 0 9408 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_80
timestamp 1698431365
transform 1 0 10304 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_99
timestamp 1698431365
transform 1 0 12432 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_131
timestamp 1698431365
transform 1 0 16016 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_135
timestamp 1698431365
transform 1 0 16464 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_137
timestamp 1698431365
transform 1 0 16688 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_171
timestamp 1698431365
transform 1 0 20496 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_179
timestamp 1698431365
transform 1 0 21392 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_183
timestamp 1698431365
transform 1 0 21840 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_186
timestamp 1698431365
transform 1 0 22176 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_194
timestamp 1698431365
transform 1 0 23072 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_212
timestamp 1698431365
transform 1 0 25088 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_228
timestamp 1698431365
transform 1 0 26880 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_242
timestamp 1698431365
transform 1 0 28448 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_246
timestamp 1698431365
transform 1 0 28896 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_254
timestamp 1698431365
transform 1 0 29792 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_258
timestamp 1698431365
transform 1 0 30240 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_260
timestamp 1698431365
transform 1 0 30464 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_271
timestamp 1698431365
transform 1 0 31696 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_275
timestamp 1698431365
transform 1 0 32144 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_277
timestamp 1698431365
transform 1 0 32368 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_282
timestamp 1698431365
transform 1 0 32928 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_292
timestamp 1698431365
transform 1 0 34048 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_298
timestamp 1698431365
transform 1 0 34720 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_340
timestamp 1698431365
transform 1 0 39424 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_344
timestamp 1698431365
transform 1 0 39872 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_348
timestamp 1698431365
transform 1 0 40320 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_352
timestamp 1698431365
transform 1 0 40768 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_416
timestamp 1698431365
transform 1 0 47936 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_2
timestamp 1698431365
transform 1 0 1568 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_34
timestamp 1698431365
transform 1 0 5152 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_37
timestamp 1698431365
transform 1 0 5488 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_69
timestamp 1698431365
transform 1 0 9072 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_88
timestamp 1698431365
transform 1 0 11200 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_104
timestamp 1698431365
transform 1 0 12992 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_107
timestamp 1698431365
transform 1 0 13328 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_139
timestamp 1698431365
transform 1 0 16912 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_147
timestamp 1698431365
transform 1 0 17808 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_151
timestamp 1698431365
transform 1 0 18256 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_156
timestamp 1698431365
transform 1 0 18816 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_172
timestamp 1698431365
transform 1 0 20608 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_177
timestamp 1698431365
transform 1 0 21168 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_190
timestamp 1698431365
transform 1 0 22624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_194
timestamp 1698431365
transform 1 0 23072 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_201
timestamp 1698431365
transform 1 0 23856 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_205
timestamp 1698431365
transform 1 0 24304 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_213
timestamp 1698431365
transform 1 0 25200 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_247
timestamp 1698431365
transform 1 0 29008 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_278
timestamp 1698431365
transform 1 0 32480 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_309
timestamp 1698431365
transform 1 0 35952 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_325
timestamp 1698431365
transform 1 0 37744 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_355
timestamp 1698431365
transform 1 0 41104 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_371
timestamp 1698431365
transform 1 0 42896 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_379
timestamp 1698431365
transform 1 0 43792 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_383
timestamp 1698431365
transform 1 0 44240 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_387
timestamp 1698431365
transform 1 0 44688 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_419
timestamp 1698431365
transform 1 0 48272 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_2
timestamp 1698431365
transform 1 0 1568 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_10
timestamp 1698431365
transform 1 0 2464 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_15
timestamp 1698431365
transform 1 0 3024 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_23
timestamp 1698431365
transform 1 0 3920 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_26
timestamp 1698431365
transform 1 0 4256 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_42
timestamp 1698431365
transform 1 0 6048 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_50
timestamp 1698431365
transform 1 0 6944 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_52
timestamp 1698431365
transform 1 0 7168 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_55
timestamp 1698431365
transform 1 0 7504 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_59
timestamp 1698431365
transform 1 0 7952 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_63
timestamp 1698431365
transform 1 0 8400 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_67
timestamp 1698431365
transform 1 0 8848 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_80
timestamp 1698431365
transform 1 0 10304 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_82
timestamp 1698431365
transform 1 0 10528 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_100
timestamp 1698431365
transform 1 0 12544 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_121
timestamp 1698431365
transform 1 0 14896 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_137
timestamp 1698431365
transform 1 0 16688 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_139
timestamp 1698431365
transform 1 0 16912 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_142
timestamp 1698431365
transform 1 0 17248 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_144
timestamp 1698431365
transform 1 0 17472 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_209
timestamp 1698431365
transform 1 0 24752 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_212
timestamp 1698431365
transform 1 0 25088 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_217
timestamp 1698431365
transform 1 0 25648 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_221
timestamp 1698431365
transform 1 0 26096 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_229
timestamp 1698431365
transform 1 0 26992 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_245
timestamp 1698431365
transform 1 0 28784 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_253
timestamp 1698431365
transform 1 0 29680 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_257
timestamp 1698431365
transform 1 0 30128 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_265
timestamp 1698431365
transform 1 0 31024 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_273
timestamp 1698431365
transform 1 0 31920 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_276
timestamp 1698431365
transform 1 0 32256 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_282
timestamp 1698431365
transform 1 0 32928 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_291
timestamp 1698431365
transform 1 0 33936 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_340
timestamp 1698431365
transform 1 0 39424 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_344
timestamp 1698431365
transform 1 0 39872 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_348
timestamp 1698431365
transform 1 0 40320 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_352
timestamp 1698431365
transform 1 0 40768 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_416
timestamp 1698431365
transform 1 0 47936 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_2
timestamp 1698431365
transform 1 0 1568 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_4
timestamp 1698431365
transform 1 0 1792 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_28
timestamp 1698431365
transform 1 0 4480 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_32
timestamp 1698431365
transform 1 0 4928 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_34
timestamp 1698431365
transform 1 0 5152 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_37
timestamp 1698431365
transform 1 0 5488 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_41
timestamp 1698431365
transform 1 0 5936 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_77
timestamp 1698431365
transform 1 0 9968 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_81
timestamp 1698431365
transform 1 0 10416 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_102
timestamp 1698431365
transform 1 0 12768 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_104
timestamp 1698431365
transform 1 0 12992 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_82_124
timestamp 1698431365
transform 1 0 15232 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_156
timestamp 1698431365
transform 1 0 18816 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_172
timestamp 1698431365
transform 1 0 20608 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_174
timestamp 1698431365
transform 1 0 20832 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_177
timestamp 1698431365
transform 1 0 21168 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_185
timestamp 1698431365
transform 1 0 22064 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_244
timestamp 1698431365
transform 1 0 28672 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_82_247
timestamp 1698431365
transform 1 0 29008 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_279
timestamp 1698431365
transform 1 0 32592 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_287
timestamp 1698431365
transform 1 0 33488 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_290
timestamp 1698431365
transform 1 0 33824 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_294
timestamp 1698431365
transform 1 0 34272 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_302
timestamp 1698431365
transform 1 0 35168 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_306
timestamp 1698431365
transform 1 0 35616 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_82_346
timestamp 1698431365
transform 1 0 40096 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_378
timestamp 1698431365
transform 1 0 43680 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_382
timestamp 1698431365
transform 1 0 44128 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_384
timestamp 1698431365
transform 1 0 44352 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_82_387
timestamp 1698431365
transform 1 0 44688 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_419
timestamp 1698431365
transform 1 0 48272 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_40
timestamp 1698431365
transform 1 0 5824 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_44
timestamp 1698431365
transform 1 0 6272 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_95
timestamp 1698431365
transform 1 0 11984 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_127
timestamp 1698431365
transform 1 0 15568 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_135
timestamp 1698431365
transform 1 0 16464 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_139
timestamp 1698431365
transform 1 0 16912 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_142
timestamp 1698431365
transform 1 0 17248 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_146
timestamp 1698431365
transform 1 0 17696 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_153
timestamp 1698431365
transform 1 0 18480 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_185
timestamp 1698431365
transform 1 0 22064 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_201
timestamp 1698431365
transform 1 0 23856 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_209
timestamp 1698431365
transform 1 0 24752 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_212
timestamp 1698431365
transform 1 0 25088 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_216
timestamp 1698431365
transform 1 0 25536 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_224
timestamp 1698431365
transform 1 0 26432 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_228
timestamp 1698431365
transform 1 0 26880 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_240
timestamp 1698431365
transform 1 0 28224 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_244
timestamp 1698431365
transform 1 0 28672 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_276
timestamp 1698431365
transform 1 0 32256 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_290
timestamp 1698431365
transform 1 0 33824 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_294
timestamp 1698431365
transform 1 0 34272 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_298
timestamp 1698431365
transform 1 0 34720 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_340
timestamp 1698431365
transform 1 0 39424 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_348
timestamp 1698431365
transform 1 0 40320 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_352
timestamp 1698431365
transform 1 0 40768 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_416
timestamp 1698431365
transform 1 0 47936 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_2
timestamp 1698431365
transform 1 0 1568 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_24
timestamp 1698431365
transform 1 0 4032 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_32
timestamp 1698431365
transform 1 0 4928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_34
timestamp 1698431365
transform 1 0 5152 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_50
timestamp 1698431365
transform 1 0 6944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_54
timestamp 1698431365
transform 1 0 7392 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_58
timestamp 1698431365
transform 1 0 7840 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_87
timestamp 1698431365
transform 1 0 11088 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_103
timestamp 1698431365
transform 1 0 12880 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_107
timestamp 1698431365
transform 1 0 13328 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_123
timestamp 1698431365
transform 1 0 15120 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_131
timestamp 1698431365
transform 1 0 16016 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_133
timestamp 1698431365
transform 1 0 16240 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_165
timestamp 1698431365
transform 1 0 19824 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_167
timestamp 1698431365
transform 1 0 20048 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_172
timestamp 1698431365
transform 1 0 20608 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_174
timestamp 1698431365
transform 1 0 20832 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_177
timestamp 1698431365
transform 1 0 21168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_181
timestamp 1698431365
transform 1 0 21616 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_189
timestamp 1698431365
transform 1 0 22512 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_191
timestamp 1698431365
transform 1 0 22736 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_194
timestamp 1698431365
transform 1 0 23072 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_198
timestamp 1698431365
transform 1 0 23520 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_230
timestamp 1698431365
transform 1 0 27104 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_238
timestamp 1698431365
transform 1 0 28000 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_242
timestamp 1698431365
transform 1 0 28448 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_244
timestamp 1698431365
transform 1 0 28672 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_247
timestamp 1698431365
transform 1 0 29008 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_263
timestamp 1698431365
transform 1 0 30800 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_267
timestamp 1698431365
transform 1 0 31248 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_300
timestamp 1698431365
transform 1 0 34944 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_308
timestamp 1698431365
transform 1 0 35840 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_312
timestamp 1698431365
transform 1 0 36288 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_314
timestamp 1698431365
transform 1 0 36512 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_317
timestamp 1698431365
transform 1 0 36848 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_381
timestamp 1698431365
transform 1 0 44016 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_387
timestamp 1698431365
transform 1 0 44688 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_419
timestamp 1698431365
transform 1 0 48272 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_2
timestamp 1698431365
transform 1 0 1568 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_6
timestamp 1698431365
transform 1 0 2016 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_8
timestamp 1698431365
transform 1 0 2240 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_21
timestamp 1698431365
transform 1 0 3696 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_53
timestamp 1698431365
transform 1 0 7280 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_69
timestamp 1698431365
transform 1 0 9072 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_72
timestamp 1698431365
transform 1 0 9408 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_88
timestamp 1698431365
transform 1 0 11200 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_92
timestamp 1698431365
transform 1 0 11648 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_94
timestamp 1698431365
transform 1 0 11872 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_97
timestamp 1698431365
transform 1 0 12208 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_129
timestamp 1698431365
transform 1 0 15792 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_137
timestamp 1698431365
transform 1 0 16688 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_139
timestamp 1698431365
transform 1 0 16912 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_142
timestamp 1698431365
transform 1 0 17248 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_158
timestamp 1698431365
transform 1 0 19040 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_166
timestamp 1698431365
transform 1 0 19936 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_190
timestamp 1698431365
transform 1 0 22624 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_196
timestamp 1698431365
transform 1 0 23296 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_202
timestamp 1698431365
transform 1 0 23968 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_206
timestamp 1698431365
transform 1 0 24416 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_212
timestamp 1698431365
transform 1 0 25088 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_216
timestamp 1698431365
transform 1 0 25536 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_220
timestamp 1698431365
transform 1 0 25984 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_265
timestamp 1698431365
transform 1 0 31024 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_273
timestamp 1698431365
transform 1 0 31920 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_277
timestamp 1698431365
transform 1 0 32368 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_279
timestamp 1698431365
transform 1 0 32592 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_288
timestamp 1698431365
transform 1 0 33600 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_308
timestamp 1698431365
transform 1 0 35840 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_340
timestamp 1698431365
transform 1 0 39424 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_348
timestamp 1698431365
transform 1 0 40320 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_352
timestamp 1698431365
transform 1 0 40768 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_416
timestamp 1698431365
transform 1 0 47936 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_2
timestamp 1698431365
transform 1 0 1568 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_18
timestamp 1698431365
transform 1 0 3360 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_26
timestamp 1698431365
transform 1 0 4256 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_28
timestamp 1698431365
transform 1 0 4480 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_31
timestamp 1698431365
transform 1 0 4816 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_41
timestamp 1698431365
transform 1 0 5936 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_45
timestamp 1698431365
transform 1 0 6384 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_49
timestamp 1698431365
transform 1 0 6832 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_65
timestamp 1698431365
transform 1 0 8624 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_69
timestamp 1698431365
transform 1 0 9072 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_71
timestamp 1698431365
transform 1 0 9296 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_74
timestamp 1698431365
transform 1 0 9632 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_78
timestamp 1698431365
transform 1 0 10080 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_86_107
timestamp 1698431365
transform 1 0 13328 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_139
timestamp 1698431365
transform 1 0 16912 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_147
timestamp 1698431365
transform 1 0 17808 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_151
timestamp 1698431365
transform 1 0 18256 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_160
timestamp 1698431365
transform 1 0 19264 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_168
timestamp 1698431365
transform 1 0 20160 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_172
timestamp 1698431365
transform 1 0 20608 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_174
timestamp 1698431365
transform 1 0 20832 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_200
timestamp 1698431365
transform 1 0 23744 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_202
timestamp 1698431365
transform 1 0 23968 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_205
timestamp 1698431365
transform 1 0 24304 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_238
timestamp 1698431365
transform 1 0 28000 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_247
timestamp 1698431365
transform 1 0 29008 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_280
timestamp 1698431365
transform 1 0 32704 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_284
timestamp 1698431365
transform 1 0 33152 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_292
timestamp 1698431365
transform 1 0 34048 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_314
timestamp 1698431365
transform 1 0 36512 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_317
timestamp 1698431365
transform 1 0 36848 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_321
timestamp 1698431365
transform 1 0 37296 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_86_387
timestamp 1698431365
transform 1 0 44688 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_419
timestamp 1698431365
transform 1 0 48272 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_2
timestamp 1698431365
transform 1 0 1568 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_18
timestamp 1698431365
transform 1 0 3360 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_20
timestamp 1698431365
transform 1 0 3584 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_72
timestamp 1698431365
transform 1 0 9408 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_120
timestamp 1698431365
transform 1 0 14784 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_136
timestamp 1698431365
transform 1 0 16576 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_142
timestamp 1698431365
transform 1 0 17248 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_87_177
timestamp 1698431365
transform 1 0 21168 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_185
timestamp 1698431365
transform 1 0 22064 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_235
timestamp 1698431365
transform 1 0 27664 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_239
timestamp 1698431365
transform 1 0 28112 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_251
timestamp 1698431365
transform 1 0 29456 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_260
timestamp 1698431365
transform 1 0 30464 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_264
timestamp 1698431365
transform 1 0 30912 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_268
timestamp 1698431365
transform 1 0 31360 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_87_272
timestamp 1698431365
transform 1 0 31808 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_282
timestamp 1698431365
transform 1 0 32928 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_286
timestamp 1698431365
transform 1 0 33376 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_290
timestamp 1698431365
transform 1 0 33824 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_87_337
timestamp 1698431365
transform 1 0 39088 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_345
timestamp 1698431365
transform 1 0 39984 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_349
timestamp 1698431365
transform 1 0 40432 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_352
timestamp 1698431365
transform 1 0 40768 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_416
timestamp 1698431365
transform 1 0 47936 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_2
timestamp 1698431365
transform 1 0 1568 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_6
timestamp 1698431365
transform 1 0 2016 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_32
timestamp 1698431365
transform 1 0 4928 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_34
timestamp 1698431365
transform 1 0 5152 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_43
timestamp 1698431365
transform 1 0 6160 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_67
timestamp 1698431365
transform 1 0 8848 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_75
timestamp 1698431365
transform 1 0 9744 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_79
timestamp 1698431365
transform 1 0 10192 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_107
timestamp 1698431365
transform 1 0 13328 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_171
timestamp 1698431365
transform 1 0 20496 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_183
timestamp 1698431365
transform 1 0 21840 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_187
timestamp 1698431365
transform 1 0 22288 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_225
timestamp 1698431365
transform 1 0 26544 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_229
timestamp 1698431365
transform 1 0 26992 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_247
timestamp 1698431365
transform 1 0 29008 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_253
timestamp 1698431365
transform 1 0 29680 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_269
timestamp 1698431365
transform 1 0 31472 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_273
timestamp 1698431365
transform 1 0 31920 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_275
timestamp 1698431365
transform 1 0 32144 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_295
timestamp 1698431365
transform 1 0 34384 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_346
timestamp 1698431365
transform 1 0 40096 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_378
timestamp 1698431365
transform 1 0 43680 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_382
timestamp 1698431365
transform 1 0 44128 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_384
timestamp 1698431365
transform 1 0 44352 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_387
timestamp 1698431365
transform 1 0 44688 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_419
timestamp 1698431365
transform 1 0 48272 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_2
timestamp 1698431365
transform 1 0 1568 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_27
timestamp 1698431365
transform 1 0 4368 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_31
timestamp 1698431365
transform 1 0 4816 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_35
timestamp 1698431365
transform 1 0 5264 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_39
timestamp 1698431365
transform 1 0 5712 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_66
timestamp 1698431365
transform 1 0 8736 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_89_95
timestamp 1698431365
transform 1 0 11984 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_127
timestamp 1698431365
transform 1 0 15568 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_135
timestamp 1698431365
transform 1 0 16464 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_139
timestamp 1698431365
transform 1 0 16912 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_142
timestamp 1698431365
transform 1 0 17248 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_158
timestamp 1698431365
transform 1 0 19040 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_166
timestamp 1698431365
transform 1 0 19936 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_168
timestamp 1698431365
transform 1 0 20160 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_209
timestamp 1698431365
transform 1 0 24752 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_212
timestamp 1698431365
transform 1 0 25088 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_214
timestamp 1698431365
transform 1 0 25312 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_219
timestamp 1698431365
transform 1 0 25872 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_89_223
timestamp 1698431365
transform 1 0 26320 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_255
timestamp 1698431365
transform 1 0 29904 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_271
timestamp 1698431365
transform 1 0 31696 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_275
timestamp 1698431365
transform 1 0 32144 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_277
timestamp 1698431365
transform 1 0 32368 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_288
timestamp 1698431365
transform 1 0 33600 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_292
timestamp 1698431365
transform 1 0 34048 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_296
timestamp 1698431365
transform 1 0 34496 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_316
timestamp 1698431365
transform 1 0 36736 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_318
timestamp 1698431365
transform 1 0 36960 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_325
timestamp 1698431365
transform 1 0 37744 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_329
timestamp 1698431365
transform 1 0 38192 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_345
timestamp 1698431365
transform 1 0 39984 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_349
timestamp 1698431365
transform 1 0 40432 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_352
timestamp 1698431365
transform 1 0 40768 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_416
timestamp 1698431365
transform 1 0 47936 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_19
timestamp 1698431365
transform 1 0 3472 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_27
timestamp 1698431365
transform 1 0 4368 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_31
timestamp 1698431365
transform 1 0 4816 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_37
timestamp 1698431365
transform 1 0 5488 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_39
timestamp 1698431365
transform 1 0 5712 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_63
timestamp 1698431365
transform 1 0 8400 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_65
timestamp 1698431365
transform 1 0 8624 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_91
timestamp 1698431365
transform 1 0 11536 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_95
timestamp 1698431365
transform 1 0 11984 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_103
timestamp 1698431365
transform 1 0 12880 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_107
timestamp 1698431365
transform 1 0 13328 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_171
timestamp 1698431365
transform 1 0 20496 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_177
timestamp 1698431365
transform 1 0 21168 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_193
timestamp 1698431365
transform 1 0 22960 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_197
timestamp 1698431365
transform 1 0 23408 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_200
timestamp 1698431365
transform 1 0 23744 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_232
timestamp 1698431365
transform 1 0 27328 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_240
timestamp 1698431365
transform 1 0 28224 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_244
timestamp 1698431365
transform 1 0 28672 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_247
timestamp 1698431365
transform 1 0 29008 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_251
timestamp 1698431365
transform 1 0 29456 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_253
timestamp 1698431365
transform 1 0 29680 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_290
timestamp 1698431365
transform 1 0 33824 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_292
timestamp 1698431365
transform 1 0 34048 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_295
timestamp 1698431365
transform 1 0 34384 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_299
timestamp 1698431365
transform 1 0 34832 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_303
timestamp 1698431365
transform 1 0 35280 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_311
timestamp 1698431365
transform 1 0 36176 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_317
timestamp 1698431365
transform 1 0 36848 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_321
timestamp 1698431365
transform 1 0 37296 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_325
timestamp 1698431365
transform 1 0 37744 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_357
timestamp 1698431365
transform 1 0 41328 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_373
timestamp 1698431365
transform 1 0 43120 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_381
timestamp 1698431365
transform 1 0 44016 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_387
timestamp 1698431365
transform 1 0 44688 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_419
timestamp 1698431365
transform 1 0 48272 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_2
timestamp 1698431365
transform 1 0 1568 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_66
timestamp 1698431365
transform 1 0 8736 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_118
timestamp 1698431365
transform 1 0 14560 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_134
timestamp 1698431365
transform 1 0 16352 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_138
timestamp 1698431365
transform 1 0 16800 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_142
timestamp 1698431365
transform 1 0 17248 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_150
timestamp 1698431365
transform 1 0 18144 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_154
timestamp 1698431365
transform 1 0 18592 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_156
timestamp 1698431365
transform 1 0 18816 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_165
timestamp 1698431365
transform 1 0 19824 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_197
timestamp 1698431365
transform 1 0 23408 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_205
timestamp 1698431365
transform 1 0 24304 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_209
timestamp 1698431365
transform 1 0 24752 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_212
timestamp 1698431365
transform 1 0 25088 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_276
timestamp 1698431365
transform 1 0 32256 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_286
timestamp 1698431365
transform 1 0 33376 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_292
timestamp 1698431365
transform 1 0 34048 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_324
timestamp 1698431365
transform 1 0 37632 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_340
timestamp 1698431365
transform 1 0 39424 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_348
timestamp 1698431365
transform 1 0 40320 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_352
timestamp 1698431365
transform 1 0 40768 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_416
timestamp 1698431365
transform 1 0 47936 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_2
timestamp 1698431365
transform 1 0 1568 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_34
timestamp 1698431365
transform 1 0 5152 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_37
timestamp 1698431365
transform 1 0 5488 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_69
timestamp 1698431365
transform 1 0 9072 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_77
timestamp 1698431365
transform 1 0 9968 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_79
timestamp 1698431365
transform 1 0 10192 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_107
timestamp 1698431365
transform 1 0 13328 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_139
timestamp 1698431365
transform 1 0 16912 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_143
timestamp 1698431365
transform 1 0 17360 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_181
timestamp 1698431365
transform 1 0 21616 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_247
timestamp 1698431365
transform 1 0 29008 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_262
timestamp 1698431365
transform 1 0 30688 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_278
timestamp 1698431365
transform 1 0 32480 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_282
timestamp 1698431365
transform 1 0 32928 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_284
timestamp 1698431365
transform 1 0 33152 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_289
timestamp 1698431365
transform 1 0 33712 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_297
timestamp 1698431365
transform 1 0 34608 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_301
timestamp 1698431365
transform 1 0 35056 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_311
timestamp 1698431365
transform 1 0 36176 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_321
timestamp 1698431365
transform 1 0 37296 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_387
timestamp 1698431365
transform 1 0 44688 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_419
timestamp 1698431365
transform 1 0 48272 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_2
timestamp 1698431365
transform 1 0 1568 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_10
timestamp 1698431365
transform 1 0 2464 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_31
timestamp 1698431365
transform 1 0 4816 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_64
timestamp 1698431365
transform 1 0 8512 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_95
timestamp 1698431365
transform 1 0 11984 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_127
timestamp 1698431365
transform 1 0 15568 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_135
timestamp 1698431365
transform 1 0 16464 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_139
timestamp 1698431365
transform 1 0 16912 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_142
timestamp 1698431365
transform 1 0 17248 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_174
timestamp 1698431365
transform 1 0 20832 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_190
timestamp 1698431365
transform 1 0 22624 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_198
timestamp 1698431365
transform 1 0 23520 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_202
timestamp 1698431365
transform 1 0 23968 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_206
timestamp 1698431365
transform 1 0 24416 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_217
timestamp 1698431365
transform 1 0 25648 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_221
timestamp 1698431365
transform 1 0 26096 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_229
timestamp 1698431365
transform 1 0 26992 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_235
timestamp 1698431365
transform 1 0 27664 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_251
timestamp 1698431365
transform 1 0 29456 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_259
timestamp 1698431365
transform 1 0 30352 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_263
timestamp 1698431365
transform 1 0 30800 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_266
timestamp 1698431365
transform 1 0 31136 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_274
timestamp 1698431365
transform 1 0 32032 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_282
timestamp 1698431365
transform 1 0 32928 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_284
timestamp 1698431365
transform 1 0 33152 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_291
timestamp 1698431365
transform 1 0 33936 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_295
timestamp 1698431365
transform 1 0 34384 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_328
timestamp 1698431365
transform 1 0 38080 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_344
timestamp 1698431365
transform 1 0 39872 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_348
timestamp 1698431365
transform 1 0 40320 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_93_352
timestamp 1698431365
transform 1 0 40768 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_416
timestamp 1698431365
transform 1 0 47936 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_94_2
timestamp 1698431365
transform 1 0 1568 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_10
timestamp 1698431365
transform 1 0 2464 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_31
timestamp 1698431365
transform 1 0 4816 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_37
timestamp 1698431365
transform 1 0 5488 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_39
timestamp 1698431365
transform 1 0 5712 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_94_65
timestamp 1698431365
transform 1 0 8624 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_98
timestamp 1698431365
transform 1 0 12320 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_100
timestamp 1698431365
transform 1 0 12544 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_103
timestamp 1698431365
transform 1 0 12880 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_94_107
timestamp 1698431365
transform 1 0 13328 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_171
timestamp 1698431365
transform 1 0 20496 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_183
timestamp 1698431365
transform 1 0 21840 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_187
timestamp 1698431365
transform 1 0 22288 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_200
timestamp 1698431365
transform 1 0 23744 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_243
timestamp 1698431365
transform 1 0 28560 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_247
timestamp 1698431365
transform 1 0 29008 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_251
timestamp 1698431365
transform 1 0 29456 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_253
timestamp 1698431365
transform 1 0 29680 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_262
timestamp 1698431365
transform 1 0 30688 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_301
timestamp 1698431365
transform 1 0 35056 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_305
timestamp 1698431365
transform 1 0 35504 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_94_309
timestamp 1698431365
transform 1 0 35952 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_94_317
timestamp 1698431365
transform 1 0 36848 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_94_381
timestamp 1698431365
transform 1 0 44016 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_94_387
timestamp 1698431365
transform 1 0 44688 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_94_419
timestamp 1698431365
transform 1 0 48272 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_2
timestamp 1698431365
transform 1 0 1568 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_67
timestamp 1698431365
transform 1 0 8848 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_69
timestamp 1698431365
transform 1 0 9072 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_72
timestamp 1698431365
transform 1 0 9408 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_76
timestamp 1698431365
transform 1 0 9856 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_95_126
timestamp 1698431365
transform 1 0 15456 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_134
timestamp 1698431365
transform 1 0 16352 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_138
timestamp 1698431365
transform 1 0 16800 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_95_142
timestamp 1698431365
transform 1 0 17248 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_95_212
timestamp 1698431365
transform 1 0 25088 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_220
timestamp 1698431365
transform 1 0 25984 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_224
timestamp 1698431365
transform 1 0 26432 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_226
timestamp 1698431365
transform 1 0 26656 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_258
timestamp 1698431365
transform 1 0 30240 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_95_266
timestamp 1698431365
transform 1 0 31136 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_274
timestamp 1698431365
transform 1 0 32032 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_278
timestamp 1698431365
transform 1 0 32480 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_282
timestamp 1698431365
transform 1 0 32928 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_95_319
timestamp 1698431365
transform 1 0 37072 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_95_335
timestamp 1698431365
transform 1 0 38864 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_343
timestamp 1698431365
transform 1 0 39760 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95_347
timestamp 1698431365
transform 1 0 40208 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_95_349
timestamp 1698431365
transform 1 0 40432 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_95_352
timestamp 1698431365
transform 1 0 40768 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95_416
timestamp 1698431365
transform 1 0 47936 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_96_19
timestamp 1698431365
transform 1 0 3472 0 1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_37
timestamp 1698431365
transform 1 0 5488 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_41
timestamp 1698431365
transform 1 0 5936 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_45
timestamp 1698431365
transform 1 0 6384 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_49
timestamp 1698431365
transform 1 0 6832 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_96_78
timestamp 1698431365
transform 1 0 10080 0 1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_96_94
timestamp 1698431365
transform 1 0 11872 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_102
timestamp 1698431365
transform 1 0 12768 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_104
timestamp 1698431365
transform 1 0 12992 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_96_107
timestamp 1698431365
transform 1 0 13328 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_171
timestamp 1698431365
transform 1 0 20496 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_177
timestamp 1698431365
transform 1 0 21168 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_96_181
timestamp 1698431365
transform 1 0 21616 0 1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_96_213
timestamp 1698431365
transform 1 0 25200 0 1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_229
timestamp 1698431365
transform 1 0 26992 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_233
timestamp 1698431365
transform 1 0 27440 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_241
timestamp 1698431365
transform 1 0 28336 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_96_247
timestamp 1698431365
transform 1 0 29008 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_255
timestamp 1698431365
transform 1 0 29904 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_257
timestamp 1698431365
transform 1 0 30128 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_96_287
timestamp 1698431365
transform 1 0 33488 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_96_291
timestamp 1698431365
transform 1 0 33936 0 1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_96_307
timestamp 1698431365
transform 1 0 35728 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_96_317
timestamp 1698431365
transform 1 0 36848 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_96_381
timestamp 1698431365
transform 1 0 44016 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_96_387
timestamp 1698431365
transform 1 0 44688 0 1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_96_419
timestamp 1698431365
transform 1 0 48272 0 1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_97_19
timestamp 1698431365
transform 1 0 3472 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_97_27
timestamp 1698431365
transform 1 0 4368 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_31
timestamp 1698431365
transform 1 0 4816 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_97_33
timestamp 1698431365
transform 1 0 5040 0 -1 78400
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_97_36
timestamp 1698431365
transform 1 0 5376 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_97_70
timestamp 1698431365
transform 1 0 9184 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_97_104
timestamp 1698431365
transform 1 0 12992 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_97_138
timestamp 1698431365
transform 1 0 16800 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_97_172
timestamp 1698431365
transform 1 0 20608 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_97_206
timestamp 1698431365
transform 1 0 24416 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_97_240
timestamp 1698431365
transform 1 0 28224 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_97_274
timestamp 1698431365
transform 1 0 32032 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_97_308
timestamp 1698431365
transform 1 0 35840 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_97_342
timestamp 1698431365
transform 1 0 39648 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_97_376
timestamp 1698431365
transform 1 0 43456 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_97_410
timestamp 1698431365
transform 1 0 47264 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_97_418
timestamp 1698431365
transform 1 0 48160 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  input2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input5
timestamp 1698431365
transform 1 0 2464 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input6
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_98 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 48608 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 48608 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_136
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_137
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_138
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_139
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_140
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_141
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_142
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_143
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_144
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_145
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_146
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_147
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_148
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_149
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_150
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_151
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_152
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_153
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_154
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_155
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 48608 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_156
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 48608 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_157
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 48608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_158
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 48608 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_159
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 48608 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_160
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 48608 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_161
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 48608 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_162
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 48608 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_163
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 48608 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_164
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 48608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_165
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 48608 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_166
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698431365
transform -1 0 48608 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_167
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698431365
transform -1 0 48608 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_168
timestamp 1698431365
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698431365
transform -1 0 48608 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_169
timestamp 1698431365
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698431365
transform -1 0 48608 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_170
timestamp 1698431365
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698431365
transform -1 0 48608 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_171
timestamp 1698431365
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1698431365
transform -1 0 48608 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_172
timestamp 1698431365
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1698431365
transform -1 0 48608 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_173
timestamp 1698431365
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1698431365
transform -1 0 48608 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_174
timestamp 1698431365
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1698431365
transform -1 0 48608 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_175
timestamp 1698431365
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1698431365
transform -1 0 48608 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_176
timestamp 1698431365
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1698431365
transform -1 0 48608 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_177
timestamp 1698431365
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1698431365
transform -1 0 48608 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_178
timestamp 1698431365
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1698431365
transform -1 0 48608 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Left_179
timestamp 1698431365
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Right_81
timestamp 1698431365
transform -1 0 48608 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Left_180
timestamp 1698431365
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Right_82
timestamp 1698431365
transform -1 0 48608 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Left_181
timestamp 1698431365
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Right_83
timestamp 1698431365
transform -1 0 48608 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Left_182
timestamp 1698431365
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Right_84
timestamp 1698431365
transform -1 0 48608 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Left_183
timestamp 1698431365
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Right_85
timestamp 1698431365
transform -1 0 48608 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Left_184
timestamp 1698431365
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Right_86
timestamp 1698431365
transform -1 0 48608 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Left_185
timestamp 1698431365
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Right_87
timestamp 1698431365
transform -1 0 48608 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Left_186
timestamp 1698431365
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Right_88
timestamp 1698431365
transform -1 0 48608 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Left_187
timestamp 1698431365
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Right_89
timestamp 1698431365
transform -1 0 48608 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Left_188
timestamp 1698431365
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Right_90
timestamp 1698431365
transform -1 0 48608 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Left_189
timestamp 1698431365
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Right_91
timestamp 1698431365
transform -1 0 48608 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Left_190
timestamp 1698431365
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Right_92
timestamp 1698431365
transform -1 0 48608 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Left_191
timestamp 1698431365
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Right_93
timestamp 1698431365
transform -1 0 48608 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_Left_192
timestamp 1698431365
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_94_Right_94
timestamp 1698431365
transform -1 0 48608 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_Left_193
timestamp 1698431365
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_95_Right_95
timestamp 1698431365
transform -1 0 48608 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_Left_194
timestamp 1698431365
transform 1 0 1344 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_96_Right_96
timestamp 1698431365
transform -1 0 48608 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_Left_195
timestamp 1698431365
transform 1 0 1344 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_97_Right_97
timestamp 1698431365
transform -1 0 48608 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  seg1._26_
timestamp 1698431365
transform -1 0 8064 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  seg1._27_
timestamp 1698431365
transform -1 0 6272 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  seg1._28_
timestamp 1698431365
transform -1 0 7280 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  seg1._29_
timestamp 1698431365
transform -1 0 5376 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  seg1._30_
timestamp 1698431365
transform -1 0 5264 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  seg1._31_
timestamp 1698431365
transform -1 0 5264 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  seg1._32_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  seg1._33_
timestamp 1698431365
transform -1 0 4928 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  seg1._34_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4928 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  seg1._35_
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  seg1._36_
timestamp 1698431365
transform 1 0 5152 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._37_
timestamp 1698431365
transform 1 0 8400 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  seg1._38_
timestamp 1698431365
transform 1 0 6720 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  seg1._39_
timestamp 1698431365
transform 1 0 6496 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._40_
timestamp 1698431365
transform 1 0 4704 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  seg1._41_
timestamp 1698431365
transform 1 0 7392 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._42_
timestamp 1698431365
transform -1 0 9968 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._43_
timestamp 1698431365
transform 1 0 7952 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  seg1._44_
timestamp 1698431365
transform -1 0 6048 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  seg1._45_ open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 8400 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  seg1._46_
timestamp 1698431365
transform -1 0 8176 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  seg1._47_
timestamp 1698431365
transform 1 0 7280 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  seg1._48_
timestamp 1698431365
transform -1 0 10080 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  seg1._49_
timestamp 1698431365
transform 1 0 6160 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._50_
timestamp 1698431365
transform 1 0 6384 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  seg1._51_
timestamp 1698431365
transform 1 0 5376 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._52_
timestamp 1698431365
transform 1 0 5824 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  seg1._53_
timestamp 1698431365
transform 1 0 9072 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  seg1._54_
timestamp 1698431365
transform 1 0 8176 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  seg1._55_
timestamp 1698431365
transform -1 0 9184 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  seg1._56_
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  seg1._57_
timestamp 1698431365
transform 1 0 5712 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  seg1._58_
timestamp 1698431365
transform 1 0 5600 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_196 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_197
timestamp 1698431365
transform 1 0 8960 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_198
timestamp 1698431365
transform 1 0 12768 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_199
timestamp 1698431365
transform 1 0 16576 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_200
timestamp 1698431365
transform 1 0 20384 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_201
timestamp 1698431365
transform 1 0 24192 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_202
timestamp 1698431365
transform 1 0 28000 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_203
timestamp 1698431365
transform 1 0 31808 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_204
timestamp 1698431365
transform 1 0 35616 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_205
timestamp 1698431365
transform 1 0 39424 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_206
timestamp 1698431365
transform 1 0 43232 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_207
timestamp 1698431365
transform 1 0 47040 0 1 1568
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_208
timestamp 1698431365
transform 1 0 9184 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_209
timestamp 1698431365
transform 1 0 17024 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_210
timestamp 1698431365
transform 1 0 24864 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_211
timestamp 1698431365
transform 1 0 32704 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_212
timestamp 1698431365
transform 1 0 40544 0 -1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_213
timestamp 1698431365
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_214
timestamp 1698431365
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_215
timestamp 1698431365
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_216
timestamp 1698431365
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_217
timestamp 1698431365
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_218
timestamp 1698431365
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_219
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_220
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_221
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_222
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_223
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_224
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_225
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_226
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_227
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_228
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_229
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_230
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_231
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_232
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_233
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_234
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_235
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_236
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_237
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_238
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_239
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_240
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_241
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_242
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_243
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_244
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_245
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_246
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_247
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_248
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_249
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_250
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_251
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_252
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_253
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_254
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_255
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_256
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_257
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_258
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_259
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_260
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_261
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_262
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_263
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_264
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_265
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_266
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_267
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_268
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_269
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_270
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_271
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_272
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_273
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_274
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_275
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_276
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_277
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_278
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_279
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_280
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_281
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_282
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_283
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_284
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_285
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_286
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_287
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_288
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_289
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_290
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_291
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_292
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_293
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_294
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_295
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_296
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_297
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_298
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_299
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_300
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_301
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_302
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_303
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_304
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_305
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_306
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_307
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_308
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_309
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_310
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_311
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_312
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_313
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_314
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_315
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_316
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_317
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_318
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_319
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_320
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_321
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_322
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_323
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_324
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_325
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_326
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_327
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_328
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_329
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_330
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_331
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_332
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_333
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_334
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_335
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_336
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_337
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_338
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_339
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_340
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_341
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_342
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_343
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_344
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_345
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_346
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_347
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_348
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_349
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_350
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_351
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_352
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_353
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_354
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_355
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_356
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_357
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_358
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_359
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_360
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_361
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_362
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_363
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_364
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_365
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_366
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_367
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_368
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_369
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_370
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_371
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_372
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_373
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_374
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_375
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_376
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_377
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_378
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_379
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_380
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_381
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_382
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_383
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_384
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_385
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_386
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_387
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_388
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_389
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_390
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_391
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_392
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_393
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_394
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_395
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_396
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_397
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_398
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_399
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_400
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_401
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_402
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_403
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_404
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_405
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_406
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_407
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_408
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_409
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_410
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_411
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_412
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_413
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_414
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_416
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_417
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_418
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_422
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_425
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_426
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_427
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_428
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_429
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_430
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_431
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_432
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_433
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_434
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_435
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_436
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_437
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_438
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_439
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_440
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_441
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_442
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_443
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_444
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_445
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_446
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_447
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_448
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_449
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_450
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_451
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_452
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_453
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_454
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_455
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_456
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_457
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_458
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_459
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_460
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_461
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_462
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_463
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_464
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_465
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_466
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_467
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_468
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_469
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_470
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_471
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_472
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_473
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_474
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_475
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_476
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_477
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_478
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_479
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_480
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_481
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_482
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_483
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_484
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_485
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_486
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_487
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_488
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_489
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_490
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_491
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_492
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_493
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_494
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_495
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_496
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_497
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_498
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_499
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_500
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_501
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_502
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_503
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_504
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_505
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_506
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_507
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_508
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_509
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_510
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_511
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_512
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_513
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_514
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_515
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_516
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_517
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_518
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_519
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_520
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_521
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_522
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_523
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_524
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_525
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_526
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_527
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_528
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_529
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_530
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_531
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_532
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_533
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_534
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_535
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_536
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_537
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_538
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_539
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_540
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_541
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_542
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_543
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_544
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_545
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_546
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_547
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_548
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_549
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_550
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_551
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_552
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_553
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_554
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_555
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_556
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_557
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_558
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_559
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_560
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_561
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_562
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_563
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_564
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_565
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_566
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_567
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_568
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_569
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_570
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_571
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_572
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_573
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_574
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_575
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_576
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_577
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_578
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_579
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_580
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_581
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_582
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_583
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_584
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_585
timestamp 1698431365
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_586
timestamp 1698431365
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_587
timestamp 1698431365
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_588
timestamp 1698431365
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_589
timestamp 1698431365
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_590
timestamp 1698431365
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_591
timestamp 1698431365
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_592
timestamp 1698431365
transform 1 0 44464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_593
timestamp 1698431365
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_594
timestamp 1698431365
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_595
timestamp 1698431365
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_596
timestamp 1698431365
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_597
timestamp 1698431365
transform 1 0 40544 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_598
timestamp 1698431365
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_599
timestamp 1698431365
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_600
timestamp 1698431365
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_601
timestamp 1698431365
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_602
timestamp 1698431365
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_603
timestamp 1698431365
transform 1 0 44464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_604
timestamp 1698431365
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_605
timestamp 1698431365
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_606
timestamp 1698431365
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_607
timestamp 1698431365
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_608
timestamp 1698431365
transform 1 0 40544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_609
timestamp 1698431365
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_610
timestamp 1698431365
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_611
timestamp 1698431365
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_612
timestamp 1698431365
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_613
timestamp 1698431365
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_614
timestamp 1698431365
transform 1 0 44464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_615
timestamp 1698431365
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_616
timestamp 1698431365
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_617
timestamp 1698431365
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_618
timestamp 1698431365
transform 1 0 32704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_619
timestamp 1698431365
transform 1 0 40544 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_620
timestamp 1698431365
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_621
timestamp 1698431365
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_622
timestamp 1698431365
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_623
timestamp 1698431365
transform 1 0 28784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_624
timestamp 1698431365
transform 1 0 36624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_625
timestamp 1698431365
transform 1 0 44464 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_626
timestamp 1698431365
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_627
timestamp 1698431365
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_628
timestamp 1698431365
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_629
timestamp 1698431365
transform 1 0 32704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_630
timestamp 1698431365
transform 1 0 40544 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_631
timestamp 1698431365
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_632
timestamp 1698431365
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_633
timestamp 1698431365
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_634
timestamp 1698431365
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_635
timestamp 1698431365
transform 1 0 36624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_636
timestamp 1698431365
transform 1 0 44464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_637
timestamp 1698431365
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_638
timestamp 1698431365
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_639
timestamp 1698431365
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_640
timestamp 1698431365
transform 1 0 32704 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_641
timestamp 1698431365
transform 1 0 40544 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_642
timestamp 1698431365
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_643
timestamp 1698431365
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_644
timestamp 1698431365
transform 1 0 20944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_645
timestamp 1698431365
transform 1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_646
timestamp 1698431365
transform 1 0 36624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_647
timestamp 1698431365
transform 1 0 44464 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_648
timestamp 1698431365
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_649
timestamp 1698431365
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_650
timestamp 1698431365
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_651
timestamp 1698431365
transform 1 0 32704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_652
timestamp 1698431365
transform 1 0 40544 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_653
timestamp 1698431365
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_654
timestamp 1698431365
transform 1 0 13104 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_655
timestamp 1698431365
transform 1 0 20944 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_656
timestamp 1698431365
transform 1 0 28784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_657
timestamp 1698431365
transform 1 0 36624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_658
timestamp 1698431365
transform 1 0 44464 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_659
timestamp 1698431365
transform 1 0 9184 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_660
timestamp 1698431365
transform 1 0 17024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_661
timestamp 1698431365
transform 1 0 24864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_662
timestamp 1698431365
transform 1 0 32704 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_663
timestamp 1698431365
transform 1 0 40544 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_664
timestamp 1698431365
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_665
timestamp 1698431365
transform 1 0 13104 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_666
timestamp 1698431365
transform 1 0 20944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_667
timestamp 1698431365
transform 1 0 28784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_668
timestamp 1698431365
transform 1 0 36624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_669
timestamp 1698431365
transform 1 0 44464 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_670
timestamp 1698431365
transform 1 0 9184 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_671
timestamp 1698431365
transform 1 0 17024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_672
timestamp 1698431365
transform 1 0 24864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_673
timestamp 1698431365
transform 1 0 32704 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_674
timestamp 1698431365
transform 1 0 40544 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_675
timestamp 1698431365
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_676
timestamp 1698431365
transform 1 0 13104 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_677
timestamp 1698431365
transform 1 0 20944 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_678
timestamp 1698431365
transform 1 0 28784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_679
timestamp 1698431365
transform 1 0 36624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_680
timestamp 1698431365
transform 1 0 44464 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_681
timestamp 1698431365
transform 1 0 9184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_682
timestamp 1698431365
transform 1 0 17024 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_683
timestamp 1698431365
transform 1 0 24864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_684
timestamp 1698431365
transform 1 0 32704 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_685
timestamp 1698431365
transform 1 0 40544 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_686
timestamp 1698431365
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_687
timestamp 1698431365
transform 1 0 13104 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_688
timestamp 1698431365
transform 1 0 20944 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_689
timestamp 1698431365
transform 1 0 28784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_690
timestamp 1698431365
transform 1 0 36624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_691
timestamp 1698431365
transform 1 0 44464 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_692
timestamp 1698431365
transform 1 0 9184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_693
timestamp 1698431365
transform 1 0 17024 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_694
timestamp 1698431365
transform 1 0 24864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_695
timestamp 1698431365
transform 1 0 32704 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_696
timestamp 1698431365
transform 1 0 40544 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_697
timestamp 1698431365
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_698
timestamp 1698431365
transform 1 0 13104 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_699
timestamp 1698431365
transform 1 0 20944 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_700
timestamp 1698431365
transform 1 0 28784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_701
timestamp 1698431365
transform 1 0 36624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_702
timestamp 1698431365
transform 1 0 44464 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_703
timestamp 1698431365
transform 1 0 9184 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_704
timestamp 1698431365
transform 1 0 17024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_705
timestamp 1698431365
transform 1 0 24864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_706
timestamp 1698431365
transform 1 0 32704 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_707
timestamp 1698431365
transform 1 0 40544 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_708
timestamp 1698431365
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_709
timestamp 1698431365
transform 1 0 13104 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_710
timestamp 1698431365
transform 1 0 20944 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_711
timestamp 1698431365
transform 1 0 28784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_712
timestamp 1698431365
transform 1 0 36624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_713
timestamp 1698431365
transform 1 0 44464 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_714
timestamp 1698431365
transform 1 0 9184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_715
timestamp 1698431365
transform 1 0 17024 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_716
timestamp 1698431365
transform 1 0 24864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_717
timestamp 1698431365
transform 1 0 32704 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_718
timestamp 1698431365
transform 1 0 40544 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_719
timestamp 1698431365
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_720
timestamp 1698431365
transform 1 0 13104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_721
timestamp 1698431365
transform 1 0 20944 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_722
timestamp 1698431365
transform 1 0 28784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_723
timestamp 1698431365
transform 1 0 36624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_94_724
timestamp 1698431365
transform 1 0 44464 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_725
timestamp 1698431365
transform 1 0 9184 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_726
timestamp 1698431365
transform 1 0 17024 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_727
timestamp 1698431365
transform 1 0 24864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_728
timestamp 1698431365
transform 1 0 32704 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_95_729
timestamp 1698431365
transform 1 0 40544 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_730
timestamp 1698431365
transform 1 0 5264 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_731
timestamp 1698431365
transform 1 0 13104 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_732
timestamp 1698431365
transform 1 0 20944 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_733
timestamp 1698431365
transform 1 0 28784 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_734
timestamp 1698431365
transform 1 0 36624 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_96_735
timestamp 1698431365
transform 1 0 44464 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_736
timestamp 1698431365
transform 1 0 5152 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_737
timestamp 1698431365
transform 1 0 8960 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_738
timestamp 1698431365
transform 1 0 12768 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_739
timestamp 1698431365
transform 1 0 16576 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_740
timestamp 1698431365
transform 1 0 20384 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_741
timestamp 1698431365
transform 1 0 24192 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_742
timestamp 1698431365
transform 1 0 28000 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_743
timestamp 1698431365
transform 1 0 31808 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_744
timestamp 1698431365
transform 1 0 35616 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_745
timestamp 1698431365
transform 1 0 39424 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_746
timestamp 1698431365
transform 1 0 43232 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_97_747
timestamp 1698431365
transform 1 0 47040 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac._4_
timestamp 1698431365
transform -1 0 4480 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  temp1.dac._5_
timestamp 1698431365
transform 1 0 3360 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[0\].vdac_batch._3_
timestamp 1698431365
transform 1 0 4816 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[0\].vdac_batch._4_
timestamp 1698431365
transform -1 0 3920 0 -1 58016
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[0\].vdac_batch._5_
timestamp 1698431365
transform 1 0 2800 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  temp1.dac.parallel_cells\[0\].vdac_batch._6_
timestamp 1698431365
transform -1 0 4816 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[0\].vdac_batch._7_
timestamp 1698431365
transform 1 0 2016 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  temp1.dac.parallel_cells\[0\].vdac_batch._8_
timestamp 1698431365
transform -1 0 2800 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].pupd open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3920 0 -1 58016
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[0\].vdac_batch.einvp_batch\[0\].vref open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 58016
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[1\].vdac_batch._3_
timestamp 1698431365
transform -1 0 4032 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[1\].vdac_batch._4_
timestamp 1698431365
transform 1 0 3584 0 1 61152
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[1\].vdac_batch._5_
timestamp 1698431365
transform -1 0 4480 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  temp1.dac.parallel_cells\[1\].vdac_batch._6_
timestamp 1698431365
transform -1 0 2912 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[1\].vdac_batch._7_
timestamp 1698431365
transform 1 0 4480 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  temp1.dac.parallel_cells\[1\].vdac_batch._8_
timestamp 1698431365
transform 1 0 5488 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1698431365
transform 1 0 1680 0 -1 62720
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform 1 0 5488 0 1 62720
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1698431365
transform 1 0 1680 0 1 61152
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[1\].vdac_batch.einvp_batch\[1\].vref
timestamp 1698431365
transform 1 0 4928 0 -1 62720
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[2\].vdac_batch._3_
timestamp 1698431365
transform 1 0 7392 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[2\].vdac_batch._4_
timestamp 1698431365
transform 1 0 5488 0 1 58016
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[2\].vdac_batch._5_
timestamp 1698431365
transform 1 0 6048 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  temp1.dac.parallel_cells\[2\].vdac_batch._6_
timestamp 1698431365
transform 1 0 6608 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[2\].vdac_batch._7_
timestamp 1698431365
transform 1 0 5712 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  temp1.dac.parallel_cells\[2\].vdac_batch._8_
timestamp 1698431365
transform 1 0 6160 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1698431365
transform 1 0 7392 0 1 61152
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform 1 0 7280 0 1 56448
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1698431365
transform 1 0 9296 0 1 61152
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[1\].vref
timestamp 1698431365
transform 1 0 9856 0 1 56448
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1698431365
transform 1 0 7280 0 -1 61152
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[2\].vref
timestamp 1698431365
transform -1 0 9184 0 1 54880
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1698431365
transform 1 0 8064 0 1 62720
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[2\].vdac_batch.einvp_batch\[3\].vref
timestamp 1698431365
transform -1 0 9184 0 -1 58016
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  temp1.dac.parallel_cells\[3\].vdac_batch._3_
timestamp 1698431365
transform -1 0 6160 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[3\].vdac_batch._4_
timestamp 1698431365
transform -1 0 6944 0 1 67424
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[3\].vdac_batch._5_
timestamp 1698431365
transform 1 0 3696 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  temp1.dac.parallel_cells\[3\].vdac_batch._6_
timestamp 1698431365
transform -1 0 4928 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[3\].vdac_batch._7_
timestamp 1698431365
transform -1 0 5936 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  temp1.dac.parallel_cells\[3\].vdac_batch._8_
timestamp 1698431365
transform -1 0 6608 0 -1 70560
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1698431365
transform 1 0 1568 0 1 72128
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform 1 0 6608 0 -1 70560
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1698431365
transform 1 0 1568 0 1 76832
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[1\].vref
timestamp 1698431365
transform 1 0 5936 0 -1 75264
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1698431365
transform 1 0 2464 0 -1 72128
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[2\].vref
timestamp 1698431365
transform 1 0 6048 0 1 75264
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1698431365
transform 1 0 2912 0 1 75264
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[3\].vref
timestamp 1698431365
transform 1 0 5824 0 1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1698431365
transform 1 0 1680 0 -1 76832
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[4\].vref
timestamp 1698431365
transform 1 0 6272 0 1 70560
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1698431365
transform 1 0 2128 0 1 70560
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[5\].vref
timestamp 1698431365
transform -1 0 6160 0 -1 76832
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1698431365
transform 1 0 1568 0 -1 78400
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_4  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[6\].vref open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6160 0 -1 76832
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1698431365
transform 1 0 2912 0 -1 75264
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[3\].vdac_batch.einvp_batch\[7\].vref
timestamp 1698431365
transform 1 0 6160 0 -1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__inv_3  temp1.dac.parallel_cells\[4\].vdac_batch._3_
timestamp 1698431365
transform 1 0 9408 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.parallel_cells\[4\].vdac_batch._4_
timestamp 1698431365
transform 1 0 6048 0 1 65856
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.parallel_cells\[4\].vdac_batch._5_
timestamp 1698431365
transform 1 0 7504 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  temp1.dac.parallel_cells\[4\].vdac_batch._6_
timestamp 1698431365
transform 1 0 8400 0 1 65856
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.parallel_cells\[4\].vdac_batch._7_
timestamp 1698431365
transform 1 0 6720 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  temp1.dac.parallel_cells\[4\].vdac_batch._8_
timestamp 1698431365
transform -1 0 9184 0 -1 67424
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].pupd
timestamp 1698431365
transform 1 0 13328 0 1 65856
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[0\].vref
timestamp 1698431365
transform 1 0 10528 0 1 73696
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].pupd
timestamp 1698431365
transform 1 0 13328 0 1 61152
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[1\].vref
timestamp 1698431365
transform 1 0 9408 0 -1 75264
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].pupd
timestamp 1698431365
transform 1 0 9296 0 1 64288
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[2\].vref
timestamp 1698431365
transform 1 0 9408 0 -1 73696
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].pupd
timestamp 1698431365
transform -1 0 12768 0 1 65856
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[3\].vref
timestamp 1698431365
transform 1 0 12880 0 -1 76832
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].pupd
timestamp 1698431365
transform 1 0 10528 0 -1 64288
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[4\].vref
timestamp 1698431365
transform 1 0 10304 0 -1 76832
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].pupd
timestamp 1698431365
transform 1 0 12656 0 -1 58016
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[5\].vref
timestamp 1698431365
transform 1 0 12208 0 -1 70560
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].pupd
timestamp 1698431365
transform 1 0 12656 0 -1 59584
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[6\].vref
timestamp 1698431365
transform 1 0 9744 0 1 75264
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].pupd
timestamp 1698431365
transform 1 0 13328 0 1 58016
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[7\].vref
timestamp 1698431365
transform 1 0 10528 0 1 70560
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].pupd
timestamp 1698431365
transform 1 0 10080 0 -1 62720
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[8\].vref
timestamp 1698431365
transform 1 0 9408 0 -1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].pupd
timestamp 1698431365
transform 1 0 10528 0 -1 59584
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[9\].vref
timestamp 1698431365
transform 1 0 8512 0 1 67424
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].pupd
timestamp 1698431365
transform 1 0 10528 0 1 58016
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[10\].vref
timestamp 1698431365
transform -1 0 10080 0 1 76832
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].pupd
timestamp 1698431365
transform 1 0 12992 0 -1 65856
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[11\].vref
timestamp 1698431365
transform -1 0 11984 0 -1 67424
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].pupd
timestamp 1698431365
transform 1 0 13328 0 1 62720
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[12\].vref
timestamp 1698431365
transform 1 0 10528 0 1 68992
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].pupd
timestamp 1698431365
transform 1 0 12880 0 -1 62720
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[13\].vref
timestamp 1698431365
transform 1 0 11984 0 -1 73696
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].pupd
timestamp 1698431365
transform 1 0 10640 0 -1 65856
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[14\].vref
timestamp 1698431365
transform 1 0 9632 0 -1 70560
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].pupd
timestamp 1698431365
transform -1 0 12432 0 -1 58016
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_3  temp1.dac.parallel_cells\[4\].vdac_batch.einvp_batch\[15\].vref
timestamp 1698431365
transform 1 0 8960 0 1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp1.dac.vdac_single._3__19 open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3248 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  temp1.dac.vdac_single._3_
timestamp 1698431365
transform 1 0 2576 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp1.dac.vdac_single._4__20
timestamp 1698431365
transform -1 0 2800 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  temp1.dac.vdac_single._4__21
timestamp 1698431365
transform -1 0 3696 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  temp1.dac.vdac_single._4_
timestamp 1698431365
transform 1 0 1904 0 1 65856
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  temp1.dac.vdac_single._5_
timestamp 1698431365
transform -1 0 3360 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  temp1.dac.vdac_single._6_
timestamp 1698431365
transform -1 0 2464 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  temp1.dac.vdac_single._7_
timestamp 1698431365
transform 1 0 3472 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  temp1.dac.vdac_single._8_
timestamp 1698431365
transform 1 0 3360 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__invz_2  temp1.dac.vdac_single.einvp_batch\[0\].pupd
timestamp 1698431365
transform 1 0 1568 0 -1 67424
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  temp1.dac.vdac_single.einvp_batch\[0\].vref open_design_environment/foundry/pdks/GF180/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3920 0 -1 67424
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__invz_1  temp1.dcdc
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  temp1.inv1_2
timestamp 1698431365
transform 1 0 1792 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  temp1.inv2_3
timestamp 1698431365
transform -1 0 4368 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  temp1.inv2_4
timestamp 1698431365
transform -1 0 3920 0 1 45472
box -86 -86 534 870
<< labels >>
flabel metal4 s 4448 1508 4768 78460 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 35168 1508 35488 78460 0 FreeSans 1280 90 0 0 VDD
port 0 nsew power bidirectional
flabel metal4 s 19808 1508 20128 78460 0 FreeSans 1280 90 0 0 VSS
port 1 nsew ground bidirectional
flabel metal3 s 0 2912 400 3024 0 FreeSans 448 0 0 0 io_in[0]
port 2 nsew signal input
flabel metal3 s 0 7840 400 7952 0 FreeSans 448 0 0 0 io_in[1]
port 3 nsew signal input
flabel metal3 s 0 12768 400 12880 0 FreeSans 448 0 0 0 io_in[2]
port 4 nsew signal input
flabel metal3 s 0 17696 400 17808 0 FreeSans 448 0 0 0 io_in[3]
port 5 nsew signal input
flabel metal3 s 0 22624 400 22736 0 FreeSans 448 0 0 0 io_in[4]
port 6 nsew signal input
flabel metal3 s 0 27552 400 27664 0 FreeSans 448 0 0 0 io_in[5]
port 7 nsew signal input
flabel metal3 s 0 32480 400 32592 0 FreeSans 448 0 0 0 io_in[6]
port 8 nsew signal input
flabel metal3 s 0 37408 400 37520 0 FreeSans 448 0 0 0 io_in[7]
port 9 nsew signal input
flabel metal3 s 0 42336 400 42448 0 FreeSans 448 0 0 0 io_out[0]
port 10 nsew signal tristate
flabel metal3 s 0 47264 400 47376 0 FreeSans 448 0 0 0 io_out[1]
port 11 nsew signal tristate
flabel metal3 s 0 52192 400 52304 0 FreeSans 448 0 0 0 io_out[2]
port 12 nsew signal tristate
flabel metal3 s 0 57120 400 57232 0 FreeSans 448 0 0 0 io_out[3]
port 13 nsew signal tristate
flabel metal3 s 0 62048 400 62160 0 FreeSans 448 0 0 0 io_out[4]
port 14 nsew signal tristate
flabel metal3 s 0 66976 400 67088 0 FreeSans 448 0 0 0 io_out[5]
port 15 nsew signal tristate
flabel metal3 s 0 71904 400 72016 0 FreeSans 448 0 0 0 io_out[6]
port 16 nsew signal tristate
flabel metal3 s 0 76832 400 76944 0 FreeSans 448 0 0 0 io_out[7]
port 17 nsew signal tristate
rlabel metal1 24976 77616 24976 77616 0 VDD
rlabel metal1 24976 78400 24976 78400 0 VSS
rlabel metal2 11592 19488 11592 19488 0 _0000_
rlabel metal2 13720 20328 13720 20328 0 _0001_
rlabel metal2 16072 23968 16072 23968 0 _0002_
rlabel metal2 15176 25984 15176 25984 0 _0003_
rlabel metal3 16744 29512 16744 29512 0 _0004_
rlabel metal2 14168 31304 14168 31304 0 _0005_
rlabel metal2 15064 53984 15064 53984 0 _0006_
rlabel metal3 17696 63224 17696 63224 0 _0007_
rlabel metal2 18144 62216 18144 62216 0 _0008_
rlabel metal2 21336 54992 21336 54992 0 _0009_
rlabel metal2 25928 53032 25928 53032 0 _0010_
rlabel metal2 30968 54208 30968 54208 0 _0011_
rlabel metal2 35224 55104 35224 55104 0 _0012_
rlabel metal2 38472 57904 38472 57904 0 _0013_
rlabel metal2 40376 61040 40376 61040 0 _0014_
rlabel metal2 41272 60424 41272 60424 0 _0015_
rlabel metal2 42168 56504 42168 56504 0 _0016_
rlabel metal2 29288 53816 29288 53816 0 _0017_
rlabel metal2 33432 60032 33432 60032 0 _0018_
rlabel metal3 35336 70056 35336 70056 0 _0019_
rlabel metal2 37800 71288 37800 71288 0 _0020_
rlabel metal3 32368 71960 32368 71960 0 _0021_
rlabel metal2 30072 72856 30072 72856 0 _0022_
rlabel metal2 26488 50120 26488 50120 0 _0023_
rlabel metal2 17976 51072 17976 51072 0 _0024_
rlabel metal2 14784 51464 14784 51464 0 _0025_
rlabel metal2 14224 47544 14224 47544 0 _0026_
rlabel metal2 15176 43876 15176 43876 0 _0027_
rlabel metal3 18480 39704 18480 39704 0 _0028_
rlabel metal2 18648 36960 18648 36960 0 _0029_
rlabel metal2 15848 33656 15848 33656 0 _0030_
rlabel metal2 15288 7896 15288 7896 0 _0031_
rlabel metal2 18200 9352 18200 9352 0 _0032_
rlabel metal2 20328 19488 20328 19488 0 _0033_
rlabel metal2 22344 25760 22344 25760 0 _0034_
rlabel metal2 23352 29288 23352 29288 0 _0035_
rlabel metal2 19208 32032 19208 32032 0 _0036_
rlabel metal2 19432 73752 19432 73752 0 _0037_
rlabel metal2 19320 76104 19320 76104 0 _0038_
rlabel metal2 22904 76048 22904 76048 0 _0039_
rlabel metal2 25592 75320 25592 75320 0 _0040_
rlabel metal2 27944 76776 27944 76776 0 _0041_
rlabel metal2 30968 76888 30968 76888 0 _0042_
rlabel metal2 34776 76048 34776 76048 0 _0043_
rlabel metal2 35784 74480 35784 74480 0 _0044_
rlabel metal2 33768 75152 33768 75152 0 _0045_
rlabel metal2 30632 73640 30632 73640 0 _0046_
rlabel metal2 28056 68936 28056 68936 0 _0047_
rlabel metal2 30464 68824 30464 68824 0 _0048_
rlabel metal2 32648 68320 32648 68320 0 _0049_
rlabel metal2 33880 64344 33880 64344 0 _0050_
rlabel metal2 30352 64792 30352 64792 0 _0051_
rlabel metal2 29176 62188 29176 62188 0 _0052_
rlabel metal2 30184 57120 30184 57120 0 _0053_
rlabel metal2 27608 11592 27608 11592 0 _0054_
rlabel metal2 25144 8372 25144 8372 0 _0055_
rlabel metal2 21560 6216 21560 6216 0 _0056_
rlabel metal2 22568 13272 22568 13272 0 _0057_
rlabel metal3 25536 18424 25536 18424 0 _0058_
rlabel metal2 24584 25816 24584 25816 0 _0059_
rlabel metal2 27384 12488 27384 12488 0 _0060_
rlabel metal2 20216 11508 20216 11508 0 _0061_
rlabel metal2 20552 7980 20552 7980 0 _0062_
rlabel metal2 21672 17304 21672 17304 0 _0063_
rlabel metal3 24808 20776 24808 20776 0 _0064_
rlabel metal2 24920 22008 24920 22008 0 _0065_
rlabel metal2 16408 21280 16408 21280 0 _0066_
rlabel metal2 15064 13216 15064 13216 0 _0067_
rlabel metal2 15512 11480 15512 11480 0 _0068_
rlabel metal2 18536 25144 18536 25144 0 _0069_
rlabel metal2 21336 30464 21336 30464 0 _0070_
rlabel metal2 23800 33600 23800 33600 0 _0071_
rlabel metal2 16296 30240 16296 30240 0 _0072_
rlabel metal2 14392 16184 14392 16184 0 _0073_
rlabel metal2 15904 17752 15904 17752 0 _0074_
rlabel metal2 18424 27328 18424 27328 0 _0075_
rlabel metal2 21784 35504 21784 35504 0 _0076_
rlabel metal2 23576 44800 23576 44800 0 _0077_
rlabel metal2 22120 47712 22120 47712 0 _0078_
rlabel metal2 19768 60984 19768 60984 0 _0079_
rlabel metal2 22008 60144 22008 60144 0 _0080_
rlabel metal2 23800 61880 23800 61880 0 _0081_
rlabel metal3 25368 60648 25368 60648 0 _0082_
rlabel metal2 26432 65688 26432 65688 0 _0083_
rlabel metal2 17976 67480 17976 67480 0 _0084_
rlabel metal2 18760 69720 18760 69720 0 _0085_
rlabel metal2 21448 71344 21448 71344 0 _0086_
rlabel metal2 23688 71064 23688 71064 0 _0087_
rlabel metal2 25704 69944 25704 69944 0 _0088_
rlabel metal2 27160 59528 27160 59528 0 _0089_
rlabel metal2 18088 59640 18088 59640 0 _0090_
rlabel metal2 16296 58912 16296 58912 0 _0091_
rlabel metal2 17080 54208 17080 54208 0 _0092_
rlabel metal2 20664 52248 20664 52248 0 _0093_
rlabel metal2 23688 50232 23688 50232 0 _0094_
rlabel metal2 26040 32872 26040 32872 0 _0095_
rlabel metal3 36680 31080 36680 31080 0 _0096_
rlabel metal2 41720 27664 41720 27664 0 _0097_
rlabel metal2 43904 24808 43904 24808 0 _0098_
rlabel metal2 45192 23576 45192 23576 0 _0099_
rlabel metal2 43064 23520 43064 23520 0 _0100_
rlabel metal2 42504 20328 42504 20328 0 _0101_
rlabel metal2 44184 17752 44184 17752 0 _0102_
rlabel metal2 42392 16128 42392 16128 0 _0103_
rlabel metal2 41720 14056 41720 14056 0 _0104_
rlabel metal2 40152 14840 40152 14840 0 _0105_
rlabel metal2 33768 16408 33768 16408 0 _0106_
rlabel metal2 23800 36736 23800 36736 0 _0107_
rlabel metal2 15400 39256 15400 39256 0 _0108_
rlabel metal2 16408 48664 16408 48664 0 _0109_
rlabel metal2 16856 46200 16856 46200 0 _0110_
rlabel metal2 18928 43624 18928 43624 0 _0111_
rlabel metal2 22120 41608 22120 41608 0 _0112_
rlabel metal3 25480 40936 25480 40936 0 _0113_
rlabel metal3 37296 43624 37296 43624 0 _0114_
rlabel metal2 40152 46368 40152 46368 0 _0115_
rlabel metal3 45080 46760 45080 46760 0 _0116_
rlabel metal2 46032 36568 46032 36568 0 _0117_
rlabel metal2 40656 28728 40656 28728 0 _0118_
rlabel metal3 38416 26488 38416 26488 0 _0119_
rlabel metal3 32704 23688 32704 23688 0 _0120_
rlabel metal2 34272 9128 34272 9128 0 _0121_
rlabel metal2 36792 7784 36792 7784 0 _0122_
rlabel metal2 39088 3640 39088 3640 0 _0123_
rlabel metal2 35784 3808 35784 3808 0 _0124_
rlabel metal3 33208 4424 33208 4424 0 _0125_
rlabel metal2 18144 4424 18144 4424 0 _0126_
rlabel metal2 13944 4648 13944 4648 0 _0127_
rlabel metal2 16072 3640 16072 3640 0 _0128_
rlabel metal2 20328 3080 20328 3080 0 _0129_
rlabel metal2 23800 4032 23800 4032 0 _0130_
rlabel metal3 25368 4424 25368 4424 0 _0131_
rlabel metal2 27160 7784 27160 7784 0 _0132_
rlabel metal2 27944 3080 27944 3080 0 _0133_
rlabel metal2 30744 3164 30744 3164 0 _0134_
rlabel metal2 30520 6944 30520 6944 0 _0135_
rlabel metal2 32312 8960 32312 8960 0 _0136_
rlabel metal2 31304 32200 31304 32200 0 _0137_
rlabel metal3 35112 34216 35112 34216 0 _0138_
rlabel metal2 36344 41216 36344 41216 0 _0139_
rlabel metal2 41720 41496 41720 41496 0 _0140_
rlabel metal2 44408 40544 44408 40544 0 _0141_
rlabel metal2 40152 38360 40152 38360 0 _0142_
rlabel metal2 36792 38668 36792 38668 0 _0143_
rlabel metal2 37912 35392 37912 35392 0 _0144_
rlabel metal2 40040 33656 40040 33656 0 _0145_
rlabel metal2 43848 32704 43848 32704 0 _0146_
rlabel metal2 45640 31892 45640 31892 0 _0147_
rlabel metal2 45752 28952 45752 28952 0 _0148_
rlabel metal2 40656 24024 40656 24024 0 _0149_
rlabel metal2 27720 20328 27720 20328 0 _0150_
rlabel metal2 28280 15260 28280 15260 0 _0151_
rlabel metal2 30408 12488 30408 12488 0 _0152_
rlabel metal2 33432 15260 33432 15260 0 _0153_
rlabel metal2 31416 17920 31416 17920 0 _0154_
rlabel metal2 31528 25760 31528 25760 0 _0155_
rlabel metal2 27888 64120 27888 64120 0 _0156_
rlabel metal2 21448 65128 21448 65128 0 _0157_
rlabel metal2 22064 64904 22064 64904 0 _0158_
rlabel metal2 23520 64792 23520 64792 0 _0159_
rlabel metal2 26040 56560 26040 56560 0 _0160_
rlabel metal2 27832 23352 27832 23352 0 _0161_
rlabel metal3 31864 20888 31864 20888 0 _0162_
rlabel metal2 34328 18368 34328 18368 0 _0163_
rlabel metal2 37576 12600 37576 12600 0 _0164_
rlabel metal2 38920 17920 38920 17920 0 _0165_
rlabel metal2 35784 22624 35784 22624 0 _0166_
rlabel metal2 34552 31024 34552 31024 0 _0167_
rlabel metal2 36344 53256 36344 53256 0 _0168_
rlabel metal2 39032 54768 39032 54768 0 _0169_
rlabel metal2 42168 54992 42168 54992 0 _0170_
rlabel metal2 43960 52584 43960 52584 0 _0171_
rlabel metal2 38696 51688 38696 51688 0 _0172_
rlabel metal2 33936 46872 33936 46872 0 _0173_
rlabel metal2 37800 47936 37800 47936 0 _0174_
rlabel metal2 38976 48104 38976 48104 0 _0175_
rlabel metal3 42560 49672 42560 49672 0 _0176_
rlabel metal2 44072 44744 44072 44744 0 _0177_
rlabel metal2 44016 35784 44016 35784 0 _0178_
rlabel metal2 33880 51016 33880 51016 0 _0179_
rlabel metal2 35840 58296 35840 58296 0 _0180_
rlabel metal3 37128 66136 37128 66136 0 _0181_
rlabel metal2 39088 63000 39088 63000 0 _0182_
rlabel metal2 37464 61376 37464 61376 0 _0183_
rlabel metal2 31640 59024 31640 59024 0 _0184_
rlabel metal2 33488 55384 33488 55384 0 _0185_
rlabel metal3 37240 22456 37240 22456 0 _0186_
rlabel metal2 39480 19600 39480 19600 0 _0187_
rlabel metal3 41608 9912 41608 9912 0 _0188_
rlabel metal2 39032 10304 39032 10304 0 _0189_
rlabel metal3 34832 11480 34832 11480 0 _0190_
rlabel metal2 34328 27216 34328 27216 0 _0191_
rlabel metal2 11480 41552 11480 41552 0 _0192_
rlabel metal2 9240 36736 9240 36736 0 _0193_
rlabel metal2 11480 43064 11480 43064 0 _0194_
rlabel metal3 11704 32648 11704 32648 0 _0195_
rlabel metal2 12600 38668 12600 38668 0 _0196_
rlabel metal2 9688 32984 9688 32984 0 _0197_
rlabel metal2 2520 41608 2520 41608 0 _0198_
rlabel metal2 11928 53088 11928 53088 0 _0199_
rlabel metal2 2576 49112 2576 49112 0 _0200_
rlabel metal2 8904 43960 8904 43960 0 _0201_
rlabel metal3 8792 45976 8792 45976 0 _0202_
rlabel metal2 8848 50456 8848 50456 0 _0203_
rlabel metal2 10360 51688 10360 51688 0 _0204_
rlabel metal2 11928 47768 11928 47768 0 _0205_
rlabel metal2 9464 42392 9464 42392 0 _0206_
rlabel metal2 2296 22400 2296 22400 0 _0207_
rlabel metal2 2576 18536 2576 18536 0 _0208_
rlabel metal2 2520 13328 2520 13328 0 _0209_
rlabel metal2 2576 3640 2576 3640 0 _0210_
rlabel metal2 2520 5040 2520 5040 0 _0211_
rlabel metal2 4200 4648 4200 4648 0 _0212_
rlabel metal2 27832 76496 27832 76496 0 _0213_
rlabel metal2 30576 75880 30576 75880 0 _0214_
rlabel metal2 28672 69384 28672 69384 0 _0215_
rlabel metal2 30688 68600 30688 68600 0 _0216_
rlabel metal2 33600 67144 33600 67144 0 _0217_
rlabel metal2 33488 64008 33488 64008 0 _0218_
rlabel metal2 30968 64792 30968 64792 0 _0219_
rlabel metal2 30072 62216 30072 62216 0 _0220_
rlabel metal2 29960 56728 29960 56728 0 _0221_
rlabel metal2 28896 15848 28896 15848 0 _0222_
rlabel metal2 24024 9352 24024 9352 0 _0223_
rlabel metal2 22176 6664 22176 6664 0 _0224_
rlabel metal2 23688 13048 23688 13048 0 _0225_
rlabel metal2 25144 18536 25144 18536 0 _0226_
rlabel metal2 25872 12936 25872 12936 0 _0227_
rlabel metal2 20944 11256 20944 11256 0 _0228_
rlabel metal2 21224 9352 21224 9352 0 _0229_
rlabel metal2 21560 16576 21560 16576 0 _0230_
rlabel metal2 22960 19432 22960 19432 0 _0231_
rlabel metal2 17752 22120 17752 22120 0 _0232_
rlabel metal2 15400 13216 15400 13216 0 _0233_
rlabel metal2 16296 12824 16296 12824 0 _0234_
rlabel metal2 18312 24024 18312 24024 0 _0235_
rlabel metal2 21000 29680 21000 29680 0 _0236_
rlabel metal2 23464 33152 23464 33152 0 _0237_
rlabel metal2 17304 31584 17304 31584 0 _0238_
rlabel metal2 14840 17808 14840 17808 0 _0239_
rlabel metal3 17584 26040 17584 26040 0 _0240_
rlabel metal2 16016 17080 16016 17080 0 _0241_
rlabel metal2 17752 26684 17752 26684 0 _0242_
rlabel metal2 21336 34160 21336 34160 0 _0243_
rlabel metal2 23016 45024 23016 45024 0 _0244_
rlabel metal2 22680 46704 22680 46704 0 _0245_
rlabel metal2 26600 65464 26600 65464 0 _0246_
rlabel metal3 22904 67032 22904 67032 0 _0247_
rlabel metal2 27496 59304 27496 59304 0 _0248_
rlabel metal2 29176 58912 29176 58912 0 _0249_
rlabel metal2 17472 57848 17472 57848 0 _0250_
rlabel metal2 17640 54768 17640 54768 0 _0251_
rlabel metal2 20160 52920 20160 52920 0 _0252_
rlabel metal2 23240 51128 23240 51128 0 _0253_
rlabel metal2 25256 33600 25256 33600 0 _0254_
rlabel metal3 23856 2744 23856 2744 0 _0255_
rlabel metal2 29736 31864 29736 31864 0 _0256_
rlabel metal2 40040 28560 40040 28560 0 _0257_
rlabel metal2 44072 26544 44072 26544 0 _0258_
rlabel metal2 44968 24192 44968 24192 0 _0259_
rlabel metal2 42224 24136 42224 24136 0 _0260_
rlabel metal2 42840 21056 42840 21056 0 _0261_
rlabel metal2 44520 18704 44520 18704 0 _0262_
rlabel metal2 24360 36344 24360 36344 0 _0263_
rlabel metal2 15736 38724 15736 38724 0 _0264_
rlabel metal2 24976 41160 24976 41160 0 _0265_
rlabel metal2 32536 41160 32536 41160 0 _0266_
rlabel metal2 39704 45976 39704 45976 0 _0267_
rlabel metal3 43568 47320 43568 47320 0 _0268_
rlabel metal2 45584 39480 45584 39480 0 _0269_
rlabel metal2 40824 35560 40824 35560 0 _0270_
rlabel metal2 37352 26628 37352 26628 0 _0271_
rlabel metal3 32816 23912 32816 23912 0 _0272_
rlabel metal2 33992 12040 33992 12040 0 _0273_
rlabel metal2 36232 8176 36232 8176 0 _0274_
rlabel metal2 37968 5096 37968 5096 0 _0275_
rlabel metal2 35560 4200 35560 4200 0 _0276_
rlabel metal2 33432 3388 33432 3388 0 _0277_
rlabel metal2 18424 4760 18424 4760 0 _0278_
rlabel metal2 14168 4032 14168 4032 0 _0279_
rlabel metal2 16632 4480 16632 4480 0 _0280_
rlabel metal2 19880 3584 19880 3584 0 _0281_
rlabel metal2 23856 2968 23856 2968 0 _0282_
rlabel metal2 24472 4704 24472 4704 0 _0283_
rlabel metal3 27272 6888 27272 6888 0 _0284_
rlabel metal2 28504 3808 28504 3808 0 _0285_
rlabel metal2 30520 3416 30520 3416 0 _0286_
rlabel metal2 31304 6328 31304 6328 0 _0287_
rlabel metal2 32424 9520 32424 9520 0 _0288_
rlabel metal2 45192 29848 45192 29848 0 _0289_
rlabel metal3 34048 34328 34048 34328 0 _0290_
rlabel metal2 37240 37968 37240 37968 0 _0291_
rlabel metal2 37576 36008 37576 36008 0 _0292_
rlabel metal2 27944 21448 27944 21448 0 _0293_
rlabel metal3 39368 65352 39368 65352 0 _0294_
rlabel metal3 28896 15288 28896 15288 0 _0295_
rlabel metal2 29400 13216 29400 13216 0 _0296_
rlabel metal2 33208 15204 33208 15204 0 _0297_
rlabel metal2 31080 17304 31080 17304 0 _0298_
rlabel metal2 31024 25368 31024 25368 0 _0299_
rlabel metal3 28504 63896 28504 63896 0 _0300_
rlabel metal2 31080 22624 31080 22624 0 _0301_
rlabel metal2 35000 19320 35000 19320 0 _0302_
rlabel metal2 37352 12824 37352 12824 0 _0303_
rlabel metal2 38416 17528 38416 17528 0 _0304_
rlabel metal2 35952 21000 35952 21000 0 _0305_
rlabel metal2 36008 52976 36008 52976 0 _0306_
rlabel metal2 34104 46928 34104 46928 0 _0307_
rlabel metal2 36456 47936 36456 47936 0 _0308_
rlabel metal2 35672 58128 35672 58128 0 _0309_
rlabel metal3 36624 64904 36624 64904 0 _0310_
rlabel metal2 38696 64456 38696 64456 0 _0311_
rlabel metal2 37016 62524 37016 62524 0 _0312_
rlabel metal2 32536 61096 32536 61096 0 _0313_
rlabel metal2 33768 56392 33768 56392 0 _0314_
rlabel metal2 38864 40600 38864 40600 0 _0315_
rlabel metal2 3864 42224 3864 42224 0 _0316_
rlabel metal2 3752 40432 3752 40432 0 _0317_
rlabel metal3 9408 37240 9408 37240 0 _0318_
rlabel metal2 12152 41160 12152 41160 0 _0319_
rlabel metal2 8568 37296 8568 37296 0 _0320_
rlabel metal2 10640 42168 10640 42168 0 _0321_
rlabel metal2 11704 34888 11704 34888 0 _0322_
rlabel metal2 11704 38024 11704 38024 0 _0323_
rlabel metal2 10136 32704 10136 32704 0 _0324_
rlabel metal2 2520 42784 2520 42784 0 _0325_
rlabel metal3 7672 42840 7672 42840 0 _0326_
rlabel metal2 6328 45528 6328 45528 0 _0327_
rlabel metal3 8232 48776 8232 48776 0 _0328_
rlabel metal2 11256 51212 11256 51212 0 _0329_
rlabel metal2 10192 47432 10192 47432 0 _0330_
rlabel metal2 11424 47320 11424 47320 0 _0331_
rlabel metal2 9688 40488 9688 40488 0 _0332_
rlabel metal2 2632 22736 2632 22736 0 _0333_
rlabel metal2 3304 19096 3304 19096 0 _0334_
rlabel metal2 2688 17528 2688 17528 0 _0335_
rlabel metal2 2296 18368 2296 18368 0 _0336_
rlabel metal2 3304 13216 3304 13216 0 _0337_
rlabel metal2 2408 10136 2408 10136 0 _0338_
rlabel metal2 3080 9016 3080 9016 0 _0339_
rlabel metal3 1904 6664 1904 6664 0 _0340_
rlabel metal3 3024 8680 3024 8680 0 _0341_
rlabel metal3 2296 6776 2296 6776 0 _0342_
rlabel metal2 3752 14224 3752 14224 0 _0343_
rlabel metal2 8232 34216 8232 34216 0 _0344_
rlabel metal2 6776 52864 6776 52864 0 _0345_
rlabel metal2 3528 52192 3528 52192 0 _0346_
rlabel metal2 2856 44632 2856 44632 0 _0347_
rlabel metal2 8232 48944 8232 48944 0 _0348_
rlabel metal2 9688 46984 9688 46984 0 _0349_
rlabel metal2 9688 40264 9688 40264 0 _0350_
rlabel metal2 2408 24472 2408 24472 0 _0351_
rlabel metal2 2520 17360 2520 17360 0 _0352_
rlabel metal2 3080 7924 3080 7924 0 _0353_
rlabel metal2 4648 7336 4648 7336 0 _0354_
rlabel metal3 25312 47432 25312 47432 0 _0355_
rlabel metal2 20384 47208 20384 47208 0 _0356_
rlabel metal2 1960 28896 1960 28896 0 _0357_
rlabel metal3 40992 30184 40992 30184 0 _0358_
rlabel metal3 23912 41888 23912 41888 0 _0359_
rlabel metal2 22568 20608 22568 20608 0 _0360_
rlabel metal2 30296 20552 30296 20552 0 _0361_
rlabel metal2 18424 42168 18424 42168 0 _0362_
rlabel metal2 24024 46704 24024 46704 0 _0363_
rlabel metal3 30464 40376 30464 40376 0 _0364_
rlabel metal3 19096 40376 19096 40376 0 _0365_
rlabel metal2 26600 46928 26600 46928 0 _0366_
rlabel metal3 32760 21784 32760 21784 0 _0367_
rlabel metal3 26264 5992 26264 5992 0 _0368_
rlabel metal3 29960 49784 29960 49784 0 _0369_
rlabel metal2 31808 18088 31808 18088 0 _0370_
rlabel metal2 29400 17948 29400 17948 0 _0371_
rlabel metal2 18984 21504 18984 21504 0 _0372_
rlabel metal2 23912 5544 23912 5544 0 _0373_
rlabel metal2 19208 14112 19208 14112 0 _0374_
rlabel metal2 19264 4872 19264 4872 0 _0375_
rlabel metal2 23352 68376 23352 68376 0 _0376_
rlabel metal2 24416 19320 24416 19320 0 _0377_
rlabel metal2 24528 41272 24528 41272 0 _0378_
rlabel metal3 25872 22904 25872 22904 0 _0379_
rlabel metal2 21784 13440 21784 13440 0 _0380_
rlabel metal2 33264 39592 33264 39592 0 _0381_
rlabel metal2 33992 40656 33992 40656 0 _0382_
rlabel metal2 19544 23016 19544 23016 0 _0383_
rlabel metal3 24248 39592 24248 39592 0 _0384_
rlabel metal2 25704 46200 25704 46200 0 _0385_
rlabel metal2 22400 20552 22400 20552 0 _0386_
rlabel metal2 21112 15288 21112 15288 0 _0387_
rlabel metal2 20216 21952 20216 21952 0 _0388_
rlabel metal3 39424 21448 39424 21448 0 _0389_
rlabel metal2 20608 39368 20608 39368 0 _0390_
rlabel metal2 41328 30296 41328 30296 0 _0391_
rlabel metal2 35168 21672 35168 21672 0 _0392_
rlabel metal2 39480 21448 39480 21448 0 _0393_
rlabel metal2 19488 41944 19488 41944 0 _0394_
rlabel metal2 38920 21224 38920 21224 0 _0395_
rlabel metal2 32536 49000 32536 49000 0 _0396_
rlabel metal2 40152 20552 40152 20552 0 _0397_
rlabel metal3 41104 17080 41104 17080 0 _0398_
rlabel metal2 36568 21280 36568 21280 0 _0399_
rlabel metal2 38136 24332 38136 24332 0 _0400_
rlabel metal2 39256 51856 39256 51856 0 _0401_
rlabel metal2 38360 66248 38360 66248 0 _0402_
rlabel metal2 31192 43008 31192 43008 0 _0403_
rlabel metal2 34720 75544 34720 75544 0 _0404_
rlabel metal2 30184 46536 30184 46536 0 _0405_
rlabel metal2 41944 38248 41944 38248 0 _0406_
rlabel metal2 34160 69160 34160 69160 0 _0407_
rlabel metal3 34888 69384 34888 69384 0 _0408_
rlabel metal2 35672 69832 35672 69832 0 _0409_
rlabel metal2 36008 67536 36008 67536 0 _0410_
rlabel metal2 37800 46256 37800 46256 0 _0411_
rlabel metal2 19992 57232 19992 57232 0 _0412_
rlabel metal2 38696 31472 38696 31472 0 _0413_
rlabel metal2 25816 49756 25816 49756 0 _0414_
rlabel metal2 18928 57512 18928 57512 0 _0415_
rlabel metal2 20104 57064 20104 57064 0 _0416_
rlabel metal3 22456 63896 22456 63896 0 _0417_
rlabel metal2 26824 55552 26824 55552 0 _0418_
rlabel metal2 23128 56504 23128 56504 0 _0419_
rlabel metal2 23352 56336 23352 56336 0 _0420_
rlabel metal2 21448 68320 21448 68320 0 _0421_
rlabel metal2 26040 70168 26040 70168 0 _0422_
rlabel metal2 21896 68992 21896 68992 0 _0423_
rlabel metal3 19376 68824 19376 68824 0 _0424_
rlabel metal3 22456 68376 22456 68376 0 _0425_
rlabel metal2 16632 47488 16632 47488 0 _0426_
rlabel metal2 20216 48776 20216 48776 0 _0427_
rlabel metal2 20664 49728 20664 49728 0 _0428_
rlabel metal2 19208 53592 19208 53592 0 _0429_
rlabel metal2 22176 56280 22176 56280 0 _0430_
rlabel metal2 38584 38584 38584 38584 0 _0431_
rlabel metal2 41272 41216 41272 41216 0 _0432_
rlabel metal2 26824 23128 26824 23128 0 _0433_
rlabel metal2 39480 40320 39480 40320 0 _0434_
rlabel metal2 39704 33376 39704 33376 0 _0435_
rlabel metal3 43008 30856 43008 30856 0 _0436_
rlabel metal2 38920 32256 38920 32256 0 _0437_
rlabel metal2 40152 33096 40152 33096 0 _0438_
rlabel metal2 38696 53424 38696 53424 0 _0439_
rlabel metal3 43960 51576 43960 51576 0 _0440_
rlabel metal2 41160 52192 41160 52192 0 _0441_
rlabel metal2 38584 56056 38584 56056 0 _0442_
rlabel metal2 39872 52360 39872 52360 0 _0443_
rlabel metal2 38864 46872 38864 46872 0 _0444_
rlabel metal2 42896 38024 42896 38024 0 _0445_
rlabel metal2 38808 44800 38808 44800 0 _0446_
rlabel metal2 38696 43148 38696 43148 0 _0447_
rlabel metal2 34776 43064 34776 43064 0 _0448_
rlabel metal2 20552 22400 20552 22400 0 _0449_
rlabel metal2 16968 23072 16968 23072 0 _0450_
rlabel metal2 7448 24080 7448 24080 0 _0451_
rlabel metal2 30576 21784 30576 21784 0 _0452_
rlabel metal2 30520 14056 30520 14056 0 _0453_
rlabel metal2 29960 10808 29960 10808 0 _0454_
rlabel metal2 23968 21448 23968 21448 0 _0455_
rlabel metal2 18984 12544 18984 12544 0 _0456_
rlabel metal2 18032 12936 18032 12936 0 _0457_
rlabel metal2 20104 13440 20104 13440 0 _0458_
rlabel metal2 19880 13384 19880 13384 0 _0459_
rlabel metal2 21672 20832 21672 20832 0 _0460_
rlabel metal2 39928 16016 39928 16016 0 _0461_
rlabel metal2 41160 16576 41160 16576 0 _0462_
rlabel metal2 39368 16576 39368 16576 0 _0463_
rlabel metal2 39536 27944 39536 27944 0 _0464_
rlabel metal3 35336 73080 35336 73080 0 _0465_
rlabel metal3 37968 71736 37968 71736 0 _0466_
rlabel metal2 36120 70112 36120 70112 0 _0467_
rlabel metal2 38584 47096 38584 47096 0 _0468_
rlabel metal2 17976 62328 17976 62328 0 _0469_
rlabel metal2 19432 57512 19432 57512 0 _0470_
rlabel metal2 19880 57400 19880 57400 0 _0471_
rlabel metal2 21896 65240 21896 65240 0 _0472_
rlabel metal3 22344 59752 22344 59752 0 _0473_
rlabel metal2 22792 58352 22792 58352 0 _0474_
rlabel metal2 21504 73976 21504 73976 0 _0475_
rlabel metal2 21000 69664 21000 69664 0 _0476_
rlabel metal2 22456 58212 22456 58212 0 _0477_
rlabel metal3 18256 48776 18256 48776 0 _0478_
rlabel metal2 19544 48496 19544 48496 0 _0479_
rlabel metal2 20776 49644 20776 49644 0 _0480_
rlabel metal2 22456 53928 22456 53928 0 _0481_
rlabel metal2 40264 42000 40264 42000 0 _0482_
rlabel metal2 41944 42952 41944 42952 0 _0483_
rlabel metal2 43288 33040 43288 33040 0 _0484_
rlabel metal2 42616 32648 42616 32648 0 _0485_
rlabel metal2 43904 38024 43904 38024 0 _0486_
rlabel metal2 42280 54376 42280 54376 0 _0487_
rlabel metal2 40768 58296 40768 58296 0 _0488_
rlabel metal2 40936 53144 40936 53144 0 _0489_
rlabel metal2 41720 48104 41720 48104 0 _0490_
rlabel metal2 40936 47712 40936 47712 0 _0491_
rlabel metal2 41160 47152 41160 47152 0 _0492_
rlabel metal2 36232 46816 36232 46816 0 _0493_
rlabel metal2 23464 20888 23464 20888 0 _0494_
rlabel metal2 18536 22064 18536 22064 0 _0495_
rlabel metal2 11256 23632 11256 23632 0 _0496_
rlabel metal2 31640 13496 31640 13496 0 _0497_
rlabel metal2 31080 11872 31080 11872 0 _0498_
rlabel metal2 24696 24136 24696 24136 0 _0499_
rlabel metal2 20720 15400 20720 15400 0 _0500_
rlabel metal2 20216 6104 20216 6104 0 _0501_
rlabel metal2 22624 15288 22624 15288 0 _0502_
rlabel metal2 19432 16408 19432 16408 0 _0503_
rlabel metal2 22904 24136 22904 24136 0 _0504_
rlabel metal2 39144 12264 39144 12264 0 _0505_
rlabel metal2 40264 13944 40264 13944 0 _0506_
rlabel metal2 38696 14616 38696 14616 0 _0507_
rlabel metal2 38920 20160 38920 20160 0 _0508_
rlabel metal2 37016 74648 37016 74648 0 _0509_
rlabel metal2 38808 71008 38808 71008 0 _0510_
rlabel metal2 36232 70224 36232 70224 0 _0511_
rlabel metal2 38472 43176 38472 43176 0 _0512_
rlabel metal2 20216 58688 20216 58688 0 _0513_
rlabel metal2 19544 54992 19544 54992 0 _0514_
rlabel metal3 23072 55160 23072 55160 0 _0515_
rlabel metal2 24584 64904 24584 64904 0 _0516_
rlabel metal2 23856 62440 23856 62440 0 _0517_
rlabel metal2 24696 57176 24696 57176 0 _0518_
rlabel metal2 23464 72912 23464 72912 0 _0519_
rlabel metal2 24472 70784 24472 70784 0 _0520_
rlabel metal2 24304 69944 24304 69944 0 _0521_
rlabel metal2 19320 45304 19320 45304 0 _0522_
rlabel metal2 20440 46368 20440 46368 0 _0523_
rlabel metal3 21448 46536 21448 46536 0 _0524_
rlabel metal2 23856 41384 23856 41384 0 _0525_
rlabel metal2 44296 41664 44296 41664 0 _0526_
rlabel metal2 43624 42672 43624 42672 0 _0527_
rlabel metal2 45080 32592 45080 32592 0 _0528_
rlabel metal2 43064 30296 43064 30296 0 _0529_
rlabel metal2 43848 32984 43848 32984 0 _0530_
rlabel metal2 44016 52136 44016 52136 0 _0531_
rlabel metal2 41384 53816 41384 53816 0 _0532_
rlabel metal2 42784 51128 42784 51128 0 _0533_
rlabel metal3 44464 44296 44464 44296 0 _0534_
rlabel metal2 41608 44576 41608 44576 0 _0535_
rlabel metal2 42840 43904 42840 43904 0 _0536_
rlabel metal2 36120 42896 36120 42896 0 _0537_
rlabel metal2 23016 24640 23016 24640 0 _0538_
rlabel metal2 12824 24640 12824 24640 0 _0539_
rlabel metal2 10808 25032 10808 25032 0 _0540_
rlabel metal2 30856 16688 30856 16688 0 _0541_
rlabel metal2 30688 16856 30688 16856 0 _0542_
rlabel metal2 23744 21224 23744 21224 0 _0543_
rlabel metal2 23072 20888 23072 20888 0 _0544_
rlabel metal3 23856 4984 23856 4984 0 _0545_
rlabel metal2 22792 22064 22792 22064 0 _0546_
rlabel metal2 22232 24136 22232 24136 0 _0547_
rlabel metal3 24976 22904 24976 22904 0 _0548_
rlabel metal3 37408 11368 37408 11368 0 _0549_
rlabel metal2 33992 16016 33992 16016 0 _0550_
rlabel metal3 36344 15960 36344 15960 0 _0551_
rlabel metal2 37912 21000 37912 21000 0 _0552_
rlabel metal2 33544 73976 33544 73976 0 _0553_
rlabel metal2 32984 72072 32984 72072 0 _0554_
rlabel metal2 33320 68992 33320 68992 0 _0555_
rlabel metal3 36960 37240 36960 37240 0 _0556_
rlabel metal3 24752 54600 24752 54600 0 _0557_
rlabel metal2 24136 53424 24136 53424 0 _0558_
rlabel metal3 25088 53592 25088 53592 0 _0559_
rlabel metal2 25536 65240 25536 65240 0 _0560_
rlabel metal2 26376 61152 26376 61152 0 _0561_
rlabel metal2 26376 55552 26376 55552 0 _0562_
rlabel metal2 25424 74984 25424 74984 0 _0563_
rlabel metal2 26152 70448 26152 70448 0 _0564_
rlabel metal2 26824 66052 26824 66052 0 _0565_
rlabel metal2 21448 42336 21448 42336 0 _0566_
rlabel metal2 20944 45080 20944 45080 0 _0567_
rlabel metal3 23352 52136 23352 52136 0 _0568_
rlabel metal2 25424 44520 25424 44520 0 _0569_
rlabel metal3 44520 39592 44520 39592 0 _0570_
rlabel metal2 44184 37856 44184 37856 0 _0571_
rlabel metal3 45920 30968 45920 30968 0 _0572_
rlabel metal2 44408 30688 44408 30688 0 _0573_
rlabel metal2 44968 37240 44968 37240 0 _0574_
rlabel metal3 42392 52192 42392 52192 0 _0575_
rlabel metal2 41720 52192 41720 52192 0 _0576_
rlabel metal2 43456 52360 43456 52360 0 _0577_
rlabel metal2 44072 38248 44072 38248 0 _0578_
rlabel metal3 43064 37800 43064 37800 0 _0579_
rlabel metal2 43064 37576 43064 37576 0 _0580_
rlabel metal2 33992 37408 33992 37408 0 _0581_
rlabel metal2 26152 22456 26152 22456 0 _0582_
rlabel metal2 11704 22456 11704 22456 0 _0583_
rlabel metal2 10920 22008 10920 22008 0 _0584_
rlabel metal3 11760 30744 11760 30744 0 _0585_
rlabel metal2 30968 45248 30968 45248 0 _0586_
rlabel metal2 29288 43904 29288 43904 0 _0587_
rlabel metal2 29624 39480 29624 39480 0 _0588_
rlabel metal2 26488 36848 26488 36848 0 _0589_
rlabel metal2 26376 38668 26376 38668 0 _0590_
rlabel metal2 26488 38864 26488 38864 0 _0591_
rlabel metal2 27496 42000 27496 42000 0 _0592_
rlabel metal2 27832 43400 27832 43400 0 _0593_
rlabel metal2 26824 38528 26824 38528 0 _0594_
rlabel metal2 26208 34328 26208 34328 0 _0595_
rlabel metal2 26152 40264 26152 40264 0 _0596_
rlabel metal2 26936 39144 26936 39144 0 _0597_
rlabel metal3 27720 38808 27720 38808 0 _0598_
rlabel metal2 30856 49896 30856 49896 0 _0599_
rlabel via2 30408 49784 30408 49784 0 _0600_
rlabel metal2 29176 46424 29176 46424 0 _0601_
rlabel metal2 28392 44632 28392 44632 0 _0602_
rlabel metal2 27272 45360 27272 45360 0 _0603_
rlabel metal3 29400 40936 29400 40936 0 _0604_
rlabel metal3 29792 41272 29792 41272 0 _0605_
rlabel metal2 29960 46424 29960 46424 0 _0606_
rlabel metal2 30184 44688 30184 44688 0 _0607_
rlabel metal2 32424 22232 32424 22232 0 _0608_
rlabel metal2 33544 30128 33544 30128 0 _0609_
rlabel metal2 37016 25508 37016 25508 0 _0610_
rlabel metal2 33376 28728 33376 28728 0 _0611_
rlabel metal2 27272 24472 27272 24472 0 _0612_
rlabel metal2 34048 49448 34048 49448 0 _0613_
rlabel metal3 32872 28840 32872 28840 0 _0614_
rlabel metal3 35672 27832 35672 27832 0 _0615_
rlabel metal3 36456 28616 36456 28616 0 _0616_
rlabel metal3 35448 28672 35448 28672 0 _0617_
rlabel metal2 47208 27272 47208 27272 0 _0618_
rlabel metal2 41720 29064 41720 29064 0 _0619_
rlabel metal2 33992 29008 33992 29008 0 _0620_
rlabel metal2 30464 27944 30464 27944 0 _0621_
rlabel metal2 25872 23352 25872 23352 0 _0622_
rlabel metal2 27048 27608 27048 27608 0 _0623_
rlabel metal2 26208 27944 26208 27944 0 _0624_
rlabel metal2 37016 42336 37016 42336 0 _0625_
rlabel metal2 35000 37128 35000 37128 0 _0626_
rlabel metal2 34608 40712 34608 40712 0 _0627_
rlabel metal3 28840 27832 28840 27832 0 _0628_
rlabel metal2 27832 27440 27832 27440 0 _0629_
rlabel metal2 27048 19768 27048 19768 0 _0630_
rlabel metal2 28280 27496 28280 27496 0 _0631_
rlabel metal2 33152 25368 33152 25368 0 _0632_
rlabel metal2 32648 26040 32648 26040 0 _0633_
rlabel metal4 30520 33152 30520 33152 0 _0634_
rlabel metal2 11480 30744 11480 30744 0 _0635_
rlabel metal2 13384 29736 13384 29736 0 _0636_
rlabel metal3 11816 29400 11816 29400 0 _0637_
rlabel metal2 9912 28840 9912 28840 0 _0638_
rlabel metal2 36232 29288 36232 29288 0 _0639_
rlabel metal2 29512 33432 29512 33432 0 _0640_
rlabel metal2 30072 32256 30072 32256 0 _0641_
rlabel metal2 30744 34048 30744 34048 0 _0642_
rlabel metal2 31528 32256 31528 32256 0 _0643_
rlabel metal2 30576 32648 30576 32648 0 _0644_
rlabel metal3 29904 33432 29904 33432 0 _0645_
rlabel metal2 30184 32424 30184 32424 0 _0646_
rlabel metal3 28784 23912 28784 23912 0 _0647_
rlabel metal3 28112 27608 28112 27608 0 _0648_
rlabel metal2 28616 32200 28616 32200 0 _0649_
rlabel metal3 27440 44072 27440 44072 0 _0650_
rlabel metal3 26880 30408 26880 30408 0 _0651_
rlabel metal2 26712 31752 26712 31752 0 _0652_
rlabel metal2 29568 26824 29568 26824 0 _0653_
rlabel metal2 29400 28336 29400 28336 0 _0654_
rlabel metal3 28448 32648 28448 32648 0 _0655_
rlabel metal2 30296 35728 30296 35728 0 _0656_
rlabel metal3 33264 42840 33264 42840 0 _0657_
rlabel metal2 35728 49224 35728 49224 0 _0658_
rlabel metal2 35000 49560 35000 49560 0 _0659_
rlabel metal2 35560 43008 35560 43008 0 _0660_
rlabel metal2 35784 40684 35784 40684 0 _0661_
rlabel metal2 36120 36960 36120 36960 0 _0662_
rlabel metal3 29064 36456 29064 36456 0 _0663_
rlabel metal2 30184 29008 30184 29008 0 _0664_
rlabel metal2 27496 36680 27496 36680 0 _0665_
rlabel metal2 27048 11480 27048 11480 0 _0666_
rlabel metal2 26936 36512 26936 36512 0 _0667_
rlabel metal2 27608 36960 27608 36960 0 _0668_
rlabel metal2 29624 36960 29624 36960 0 _0669_
rlabel metal2 15624 27944 15624 27944 0 _0670_
rlabel metal2 11928 28280 11928 28280 0 _0671_
rlabel metal2 6440 52472 6440 52472 0 _0672_
rlabel metal2 3752 50624 3752 50624 0 _0673_
rlabel metal2 3248 23800 3248 23800 0 _0674_
rlabel metal2 4312 19656 4312 19656 0 _0675_
rlabel metal2 3192 16632 3192 16632 0 _0676_
rlabel metal2 3192 29624 3192 29624 0 _0677_
rlabel metal3 3472 51240 3472 51240 0 _0678_
rlabel metal2 7616 51352 7616 51352 0 _0679_
rlabel metal2 3752 53256 3752 53256 0 _0680_
rlabel metal2 2968 30632 2968 30632 0 _0681_
rlabel metal2 2184 26992 2184 26992 0 _0682_
rlabel metal2 2856 34608 2856 34608 0 _0683_
rlabel metal2 2352 35112 2352 35112 0 _0684_
rlabel metal2 1960 43400 1960 43400 0 _0685_
rlabel metal2 2968 27832 2968 27832 0 _0686_
rlabel metal2 2296 37576 2296 37576 0 _0687_
rlabel metal3 4256 34216 4256 34216 0 _0688_
rlabel metal3 2828 23912 2828 23912 0 _0689_
rlabel metal3 6552 24808 6552 24808 0 _0690_
rlabel metal2 2744 27888 2744 27888 0 _0691_
rlabel metal2 5992 27440 5992 27440 0 _0692_
rlabel metal2 3752 26572 3752 26572 0 _0693_
rlabel metal2 5264 27832 5264 27832 0 _0694_
rlabel metal2 5320 28672 5320 28672 0 _0695_
rlabel metal2 7448 43008 7448 43008 0 _0696_
rlabel metal2 6048 23352 6048 23352 0 _0697_
rlabel metal2 4984 29400 4984 29400 0 _0698_
rlabel metal2 5656 29848 5656 29848 0 _0699_
rlabel metal2 4872 35840 4872 35840 0 _0700_
rlabel metal2 3528 38724 3528 38724 0 _0701_
rlabel metal2 3192 39312 3192 39312 0 _0702_
rlabel metal2 2968 36512 2968 36512 0 _0703_
rlabel metal2 2800 38024 2800 38024 0 _0704_
rlabel metal2 4760 42504 4760 42504 0 _0705_
rlabel metal2 5152 39816 5152 39816 0 _0706_
rlabel metal2 3192 40880 3192 40880 0 _0707_
rlabel metal2 3192 47152 3192 47152 0 _0708_
rlabel metal2 4088 52752 4088 52752 0 _0709_
rlabel metal2 2520 47712 2520 47712 0 _0710_
rlabel metal2 9800 24248 9800 24248 0 _0711_
rlabel metal2 8568 23408 8568 23408 0 _0712_
rlabel metal3 8512 24696 8512 24696 0 _0713_
rlabel metal3 9688 25816 9688 25816 0 _0714_
rlabel metal2 3976 24360 3976 24360 0 _0715_
rlabel metal2 4424 32312 4424 32312 0 _0716_
rlabel metal2 4312 34496 4312 34496 0 _0717_
rlabel metal2 3304 37912 3304 37912 0 _0718_
rlabel metal3 2856 47320 2856 47320 0 _0719_
rlabel metal2 7672 23128 7672 23128 0 _0720_
rlabel metal2 6440 23408 6440 23408 0 _0721_
rlabel metal3 6440 23240 6440 23240 0 _0722_
rlabel metal2 8120 24696 8120 24696 0 _0723_
rlabel metal3 6160 23128 6160 23128 0 _0724_
rlabel metal2 5040 24920 5040 24920 0 _0725_
rlabel metal2 5936 34328 5936 34328 0 _0726_
rlabel metal2 6104 36568 6104 36568 0 _0727_
rlabel metal2 5600 44520 5600 44520 0 _0728_
rlabel metal2 5096 53144 5096 53144 0 _0729_
rlabel metal2 4816 52360 4816 52360 0 _0730_
rlabel metal2 5992 53536 5992 53536 0 _0731_
rlabel metal2 2744 10696 2744 10696 0 _0733_
rlabel metal3 9128 25256 9128 25256 0 _0734_
rlabel metal2 8232 23184 8232 23184 0 _0735_
rlabel metal2 8848 24472 8848 24472 0 _0736_
rlabel metal2 8568 26152 8568 26152 0 _0737_
rlabel metal3 7784 25480 7784 25480 0 _0738_
rlabel metal2 8232 26544 8232 26544 0 _0739_
rlabel metal2 6888 34216 6888 34216 0 _0740_
rlabel metal2 7672 39508 7672 39508 0 _0741_
rlabel metal2 7056 53704 7056 53704 0 _0742_
rlabel metal2 7224 54488 7224 54488 0 _0743_
rlabel metal3 6832 23800 6832 23800 0 _0744_
rlabel metal3 8344 23912 8344 23912 0 _0745_
rlabel metal2 5600 22904 5600 22904 0 _0746_
rlabel metal2 6328 23632 6328 23632 0 _0747_
rlabel metal2 6776 24248 6776 24248 0 _0748_
rlabel metal2 6608 24920 6608 24920 0 _0749_
rlabel metal2 6160 33320 6160 33320 0 _0750_
rlabel metal3 7224 35896 7224 35896 0 _0751_
rlabel metal2 3920 49896 3920 49896 0 _0752_
rlabel metal2 3640 53760 3640 53760 0 _0753_
rlabel metal2 8904 21000 8904 21000 0 _0754_
rlabel metal2 11032 29680 11032 29680 0 _0755_
rlabel metal2 8568 29512 8568 29512 0 _0756_
rlabel metal3 7952 30072 7952 30072 0 _0757_
rlabel metal2 7168 29624 7168 29624 0 _0758_
rlabel metal3 7000 30184 7000 30184 0 _0759_
rlabel metal2 7448 30296 7448 30296 0 _0760_
rlabel metal3 6832 32536 6832 32536 0 _0761_
rlabel metal2 7392 37016 7392 37016 0 _0762_
rlabel metal2 3640 42504 3640 42504 0 _0763_
rlabel metal2 4536 47040 4536 47040 0 _0764_
rlabel metal2 10248 27552 10248 27552 0 _0765_
rlabel metal2 6328 29120 6328 29120 0 _0766_
rlabel metal2 5656 30688 5656 30688 0 _0767_
rlabel metal2 6440 34160 6440 34160 0 _0768_
rlabel metal2 6328 37128 6328 37128 0 _0769_
rlabel metal2 3024 53816 3024 53816 0 _0770_
rlabel metal2 4200 53424 4200 53424 0 _0771_
rlabel metal2 2856 28056 2856 28056 0 _0772_
rlabel metal2 3640 29680 3640 29680 0 _0773_
rlabel metal3 2520 36960 2520 36960 0 _0774_
rlabel metal3 3416 37912 3416 37912 0 _0775_
rlabel metal2 1736 38388 1736 38388 0 _0776_
rlabel metal2 2408 39984 2408 39984 0 _0777_
rlabel metal2 2856 45864 2856 45864 0 _0778_
rlabel metal2 15512 6160 15512 6160 0 _0779_
rlabel metal3 41720 50456 41720 50456 0 _0780_
rlabel metal2 11368 18928 11368 18928 0 _0781_
rlabel metal2 38920 39368 38920 39368 0 _0782_
rlabel metal2 1848 6664 1848 6664 0 _0783_
rlabel metal2 14336 20776 14336 20776 0 _0784_
rlabel metal2 15064 23576 15064 23576 0 _0785_
rlabel metal2 15232 24136 15232 24136 0 _0786_
rlabel metal2 16632 29120 16632 29120 0 _0787_
rlabel metal2 13496 31024 13496 31024 0 _0788_
rlabel metal2 14952 52248 14952 52248 0 _0789_
rlabel metal2 26376 71400 26376 71400 0 _0790_
rlabel metal2 25368 23128 25368 23128 0 _0791_
rlabel metal3 29960 53928 29960 53928 0 _0792_
rlabel metal2 34216 54208 34216 54208 0 _0793_
rlabel metal2 28952 54432 28952 54432 0 _0794_
rlabel metal2 32368 53144 32368 53144 0 _0795_
rlabel metal2 26936 50512 26936 50512 0 _0796_
rlabel metal2 26824 50288 26824 50288 0 _0797_
rlabel metal2 14000 50792 14000 50792 0 _0798_
rlabel metal2 14392 48496 14392 48496 0 _0799_
rlabel metal2 15792 44184 15792 44184 0 _0800_
rlabel metal2 19208 41048 19208 41048 0 _0801_
rlabel metal2 22792 23632 22792 23632 0 _0802_
rlabel metal2 19432 37576 19432 37576 0 _0803_
rlabel metal3 17976 35112 17976 35112 0 _0804_
rlabel metal2 22176 8344 22176 8344 0 _0805_
rlabel metal2 15624 7980 15624 7980 0 _0806_
rlabel metal2 18312 9072 18312 9072 0 _0807_
rlabel metal2 20216 18816 20216 18816 0 _0808_
rlabel metal2 21784 24752 21784 24752 0 _0809_
rlabel metal2 23576 27944 23576 27944 0 _0810_
rlabel metal2 19096 31248 19096 31248 0 _0811_
rlabel metal2 42840 24192 42840 24192 0 cal_lut\[100\]
rlabel metal3 41496 23016 41496 23016 0 cal_lut\[101\]
rlabel metal2 44408 19600 44408 19600 0 cal_lut\[102\]
rlabel metal2 46312 17136 46312 17136 0 cal_lut\[103\]
rlabel metal2 44520 15568 44520 15568 0 cal_lut\[104\]
rlabel metal2 43848 14000 43848 14000 0 cal_lut\[105\]
rlabel metal2 42280 14840 42280 14840 0 cal_lut\[106\]
rlabel metal2 26712 25368 26712 25368 0 cal_lut\[107\]
rlabel metal3 19264 37128 19264 37128 0 cal_lut\[108\]
rlabel metal2 16800 39704 16800 39704 0 cal_lut\[109\]
rlabel metal2 23744 54376 23744 54376 0 cal_lut\[10\]
rlabel metal2 18592 49112 18592 49112 0 cal_lut\[110\]
rlabel metal2 19040 45192 19040 45192 0 cal_lut\[111\]
rlabel metal2 21336 43120 21336 43120 0 cal_lut\[112\]
rlabel metal3 25032 41272 25032 41272 0 cal_lut\[113\]
rlabel metal2 28168 41160 28168 41160 0 cal_lut\[114\]
rlabel metal2 39144 44408 39144 44408 0 cal_lut\[115\]
rlabel metal2 42728 47880 42728 47880 0 cal_lut\[116\]
rlabel metal2 42392 45136 42392 45136 0 cal_lut\[117\]
rlabel metal2 42392 37184 42392 37184 0 cal_lut\[118\]
rlabel metal3 37856 28392 37856 28392 0 cal_lut\[119\]
rlabel metal2 29232 46984 29232 46984 0 cal_lut\[11\]
rlabel metal2 32032 24024 32032 24024 0 cal_lut\[120\]
rlabel metal2 34664 22008 34664 22008 0 cal_lut\[121\]
rlabel metal2 37128 15596 37128 15596 0 cal_lut\[122\]
rlabel metal2 38920 7168 38920 7168 0 cal_lut\[123\]
rlabel metal2 37016 4312 37016 4312 0 cal_lut\[124\]
rlabel metal3 33992 16968 33992 16968 0 cal_lut\[125\]
rlabel metal2 36064 4200 36064 4200 0 cal_lut\[126\]
rlabel metal2 19096 4592 19096 4592 0 cal_lut\[127\]
rlabel metal3 16632 5208 16632 5208 0 cal_lut\[128\]
rlabel metal2 18984 4872 18984 4872 0 cal_lut\[129\]
rlabel metal2 32816 44520 32816 44520 0 cal_lut\[12\]
rlabel metal2 22456 3808 22456 3808 0 cal_lut\[130\]
rlabel metal2 25984 5096 25984 5096 0 cal_lut\[131\]
rlabel metal2 27440 6776 27440 6776 0 cal_lut\[132\]
rlabel metal2 29288 5880 29288 5880 0 cal_lut\[133\]
rlabel metal2 30016 2632 30016 2632 0 cal_lut\[134\]
rlabel metal2 30744 7784 30744 7784 0 cal_lut\[135\]
rlabel metal2 31864 8120 31864 8120 0 cal_lut\[136\]
rlabel metal3 33992 8344 33992 8344 0 cal_lut\[137\]
rlabel metal2 33096 34944 33096 34944 0 cal_lut\[138\]
rlabel metal2 37576 34384 37576 34384 0 cal_lut\[139\]
rlabel metal2 38248 56336 38248 56336 0 cal_lut\[13\]
rlabel metal2 40432 40488 40432 40488 0 cal_lut\[140\]
rlabel metal2 44016 41272 44016 41272 0 cal_lut\[141\]
rlabel metal2 46536 39984 46536 39984 0 cal_lut\[142\]
rlabel metal2 35896 38360 35896 38360 0 cal_lut\[143\]
rlabel metal2 35336 36568 35336 36568 0 cal_lut\[144\]
rlabel metal2 40264 34608 40264 34608 0 cal_lut\[145\]
rlabel metal2 42392 33040 42392 33040 0 cal_lut\[146\]
rlabel metal2 45976 32480 45976 32480 0 cal_lut\[147\]
rlabel metal2 46424 31472 46424 31472 0 cal_lut\[148\]
rlabel metal2 47320 28336 47320 28336 0 cal_lut\[149\]
rlabel metal2 40936 58520 40936 58520 0 cal_lut\[14\]
rlabel metal2 27832 23968 27832 23968 0 cal_lut\[150\]
rlabel metal2 29848 18032 29848 18032 0 cal_lut\[151\]
rlabel metal2 29400 14448 29400 14448 0 cal_lut\[152\]
rlabel via2 32536 12824 32536 12824 0 cal_lut\[153\]
rlabel metal3 31248 15848 31248 15848 0 cal_lut\[154\]
rlabel metal2 30072 23688 30072 23688 0 cal_lut\[155\]
rlabel metal2 29680 26152 29680 26152 0 cal_lut\[156\]
rlabel metal3 24304 64008 24304 64008 0 cal_lut\[157\]
rlabel metal2 20888 65800 20888 65800 0 cal_lut\[158\]
rlabel metal2 24304 65352 24304 65352 0 cal_lut\[159\]
rlabel metal2 42392 60872 42392 60872 0 cal_lut\[15\]
rlabel metal2 25312 65576 25312 65576 0 cal_lut\[160\]
rlabel metal2 27776 44520 27776 44520 0 cal_lut\[161\]
rlabel metal3 30184 23128 30184 23128 0 cal_lut\[162\]
rlabel metal2 34440 21112 34440 21112 0 cal_lut\[163\]
rlabel metal2 39704 16016 39704 16016 0 cal_lut\[164\]
rlabel metal3 39256 16856 39256 16856 0 cal_lut\[165\]
rlabel metal2 37016 18200 37016 18200 0 cal_lut\[166\]
rlabel metal2 37576 23408 37576 23408 0 cal_lut\[167\]
rlabel metal2 35000 46032 35000 46032 0 cal_lut\[168\]
rlabel metal2 38472 53200 38472 53200 0 cal_lut\[169\]
rlabel metal2 42840 60368 42840 60368 0 cal_lut\[16\]
rlabel metal3 41832 55384 41832 55384 0 cal_lut\[170\]
rlabel metal2 44072 54096 44072 54096 0 cal_lut\[171\]
rlabel metal2 45192 52528 45192 52528 0 cal_lut\[172\]
rlabel metal2 34664 47264 34664 47264 0 cal_lut\[173\]
rlabel metal2 35896 46144 35896 46144 0 cal_lut\[174\]
rlabel metal2 39032 46984 39032 46984 0 cal_lut\[175\]
rlabel metal2 41384 49112 41384 49112 0 cal_lut\[176\]
rlabel metal2 44968 49392 44968 49392 0 cal_lut\[177\]
rlabel metal2 45976 44296 45976 44296 0 cal_lut\[178\]
rlabel metal2 46032 35560 46032 35560 0 cal_lut\[179\]
rlabel metal2 41384 55832 41384 55832 0 cal_lut\[17\]
rlabel metal2 35056 50568 35056 50568 0 cal_lut\[180\]
rlabel metal2 37520 64680 37520 64680 0 cal_lut\[181\]
rlabel metal3 39592 66360 39592 66360 0 cal_lut\[182\]
rlabel metal2 37800 64344 37800 64344 0 cal_lut\[183\]
rlabel metal3 34440 63000 34440 63000 0 cal_lut\[184\]
rlabel metal3 34160 58520 34160 58520 0 cal_lut\[185\]
rlabel metal2 38808 46088 38808 46088 0 cal_lut\[186\]
rlabel metal2 40152 22456 40152 22456 0 cal_lut\[187\]
rlabel metal2 41048 18928 41048 18928 0 cal_lut\[188\]
rlabel metal2 40992 9912 40992 9912 0 cal_lut\[189\]
rlabel metal2 31528 52808 31528 52808 0 cal_lut\[18\]
rlabel metal2 40600 9968 40600 9968 0 cal_lut\[190\]
rlabel metal2 36680 12488 36680 12488 0 cal_lut\[191\]
rlabel metal2 36400 27160 36400 27160 0 cal_lut\[192\]
rlabel metal2 35784 68488 35784 68488 0 cal_lut\[19\]
rlabel metal2 17528 21784 17528 21784 0 cal_lut\[1\]
rlabel metal2 38024 70112 38024 70112 0 cal_lut\[20\]
rlabel metal2 38920 70672 38920 70672 0 cal_lut\[21\]
rlabel metal2 33656 72912 33656 72912 0 cal_lut\[22\]
rlabel metal2 28280 51856 28280 51856 0 cal_lut\[23\]
rlabel metal2 28616 49784 28616 49784 0 cal_lut\[24\]
rlabel metal3 19264 50680 19264 50680 0 cal_lut\[25\]
rlabel metal2 18816 48328 18816 48328 0 cal_lut\[26\]
rlabel metal2 16632 45080 16632 45080 0 cal_lut\[27\]
rlabel metal2 17528 42336 17528 42336 0 cal_lut\[28\]
rlabel metal2 20160 39704 20160 39704 0 cal_lut\[29\]
rlabel metal3 17248 21448 17248 21448 0 cal_lut\[2\]
rlabel metal2 20776 36680 20776 36680 0 cal_lut\[30\]
rlabel metal2 18088 14448 18088 14448 0 cal_lut\[31\]
rlabel metal2 17192 8372 17192 8372 0 cal_lut\[32\]
rlabel metal2 20216 15792 20216 15792 0 cal_lut\[33\]
rlabel metal2 22288 20664 22288 20664 0 cal_lut\[34\]
rlabel metal2 24248 26516 24248 26516 0 cal_lut\[35\]
rlabel metal2 25256 30576 25256 30576 0 cal_lut\[36\]
rlabel metal2 20944 67704 20944 67704 0 cal_lut\[37\]
rlabel metal2 21056 74200 21056 74200 0 cal_lut\[38\]
rlabel metal2 23576 76048 23576 76048 0 cal_lut\[39\]
rlabel metal3 17920 24584 17920 24584 0 cal_lut\[3\]
rlabel metal2 24136 76048 24136 76048 0 cal_lut\[40\]
rlabel metal2 27552 75768 27552 75768 0 cal_lut\[41\]
rlabel metal2 30968 74368 30968 74368 0 cal_lut\[42\]
rlabel metal2 33544 76944 33544 76944 0 cal_lut\[43\]
rlabel metal2 36456 76048 36456 76048 0 cal_lut\[44\]
rlabel metal2 37128 74480 37128 74480 0 cal_lut\[45\]
rlabel metal2 33544 74984 33544 74984 0 cal_lut\[46\]
rlabel metal2 29680 48328 29680 48328 0 cal_lut\[47\]
rlabel metal3 30520 43624 30520 43624 0 cal_lut\[48\]
rlabel metal2 33040 66920 33040 66920 0 cal_lut\[49\]
rlabel metal2 22120 24864 22120 24864 0 cal_lut\[4\]
rlabel metal3 34552 67032 34552 67032 0 cal_lut\[50\]
rlabel metal3 33432 63896 33432 63896 0 cal_lut\[51\]
rlabel metal2 32424 63952 32424 63952 0 cal_lut\[52\]
rlabel metal2 31304 62188 31304 62188 0 cal_lut\[53\]
rlabel metal3 29288 16968 29288 16968 0 cal_lut\[54\]
rlabel metal2 24472 11088 24472 11088 0 cal_lut\[55\]
rlabel metal2 22680 8372 22680 8372 0 cal_lut\[56\]
rlabel metal2 23128 11256 23128 11256 0 cal_lut\[57\]
rlabel metal2 24584 15288 24584 15288 0 cal_lut\[58\]
rlabel metal2 28168 18704 28168 18704 0 cal_lut\[59\]
rlabel metal3 13104 30072 13104 30072 0 cal_lut\[5\]
rlabel metal2 26600 25592 26600 25592 0 cal_lut\[60\]
rlabel metal3 22512 12152 22512 12152 0 cal_lut\[61\]
rlabel metal2 22008 12880 22008 12880 0 cal_lut\[62\]
rlabel metal2 22624 7336 22624 7336 0 cal_lut\[63\]
rlabel metal3 23912 18424 23912 18424 0 cal_lut\[64\]
rlabel metal2 25928 22232 25928 22232 0 cal_lut\[65\]
rlabel metal2 19208 22848 19208 22848 0 cal_lut\[66\]
rlabel metal2 18424 17136 18424 17136 0 cal_lut\[67\]
rlabel metal2 16856 14112 16856 14112 0 cal_lut\[68\]
rlabel metal2 17528 23016 17528 23016 0 cal_lut\[69\]
rlabel metal2 12040 32032 12040 32032 0 cal_lut\[6\]
rlabel metal2 20664 26236 20664 26236 0 cal_lut\[70\]
rlabel metal2 22568 35616 22568 35616 0 cal_lut\[71\]
rlabel metal3 23912 33992 23912 33992 0 cal_lut\[72\]
rlabel metal2 18368 26376 18368 26376 0 cal_lut\[73\]
rlabel metal2 16408 16128 16408 16128 0 cal_lut\[74\]
rlabel metal2 18256 26152 18256 26152 0 cal_lut\[75\]
rlabel metal2 22232 26992 22232 26992 0 cal_lut\[76\]
rlabel metal2 24192 44968 24192 44968 0 cal_lut\[77\]
rlabel metal2 25704 44520 25704 44520 0 cal_lut\[78\]
rlabel metal3 23184 52024 23184 52024 0 cal_lut\[79\]
rlabel metal2 16632 54768 16632 54768 0 cal_lut\[7\]
rlabel metal2 21224 61656 21224 61656 0 cal_lut\[80\]
rlabel metal2 23912 60368 23912 60368 0 cal_lut\[81\]
rlabel metal2 26096 61656 26096 61656 0 cal_lut\[82\]
rlabel metal2 27104 45304 27104 45304 0 cal_lut\[83\]
rlabel metal2 28728 43624 28728 43624 0 cal_lut\[84\]
rlabel metal2 19656 68208 19656 68208 0 cal_lut\[85\]
rlabel metal2 20720 70056 20720 70056 0 cal_lut\[86\]
rlabel via1 23576 71610 23576 71610 0 cal_lut\[87\]
rlabel metal2 25648 71064 25648 71064 0 cal_lut\[88\]
rlabel metal2 28000 65800 28000 65800 0 cal_lut\[89\]
rlabel metal2 18536 63896 18536 63896 0 cal_lut\[8\]
rlabel metal2 29736 57904 29736 57904 0 cal_lut\[90\]
rlabel metal2 17976 58912 17976 58912 0 cal_lut\[91\]
rlabel metal2 18424 56952 18424 56952 0 cal_lut\[92\]
rlabel metal2 19208 54208 19208 54208 0 cal_lut\[93\]
rlabel metal2 23688 52136 23688 52136 0 cal_lut\[94\]
rlabel metal2 26376 39312 26376 39312 0 cal_lut\[95\]
rlabel metal2 28168 31696 28168 31696 0 cal_lut\[96\]
rlabel metal2 39592 30184 39592 30184 0 cal_lut\[97\]
rlabel metal3 43064 27160 43064 27160 0 cal_lut\[98\]
rlabel metal2 45416 26432 45416 26432 0 cal_lut\[99\]
rlabel metal2 20328 63112 20328 63112 0 cal_lut\[9\]
rlabel metal2 7560 40320 7560 40320 0 clknet_0__0316_
rlabel metal2 15288 39536 15288 39536 0 clknet_0__0318_
rlabel metal3 10192 20888 10192 20888 0 clknet_0_io_in[0]
rlabel metal2 8120 45640 8120 45640 0 clknet_0_net23
rlabel metal2 6328 53256 6328 53256 0 clknet_0_temp1.i_precharge_n
rlabel metal2 3920 40152 3920 40152 0 clknet_1_0__leaf__0316_
rlabel metal2 9352 37352 9352 37352 0 clknet_1_0__leaf__0318_
rlabel metal2 1736 5768 1736 5768 0 clknet_1_0__leaf_io_in[0]
rlabel metal3 6328 42616 6328 42616 0 clknet_1_0__leaf_net23
rlabel metal3 5992 53032 5992 53032 0 clknet_1_0__leaf_temp1.i_precharge_n
rlabel metal2 2744 43064 2744 43064 0 clknet_1_1__leaf__0316_
rlabel metal2 12264 40712 12264 40712 0 clknet_1_1__leaf__0318_
rlabel metal2 7896 50512 7896 50512 0 clknet_1_1__leaf_io_in[0]
rlabel metal2 3808 45864 3808 45864 0 clknet_1_1__leaf_net23
rlabel metal2 3192 55216 3192 55216 0 clknet_1_1__leaf_temp1.i_precharge_n
rlabel metal2 14056 53256 14056 53256 0 ctr\[0\]
rlabel metal2 3864 14000 3864 14000 0 ctr\[10\]
rlabel metal2 3528 15288 3528 15288 0 ctr\[11\]
rlabel metal2 2968 6608 2968 6608 0 ctr\[12\]
rlabel metal2 4424 43848 4424 43848 0 ctr\[1\]
rlabel metal2 7560 42896 7560 42896 0 ctr\[2\]
rlabel metal3 6832 50568 6832 50568 0 ctr\[3\]
rlabel metal2 7560 50568 7560 50568 0 ctr\[4\]
rlabel metal2 12488 51296 12488 51296 0 ctr\[5\]
rlabel metal3 10920 38808 10920 38808 0 ctr\[6\]
rlabel metal2 9016 47768 9016 47768 0 ctr\[7\]
rlabel metal2 3304 16296 3304 16296 0 ctr\[8\]
rlabel metal2 4648 18256 4648 18256 0 ctr\[9\]
rlabel metal2 13944 42280 13944 42280 0 dbg3\[0\]
rlabel metal2 11368 36120 11368 36120 0 dbg3\[1\]
rlabel metal2 12936 44744 12936 44744 0 dbg3\[2\]
rlabel metal2 14336 32424 14336 32424 0 dbg3\[3\]
rlabel metal2 14728 38360 14728 38360 0 dbg3\[4\]
rlabel metal2 10696 30912 10696 30912 0 dbg3\[5\]
rlabel metal3 6272 9016 6272 9016 0 dec1._000_
rlabel metal3 5544 6552 5544 6552 0 dec1._001_
rlabel metal3 8232 6440 8232 6440 0 dec1._002_
rlabel metal2 11704 11984 11704 11984 0 dec1._003_
rlabel metal3 12488 15064 12488 15064 0 dec1._004_
rlabel metal2 12600 14000 12600 14000 0 dec1._005_
rlabel metal2 11928 13552 11928 13552 0 dec1._006_
rlabel metal3 13384 6552 13384 6552 0 dec1._007_
rlabel metal2 11592 12880 11592 12880 0 dec1._008_
rlabel metal2 13608 12992 13608 12992 0 dec1._009_
rlabel metal2 13608 10192 13608 10192 0 dec1._010_
rlabel metal3 15204 9912 15204 9912 0 dec1._011_
rlabel metal2 12600 10136 12600 10136 0 dec1._012_
rlabel metal2 14280 6608 14280 6608 0 dec1._013_
rlabel metal2 14056 7784 14056 7784 0 dec1._014_
rlabel metal2 13832 5096 13832 5096 0 dec1._015_
rlabel metal3 12152 6664 12152 6664 0 dec1._016_
rlabel metal2 13384 9688 13384 9688 0 dec1._017_
rlabel metal2 10472 9296 10472 9296 0 dec1._018_
rlabel metal2 14952 8512 14952 8512 0 dec1._019_
rlabel metal2 10248 14224 10248 14224 0 dec1._020_
rlabel metal2 11480 12992 11480 12992 0 dec1._021_
rlabel metal2 11704 15540 11704 15540 0 dec1._022_
rlabel metal2 12712 10248 12712 10248 0 dec1._023_
rlabel metal2 11928 12264 11928 12264 0 dec1._024_
rlabel metal2 11368 7280 11368 7280 0 dec1._025_
rlabel metal2 10360 2576 10360 2576 0 dec1._026_
rlabel metal2 12040 3304 12040 3304 0 dec1._027_
rlabel metal2 10752 5880 10752 5880 0 dec1._028_
rlabel metal2 12040 11928 12040 11928 0 dec1._029_
rlabel metal3 15288 7784 15288 7784 0 dec1._030_
rlabel metal2 12264 4760 12264 4760 0 dec1._031_
rlabel metal2 8456 4088 8456 4088 0 dec1._032_
rlabel metal2 8904 4312 8904 4312 0 dec1._033_
rlabel metal3 13832 5992 13832 5992 0 dec1._034_
rlabel metal3 13048 5768 13048 5768 0 dec1._035_
rlabel metal2 11032 5320 11032 5320 0 dec1._036_
rlabel metal2 10528 5656 10528 5656 0 dec1._037_
rlabel metal2 11032 3640 11032 3640 0 dec1._038_
rlabel metal2 11256 5544 11256 5544 0 dec1._039_
rlabel metal2 7560 4984 7560 4984 0 dec1._040_
rlabel metal2 7448 8624 7448 8624 0 dec1._041_
rlabel metal2 10136 12992 10136 12992 0 dec1._042_
rlabel metal2 9912 11816 9912 11816 0 dec1._043_
rlabel metal2 9576 13216 9576 13216 0 dec1._044_
rlabel metal2 10024 12432 10024 12432 0 dec1._045_
rlabel metal2 8344 12600 8344 12600 0 dec1._046_
rlabel metal2 8064 2744 8064 2744 0 dec1._047_
rlabel metal2 9800 5096 9800 5096 0 dec1._048_
rlabel metal2 10584 3052 10584 3052 0 dec1._049_
rlabel metal3 8736 2520 8736 2520 0 dec1._050_
rlabel metal2 6104 4928 6104 4928 0 dec1._051_
rlabel metal2 9016 8568 9016 8568 0 dec1._052_
rlabel metal3 7560 7448 7560 7448 0 dec1._053_
rlabel metal3 7840 7672 7840 7672 0 dec1._054_
rlabel metal2 8008 7784 8008 7784 0 dec1._055_
rlabel metal2 10248 11648 10248 11648 0 dec1._056_
rlabel metal2 6888 4592 6888 4592 0 dec1._057_
rlabel metal2 6944 2968 6944 2968 0 dec1._058_
rlabel metal4 7448 7560 7448 7560 0 dec1._059_
rlabel metal2 7224 24136 7224 24136 0 dec1.i_bin\[0\]
rlabel metal2 10864 18536 10864 18536 0 dec1.i_bin\[1\]
rlabel metal2 12040 9576 12040 9576 0 dec1.i_bin\[2\]
rlabel metal2 15176 7056 15176 7056 0 dec1.i_bin\[3\]
rlabel metal2 11480 16856 11480 16856 0 dec1.i_bin\[4\]
rlabel metal2 11984 16856 11984 16856 0 dec1.i_bin\[5\]
rlabel metal2 15288 23912 15288 23912 0 dec1.i_bin\[6\]
rlabel metal2 6552 2968 6552 2968 0 dec1.i_ones
rlabel metal3 2688 27832 2688 27832 0 dec1.i_tens
rlabel metal3 5600 17528 5600 17528 0 dec1.o_dec\[0\]
rlabel metal3 6384 16856 6384 16856 0 dec1.o_dec\[1\]
rlabel metal2 7000 11032 7000 11032 0 dec1.o_dec\[2\]
rlabel metal3 8288 11480 8288 11480 0 dec1.o_dec\[3\]
rlabel metal3 3094 2968 3094 2968 0 io_in[0]
rlabel metal2 1848 7952 1848 7952 0 io_in[1]
rlabel metal3 1022 12824 1022 12824 0 io_in[2]
rlabel metal2 1736 17696 1736 17696 0 io_in[3]
rlabel metal2 1736 22176 1736 22176 0 io_in[4]
rlabel metal2 2632 27048 2632 27048 0 io_in[5]
rlabel metal2 1848 31892 1848 31892 0 io_in[6]
rlabel metal3 1134 37464 1134 37464 0 io_in[7]
rlabel metal2 3416 41328 3416 41328 0 io_out[0]
rlabel metal3 1358 47320 1358 47320 0 io_out[1]
rlabel metal3 2814 52248 2814 52248 0 io_out[2]
rlabel metal2 6776 53816 6776 53816 0 io_out[3]
rlabel metal2 3808 53816 3808 53816 0 io_out[4]
rlabel metal2 4088 51016 4088 51016 0 io_out[5]
rlabel metal2 2632 54264 2632 54264 0 io_out[6]
rlabel metal2 3528 52360 3528 52360 0 io_out[7]
rlabel metal2 2072 7952 2072 7952 0 net1
rlabel metal2 43736 9520 43736 9520 0 net10
rlabel metal2 23968 25480 23968 25480 0 net11
rlabel metal3 44632 28616 44632 28616 0 net12
rlabel metal3 44576 31976 44576 31976 0 net13
rlabel metal2 40936 39760 40936 39760 0 net14
rlabel metal2 13832 54432 13832 54432 0 net15
rlabel metal3 25424 73192 25424 73192 0 net16
rlabel metal2 31304 76440 31304 76440 0 net17
rlabel metal2 25032 68936 25032 68936 0 net18
rlabel metal2 2912 68712 2912 68712 0 net19
rlabel metal2 42224 50680 42224 50680 0 net2
rlabel metal2 2632 68712 2632 68712 0 net20
rlabel metal2 3136 66584 3136 66584 0 net21
rlabel metal3 7616 53480 7616 53480 0 net22
rlabel metal2 2072 52248 2072 52248 0 net23
rlabel metal2 3752 42728 3752 42728 0 net24
rlabel metal3 3472 45864 3472 45864 0 net25
rlabel metal2 2072 17696 2072 17696 0 net3
rlabel metal2 2072 22064 2072 22064 0 net4
rlabel metal2 3080 29008 3080 29008 0 net5
rlabel metal2 2296 30184 2296 30184 0 net6
rlabel metal2 2128 37240 2128 37240 0 net7
rlabel metal2 20776 6216 20776 6216 0 net8
rlabel metal2 25144 13328 25144 13328 0 net9
rlabel metal2 5208 12208 5208 12208 0 seg1._00_
rlabel metal2 5544 12376 5544 12376 0 seg1._01_
rlabel metal2 5656 11760 5656 11760 0 seg1._02_
rlabel metal2 5656 17248 5656 17248 0 seg1._03_
rlabel metal3 5544 12936 5544 12936 0 seg1._04_
rlabel metal2 4872 11928 4872 11928 0 seg1._05_
rlabel metal2 5768 12320 5768 12320 0 seg1._06_
rlabel metal3 4872 12040 4872 12040 0 seg1._07_
rlabel metal3 5600 17752 5600 17752 0 seg1._08_
rlabel metal2 8120 17864 8120 17864 0 seg1._09_
rlabel metal2 8400 19208 8400 19208 0 seg1._10_
rlabel metal2 7896 18088 7896 18088 0 seg1._11_
rlabel metal2 7448 18424 7448 18424 0 seg1._12_
rlabel metal3 5768 18424 5768 18424 0 seg1._13_
rlabel metal2 8120 16912 8120 16912 0 seg1._14_
rlabel metal2 9464 18536 9464 18536 0 seg1._15_
rlabel metal2 7448 18928 7448 18928 0 seg1._16_
rlabel metal2 7560 17864 7560 17864 0 seg1._17_
rlabel metal2 8008 20496 8008 20496 0 seg1._18_
rlabel metal2 6440 18872 6440 18872 0 seg1._19_
rlabel metal3 6496 18984 6496 18984 0 seg1._20_
rlabel metal2 5992 18592 5992 18592 0 seg1._21_
rlabel metal2 8568 17304 8568 17304 0 seg1._22_
rlabel metal2 8960 17864 8960 17864 0 seg1._23_
rlabel metal2 5768 16520 5768 16520 0 seg1._24_
rlabel metal2 6104 12712 6104 12712 0 seg1._25_
rlabel metal2 6608 19432 6608 19432 0 seg1.o_segments\[0\]
rlabel metal2 8232 21448 8232 21448 0 seg1.o_segments\[1\]
rlabel metal2 5768 19040 5768 19040 0 seg1.o_segments\[2\]
rlabel metal3 8792 21784 8792 21784 0 seg1.o_segments\[3\]
rlabel metal2 6104 19656 6104 19656 0 seg1.o_segments\[4\]
rlabel metal2 8904 19992 8904 19992 0 seg1.o_segments\[5\]
rlabel metal2 5880 17024 5880 17024 0 seg1.o_segments\[6\]
rlabel metal2 3192 67480 3192 67480 0 temp1.dac._0_
rlabel metal3 3976 66024 3976 66024 0 temp1.dac._1_
rlabel metal2 4872 52696 4872 52696 0 temp1.dac.i_data\[0\]
rlabel metal2 4368 52696 4368 52696 0 temp1.dac.i_data\[1\]
rlabel metal2 4872 53424 4872 53424 0 temp1.dac.i_data\[2\]
rlabel metal2 5992 54824 5992 54824 0 temp1.dac.i_data\[3\]
rlabel metal2 7784 54460 7784 54460 0 temp1.dac.i_data\[4\]
rlabel metal2 7280 51576 7280 51576 0 temp1.dac.i_data\[5\]
rlabel metal2 2632 7840 2632 7840 0 temp1.dac.i_enable
rlabel metal2 2352 57848 2352 57848 0 temp1.dac.parallel_cells\[0\].vdac_batch._0_
rlabel metal2 2632 58352 2632 58352 0 temp1.dac.parallel_cells\[0\].vdac_batch._1_
rlabel metal2 3528 57232 3528 57232 0 temp1.dac.parallel_cells\[0\].vdac_batch._2_
rlabel metal2 4256 57624 4256 57624 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_pupd
rlabel metal2 1848 58688 1848 58688 0 temp1.dac.parallel_cells\[0\].vdac_batch.en_vref
rlabel metal2 5096 57120 5096 57120 0 temp1.dac.parallel_cells\[0\].vdac_batch.npu_pd
rlabel metal3 5656 55272 5656 55272 0 temp1.dac.parallel_cells\[0\].vdac_batch.vout_notouch_
rlabel metal2 5880 61768 5880 61768 0 temp1.dac.parallel_cells\[1\].vdac_batch._0_
rlabel metal2 4256 61768 4256 61768 0 temp1.dac.parallel_cells\[1\].vdac_batch._1_
rlabel metal2 3752 62776 3752 62776 0 temp1.dac.parallel_cells\[1\].vdac_batch._2_
rlabel metal2 1960 62608 1960 62608 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_pupd
rlabel metal2 5488 61656 5488 61656 0 temp1.dac.parallel_cells\[1\].vdac_batch.en_vref
rlabel metal2 3304 61096 3304 61096 0 temp1.dac.parallel_cells\[1\].vdac_batch.npu_pd
rlabel metal2 5992 56784 5992 56784 0 temp1.dac.parallel_cells\[2\].vdac_batch._0_
rlabel metal2 6664 57736 6664 57736 0 temp1.dac.parallel_cells\[2\].vdac_batch._1_
rlabel metal2 6776 59584 6776 59584 0 temp1.dac.parallel_cells\[2\].vdac_batch._2_
rlabel metal3 8008 61544 8008 61544 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_pupd
rlabel metal3 7336 56840 7336 56840 0 temp1.dac.parallel_cells\[2\].vdac_batch.en_vref
rlabel metal2 7672 60480 7672 60480 0 temp1.dac.parallel_cells\[2\].vdac_batch.npu_pd
rlabel metal2 5656 69888 5656 69888 0 temp1.dac.parallel_cells\[3\].vdac_batch._0_
rlabel metal2 4984 69160 4984 69160 0 temp1.dac.parallel_cells\[3\].vdac_batch._1_
rlabel metal2 4424 70672 4424 70672 0 temp1.dac.parallel_cells\[3\].vdac_batch._2_
rlabel metal2 2744 71344 2744 71344 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_pupd
rlabel metal2 6216 75264 6216 75264 0 temp1.dac.parallel_cells\[3\].vdac_batch.en_vref
rlabel metal2 3192 72464 3192 72464 0 temp1.dac.parallel_cells\[3\].vdac_batch.npu_pd
rlabel metal3 7280 66808 7280 66808 0 temp1.dac.parallel_cells\[4\].vdac_batch._0_
rlabel metal2 7224 66752 7224 66752 0 temp1.dac.parallel_cells\[4\].vdac_batch._1_
rlabel metal2 8400 66136 8400 66136 0 temp1.dac.parallel_cells\[4\].vdac_batch._2_
rlabel metal2 10640 59192 10640 59192 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_pupd
rlabel metal2 10696 74032 10696 74032 0 temp1.dac.parallel_cells\[4\].vdac_batch.en_vref
rlabel metal2 11984 59304 11984 59304 0 temp1.dac.parallel_cells\[4\].vdac_batch.npu_pd
rlabel metal2 3752 67424 3752 67424 0 temp1.dac.vdac_single._0_
rlabel metal3 2800 67480 2800 67480 0 temp1.dac.vdac_single._1_
rlabel metal2 2464 67704 2464 67704 0 temp1.dac.vdac_single._2_
rlabel metal2 1960 67396 1960 67396 0 temp1.dac.vdac_single.en_pupd
rlabel metal2 4088 67536 4088 67536 0 temp1.dac.vdac_single.en_vref
rlabel metal2 2688 65240 2688 65240 0 temp1.dac.vdac_single.npu_pd
rlabel metal2 1960 54040 1960 54040 0 temp1.dcdel_capnode_notouch_
rlabel metal2 3304 53816 3304 53816 0 temp1.i_precharge_n
rlabel metal2 2632 41048 2632 41048 0 temp_delay_last
<< properties >>
string FIXED_BBOX 0 0 50000 80000
<< end >>
