VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_wrapper
  CLASS BLOCK ;
  FOREIGN analog_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2550.000 BY 1750.000 ;
  PIN in1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.519000 ;
    PORT
      LAYER Metal2 ;
        RECT 1273.440 0.000 1274.000 4.000 ;
    END
  END in1
  PIN in2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.519000 ;
    PORT
      LAYER Metal2 ;
        RECT 1270.080 0.000 1270.640 4.000 ;
    END
  END in2
  PIN out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.893200 ;
    PORT
      LAYER Metal2 ;
        RECT 1273.440 1746.000 1274.000 1750.000 ;
    END
  END out
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 19.940 15.380 26.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 119.940 15.380 126.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 219.940 15.380 226.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 319.940 15.380 326.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 419.940 15.380 426.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 519.940 15.380 526.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 619.940 15.380 626.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 719.940 15.380 726.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 819.940 15.380 826.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 919.940 15.380 926.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1019.940 15.380 1026.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1119.940 15.380 1126.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1219.940 15.380 1226.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1319.940 15.380 1326.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1419.940 15.380 1426.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1519.940 15.380 1526.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1619.940 15.380 1626.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1719.940 15.380 1726.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1819.940 15.380 1826.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1919.940 15.380 1926.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.940 15.380 2026.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2119.940 15.380 2126.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2219.940 15.380 2226.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2319.940 15.380 2326.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2419.940 15.380 2426.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2519.940 15.380 2526.140 1732.940 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 69.940 15.380 76.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 169.940 15.380 176.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 269.940 15.380 276.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 369.940 15.380 376.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 469.940 15.380 476.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 569.940 15.380 576.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 669.940 15.380 676.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 769.940 15.380 776.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 869.940 15.380 876.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 969.940 15.380 976.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1069.940 15.380 1076.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1169.940 15.380 1176.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1269.940 15.380 1276.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1369.940 15.380 1376.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1469.940 15.380 1476.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1569.940 15.380 1576.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1669.940 15.380 1676.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1769.940 15.380 1776.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1869.940 15.380 1876.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1969.940 15.380 1976.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2069.940 15.380 2076.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2169.940 15.380 2176.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2269.940 15.380 2276.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2369.940 15.380 2376.140 1732.940 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2469.940 15.380 2476.140 1732.940 ;
    END
  END vss
  OBS
      LAYER Pwell ;
        RECT 6.290 1730.880 2543.390 1733.070 ;
      LAYER Nwell ;
        RECT 6.290 1726.560 2543.390 1730.880 ;
      LAYER Pwell ;
        RECT 6.290 1723.040 2543.390 1726.560 ;
      LAYER Nwell ;
        RECT 6.290 1718.720 2543.390 1723.040 ;
      LAYER Pwell ;
        RECT 6.290 1715.200 2543.390 1718.720 ;
      LAYER Nwell ;
        RECT 6.290 1710.880 2543.390 1715.200 ;
      LAYER Pwell ;
        RECT 6.290 1707.360 2543.390 1710.880 ;
      LAYER Nwell ;
        RECT 6.290 1703.040 2543.390 1707.360 ;
      LAYER Pwell ;
        RECT 6.290 1699.520 2543.390 1703.040 ;
      LAYER Nwell ;
        RECT 6.290 1695.200 2543.390 1699.520 ;
      LAYER Pwell ;
        RECT 6.290 1691.680 2543.390 1695.200 ;
      LAYER Nwell ;
        RECT 6.290 1687.360 2543.390 1691.680 ;
      LAYER Pwell ;
        RECT 6.290 1683.840 2543.390 1687.360 ;
      LAYER Nwell ;
        RECT 6.290 1679.520 2543.390 1683.840 ;
      LAYER Pwell ;
        RECT 6.290 1676.000 2543.390 1679.520 ;
      LAYER Nwell ;
        RECT 6.290 1671.680 2543.390 1676.000 ;
      LAYER Pwell ;
        RECT 6.290 1668.160 2543.390 1671.680 ;
      LAYER Nwell ;
        RECT 6.290 1663.840 2543.390 1668.160 ;
      LAYER Pwell ;
        RECT 6.290 1660.320 2543.390 1663.840 ;
      LAYER Nwell ;
        RECT 6.290 1656.000 2543.390 1660.320 ;
      LAYER Pwell ;
        RECT 6.290 1652.480 2543.390 1656.000 ;
      LAYER Nwell ;
        RECT 6.290 1648.160 2543.390 1652.480 ;
      LAYER Pwell ;
        RECT 6.290 1644.640 2543.390 1648.160 ;
      LAYER Nwell ;
        RECT 6.290 1640.320 2543.390 1644.640 ;
      LAYER Pwell ;
        RECT 6.290 1636.800 2543.390 1640.320 ;
      LAYER Nwell ;
        RECT 6.290 1632.480 2543.390 1636.800 ;
      LAYER Pwell ;
        RECT 6.290 1628.960 2543.390 1632.480 ;
      LAYER Nwell ;
        RECT 6.290 1624.640 2543.390 1628.960 ;
      LAYER Pwell ;
        RECT 6.290 1621.120 2543.390 1624.640 ;
      LAYER Nwell ;
        RECT 6.290 1616.800 2543.390 1621.120 ;
      LAYER Pwell ;
        RECT 6.290 1613.280 2543.390 1616.800 ;
      LAYER Nwell ;
        RECT 6.290 1608.960 2543.390 1613.280 ;
      LAYER Pwell ;
        RECT 6.290 1605.440 2543.390 1608.960 ;
      LAYER Nwell ;
        RECT 6.290 1601.120 2543.390 1605.440 ;
      LAYER Pwell ;
        RECT 6.290 1597.600 2543.390 1601.120 ;
      LAYER Nwell ;
        RECT 6.290 1593.280 2543.390 1597.600 ;
      LAYER Pwell ;
        RECT 6.290 1589.760 2543.390 1593.280 ;
      LAYER Nwell ;
        RECT 6.290 1585.440 2543.390 1589.760 ;
      LAYER Pwell ;
        RECT 6.290 1581.920 2543.390 1585.440 ;
      LAYER Nwell ;
        RECT 6.290 1577.600 2543.390 1581.920 ;
      LAYER Pwell ;
        RECT 6.290 1574.080 2543.390 1577.600 ;
      LAYER Nwell ;
        RECT 6.290 1569.760 2543.390 1574.080 ;
      LAYER Pwell ;
        RECT 6.290 1566.240 2543.390 1569.760 ;
      LAYER Nwell ;
        RECT 6.290 1561.920 2543.390 1566.240 ;
      LAYER Pwell ;
        RECT 6.290 1558.400 2543.390 1561.920 ;
      LAYER Nwell ;
        RECT 6.290 1554.080 2543.390 1558.400 ;
      LAYER Pwell ;
        RECT 6.290 1550.560 2543.390 1554.080 ;
      LAYER Nwell ;
        RECT 6.290 1546.240 2543.390 1550.560 ;
      LAYER Pwell ;
        RECT 6.290 1542.720 2543.390 1546.240 ;
      LAYER Nwell ;
        RECT 6.290 1538.400 2543.390 1542.720 ;
      LAYER Pwell ;
        RECT 6.290 1534.880 2543.390 1538.400 ;
      LAYER Nwell ;
        RECT 6.290 1530.560 2543.390 1534.880 ;
      LAYER Pwell ;
        RECT 6.290 1527.040 2543.390 1530.560 ;
      LAYER Nwell ;
        RECT 6.290 1522.720 2543.390 1527.040 ;
      LAYER Pwell ;
        RECT 6.290 1519.200 2543.390 1522.720 ;
      LAYER Nwell ;
        RECT 6.290 1514.880 2543.390 1519.200 ;
      LAYER Pwell ;
        RECT 6.290 1511.360 2543.390 1514.880 ;
      LAYER Nwell ;
        RECT 6.290 1507.040 2543.390 1511.360 ;
      LAYER Pwell ;
        RECT 6.290 1503.520 2543.390 1507.040 ;
      LAYER Nwell ;
        RECT 6.290 1499.200 2543.390 1503.520 ;
      LAYER Pwell ;
        RECT 6.290 1495.680 2543.390 1499.200 ;
      LAYER Nwell ;
        RECT 6.290 1491.360 2543.390 1495.680 ;
      LAYER Pwell ;
        RECT 6.290 1487.840 2543.390 1491.360 ;
      LAYER Nwell ;
        RECT 6.290 1483.520 2543.390 1487.840 ;
      LAYER Pwell ;
        RECT 6.290 1480.000 2543.390 1483.520 ;
      LAYER Nwell ;
        RECT 6.290 1475.680 2543.390 1480.000 ;
      LAYER Pwell ;
        RECT 6.290 1472.160 2543.390 1475.680 ;
      LAYER Nwell ;
        RECT 6.290 1467.840 2543.390 1472.160 ;
      LAYER Pwell ;
        RECT 6.290 1464.320 2543.390 1467.840 ;
      LAYER Nwell ;
        RECT 6.290 1460.000 2543.390 1464.320 ;
      LAYER Pwell ;
        RECT 6.290 1456.480 2543.390 1460.000 ;
      LAYER Nwell ;
        RECT 6.290 1452.160 2543.390 1456.480 ;
      LAYER Pwell ;
        RECT 6.290 1448.640 2543.390 1452.160 ;
      LAYER Nwell ;
        RECT 6.290 1444.320 2543.390 1448.640 ;
      LAYER Pwell ;
        RECT 6.290 1440.800 2543.390 1444.320 ;
      LAYER Nwell ;
        RECT 6.290 1436.480 2543.390 1440.800 ;
      LAYER Pwell ;
        RECT 6.290 1432.960 2543.390 1436.480 ;
      LAYER Nwell ;
        RECT 6.290 1428.640 2543.390 1432.960 ;
      LAYER Pwell ;
        RECT 6.290 1425.120 2543.390 1428.640 ;
      LAYER Nwell ;
        RECT 6.290 1420.800 2543.390 1425.120 ;
      LAYER Pwell ;
        RECT 6.290 1417.280 2543.390 1420.800 ;
      LAYER Nwell ;
        RECT 6.290 1412.960 2543.390 1417.280 ;
      LAYER Pwell ;
        RECT 6.290 1409.440 2543.390 1412.960 ;
      LAYER Nwell ;
        RECT 6.290 1405.120 2543.390 1409.440 ;
      LAYER Pwell ;
        RECT 6.290 1401.600 2543.390 1405.120 ;
      LAYER Nwell ;
        RECT 6.290 1397.280 2543.390 1401.600 ;
      LAYER Pwell ;
        RECT 6.290 1393.760 2543.390 1397.280 ;
      LAYER Nwell ;
        RECT 6.290 1389.440 2543.390 1393.760 ;
      LAYER Pwell ;
        RECT 6.290 1385.920 2543.390 1389.440 ;
      LAYER Nwell ;
        RECT 6.290 1381.600 2543.390 1385.920 ;
      LAYER Pwell ;
        RECT 6.290 1378.080 2543.390 1381.600 ;
      LAYER Nwell ;
        RECT 6.290 1373.760 2543.390 1378.080 ;
      LAYER Pwell ;
        RECT 6.290 1370.240 2543.390 1373.760 ;
      LAYER Nwell ;
        RECT 6.290 1365.920 2543.390 1370.240 ;
      LAYER Pwell ;
        RECT 6.290 1362.400 2543.390 1365.920 ;
      LAYER Nwell ;
        RECT 6.290 1358.080 2543.390 1362.400 ;
      LAYER Pwell ;
        RECT 6.290 1354.560 2543.390 1358.080 ;
      LAYER Nwell ;
        RECT 6.290 1350.240 2543.390 1354.560 ;
      LAYER Pwell ;
        RECT 6.290 1346.720 2543.390 1350.240 ;
      LAYER Nwell ;
        RECT 6.290 1342.400 2543.390 1346.720 ;
      LAYER Pwell ;
        RECT 6.290 1338.880 2543.390 1342.400 ;
      LAYER Nwell ;
        RECT 6.290 1334.560 2543.390 1338.880 ;
      LAYER Pwell ;
        RECT 6.290 1331.040 2543.390 1334.560 ;
      LAYER Nwell ;
        RECT 6.290 1326.720 2543.390 1331.040 ;
      LAYER Pwell ;
        RECT 6.290 1323.200 2543.390 1326.720 ;
      LAYER Nwell ;
        RECT 6.290 1318.880 2543.390 1323.200 ;
      LAYER Pwell ;
        RECT 6.290 1315.360 2543.390 1318.880 ;
      LAYER Nwell ;
        RECT 6.290 1311.040 2543.390 1315.360 ;
      LAYER Pwell ;
        RECT 6.290 1307.520 2543.390 1311.040 ;
      LAYER Nwell ;
        RECT 6.290 1303.200 2543.390 1307.520 ;
      LAYER Pwell ;
        RECT 6.290 1299.680 2543.390 1303.200 ;
      LAYER Nwell ;
        RECT 6.290 1295.360 2543.390 1299.680 ;
      LAYER Pwell ;
        RECT 6.290 1291.840 2543.390 1295.360 ;
      LAYER Nwell ;
        RECT 6.290 1287.520 2543.390 1291.840 ;
      LAYER Pwell ;
        RECT 6.290 1284.000 2543.390 1287.520 ;
      LAYER Nwell ;
        RECT 6.290 1279.680 2543.390 1284.000 ;
      LAYER Pwell ;
        RECT 6.290 1276.160 2543.390 1279.680 ;
      LAYER Nwell ;
        RECT 6.290 1271.840 2543.390 1276.160 ;
      LAYER Pwell ;
        RECT 6.290 1268.320 2543.390 1271.840 ;
      LAYER Nwell ;
        RECT 6.290 1264.000 2543.390 1268.320 ;
      LAYER Pwell ;
        RECT 6.290 1260.480 2543.390 1264.000 ;
      LAYER Nwell ;
        RECT 6.290 1256.160 2543.390 1260.480 ;
      LAYER Pwell ;
        RECT 6.290 1252.640 2543.390 1256.160 ;
      LAYER Nwell ;
        RECT 6.290 1248.320 2543.390 1252.640 ;
      LAYER Pwell ;
        RECT 6.290 1244.800 2543.390 1248.320 ;
      LAYER Nwell ;
        RECT 6.290 1240.480 2543.390 1244.800 ;
      LAYER Pwell ;
        RECT 6.290 1236.960 2543.390 1240.480 ;
      LAYER Nwell ;
        RECT 6.290 1232.640 2543.390 1236.960 ;
      LAYER Pwell ;
        RECT 6.290 1229.120 2543.390 1232.640 ;
      LAYER Nwell ;
        RECT 6.290 1224.800 2543.390 1229.120 ;
      LAYER Pwell ;
        RECT 6.290 1221.280 2543.390 1224.800 ;
      LAYER Nwell ;
        RECT 6.290 1216.960 2543.390 1221.280 ;
      LAYER Pwell ;
        RECT 6.290 1213.440 2543.390 1216.960 ;
      LAYER Nwell ;
        RECT 6.290 1209.120 2543.390 1213.440 ;
      LAYER Pwell ;
        RECT 6.290 1205.600 2543.390 1209.120 ;
      LAYER Nwell ;
        RECT 6.290 1201.280 2543.390 1205.600 ;
      LAYER Pwell ;
        RECT 6.290 1197.760 2543.390 1201.280 ;
      LAYER Nwell ;
        RECT 6.290 1193.440 2543.390 1197.760 ;
      LAYER Pwell ;
        RECT 6.290 1189.920 2543.390 1193.440 ;
      LAYER Nwell ;
        RECT 6.290 1185.600 2543.390 1189.920 ;
      LAYER Pwell ;
        RECT 6.290 1182.080 2543.390 1185.600 ;
      LAYER Nwell ;
        RECT 6.290 1177.760 2543.390 1182.080 ;
      LAYER Pwell ;
        RECT 6.290 1174.240 2543.390 1177.760 ;
      LAYER Nwell ;
        RECT 6.290 1169.920 2543.390 1174.240 ;
      LAYER Pwell ;
        RECT 6.290 1166.400 2543.390 1169.920 ;
      LAYER Nwell ;
        RECT 6.290 1162.080 2543.390 1166.400 ;
      LAYER Pwell ;
        RECT 6.290 1158.560 2543.390 1162.080 ;
      LAYER Nwell ;
        RECT 6.290 1154.240 2543.390 1158.560 ;
      LAYER Pwell ;
        RECT 6.290 1150.720 2543.390 1154.240 ;
      LAYER Nwell ;
        RECT 6.290 1146.400 2543.390 1150.720 ;
      LAYER Pwell ;
        RECT 6.290 1142.880 2543.390 1146.400 ;
      LAYER Nwell ;
        RECT 6.290 1138.560 2543.390 1142.880 ;
      LAYER Pwell ;
        RECT 6.290 1135.040 2543.390 1138.560 ;
      LAYER Nwell ;
        RECT 6.290 1130.720 2543.390 1135.040 ;
      LAYER Pwell ;
        RECT 6.290 1127.200 2543.390 1130.720 ;
      LAYER Nwell ;
        RECT 6.290 1122.880 2543.390 1127.200 ;
      LAYER Pwell ;
        RECT 6.290 1119.360 2543.390 1122.880 ;
      LAYER Nwell ;
        RECT 6.290 1115.040 2543.390 1119.360 ;
      LAYER Pwell ;
        RECT 6.290 1111.520 2543.390 1115.040 ;
      LAYER Nwell ;
        RECT 6.290 1107.200 2543.390 1111.520 ;
      LAYER Pwell ;
        RECT 6.290 1103.680 2543.390 1107.200 ;
      LAYER Nwell ;
        RECT 6.290 1099.360 2543.390 1103.680 ;
      LAYER Pwell ;
        RECT 6.290 1095.840 2543.390 1099.360 ;
      LAYER Nwell ;
        RECT 6.290 1091.520 2543.390 1095.840 ;
      LAYER Pwell ;
        RECT 6.290 1088.000 2543.390 1091.520 ;
      LAYER Nwell ;
        RECT 6.290 1083.680 2543.390 1088.000 ;
      LAYER Pwell ;
        RECT 6.290 1080.160 2543.390 1083.680 ;
      LAYER Nwell ;
        RECT 6.290 1075.840 2543.390 1080.160 ;
      LAYER Pwell ;
        RECT 6.290 1072.320 2543.390 1075.840 ;
      LAYER Nwell ;
        RECT 6.290 1068.000 2543.390 1072.320 ;
      LAYER Pwell ;
        RECT 6.290 1064.480 2543.390 1068.000 ;
      LAYER Nwell ;
        RECT 6.290 1060.160 2543.390 1064.480 ;
      LAYER Pwell ;
        RECT 6.290 1056.640 2543.390 1060.160 ;
      LAYER Nwell ;
        RECT 6.290 1052.320 2543.390 1056.640 ;
      LAYER Pwell ;
        RECT 6.290 1048.800 2543.390 1052.320 ;
      LAYER Nwell ;
        RECT 6.290 1044.480 2543.390 1048.800 ;
      LAYER Pwell ;
        RECT 6.290 1040.960 2543.390 1044.480 ;
      LAYER Nwell ;
        RECT 6.290 1036.640 2543.390 1040.960 ;
      LAYER Pwell ;
        RECT 6.290 1033.120 2543.390 1036.640 ;
      LAYER Nwell ;
        RECT 6.290 1028.800 2543.390 1033.120 ;
      LAYER Pwell ;
        RECT 6.290 1025.280 2543.390 1028.800 ;
      LAYER Nwell ;
        RECT 6.290 1020.960 2543.390 1025.280 ;
      LAYER Pwell ;
        RECT 6.290 1017.440 2543.390 1020.960 ;
      LAYER Nwell ;
        RECT 6.290 1013.120 2543.390 1017.440 ;
      LAYER Pwell ;
        RECT 6.290 1009.600 2543.390 1013.120 ;
      LAYER Nwell ;
        RECT 6.290 1005.280 2543.390 1009.600 ;
      LAYER Pwell ;
        RECT 6.290 1001.760 2543.390 1005.280 ;
      LAYER Nwell ;
        RECT 6.290 997.440 2543.390 1001.760 ;
      LAYER Pwell ;
        RECT 6.290 993.920 2543.390 997.440 ;
      LAYER Nwell ;
        RECT 6.290 989.600 2543.390 993.920 ;
      LAYER Pwell ;
        RECT 6.290 986.080 2543.390 989.600 ;
      LAYER Nwell ;
        RECT 6.290 981.760 2543.390 986.080 ;
      LAYER Pwell ;
        RECT 6.290 978.240 2543.390 981.760 ;
      LAYER Nwell ;
        RECT 6.290 973.920 2543.390 978.240 ;
      LAYER Pwell ;
        RECT 6.290 970.400 2543.390 973.920 ;
      LAYER Nwell ;
        RECT 6.290 966.080 2543.390 970.400 ;
      LAYER Pwell ;
        RECT 6.290 962.560 2543.390 966.080 ;
      LAYER Nwell ;
        RECT 6.290 958.240 2543.390 962.560 ;
      LAYER Pwell ;
        RECT 6.290 954.720 2543.390 958.240 ;
      LAYER Nwell ;
        RECT 6.290 950.400 2543.390 954.720 ;
      LAYER Pwell ;
        RECT 6.290 946.880 2543.390 950.400 ;
      LAYER Nwell ;
        RECT 6.290 942.560 2543.390 946.880 ;
      LAYER Pwell ;
        RECT 6.290 939.040 2543.390 942.560 ;
      LAYER Nwell ;
        RECT 6.290 934.720 2543.390 939.040 ;
      LAYER Pwell ;
        RECT 6.290 931.200 2543.390 934.720 ;
      LAYER Nwell ;
        RECT 6.290 926.880 2543.390 931.200 ;
      LAYER Pwell ;
        RECT 6.290 923.360 2543.390 926.880 ;
      LAYER Nwell ;
        RECT 6.290 919.040 2543.390 923.360 ;
      LAYER Pwell ;
        RECT 6.290 915.520 2543.390 919.040 ;
      LAYER Nwell ;
        RECT 6.290 911.200 2543.390 915.520 ;
      LAYER Pwell ;
        RECT 6.290 907.680 2543.390 911.200 ;
      LAYER Nwell ;
        RECT 6.290 903.360 2543.390 907.680 ;
      LAYER Pwell ;
        RECT 6.290 899.840 2543.390 903.360 ;
      LAYER Nwell ;
        RECT 6.290 895.520 2543.390 899.840 ;
      LAYER Pwell ;
        RECT 6.290 892.000 2543.390 895.520 ;
      LAYER Nwell ;
        RECT 6.290 887.680 2543.390 892.000 ;
      LAYER Pwell ;
        RECT 6.290 884.160 2543.390 887.680 ;
      LAYER Nwell ;
        RECT 6.290 879.840 2543.390 884.160 ;
      LAYER Pwell ;
        RECT 6.290 876.320 2543.390 879.840 ;
      LAYER Nwell ;
        RECT 6.290 872.000 2543.390 876.320 ;
      LAYER Pwell ;
        RECT 6.290 868.480 2543.390 872.000 ;
      LAYER Nwell ;
        RECT 6.290 864.160 2543.390 868.480 ;
      LAYER Pwell ;
        RECT 6.290 860.640 2543.390 864.160 ;
      LAYER Nwell ;
        RECT 6.290 856.320 2543.390 860.640 ;
      LAYER Pwell ;
        RECT 6.290 852.800 2543.390 856.320 ;
      LAYER Nwell ;
        RECT 6.290 848.480 2543.390 852.800 ;
      LAYER Pwell ;
        RECT 6.290 844.960 2543.390 848.480 ;
      LAYER Nwell ;
        RECT 6.290 840.640 2543.390 844.960 ;
      LAYER Pwell ;
        RECT 6.290 837.120 2543.390 840.640 ;
      LAYER Nwell ;
        RECT 6.290 832.800 2543.390 837.120 ;
      LAYER Pwell ;
        RECT 6.290 829.280 2543.390 832.800 ;
      LAYER Nwell ;
        RECT 6.290 824.960 2543.390 829.280 ;
      LAYER Pwell ;
        RECT 6.290 821.440 2543.390 824.960 ;
      LAYER Nwell ;
        RECT 6.290 817.120 2543.390 821.440 ;
      LAYER Pwell ;
        RECT 6.290 813.600 2543.390 817.120 ;
      LAYER Nwell ;
        RECT 6.290 809.280 2543.390 813.600 ;
      LAYER Pwell ;
        RECT 6.290 805.760 2543.390 809.280 ;
      LAYER Nwell ;
        RECT 6.290 801.440 2543.390 805.760 ;
      LAYER Pwell ;
        RECT 6.290 797.920 2543.390 801.440 ;
      LAYER Nwell ;
        RECT 6.290 793.600 2543.390 797.920 ;
      LAYER Pwell ;
        RECT 6.290 790.080 2543.390 793.600 ;
      LAYER Nwell ;
        RECT 6.290 785.760 2543.390 790.080 ;
      LAYER Pwell ;
        RECT 6.290 782.240 2543.390 785.760 ;
      LAYER Nwell ;
        RECT 6.290 777.920 2543.390 782.240 ;
      LAYER Pwell ;
        RECT 6.290 774.400 2543.390 777.920 ;
      LAYER Nwell ;
        RECT 6.290 770.080 2543.390 774.400 ;
      LAYER Pwell ;
        RECT 6.290 766.560 2543.390 770.080 ;
      LAYER Nwell ;
        RECT 6.290 762.240 2543.390 766.560 ;
      LAYER Pwell ;
        RECT 6.290 758.720 2543.390 762.240 ;
      LAYER Nwell ;
        RECT 6.290 754.400 2543.390 758.720 ;
      LAYER Pwell ;
        RECT 6.290 750.880 2543.390 754.400 ;
      LAYER Nwell ;
        RECT 6.290 746.560 2543.390 750.880 ;
      LAYER Pwell ;
        RECT 6.290 743.040 2543.390 746.560 ;
      LAYER Nwell ;
        RECT 6.290 738.720 2543.390 743.040 ;
      LAYER Pwell ;
        RECT 6.290 735.200 2543.390 738.720 ;
      LAYER Nwell ;
        RECT 6.290 730.880 2543.390 735.200 ;
      LAYER Pwell ;
        RECT 6.290 727.360 2543.390 730.880 ;
      LAYER Nwell ;
        RECT 6.290 723.040 2543.390 727.360 ;
      LAYER Pwell ;
        RECT 6.290 719.520 2543.390 723.040 ;
      LAYER Nwell ;
        RECT 6.290 715.200 2543.390 719.520 ;
      LAYER Pwell ;
        RECT 6.290 711.680 2543.390 715.200 ;
      LAYER Nwell ;
        RECT 6.290 707.360 2543.390 711.680 ;
      LAYER Pwell ;
        RECT 6.290 703.840 2543.390 707.360 ;
      LAYER Nwell ;
        RECT 6.290 699.520 2543.390 703.840 ;
      LAYER Pwell ;
        RECT 6.290 696.000 2543.390 699.520 ;
      LAYER Nwell ;
        RECT 6.290 691.680 2543.390 696.000 ;
      LAYER Pwell ;
        RECT 6.290 688.160 2543.390 691.680 ;
      LAYER Nwell ;
        RECT 6.290 683.840 2543.390 688.160 ;
      LAYER Pwell ;
        RECT 6.290 680.320 2543.390 683.840 ;
      LAYER Nwell ;
        RECT 6.290 676.000 2543.390 680.320 ;
      LAYER Pwell ;
        RECT 6.290 672.480 2543.390 676.000 ;
      LAYER Nwell ;
        RECT 6.290 668.160 2543.390 672.480 ;
      LAYER Pwell ;
        RECT 6.290 664.640 2543.390 668.160 ;
      LAYER Nwell ;
        RECT 6.290 660.320 2543.390 664.640 ;
      LAYER Pwell ;
        RECT 6.290 656.800 2543.390 660.320 ;
      LAYER Nwell ;
        RECT 6.290 652.480 2543.390 656.800 ;
      LAYER Pwell ;
        RECT 6.290 648.960 2543.390 652.480 ;
      LAYER Nwell ;
        RECT 6.290 644.640 2543.390 648.960 ;
      LAYER Pwell ;
        RECT 6.290 641.120 2543.390 644.640 ;
      LAYER Nwell ;
        RECT 6.290 636.800 2543.390 641.120 ;
      LAYER Pwell ;
        RECT 6.290 633.280 2543.390 636.800 ;
      LAYER Nwell ;
        RECT 6.290 628.960 2543.390 633.280 ;
      LAYER Pwell ;
        RECT 6.290 625.440 2543.390 628.960 ;
      LAYER Nwell ;
        RECT 6.290 621.120 2543.390 625.440 ;
      LAYER Pwell ;
        RECT 6.290 617.600 2543.390 621.120 ;
      LAYER Nwell ;
        RECT 6.290 613.280 2543.390 617.600 ;
      LAYER Pwell ;
        RECT 6.290 609.760 2543.390 613.280 ;
      LAYER Nwell ;
        RECT 6.290 605.440 2543.390 609.760 ;
      LAYER Pwell ;
        RECT 6.290 601.920 2543.390 605.440 ;
      LAYER Nwell ;
        RECT 6.290 597.600 2543.390 601.920 ;
      LAYER Pwell ;
        RECT 6.290 594.080 2543.390 597.600 ;
      LAYER Nwell ;
        RECT 6.290 589.760 2543.390 594.080 ;
      LAYER Pwell ;
        RECT 6.290 586.240 2543.390 589.760 ;
      LAYER Nwell ;
        RECT 6.290 581.920 2543.390 586.240 ;
      LAYER Pwell ;
        RECT 6.290 578.400 2543.390 581.920 ;
      LAYER Nwell ;
        RECT 6.290 574.080 2543.390 578.400 ;
      LAYER Pwell ;
        RECT 6.290 570.560 2543.390 574.080 ;
      LAYER Nwell ;
        RECT 6.290 566.240 2543.390 570.560 ;
      LAYER Pwell ;
        RECT 6.290 562.720 2543.390 566.240 ;
      LAYER Nwell ;
        RECT 6.290 558.400 2543.390 562.720 ;
      LAYER Pwell ;
        RECT 6.290 554.880 2543.390 558.400 ;
      LAYER Nwell ;
        RECT 6.290 550.560 2543.390 554.880 ;
      LAYER Pwell ;
        RECT 6.290 547.040 2543.390 550.560 ;
      LAYER Nwell ;
        RECT 6.290 542.720 2543.390 547.040 ;
      LAYER Pwell ;
        RECT 6.290 539.200 2543.390 542.720 ;
      LAYER Nwell ;
        RECT 6.290 534.880 2543.390 539.200 ;
      LAYER Pwell ;
        RECT 6.290 531.360 2543.390 534.880 ;
      LAYER Nwell ;
        RECT 6.290 527.040 2543.390 531.360 ;
      LAYER Pwell ;
        RECT 6.290 523.520 2543.390 527.040 ;
      LAYER Nwell ;
        RECT 6.290 519.200 2543.390 523.520 ;
      LAYER Pwell ;
        RECT 6.290 515.680 2543.390 519.200 ;
      LAYER Nwell ;
        RECT 6.290 511.360 2543.390 515.680 ;
      LAYER Pwell ;
        RECT 6.290 507.840 2543.390 511.360 ;
      LAYER Nwell ;
        RECT 6.290 503.520 2543.390 507.840 ;
      LAYER Pwell ;
        RECT 6.290 500.000 2543.390 503.520 ;
      LAYER Nwell ;
        RECT 6.290 495.680 2543.390 500.000 ;
      LAYER Pwell ;
        RECT 6.290 492.160 2543.390 495.680 ;
      LAYER Nwell ;
        RECT 6.290 487.840 2543.390 492.160 ;
      LAYER Pwell ;
        RECT 6.290 484.320 2543.390 487.840 ;
      LAYER Nwell ;
        RECT 6.290 480.000 2543.390 484.320 ;
      LAYER Pwell ;
        RECT 6.290 476.480 2543.390 480.000 ;
      LAYER Nwell ;
        RECT 6.290 472.160 2543.390 476.480 ;
      LAYER Pwell ;
        RECT 6.290 468.640 2543.390 472.160 ;
      LAYER Nwell ;
        RECT 6.290 464.320 2543.390 468.640 ;
      LAYER Pwell ;
        RECT 6.290 460.800 2543.390 464.320 ;
      LAYER Nwell ;
        RECT 6.290 456.480 2543.390 460.800 ;
      LAYER Pwell ;
        RECT 6.290 452.960 2543.390 456.480 ;
      LAYER Nwell ;
        RECT 6.290 448.640 2543.390 452.960 ;
      LAYER Pwell ;
        RECT 6.290 445.120 2543.390 448.640 ;
      LAYER Nwell ;
        RECT 6.290 440.800 2543.390 445.120 ;
      LAYER Pwell ;
        RECT 6.290 437.280 2543.390 440.800 ;
      LAYER Nwell ;
        RECT 6.290 432.960 2543.390 437.280 ;
      LAYER Pwell ;
        RECT 6.290 429.440 2543.390 432.960 ;
      LAYER Nwell ;
        RECT 6.290 425.120 2543.390 429.440 ;
      LAYER Pwell ;
        RECT 6.290 421.600 2543.390 425.120 ;
      LAYER Nwell ;
        RECT 6.290 417.280 2543.390 421.600 ;
      LAYER Pwell ;
        RECT 6.290 413.760 2543.390 417.280 ;
      LAYER Nwell ;
        RECT 6.290 409.440 2543.390 413.760 ;
      LAYER Pwell ;
        RECT 6.290 405.920 2543.390 409.440 ;
      LAYER Nwell ;
        RECT 6.290 401.600 2543.390 405.920 ;
      LAYER Pwell ;
        RECT 6.290 398.080 2543.390 401.600 ;
      LAYER Nwell ;
        RECT 6.290 393.760 2543.390 398.080 ;
      LAYER Pwell ;
        RECT 6.290 390.240 2543.390 393.760 ;
      LAYER Nwell ;
        RECT 6.290 385.920 2543.390 390.240 ;
      LAYER Pwell ;
        RECT 6.290 382.400 2543.390 385.920 ;
      LAYER Nwell ;
        RECT 6.290 378.080 2543.390 382.400 ;
      LAYER Pwell ;
        RECT 6.290 374.560 2543.390 378.080 ;
      LAYER Nwell ;
        RECT 6.290 370.240 2543.390 374.560 ;
      LAYER Pwell ;
        RECT 6.290 366.720 2543.390 370.240 ;
      LAYER Nwell ;
        RECT 6.290 362.400 2543.390 366.720 ;
      LAYER Pwell ;
        RECT 6.290 358.880 2543.390 362.400 ;
      LAYER Nwell ;
        RECT 6.290 354.560 2543.390 358.880 ;
      LAYER Pwell ;
        RECT 6.290 351.040 2543.390 354.560 ;
      LAYER Nwell ;
        RECT 6.290 346.720 2543.390 351.040 ;
      LAYER Pwell ;
        RECT 6.290 343.200 2543.390 346.720 ;
      LAYER Nwell ;
        RECT 6.290 338.880 2543.390 343.200 ;
      LAYER Pwell ;
        RECT 6.290 335.360 2543.390 338.880 ;
      LAYER Nwell ;
        RECT 6.290 331.040 2543.390 335.360 ;
      LAYER Pwell ;
        RECT 6.290 327.520 2543.390 331.040 ;
      LAYER Nwell ;
        RECT 6.290 323.200 2543.390 327.520 ;
      LAYER Pwell ;
        RECT 6.290 319.680 2543.390 323.200 ;
      LAYER Nwell ;
        RECT 6.290 315.360 2543.390 319.680 ;
      LAYER Pwell ;
        RECT 6.290 311.840 2543.390 315.360 ;
      LAYER Nwell ;
        RECT 6.290 307.520 2543.390 311.840 ;
      LAYER Pwell ;
        RECT 6.290 304.000 2543.390 307.520 ;
      LAYER Nwell ;
        RECT 6.290 299.680 2543.390 304.000 ;
      LAYER Pwell ;
        RECT 6.290 296.160 2543.390 299.680 ;
      LAYER Nwell ;
        RECT 6.290 291.840 2543.390 296.160 ;
      LAYER Pwell ;
        RECT 6.290 288.320 2543.390 291.840 ;
      LAYER Nwell ;
        RECT 6.290 284.000 2543.390 288.320 ;
      LAYER Pwell ;
        RECT 6.290 280.480 2543.390 284.000 ;
      LAYER Nwell ;
        RECT 6.290 276.160 2543.390 280.480 ;
      LAYER Pwell ;
        RECT 6.290 272.640 2543.390 276.160 ;
      LAYER Nwell ;
        RECT 6.290 268.320 2543.390 272.640 ;
      LAYER Pwell ;
        RECT 6.290 264.800 2543.390 268.320 ;
      LAYER Nwell ;
        RECT 6.290 260.480 2543.390 264.800 ;
      LAYER Pwell ;
        RECT 6.290 256.960 2543.390 260.480 ;
      LAYER Nwell ;
        RECT 6.290 252.640 2543.390 256.960 ;
      LAYER Pwell ;
        RECT 6.290 249.120 2543.390 252.640 ;
      LAYER Nwell ;
        RECT 6.290 244.800 2543.390 249.120 ;
      LAYER Pwell ;
        RECT 6.290 241.280 2543.390 244.800 ;
      LAYER Nwell ;
        RECT 6.290 236.960 2543.390 241.280 ;
      LAYER Pwell ;
        RECT 6.290 233.440 2543.390 236.960 ;
      LAYER Nwell ;
        RECT 6.290 229.120 2543.390 233.440 ;
      LAYER Pwell ;
        RECT 6.290 225.600 2543.390 229.120 ;
      LAYER Nwell ;
        RECT 6.290 221.280 2543.390 225.600 ;
      LAYER Pwell ;
        RECT 6.290 217.760 2543.390 221.280 ;
      LAYER Nwell ;
        RECT 6.290 213.440 2543.390 217.760 ;
      LAYER Pwell ;
        RECT 6.290 209.920 2543.390 213.440 ;
      LAYER Nwell ;
        RECT 6.290 205.600 2543.390 209.920 ;
      LAYER Pwell ;
        RECT 6.290 202.080 2543.390 205.600 ;
      LAYER Nwell ;
        RECT 6.290 197.760 2543.390 202.080 ;
      LAYER Pwell ;
        RECT 6.290 194.240 2543.390 197.760 ;
      LAYER Nwell ;
        RECT 6.290 189.920 2543.390 194.240 ;
      LAYER Pwell ;
        RECT 6.290 186.400 2543.390 189.920 ;
      LAYER Nwell ;
        RECT 6.290 182.080 2543.390 186.400 ;
      LAYER Pwell ;
        RECT 6.290 178.560 2543.390 182.080 ;
      LAYER Nwell ;
        RECT 6.290 174.240 2543.390 178.560 ;
      LAYER Pwell ;
        RECT 6.290 170.720 2543.390 174.240 ;
      LAYER Nwell ;
        RECT 6.290 166.400 2543.390 170.720 ;
      LAYER Pwell ;
        RECT 6.290 162.880 2543.390 166.400 ;
      LAYER Nwell ;
        RECT 6.290 158.560 2543.390 162.880 ;
      LAYER Pwell ;
        RECT 6.290 155.040 2543.390 158.560 ;
      LAYER Nwell ;
        RECT 6.290 150.720 2543.390 155.040 ;
      LAYER Pwell ;
        RECT 6.290 147.200 2543.390 150.720 ;
      LAYER Nwell ;
        RECT 6.290 142.880 2543.390 147.200 ;
      LAYER Pwell ;
        RECT 6.290 139.360 2543.390 142.880 ;
      LAYER Nwell ;
        RECT 6.290 135.040 2543.390 139.360 ;
      LAYER Pwell ;
        RECT 6.290 131.520 2543.390 135.040 ;
      LAYER Nwell ;
        RECT 6.290 127.200 2543.390 131.520 ;
      LAYER Pwell ;
        RECT 6.290 123.680 2543.390 127.200 ;
      LAYER Nwell ;
        RECT 6.290 119.360 2543.390 123.680 ;
      LAYER Pwell ;
        RECT 6.290 115.840 2543.390 119.360 ;
      LAYER Nwell ;
        RECT 6.290 111.520 2543.390 115.840 ;
      LAYER Pwell ;
        RECT 6.290 108.000 2543.390 111.520 ;
      LAYER Nwell ;
        RECT 6.290 103.680 2543.390 108.000 ;
      LAYER Pwell ;
        RECT 6.290 100.160 2543.390 103.680 ;
      LAYER Nwell ;
        RECT 6.290 95.840 2543.390 100.160 ;
      LAYER Pwell ;
        RECT 6.290 92.320 2543.390 95.840 ;
      LAYER Nwell ;
        RECT 6.290 88.000 2543.390 92.320 ;
      LAYER Pwell ;
        RECT 6.290 84.480 2543.390 88.000 ;
      LAYER Nwell ;
        RECT 6.290 80.160 2543.390 84.480 ;
      LAYER Pwell ;
        RECT 6.290 76.640 2543.390 80.160 ;
      LAYER Nwell ;
        RECT 6.290 72.320 2543.390 76.640 ;
      LAYER Pwell ;
        RECT 6.290 68.800 2543.390 72.320 ;
      LAYER Nwell ;
        RECT 6.290 64.480 2543.390 68.800 ;
      LAYER Pwell ;
        RECT 6.290 60.960 2543.390 64.480 ;
      LAYER Nwell ;
        RECT 6.290 56.640 2543.390 60.960 ;
      LAYER Pwell ;
        RECT 6.290 53.120 2543.390 56.640 ;
      LAYER Nwell ;
        RECT 6.290 48.800 2543.390 53.120 ;
      LAYER Pwell ;
        RECT 6.290 45.280 2543.390 48.800 ;
      LAYER Nwell ;
        RECT 6.290 40.960 2543.390 45.280 ;
      LAYER Pwell ;
        RECT 6.290 37.440 2543.390 40.960 ;
      LAYER Nwell ;
        RECT 6.290 33.120 2543.390 37.440 ;
      LAYER Pwell ;
        RECT 6.290 29.600 2543.390 33.120 ;
      LAYER Nwell ;
        RECT 6.290 25.280 2543.390 29.600 ;
      LAYER Pwell ;
        RECT 6.290 21.760 2543.390 25.280 ;
      LAYER Nwell ;
        RECT 6.290 17.440 2543.390 21.760 ;
      LAYER Pwell ;
        RECT 6.290 15.250 2543.390 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 2542.960 1732.940 ;
      LAYER Metal2 ;
        RECT 20.040 1745.700 1273.140 1746.000 ;
        RECT 1274.300 1745.700 2526.040 1746.000 ;
        RECT 20.040 4.300 2526.040 1745.700 ;
        RECT 20.040 4.000 1269.780 4.300 ;
        RECT 1270.940 4.000 1273.140 4.300 ;
        RECT 1274.300 4.000 2526.040 4.300 ;
      LAYER Metal3 ;
        RECT 19.990 4.620 2526.090 1732.780 ;
  END
END analog_wrapper
END LIBRARY

