* NGSPICE file created from serv_rf_top.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 ZN VSS VDD C2 C1 B2 B1 A2 VNW VPW
X0 ZN A2 a_1812_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X1 a_224_472# C2 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X2 ZN A1 a_4876_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
X3 a_1812_472# A1 ZN VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X4 a_2010_68# B1 ZN VPW nfet_06v0 ad=0.152p pd=1.19u as=0.488p ps=2.01u w=0.82u l=0.6u
X5 VSS A2 a_3652_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X6 a_3652_68# A1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X7 VDD C1 a_224_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X8 a_244_68# C1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
X9 VSS C2 a_244_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X10 a_1812_472# B2 a_224_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X11 a_1468_68# C2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X12 a_2428_68# B2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X13 a_224_472# C1 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X14 a_4468_68# A1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X15 a_224_472# B2 a_1812_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X16 a_224_472# B1 a_1812_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.537p ps=3.32u w=1.22u l=0.5u
X17 a_4060_68# A2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X18 a_1812_472# B1 a_224_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X19 a_652_68# C2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X20 ZN C1 a_652_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X21 VDD C2 a_224_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X22 a_2836_68# B1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X23 a_224_472# B2 a_1812_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X24 a_224_472# B1 a_1812_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X25 VSS C2 a_1060_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X26 a_224_472# C2 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X27 VSS B2 a_2010_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.152p ps=1.19u w=0.82u l=0.6u
X28 a_4876_68# A2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X29 a_1812_472# B1 a_224_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X30 a_1812_472# B2 a_224_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X31 a_1060_68# C1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X32 ZN A1 a_4060_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X33 VDD C1 a_224_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X34 ZN A1 a_1812_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X35 a_1812_472# A1 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X36 ZN C1 a_1468_68# VPW nfet_06v0 ad=0.488p pd=2.01u as=0.131p ps=1.14u w=0.82u l=0.6u
X37 a_1812_472# A2 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X38 ZN B1 a_2428_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X39 ZN A2 a_1812_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X40 ZN A1 a_1812_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X41 VSS A2 a_4468_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X42 a_224_472# C1 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.537p ps=3.32u w=1.22u l=0.5u
X43 a_1812_472# A2 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X44 ZN B1 a_3244_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X45 a_3244_68# B2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X46 VDD C2 a_224_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X47 VSS B2 a_2836_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__antenna VSS I VDD VNW VPW
D0 VPW I diode_nd2ps_06v0 pj=1.86u area=0.205p
D1 I VNW diode_pd2nw_06v0 pj=1.86u area=0.205p
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS VNW VPW
X0 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X1 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A2 VDD VNW pfet_06v0 ad=0.294p pd=1.65u as=0.497p ps=3.14u w=1.13u l=0.5u
X1 ZN A1 a_245_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
X2 VDD A1 ZN VNW pfet_06v0 ad=0.497p pd=3.14u as=0.294p ps=1.65u w=1.13u l=0.5u
X3 a_245_68# A2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 VDD VSS ZN A1 A2 VNW VPW
X0 a_1140_472# A2 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
X1 ZN A1 VSS VPW nfet_06v0 ad=0.147p pd=1.09u as=0.147p ps=1.09u w=0.565u l=0.6u
X2 ZN A1 a_1140_472# VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X3 ZN A2 VSS VPW nfet_06v0 ad=0.147p pd=1.09u as=0.249p ps=2.01u w=0.565u l=0.6u
X4 a_1588_472# A1 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
X5 VDD A2 a_1588_472# VNW pfet_06v0 ad=0.598p pd=3.42u as=0.317p ps=1.74u w=1.22u l=0.5u
X6 ZN A1 VSS VPW nfet_06v0 ad=0.147p pd=1.09u as=0.147p ps=1.09u w=0.565u l=0.6u
X7 a_244_472# A2 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.598p ps=3.42u w=1.22u l=0.5u
X8 ZN A1 a_244_472# VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X9 a_692_472# A1 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
X10 VSS A2 ZN VPW nfet_06v0 ad=0.249p pd=2.01u as=0.147p ps=1.09u w=0.565u l=0.6u
X11 VDD A2 a_692_472# VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X12 VSS A1 ZN VPW nfet_06v0 ad=0.147p pd=1.09u as=0.147p ps=1.09u w=0.565u l=0.6u
X13 VSS A2 ZN VPW nfet_06v0 ad=0.147p pd=1.09u as=0.147p ps=1.09u w=0.565u l=0.6u
X14 VSS A1 ZN VPW nfet_06v0 ad=0.147p pd=1.09u as=0.147p ps=1.09u w=0.565u l=0.6u
X15 ZN A2 VSS VPW nfet_06v0 ad=0.147p pd=1.09u as=0.147p ps=1.09u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 VDD B A2 ZN A1 VSS VNW VPW
X0 VSS B a_36_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X2 VDD B ZN VNW pfet_06v0 ad=0.497p pd=3.14u as=0.425p ps=1.94u w=1.13u l=0.5u
X3 a_244_472# A2 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.598p ps=3.42u w=1.22u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.425p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 B1 B2 VDD VSS ZN A1 A2 C VNW VPW
X0 a_56_492# A2 ZN VNW pfet_06v0 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.5u
X1 a_512_68# B2 VSS VPW nfet_06v0 ad=0.164p pd=1.17u as=0.218p ps=1.45u w=0.715u l=0.6u
X2 ZN C VSS VPW nfet_06v0 ad=0.234p pd=1.43u as=0.652p ps=2.69u w=0.575u l=0.6u
X3 a_244_492# B2 VDD VNW pfet_06v0 ad=0.706p pd=2.38u as=0.566p ps=2.24u w=1.12u l=0.5u
X4 a_948_68# B1 ZN VPW nfet_06v0 ad=0.107p pd=1.01u as=0.186p ps=1.24u w=0.715u l=0.6u
X5 VSS B2 a_948_68# VPW nfet_06v0 ad=0.652p pd=2.69u as=0.107p ps=1.01u w=0.715u l=0.6u
X6 a_56_492# C a_244_492# VNW pfet_06v0 ad=0.311p pd=1.67u as=0.706p ps=2.38u w=1.12u l=0.5u
X7 VSS C ZN VPW nfet_06v0 ad=0.218p pd=1.45u as=0.178p ps=1.69u w=0.405u l=0.6u
X8 VDD B1 a_244_492# VNW pfet_06v0 ad=0.566p pd=2.24u as=0.302p ps=1.66u w=1.12u l=0.5u
X9 a_2267_68# A2 VSS VPW nfet_06v0 ad=85.8f pd=0.955u as=0.186p ps=1.24u w=0.715u l=0.6u
X10 a_1875_68# A1 ZN VPW nfet_06v0 ad=85.8f pd=0.955u as=0.234p ps=1.43u w=0.715u l=0.6u
X11 VSS A2 a_1875_68# VPW nfet_06v0 ad=0.186p pd=1.24u as=85.8f ps=0.955u w=0.715u l=0.6u
X12 ZN A1 a_2267_68# VPW nfet_06v0 ad=0.315p pd=2.31u as=85.8f ps=0.955u w=0.715u l=0.6u
X13 a_244_492# B1 VDD VNW pfet_06v0 ad=0.302p pd=1.66u as=0.566p ps=2.24u w=1.12u l=0.5u
X14 ZN B1 a_512_68# VPW nfet_06v0 ad=0.186p pd=1.24u as=0.164p ps=1.17u w=0.715u l=0.6u
X15 a_244_492# C a_56_492# VNW pfet_06v0 ad=0.291p pd=1.64u as=0.493p ps=3.12u w=1.12u l=0.5u
X16 ZN A2 a_56_492# VNW pfet_06v0 ad=0.291p pd=1.64u as=0.291p ps=1.64u w=1.12u l=0.5u
X17 VDD B2 a_244_492# VNW pfet_06v0 ad=0.566p pd=2.24u as=0.291p ps=1.64u w=1.12u l=0.5u
X18 ZN A1 a_56_492# VNW pfet_06v0 ad=0.291p pd=1.64u as=0.311p ps=1.67u w=1.12u l=0.5u
X19 a_56_492# A1 ZN VNW pfet_06v0 ad=0.493p pd=3.12u as=0.291p ps=1.64u w=1.12u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 B2 B1 A2 A1 ZN VSS VDD C2 C1 VNW VPW
X0 VSS C2 a_251_68# VPW nfet_06v0 ad=0.316p pd=1.59u as=96f ps=1.04u w=0.8u l=0.6u
X1 ZN C1 a_697_68# VPW nfet_06v0 ad=0.384p pd=1.76u as=0.124p ps=1.11u w=0.8u l=0.6u
X2 a_231_472# C1 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.537p ps=3.32u w=1.22u l=0.5u
X3 a_1003_472# B2 a_231_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X4 ZN A2 a_1003_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X5 ZN A1 a_1003_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.326p ps=1.75u w=1.22u l=0.5u
X6 VSS B2 a_1191_68# VPW nfet_06v0 ad=0.208p pd=1.32u as=0.168p ps=1.22u w=0.8u l=0.6u
X7 a_231_472# B2 a_1003_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X8 a_1003_472# A1 ZN VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X9 VDD C2 a_231_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X10 a_231_472# C2 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X11 ZN B1 a_1619_68# VPW nfet_06v0 ad=0.214p pd=1.34u as=0.128p ps=1.12u w=0.8u l=0.6u
X12 VDD C1 a_231_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X13 a_2438_68# A2 VSS VPW nfet_06v0 ad=0.128p pd=1.12u as=0.208p ps=1.32u w=0.8u l=0.6u
X14 a_2030_68# A1 ZN VPW nfet_06v0 ad=0.128p pd=1.12u as=0.214p ps=1.34u w=0.8u l=0.6u
X15 a_251_68# C1 ZN VPW nfet_06v0 ad=96f pd=1.04u as=0.352p ps=2.48u w=0.8u l=0.6u
X16 a_1003_472# B1 a_231_472# VNW pfet_06v0 ad=0.326p pd=1.75u as=0.317p ps=1.74u w=1.22u l=0.5u
X17 VSS A2 a_2030_68# VPW nfet_06v0 ad=0.208p pd=1.32u as=0.128p ps=1.12u w=0.8u l=0.6u
X18 a_1191_68# B1 ZN VPW nfet_06v0 ad=0.168p pd=1.22u as=0.384p ps=1.76u w=0.8u l=0.6u
X19 a_1619_68# B2 VSS VPW nfet_06v0 ad=0.128p pd=1.12u as=0.208p ps=1.32u w=0.8u l=0.6u
X20 ZN A1 a_2438_68# VPW nfet_06v0 ad=0.352p pd=2.48u as=0.128p ps=1.12u w=0.8u l=0.6u
X21 a_231_472# B1 a_1003_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.537p ps=3.32u w=1.22u l=0.5u
X22 a_697_68# C2 VSS VPW nfet_06v0 ad=0.124p pd=1.11u as=0.316p ps=1.59u w=0.8u l=0.6u
X23 a_1003_472# A2 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X3 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X4 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X5 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X6 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X7 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X1 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X2 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X3 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X4 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X5 a_1916_375# a_1828_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X6 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X7 a_2812_375# a_2724_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X8 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X9 a_2364_375# a_2276_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X10 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X11 a_3260_375# a_3172_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X12 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X13 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X14 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X15 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS VNW VPW
X0 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X1 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X2 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X3 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 B VDD VSS ZN A1 A2 VNW VPW
X0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.257p pd=1.56u as=0.131p ps=1.14u w=0.82u l=0.6u
X2 VDD B a_36_472# VNW pfet_06v0 ad=0.535p pd=3.31u as=0.45p ps=1.96u w=1.22u l=0.5u
X3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.535p ps=3.31u w=1.22u l=0.5u
X4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.45p pd=1.96u as=0.316p ps=1.74u w=1.22u l=0.5u
X5 VSS B ZN VPW nfet_06v0 ad=0.224p pd=1.9u as=0.257p ps=1.56u w=0.51u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 B VDD VSS ZN A1 A2 VNW VPW
X0 VSS A2 a_1133_69# VPW nfet_06v0 ad=0.341p pd=2.43u as=93f ps=1.01u w=0.775u l=0.6u
X1 VDD B a_49_472# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.535p ps=3.31u w=1.22u l=0.5u
X2 ZN A1 a_49_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.328p ps=1.75u w=1.22u l=0.5u
X3 a_741_69# A2 VSS VPW nfet_06v0 ad=93f pd=1.01u as=0.24p ps=1.48u w=0.775u l=0.6u
X4 a_49_472# A1 ZN VNW pfet_06v0 ad=0.328p pd=1.75u as=0.377p ps=1.83u w=1.22u l=0.5u
X5 ZN B VSS VPW nfet_06v0 ad=0.147p pd=1.09u as=0.249p ps=2.01u w=0.565u l=0.6u
X6 a_49_472# A2 ZN VNW pfet_06v0 ad=0.535p pd=3.31u as=0.316p ps=1.74u w=1.22u l=0.5u
X7 a_49_472# B VDD VNW pfet_06v0 ad=0.316p pd=1.74u as=0.377p ps=1.83u w=1.22u l=0.5u
X8 ZN A2 a_49_472# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.316p ps=1.74u w=1.22u l=0.5u
X9 VSS B ZN VPW nfet_06v0 ad=0.24p pd=1.48u as=0.147p ps=1.09u w=0.565u l=0.6u
X10 ZN A1 a_741_69# VPW nfet_06v0 ad=0.201p pd=1.29u as=93f ps=1.01u w=0.775u l=0.6u
X11 a_1133_69# A1 ZN VPW nfet_06v0 ad=93f pd=1.01u as=0.201p ps=1.29u w=0.775u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A2 B1 B2 C VDD VSS ZN A1 VNW VPW
X0 VSS B2 a_1070_69# VPW nfet_06v0 ad=0.2p pd=1.29u as=0.123p ps=1.09u w=0.77u l=0.6u
X1 VDD B2 a_234_508# VNW pfet_06v0 ad=0.269p pd=1.55u as=0.269p ps=1.55u w=1.03u l=0.5u
X2 VSS A2 a_3728_69# VPW nfet_06v0 ad=0.2p pd=1.29u as=0.123p ps=1.09u w=0.77u l=0.6u
X3 a_234_508# C a_1822_472# VNW pfet_06v0 ad=0.346p pd=1.78u as=0.316p ps=1.74u w=1.22u l=0.5u
X4 a_1822_472# A1 ZN VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X5 a_234_508# C a_1822_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.535p ps=3.31u w=1.22u l=0.5u
X6 ZN A2 a_1822_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X7 a_1070_69# B1 ZN VPW nfet_06v0 ad=0.123p pd=1.09u as=0.2p ps=1.29u w=0.77u l=0.6u
X8 a_234_508# B2 VDD VNW pfet_06v0 ad=0.269p pd=1.55u as=0.269p ps=1.55u w=1.03u l=0.5u
X9 ZN A1 a_1822_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X10 a_1822_472# A1 ZN VNW pfet_06v0 ad=0.535p pd=3.31u as=0.316p ps=1.74u w=1.22u l=0.5u
X11 VDD B1 a_234_508# VNW pfet_06v0 ad=0.455p pd=2.95u as=0.269p ps=1.55u w=1.03u l=0.5u
X12 a_1822_472# A2 ZN VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X13 a_2912_69# A1 ZN VPW nfet_06v0 ad=0.123p pd=1.09u as=0.226p ps=1.47u w=0.77u l=0.6u
X14 VSS A2 a_2912_69# VPW nfet_06v0 ad=0.2p pd=1.29u as=0.123p ps=1.09u w=0.77u l=0.6u
X15 a_234_508# B1 VDD VNW pfet_06v0 ad=0.269p pd=1.55u as=0.455p ps=2.95u w=1.03u l=0.5u
X16 a_3728_69# A1 ZN VPW nfet_06v0 ad=0.123p pd=1.09u as=0.2p ps=1.29u w=0.77u l=0.6u
X17 ZN A1 a_4136_69# VPW nfet_06v0 ad=0.339p pd=2.42u as=0.123p ps=1.09u w=0.77u l=0.6u
X18 a_244_69# B1 ZN VPW nfet_06v0 ad=0.142p pd=1.14u as=0.339p ps=2.42u w=0.77u l=0.6u
X19 VSS C ZN VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
X20 VDD B2 a_234_508# VNW pfet_06v0 ad=0.269p pd=1.55u as=0.269p ps=1.55u w=1.03u l=0.5u
X21 ZN B1 a_1478_69# VPW nfet_06v0 ad=0.299p pd=1.66u as=0.162p ps=1.19u w=0.77u l=0.6u
X22 a_234_508# B2 VDD VNW pfet_06v0 ad=0.269p pd=1.55u as=0.269p ps=1.55u w=1.03u l=0.5u
X23 VSS B2 a_244_69# VPW nfet_06v0 ad=0.2p pd=1.29u as=0.142p ps=1.14u w=0.77u l=0.6u
X24 a_1478_69# B2 VSS VPW nfet_06v0 ad=0.162p pd=1.19u as=0.2p ps=1.29u w=0.77u l=0.6u
X25 VDD B1 a_234_508# VNW pfet_06v0 ad=0.269p pd=1.55u as=0.269p ps=1.55u w=1.03u l=0.5u
X26 ZN A1 a_1822_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.486p ps=2.02u w=1.22u l=0.5u
X27 ZN C VSS VPW nfet_06v0 ad=0.226p pd=1.47u as=0.125p ps=1u w=0.48u l=0.6u
X28 a_3320_69# A2 VSS VPW nfet_06v0 ad=0.123p pd=1.09u as=0.2p ps=1.29u w=0.77u l=0.6u
X29 ZN A1 a_3320_69# VPW nfet_06v0 ad=0.2p pd=1.29u as=0.123p ps=1.09u w=0.77u l=0.6u
X30 a_234_508# B1 VDD VNW pfet_06v0 ad=0.269p pd=1.55u as=0.269p ps=1.55u w=1.03u l=0.5u
X31 ZN C VSS VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
X32 a_1822_472# C a_234_508# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.346p ps=1.78u w=1.22u l=0.5u
X33 a_1822_472# A2 ZN VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X34 ZN B1 a_662_69# VPW nfet_06v0 ad=0.2p pd=1.29u as=0.123p ps=1.09u w=0.77u l=0.6u
X35 a_662_69# B2 VSS VPW nfet_06v0 ad=0.123p pd=1.09u as=0.2p ps=1.29u w=0.77u l=0.6u
X36 VSS C ZN VPW nfet_06v0 ad=0.125p pd=1u as=0.299p ps=1.66u w=0.48u l=0.6u
X37 a_1822_472# C a_234_508# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X38 ZN A2 a_1822_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X39 a_4136_69# A2 VSS VPW nfet_06v0 ad=0.123p pd=1.09u as=0.2p ps=1.29u w=0.77u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 VDD Q CLK VSS D VNW VPW
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.105p pd=0.925u as=0.178p ps=1.69u w=0.405u l=0.6u
X1 Q a_2304_115# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=0.6u
X2 a_2304_115# a_2011_527# VSS VPW nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X3 a_1004_159# D a_836_159# VPW nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X4 a_1004_159# D a_880_527# VNW pfet_06v0 ad=0.187p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X5 a_2011_527# a_36_151# a_1376_115# VNW pfet_06v0 ad=0.166p pd=1.28u as=0.179p ps=1.36u w=0.36u l=0.5u
X6 a_2296_527# a_448_472# a_2011_527# VNW pfet_06v0 ad=50.4f pd=0.64u as=0.166p ps=1.28u w=0.36u l=0.5u
X7 a_1376_115# a_1004_159# VDD VNW pfet_06v0 ad=0.179p pd=1.36u as=0.104p ps=0.94u w=0.36u l=0.5u
X8 VDD CLK a_36_151# VNW pfet_06v0 ad=0.225p pd=1.38u as=0.381p ps=2.61u w=0.865u l=0.5u
X9 VSS a_1376_115# a_1328_159# VPW nfet_06v0 ad=0.264p pd=1.82u as=43.2f ps=0.6u w=0.36u l=0.6u
X10 a_2011_527# a_448_472# a_1376_115# VPW nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X11 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.381p pd=2.61u as=0.225p ps=1.38u w=0.865u l=0.5u
X12 Q a_2304_115# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=0.5u
X13 a_1376_115# a_1004_159# VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.264p ps=1.82u w=0.36u l=0.6u
X14 VSS a_2304_115# a_2256_159# VPW nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X15 a_836_159# a_36_151# VSS VPW nfet_06v0 ad=43.2f pd=0.6u as=0.158p ps=1.6u w=0.36u l=0.6u
X16 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.178p pd=1.69u as=0.105p ps=0.925u w=0.405u l=0.6u
X17 a_2256_159# a_36_151# a_2011_527# VPW nfet_06v0 ad=43.2f pd=0.6u as=93.6f ps=0.88u w=0.36u l=0.6u
X18 a_880_527# a_448_472# VDD VNW pfet_06v0 ad=54f pd=0.66u as=0.455p ps=3.25u w=0.36u l=0.5u
X19 a_1348_527# a_36_151# a_1004_159# VNW pfet_06v0 ad=43.2f pd=0.6u as=0.187p ps=1.4u w=0.36u l=0.5u
X20 a_1328_159# a_448_472# a_1004_159# VPW nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X21 VDD a_1376_115# a_1348_527# VNW pfet_06v0 ad=0.104p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X22 VDD a_2304_115# a_2296_527# VNW pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X23 a_2304_115# a_2011_527# VDD VNW pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS VNW VPW
X0 a_4604_375# a_4516_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X1 VDD a_572_375# a_484_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X2 VDD a_2364_375# a_2276_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X3 a_4156_375# a_4068_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X4 a_5500_375# a_5412_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X5 a_572_375# a_484_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X6 VDD a_5052_375# a_4964_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X7 VDD a_6844_375# a_6756_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X8 VDD a_1916_375# a_1828_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X9 a_124_375# a_36_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X10 a_5052_375# a_4964_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X11 a_1916_375# a_1828_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X12 VDD a_4604_375# a_4516_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X13 a_1468_375# a_1380_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X14 a_2812_375# a_2724_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X15 VDD a_3260_375# a_3172_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X16 a_2364_375# a_2276_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X17 a_5948_375# a_5860_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X18 VDD a_2812_375# a_2724_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X19 a_3260_375# a_3172_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X20 VDD a_1020_375# a_932_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X21 VDD a_5500_375# a_5412_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X22 a_6844_375# a_6756_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X23 a_6396_375# a_6308_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X24 VDD a_6396_375# a_6308_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X25 VDD a_1468_375# a_1380_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X26 VDD a_4156_375# a_4068_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X27 VDD a_5948_375# a_5860_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X28 VDD a_124_375# a_36_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X29 a_3708_375# a_3620_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
X30 VDD a_3708_375# a_3620_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=1u
X31 a_1020_375# a_932_472# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=1u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 Z I VDD VSS VNW VPW
X0 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 VDD a_224_472# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X3 a_224_472# I VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X4 VDD I a_224_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X6 VDD a_224_472# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X7 VSS a_224_472# Z VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X8 VSS a_224_472# Z VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X9 a_224_472# I VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
X10 VSS I a_224_472# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X11 Z a_224_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 Z I VDD VSS VNW VPW
X0 a_224_472# I VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X1 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X2 a_224_472# I VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X3 VSS a_224_472# Z VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X4 VDD a_224_472# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X5 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X6 a_224_472# I VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X7 Z a_224_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X8 VDD a_224_472# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X9 Z a_224_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X10 Z a_224_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X11 VDD I a_224_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X12 VDD a_224_472# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X13 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X14 VSS a_224_472# Z VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X15 VDD I a_224_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X16 VSS a_224_472# Z VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X17 VDD a_224_472# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X18 VSS a_224_472# Z VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X19 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X20 VSS I a_224_472# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X21 a_224_472# I VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
X22 VSS I a_224_472# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X23 Z a_224_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.211p pd=1.84u as=0.211p ps=1.84u w=0.48u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 B C VDD VSS ZN A1 A2 VNW VPW
X0 a_692_68# B a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X1 ZN A2 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# A2 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.598p ps=3.42u w=1.22u l=0.5u
X3 VDD B ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.402p ps=1.94u w=0.985u l=0.5u
X4 ZN A1 a_244_472# VNW pfet_06v0 ad=0.402p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X5 ZN C VDD VNW pfet_06v0 ad=0.443p pd=2.87u as=0.256p ps=1.5u w=0.985u l=0.5u
X6 VSS C a_692_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X7 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 Z VSS VDD I VNW VPW
X0 Z a_224_552# VSS VPW nfet_06v0 ad=0.112p pd=0.95u as=0.189p ps=1.74u w=0.43u l=0.6u
X1 VSS a_224_552# Z VPW nfet_06v0 ad=0.112p pd=0.95u as=0.112p ps=0.95u w=0.43u l=0.6u
X2 VDD a_224_552# Z VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
X3 a_224_552# I VDD VNW pfet_06v0 ad=0.295p pd=1.54u as=0.361p ps=2.52u w=0.82u l=0.5u
X4 VDD I a_224_552# VNW pfet_06v0 ad=0.213p pd=1.34u as=0.295p ps=1.54u w=0.82u l=0.5u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X6 VDD a_224_552# Z VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
X7 VSS I a_224_552# VPW nfet_06v0 ad=0.105p pd=0.925u as=0.105p ps=0.925u w=0.405u l=0.6u
X8 a_224_552# I VDD VNW pfet_06v0 ad=0.295p pd=1.54u as=0.213p ps=1.34u w=0.82u l=0.5u
X9 VDD a_224_552# Z VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
X10 VSS a_224_552# Z VPW nfet_06v0 ad=0.189p pd=1.74u as=0.112p ps=0.95u w=0.43u l=0.6u
X11 Z a_224_552# VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X12 Z a_224_552# VSS VPW nfet_06v0 ad=0.112p pd=0.95u as=0.112p ps=0.95u w=0.43u l=0.6u
X13 VSS a_224_552# Z VPW nfet_06v0 ad=0.112p pd=0.95u as=0.112p ps=0.95u w=0.43u l=0.6u
X14 Z a_224_552# VSS VPW nfet_06v0 ad=0.112p pd=0.95u as=0.112p ps=0.95u w=0.43u l=0.6u
X15 Z a_224_552# VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X16 VDD I a_224_552# VNW pfet_06v0 ad=0.367p pd=1.92u as=0.295p ps=1.54u w=0.82u l=0.5u
X17 VDD a_224_552# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.439p ps=1.94u w=1.22u l=0.5u
X18 a_224_552# I VSS VPW nfet_06v0 ad=0.105p pd=0.925u as=0.178p ps=1.69u w=0.405u l=0.6u
X19 Z a_224_552# VSS VPW nfet_06v0 ad=0.112p pd=0.95u as=0.112p ps=0.95u w=0.43u l=0.6u
X20 Z a_224_552# VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.367p ps=1.92u w=1.22u l=0.5u
X21 a_224_552# I VSS VPW nfet_06v0 ad=0.178p pd=1.69u as=0.105p ps=0.925u w=0.405u l=0.6u
X22 VSS a_224_552# Z VPW nfet_06v0 ad=0.112p pd=0.95u as=0.112p ps=0.95u w=0.43u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 VDD VSS ZN A1 A2 VNW VPW
X0 a_672_472# A1 ZN VNW pfet_06v0 ad=0.409p pd=1.89u as=0.348p ps=1.79u w=1.22u l=0.5u
X1 ZN A1 VSS VPW nfet_06v0 ad=0.147p pd=1.09u as=0.147p ps=1.09u w=0.565u l=0.6u
X2 ZN A1 a_234_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.378p ps=1.84u w=1.22u l=0.5u
X3 VSS A1 ZN VPW nfet_06v0 ad=0.147p pd=1.09u as=0.147p ps=1.09u w=0.565u l=0.6u
X4 a_234_472# A2 VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
X5 VDD A2 a_672_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.409p ps=1.89u w=1.22u l=0.5u
X6 VSS A2 ZN VPW nfet_06v0 ad=0.249p pd=2.01u as=0.147p ps=1.09u w=0.565u l=0.6u
X7 ZN A2 VSS VPW nfet_06v0 ad=0.147p pd=1.09u as=0.249p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A3 VDD VSS ZN A1 A2 VNW VPW
X0 VDD A1 ZN VNW pfet_06v0 ad=0.433p pd=2.85u as=0.522p ps=2.05u w=0.985u l=0.5u
X1 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.416p ps=1.9u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.305p ps=1.61u w=0.985u l=0.5u
X3 a_36_68# A2 a_672_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.172p ps=1.24u w=0.82u l=0.6u
X4 a_1732_68# A2 a_1528_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.172p ps=1.24u w=0.82u l=0.6u
X5 ZN A3 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.305p ps=1.61u w=0.985u l=0.5u
X6 a_244_68# A2 a_36_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.361p ps=2.52u w=0.82u l=0.6u
X7 a_1528_68# A3 VSS VPW nfet_06v0 ad=0.172p pd=1.24u as=0.213p ps=1.34u w=0.82u l=0.6u
X8 VDD A2 ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X9 ZN A1 a_36_68# VPW nfet_06v0 ad=0.416p pd=1.9u as=0.213p ps=1.34u w=0.82u l=0.6u
X10 VDD A3 ZN VNW pfet_06v0 ad=0.305p pd=1.61u as=0.256p ps=1.5u w=0.985u l=0.5u
X11 VDD A1 ZN VNW pfet_06v0 ad=0.305p pd=1.61u as=0.522p ps=2.05u w=0.985u l=0.5u
X12 a_1100_68# A2 a_36_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.213p ps=1.34u w=0.82u l=0.6u
X13 ZN A1 VDD VNW pfet_06v0 ad=0.522p pd=2.05u as=0.256p ps=1.5u w=0.985u l=0.5u
X14 ZN A3 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.305p ps=1.61u w=0.985u l=0.5u
X15 ZN A1 a_1732_68# VPW nfet_06v0 ad=0.416p pd=1.9u as=0.172p ps=1.24u w=0.82u l=0.6u
X16 VSS A3 a_244_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.172p ps=1.24u w=0.82u l=0.6u
X17 VDD A2 ZN VNW pfet_06v0 ad=0.305p pd=1.61u as=0.256p ps=1.5u w=0.985u l=0.5u
X18 VSS A3 a_1100_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.172p ps=1.24u w=0.82u l=0.6u
X19 a_36_68# A1 ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.416p ps=1.9u w=0.82u l=0.6u
X20 ZN A2 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.433p ps=2.85u w=0.985u l=0.5u
X21 a_672_68# A3 VSS VPW nfet_06v0 ad=0.172p pd=1.24u as=0.213p ps=1.34u w=0.82u l=0.6u
X22 VDD A3 ZN VNW pfet_06v0 ad=0.305p pd=1.61u as=0.256p ps=1.5u w=0.985u l=0.5u
X23 ZN A1 VDD VNW pfet_06v0 ad=0.522p pd=2.05u as=0.305p ps=1.61u w=0.985u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 B1 B2 VDD VSS ZN A1 A2 VNW VPW
X0 ZN B1 a_257_69# VPW nfet_06v0 ad=0.212p pd=1.34u as=0.13p ps=1.13u w=0.815u l=0.6u
X1 VDD B2 a_49_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.535p ps=3.31u w=1.22u l=0.5u
X2 a_49_472# B1 VDD VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X3 ZN A1 a_49_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X4 a_49_472# A2 ZN VNW pfet_06v0 ad=0.535p pd=3.31u as=0.316p ps=1.74u w=1.22u l=0.5u
X5 a_257_69# B2 VSS VPW nfet_06v0 ad=0.13p pd=1.13u as=0.359p ps=2.51u w=0.815u l=0.6u
X6 a_665_69# A1 ZN VPW nfet_06v0 ad=0.13p pd=1.13u as=0.212p ps=1.34u w=0.815u l=0.6u
X7 VSS A2 a_665_69# VPW nfet_06v0 ad=0.359p pd=2.51u as=0.13p ps=1.13u w=0.815u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A3 VDD VSS ZN A1 A2 VNW VPW
X0 VDD A3 a_1130_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.348p ps=1.79u w=1.22u l=0.5u
X1 a_1130_472# A2 a_906_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.378p ps=1.84u w=1.22u l=0.5u
X2 ZN A3 VSS VPW nfet_06v0 ad=0.205p pd=1.81u as=0.121p ps=0.985u w=0.465u l=0.6u
X3 a_244_472# A3 VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
X4 ZN A1 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X5 ZN A2 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X6 VSS A2 ZN VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X7 a_906_472# A1 ZN VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X8 ZN A1 a_468_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.348p ps=1.79u w=1.22u l=0.5u
X9 VSS A1 ZN VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X10 VSS A3 ZN VPW nfet_06v0 ad=0.121p pd=0.985u as=0.205p ps=1.81u w=0.465u l=0.6u
X11 a_468_472# A2 a_244_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.378p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 VDD VSS Z I VNW VPW
X0 VSS I a_224_552# VPW nfet_06v0 ad=94.9f pd=0.885u as=94.9f ps=0.885u w=0.365u l=0.6u
X1 VSS a_224_552# Z VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
X2 a_224_552# I VSS VPW nfet_06v0 ad=0.161p pd=1.61u as=94.9f ps=0.885u w=0.365u l=0.6u
X3 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X4 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X5 VSS I a_224_552# VPW nfet_06v0 ad=94.9f pd=0.885u as=94.9f ps=0.885u w=0.365u l=0.6u
X6 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.361p ps=2.52u w=0.82u l=0.5u
X7 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X8 VSS a_224_552# Z VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
X9 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.408p ps=2.02u w=1.22u l=0.5u
X10 Z a_224_552# VSS VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
X11 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X12 VSS a_224_552# Z VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
X13 a_224_552# I VSS VPW nfet_06v0 ad=94.9f pd=0.885u as=0.161p ps=1.61u w=0.365u l=0.6u
X14 Z a_224_552# VSS VPW nfet_06v0 ad=0.125p pd=1u as=0.211p ps=1.84u w=0.48u l=0.6u
X15 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X16 VDD I a_224_552# VNW pfet_06v0 ad=0.408p pd=2.02u as=0.254p ps=1.44u w=0.82u l=0.5u
X17 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X18 a_224_552# I VSS VPW nfet_06v0 ad=94.9f pd=0.885u as=94.9f ps=0.885u w=0.365u l=0.6u
X19 Z a_224_552# VSS VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
X20 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X21 VSS a_224_552# Z VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
X22 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X23 Z a_224_552# VSS VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
X24 VDD I a_224_552# VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X25 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X26 VDD a_224_552# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X27 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X28 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X29 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X30 Z a_224_552# VSS VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
X31 VSS a_224_552# Z VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
X32 VSS a_224_552# Z VPW nfet_06v0 ad=0.211p pd=1.84u as=0.125p ps=1u w=0.48u l=0.6u
X33 VDD I a_224_552# VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X34 Z a_224_552# VSS VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 B2 C VDD VSS ZN A1 A2 B1 VNW VPW
X0 a_672_472# C a_56_472# VNW pfet_06v0 ad=0.34p pd=1.77u as=0.377p ps=1.83u w=1.22u l=0.5u
X1 VDD B2 a_56_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.535p ps=3.31u w=1.22u l=0.5u
X2 ZN A1 a_940_90# VPW nfet_06v0 ad=0.312p pd=2.3u as=85.2f ps=0.95u w=0.71u l=0.6u
X3 a_56_472# B1 VDD VNW pfet_06v0 ad=0.377p pd=1.83u as=0.316p ps=1.74u w=1.22u l=0.5u
X4 a_672_472# A1 ZN VNW pfet_06v0 ad=0.535p pd=3.31u as=0.377p ps=1.83u w=1.22u l=0.5u
X5 ZN A2 a_672_472# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.34p ps=1.77u w=1.22u l=0.5u
X6 a_244_90# B2 VSS VPW nfet_06v0 ad=85.2f pd=0.95u as=0.312p ps=2.3u w=0.71u l=0.6u
X7 ZN B1 a_244_90# VPW nfet_06v0 ad=0.212p pd=1.41u as=85.2f ps=0.95u w=0.71u l=0.6u
X8 a_940_90# A2 VSS VPW nfet_06v0 ad=85.2f pd=0.95u as=0.226p ps=1.45u w=0.71u l=0.6u
X9 VSS C ZN VPW nfet_06v0 ad=0.226p pd=1.45u as=0.212p ps=1.41u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 VSS Z I VDD VNW VPW
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.494p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VPW nfet_06v0 ad=0.291p pd=1.53u as=0.361p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.291p ps=1.53u w=0.82u l=0.6u
X3 VDD I a_36_68# VNW pfet_06v0 ad=0.494p pd=2.03u as=0.537p ps=3.32u w=1.22u l=0.5u
X4 VSS a_36_68# Z VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X5 VDD a_36_68# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 VDD VSS ZN A1 A2 VNW VPW
X0 a_244_68# A2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
X1 ZN A1 a_244_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.294p pd=1.65u as=0.497p ps=3.14u w=1.13u l=0.5u
X3 VDD A1 ZN VNW pfet_06v0 ad=0.294p pd=1.65u as=0.294p ps=1.65u w=1.13u l=0.5u
X4 a_652_68# A1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X5 VSS A2 a_652_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
X6 ZN A1 VDD VNW pfet_06v0 ad=0.294p pd=1.65u as=0.294p ps=1.65u w=1.13u l=0.5u
X7 VDD A2 ZN VNW pfet_06v0 ad=0.497p pd=3.14u as=0.294p ps=1.65u w=1.13u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 VDD VSS Z A1 A2 VNW VPW
X0 a_255_603# A1 a_67_603# VNW pfet_06v0 ad=0.147p pd=1.09u as=0.249p ps=2.01u w=0.565u l=0.5u
X1 Z a_67_603# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.229p ps=1.58u w=0.82u l=0.6u
X2 VDD A2 a_255_603# VNW pfet_06v0 ad=0.387p pd=2.08u as=0.147p ps=1.09u w=0.565u l=0.5u
X3 VSS A2 a_67_603# VPW nfet_06v0 ad=0.229p pd=1.58u as=93.6f ps=0.88u w=0.36u l=0.6u
X4 Z a_67_603# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.387p ps=2.08u w=1.22u l=0.5u
X5 a_67_603# A1 VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 VSS Z I VDD VNW VPW
X0 VDD I a_36_113# VNW pfet_06v0 ad=0.401p pd=1.92u as=0.462p ps=2.98u w=1.05u l=0.5u
X1 Z a_36_113# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.401p ps=1.92u w=1.22u l=0.5u
X2 Z a_36_113# VSS VPW nfet_06v0 ad=0.218p pd=1.87u as=0.153p ps=1.19u w=0.495u l=0.6u
X3 VSS I a_36_113# VPW nfet_06v0 ad=0.153p pd=1.19u as=0.158p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D VDD VSS CLK Q VNW VPW
X0 VSS a_2304_115# Q VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X1 VSS CLK a_36_151# VPW nfet_06v0 ad=0.105p pd=0.925u as=0.178p ps=1.69u w=0.405u l=0.6u
X2 Q a_2304_115# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X3 a_2304_115# a_2011_527# VSS VPW nfet_06v0 ad=0.176p pd=1.68u as=0.142p ps=1.14u w=0.4u l=0.6u
X4 a_1004_159# D a_836_159# VPW nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X5 a_1004_159# D a_880_527# VNW pfet_06v0 ad=0.187p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X6 a_2011_527# a_36_151# a_1376_115# VNW pfet_06v0 ad=0.166p pd=1.28u as=0.179p ps=1.36u w=0.36u l=0.5u
X7 a_2296_527# a_448_472# a_2011_527# VNW pfet_06v0 ad=50.4f pd=0.64u as=0.166p ps=1.28u w=0.36u l=0.5u
X8 a_1376_115# a_1004_159# VDD VNW pfet_06v0 ad=0.179p pd=1.36u as=0.104p ps=0.94u w=0.36u l=0.5u
X9 VDD CLK a_36_151# VNW pfet_06v0 ad=0.225p pd=1.38u as=0.381p ps=2.61u w=0.865u l=0.5u
X10 VDD a_2304_115# Q VNW pfet_06v0 ad=0.854p pd=3.84u as=0.317p ps=1.74u w=1.22u l=0.5u
X11 VSS a_1376_115# a_1328_159# VPW nfet_06v0 ad=0.264p pd=1.82u as=43.2f ps=0.6u w=0.36u l=0.6u
X12 a_2011_527# a_448_472# a_1376_115# VPW nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X13 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.381p pd=2.61u as=0.225p ps=1.38u w=0.865u l=0.5u
X14 Q a_2304_115# VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.537p ps=3.32u w=1.22u l=0.5u
X15 a_1376_115# a_1004_159# VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.264p ps=1.82u w=0.36u l=0.6u
X16 VSS a_2304_115# a_2256_159# VPW nfet_06v0 ad=0.142p pd=1.14u as=43.2f ps=0.6u w=0.36u l=0.6u
X17 a_836_159# a_36_151# VSS VPW nfet_06v0 ad=43.2f pd=0.6u as=0.158p ps=1.6u w=0.36u l=0.6u
X18 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.178p pd=1.69u as=0.105p ps=0.925u w=0.405u l=0.6u
X19 a_2256_159# a_36_151# a_2011_527# VPW nfet_06v0 ad=43.2f pd=0.6u as=93.6f ps=0.88u w=0.36u l=0.6u
X20 a_880_527# a_448_472# VDD VNW pfet_06v0 ad=54f pd=0.66u as=0.455p ps=3.25u w=0.36u l=0.5u
X21 a_1348_527# a_36_151# a_1004_159# VNW pfet_06v0 ad=43.2f pd=0.6u as=0.187p ps=1.4u w=0.36u l=0.5u
X22 a_1328_159# a_448_472# a_1004_159# VPW nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X23 VDD a_1376_115# a_1348_527# VNW pfet_06v0 ad=0.104p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X24 VDD a_2304_115# a_2296_527# VNW pfet_06v0 ad=0.23p pd=1.54u as=50.4f ps=0.64u w=0.36u l=0.5u
X25 a_2304_115# a_2011_527# VDD VNW pfet_06v0 ad=0.352p pd=2.48u as=0.23p ps=1.54u w=0.8u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 VSS Z I VDD VNW VPW
X0 Z a_36_160# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.234p ps=1.56u w=0.82u l=0.6u
X1 Z a_36_160# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.353p ps=1.96u w=1.22u l=0.5u
X2 VDD I a_36_160# VNW pfet_06v0 ad=0.353p pd=1.96u as=0.249p ps=2.01u w=0.565u l=0.5u
X3 VSS I a_36_160# VPW nfet_06v0 ad=0.234p pd=1.56u as=0.158p ps=1.6u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 VDD VSS I ZN VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.125p pd=1u as=0.211p ps=1.84u w=0.48u l=0.6u
X1 VDD I ZN VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X2 ZN I VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
X3 VSS I ZN VPW nfet_06v0 ad=0.211p pd=1.84u as=0.125p ps=1u w=0.48u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 VSS ZN I VDD VNW VPW
X0 VDD I ZN VNW pfet_06v0 ad=0.537p pd=3.32u as=0.457p ps=1.97u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.225p pd=1.37u as=0.361p ps=2.52u w=0.82u l=0.6u
X2 VSS I ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.225p ps=1.37u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.457p pd=1.97u as=0.537p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 VDD VSS Z I VNW VPW
X0 VSS I a_224_552# VPW nfet_06v0 ad=0.105p pd=0.925u as=0.105p ps=0.925u w=0.405u l=0.6u
X1 VSS a_224_552# Z VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X2 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X3 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X4 Z a_224_552# VSS VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X5 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X6 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X7 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X8 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.361p ps=2.52u w=0.82u l=0.5u
X9 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X10 Z a_224_552# VSS VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X11 VSS a_224_552# Z VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X12 VSS a_224_552# Z VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X13 VDD a_224_552# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X14 Z a_224_552# VSS VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X15 VSS I a_224_552# VPW nfet_06v0 ad=0.105p pd=0.925u as=0.178p ps=1.69u w=0.405u l=0.6u
X16 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X17 a_224_552# I VSS VPW nfet_06v0 ad=0.105p pd=0.925u as=0.105p ps=0.925u w=0.405u l=0.6u
X18 VSS a_224_552# Z VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X19 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X20 VDD I a_224_552# VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X21 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X22 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X23 VSS I a_224_552# VPW nfet_06v0 ad=0.105p pd=0.925u as=0.105p ps=0.925u w=0.405u l=0.6u
X24 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X25 Z a_224_552# VSS VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X26 VSS a_224_552# Z VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X27 VSS a_224_552# Z VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X28 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.254p ps=1.44u w=0.82u l=0.5u
X29 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X30 a_224_552# I VSS VPW nfet_06v0 ad=0.178p pd=1.69u as=0.105p ps=0.925u w=0.405u l=0.6u
X31 Z a_224_552# VSS VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X32 VSS a_224_552# Z VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X33 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X34 VSS a_224_552# Z VPW nfet_06v0 ad=0.213p pd=1.85u as=0.126p ps=1u w=0.485u l=0.6u
X35 VDD I a_224_552# VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X36 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X37 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X38 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X39 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X40 a_224_552# I VSS VPW nfet_06v0 ad=0.105p pd=0.925u as=0.105p ps=0.925u w=0.405u l=0.6u
X41 Z a_224_552# VSS VPW nfet_06v0 ad=0.126p pd=1u as=0.213p ps=1.85u w=0.485u l=0.6u
X42 VDD I a_224_552# VNW pfet_06v0 ad=0.254p pd=1.44u as=0.254p ps=1.44u w=0.82u l=0.5u
X43 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X44 Z a_224_552# VSS VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
X45 Z a_224_552# VSS VPW nfet_06v0 ad=0.126p pd=1u as=0.126p ps=1u w=0.485u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A3 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_455_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.172p ps=1.24u w=0.82u l=0.6u
X1 ZN A3 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.433p ps=2.85u w=0.985u l=0.5u
X2 VDD A2 ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X3 ZN A1 VDD VNW pfet_06v0 ad=0.433p pd=2.85u as=0.256p ps=1.5u w=0.985u l=0.5u
X4 a_271_68# A3 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
X5 a_455_68# A2 a_271_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.131p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 VDD VNW pfet_06v0 ad=0.294p pd=1.65u as=0.294p ps=1.65u w=1.13u l=0.5u
X1 VSS A2 a_661_68# VPW nfet_06v0 ad=0.228p pd=1.38u as=98.4f ps=1.06u w=0.82u l=0.6u
X2 VDD A2 ZN VNW pfet_06v0 ad=0.294p pd=1.65u as=0.294p ps=1.65u w=1.13u l=0.5u
X3 ZN A1 a_260_68# VPW nfet_06v0 ad=0.232p pd=1.38u as=98.4f ps=1.06u w=0.82u l=0.6u
X4 a_1468_68# A1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X5 ZN A2 VDD VNW pfet_06v0 ad=0.294p pd=1.65u as=0.294p ps=1.65u w=1.13u l=0.5u
X6 VDD A1 ZN VNW pfet_06v0 ad=0.294p pd=1.65u as=0.294p ps=1.65u w=1.13u l=0.5u
X7 ZN A1 a_1060_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X8 ZN A1 VDD VNW pfet_06v0 ad=0.294p pd=1.65u as=0.294p ps=1.65u w=1.13u l=0.5u
X9 a_661_68# A1 ZN VPW nfet_06v0 ad=98.4f pd=1.06u as=0.232p ps=1.38u w=0.82u l=0.6u
X10 a_1060_68# A2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.228p ps=1.38u w=0.82u l=0.6u
X11 VDD A2 ZN VNW pfet_06v0 ad=0.497p pd=3.14u as=0.294p ps=1.65u w=1.13u l=0.5u
X12 a_260_68# A2 VSS VPW nfet_06v0 ad=98.4f pd=1.06u as=0.361p ps=2.52u w=0.82u l=0.6u
X13 VSS A2 a_1468_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
X14 ZN A2 VDD VNW pfet_06v0 ad=0.294p pd=1.65u as=0.497p ps=3.14u w=1.13u l=0.5u
X15 VDD A1 ZN VNW pfet_06v0 ad=0.294p pd=1.65u as=0.294p ps=1.65u w=1.13u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 VSS Z I VDD VNW VPW
X0 Z a_36_68# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.494p ps=2.03u w=1.22u l=0.5u
X1 VSS I a_36_68# VPW nfet_06v0 ad=0.291p pd=1.53u as=0.361p ps=2.52u w=0.82u l=0.6u
X2 Z a_36_68# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_68# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X4 Z a_36_68# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.291p ps=1.53u w=0.82u l=0.6u
X5 VDD I a_36_68# VNW pfet_06v0 ad=0.494p pd=2.03u as=0.537p ps=3.32u w=1.22u l=0.5u
X6 VSS a_36_68# Z VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X7 VDD a_36_68# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 B C VDD VSS ZN A1 A2 VNW VPW
X0 VDD A2 a_1612_497# VNW pfet_06v0 ad=0.377p pd=1.81u as=0.46p ps=1.93u w=1.1u l=0.5u
X1 VDD C ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.394p pd=1.81u as=0.285p ps=1.62u w=1.1u l=0.5u
X4 VDD A2 a_716_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.394p ps=1.81u w=1.1u l=0.5u
X5 ZN C VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X6 a_2124_68# B a_36_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.213p ps=1.34u w=0.82u l=0.6u
X7 VDD C ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X8 ZN A2 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.361p ps=2.52u w=0.82u l=0.6u
X9 a_36_68# A2 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.31p ps=1.68u w=0.82u l=0.6u
X10 VSS C a_2960_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X11 VDD B ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X12 ZN C VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X13 a_36_68# A2 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X14 a_1164_497# A2 VDD VNW pfet_06v0 ad=0.394p pd=1.81u as=0.285p ps=1.62u w=1.1u l=0.5u
X15 ZN B VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X16 VDD B ZN VNW pfet_06v0 ad=0.433p pd=2.85u as=0.256p ps=1.5u w=0.985u l=0.5u
X17 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.31p ps=1.68u w=0.82u l=0.6u
X18 a_36_68# B a_3368_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
X19 a_244_497# A2 VDD VNW pfet_06v0 ad=0.46p pd=1.93u as=0.482p ps=3.07u w=1.1u l=0.5u
X20 VSS C a_2124_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.172p ps=1.24u w=0.82u l=0.6u
X21 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X22 ZN A1 a_1164_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.394p ps=1.81u w=1.1u l=0.5u
X23 a_36_68# B a_2552_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X24 a_2552_68# C VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X25 a_1612_497# A1 ZN VNW pfet_06v0 ad=0.46p pd=1.93u as=0.285p ps=1.62u w=1.1u l=0.5u
X26 ZN A1 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u
X27 ZN A2 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X28 a_3368_68# C VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X29 ZN B VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.377p ps=1.81u w=0.985u l=0.5u
X30 a_2960_68# B a_36_68# VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X31 ZN A1 a_244_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.46p ps=1.93u w=1.1u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A2 B C VDD VSS ZN A1 VNW VPW
X0 a_170_472# B a_3662_472# VNW pfet_06v0 ad=0.598p pd=3.42u as=0.317p ps=1.74u w=1.22u l=0.5u
X1 a_1194_69# A2 VSS VPW nfet_06v0 ad=0.123p pd=1.09u as=0.2p ps=1.29u w=0.77u l=0.6u
X2 ZN A1 a_1194_69# VPW nfet_06v0 ad=0.2p pd=1.29u as=0.123p ps=1.09u w=0.77u l=0.6u
X3 VSS C ZN VPW nfet_06v0 ad=0.254p pd=1.61u as=0.12p ps=0.98u w=0.46u l=0.6u
X4 a_170_472# A1 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X5 ZN B VSS VPW nfet_06v0 ad=0.12p pd=0.98u as=0.238p ps=1.51u w=0.46u l=0.6u
X6 a_3126_472# B a_170_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.708p ps=2.38u w=1.22u l=0.5u
X7 ZN A1 a_170_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X8 ZN A1 a_358_69# VPW nfet_06v0 ad=0.2p pd=1.29u as=0.162p ps=1.19u w=0.77u l=0.6u
X9 ZN C VSS VPW nfet_06v0 ad=0.12p pd=0.98u as=0.254p ps=1.61u w=0.46u l=0.6u
X10 VDD C a_3126_472# VNW pfet_06v0 ad=0.708p pd=2.38u as=0.317p ps=1.74u w=1.22u l=0.5u
X11 VSS A2 a_1602_69# VPW nfet_06v0 ad=0.238p pd=1.51u as=0.123p ps=1.09u w=0.77u l=0.6u
X12 VSS B ZN VPW nfet_06v0 ad=0.254p pd=1.61u as=0.12p ps=0.98u w=0.46u l=0.6u
X13 a_1602_69# A1 ZN VPW nfet_06v0 ad=0.123p pd=1.09u as=0.2p ps=1.29u w=0.77u l=0.6u
X14 a_170_472# A2 ZN VNW pfet_06v0 ad=0.451p pd=1.96u as=0.317p ps=1.74u w=1.22u l=0.5u
X15 a_2034_472# B a_170_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.451p ps=1.96u w=1.22u l=0.5u
X16 a_2590_472# C VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.708p ps=2.38u w=1.22u l=0.5u
X17 a_358_69# A2 VSS VPW nfet_06v0 ad=0.162p pd=1.19u as=0.447p ps=2.7u w=0.77u l=0.6u
X18 VSS A2 a_786_69# VPW nfet_06v0 ad=0.2p pd=1.29u as=0.123p ps=1.09u w=0.77u l=0.6u
X19 a_170_472# B a_2590_472# VNW pfet_06v0 ad=0.708p pd=2.38u as=0.317p ps=1.74u w=1.22u l=0.5u
X20 VSS C ZN VPW nfet_06v0 ad=0.264p pd=1.66u as=0.12p ps=0.98u w=0.46u l=0.6u
X21 ZN B VSS VPW nfet_06v0 ad=0.12p pd=0.98u as=0.254p ps=1.61u w=0.46u l=0.6u
X22 ZN A2 a_170_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.537p ps=3.32u w=1.22u l=0.5u
X23 a_170_472# A1 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X24 ZN C VSS VPW nfet_06v0 ad=0.12p pd=0.98u as=0.264p ps=1.66u w=0.46u l=0.6u
X25 VDD C a_2034_472# VNW pfet_06v0 ad=0.708p pd=2.38u as=0.378p ps=1.84u w=1.22u l=0.5u
X26 ZN A1 a_170_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X27 a_170_472# A2 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X28 VSS B ZN VPW nfet_06v0 ad=0.202p pd=1.8u as=0.12p ps=0.98u w=0.46u l=0.6u
X29 a_786_69# A1 ZN VPW nfet_06v0 ad=0.123p pd=1.09u as=0.2p ps=1.29u w=0.77u l=0.6u
X30 a_3662_472# C VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.708p ps=2.38u w=1.22u l=0.5u
X31 ZN A2 a_170_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 VDD VSS Z A1 A2 VNW VPW
X0 VDD A2 a_36_159# VNW pfet_06v0 ad=0.406p pd=2.05u as=0.156p ps=1.12u w=0.6u l=0.5u
X1 Z a_36_159# VDD VNW pfet_06v0 ad=0.535p pd=3.31u as=0.406p ps=2.05u w=1.22u l=0.5u
X2 Z a_36_159# VSS VPW nfet_06v0 ad=0.359p pd=2.51u as=0.234p ps=1.55u w=0.815u l=0.6u
X3 VSS A2 a_244_159# VPW nfet_06v0 ad=0.234p pd=1.55u as=58.4f ps=0.685u w=0.365u l=0.6u
X4 a_244_159# A1 a_36_159# VPW nfet_06v0 ad=58.4f pd=0.685u as=0.161p ps=1.61u w=0.365u l=0.6u
X5 a_36_159# A1 VDD VNW pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 S VDD VSS Z I0 I1 VNW VPW
X0 a_1152_472# S a_124_24# VNW pfet_06v0 ad=0.146p pd=1.46u as=0.317p ps=1.74u w=1.22u l=0.5u
X1 a_692_68# I1 VSS VPW nfet_06v0 ad=98.4f pd=1.06u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 a_124_24# S a_692_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=98.4f ps=1.06u w=0.82u l=0.6u
X3 Z a_124_24# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X4 a_848_380# S VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X5 VDD a_124_24# Z VNW pfet_06v0 ad=0.439p pd=1.94u as=0.348p ps=1.79u w=1.22u l=0.5u
X6 VDD I0 a_1152_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.146p ps=1.46u w=1.22u l=0.5u
X7 a_692_472# I1 VDD VNW pfet_06v0 ad=0.476p pd=2u as=0.439p ps=1.94u w=1.22u l=0.5u
X8 a_848_380# S VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X9 Z a_124_24# VDD VNW pfet_06v0 ad=0.348p pd=1.79u as=0.537p ps=3.32u w=1.22u l=0.5u
X10 VSS I0 a_1084_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.197p ps=1.3u w=0.82u l=0.6u
X11 a_1084_68# a_848_380# a_124_24# VPW nfet_06v0 ad=0.197p pd=1.3u as=0.213p ps=1.34u w=0.82u l=0.6u
X12 VSS a_124_24# Z VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X13 a_124_24# a_848_380# a_692_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.476p ps=2u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 B1 C VDD VSS ZN A1 A2 B2 VNW VPW
X0 a_692_68# C a_36_68# VPW nfet_06v0 ad=0.246p pd=1.42u as=0.213p ps=1.34u w=0.82u l=0.6u
X1 a_932_472# A2 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.386p ps=1.92u w=1.22u l=0.5u
X2 VSS B2 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X3 ZN A2 a_692_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.246p ps=1.42u w=0.82u l=0.6u
X4 a_244_472# B2 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.659p ps=3.52u w=1.22u l=0.5u
X5 ZN A1 a_932_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X6 VDD C ZN VNW pfet_06v0 ad=0.386p pd=1.92u as=0.395p ps=1.94u w=0.945u l=0.5u
X7 ZN B1 a_244_472# VNW pfet_06v0 ad=0.395p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X8 a_36_68# B1 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X9 a_692_68# A1 ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 Z VSS VDD I VNW VPW
X0 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X1 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.361p ps=2.52u w=0.82u l=0.5u
X2 VSS a_224_552# Z VPW nfet_06v0 ad=0.118p pd=0.975u as=0.118p ps=0.975u w=0.455u l=0.6u
X3 VDD a_224_552# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X4 VSS a_224_552# Z VPW nfet_06v0 ad=0.2p pd=1.79u as=0.118p ps=0.975u w=0.455u l=0.6u
X5 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X6 Z a_224_552# VSS VPW nfet_06v0 ad=0.118p pd=0.975u as=0.234p ps=1.94u w=0.455u l=0.6u
X7 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.254p ps=1.44u w=0.82u l=0.5u
X8 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X9 a_224_552# I VSS VPW nfet_06v0 ad=0.514p pd=2.91u as=0.266p ps=2.09u w=0.605u l=0.6u
X10 Z a_224_552# VSS VPW nfet_06v0 ad=0.118p pd=0.975u as=0.118p ps=0.975u w=0.455u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A2 B1 B2 VDD VSS ZN A1 VNW VPW
X0 ZN A1 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X1 VSS B2 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# B2 VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.659p ps=3.52u w=1.22u l=0.5u
X3 a_692_472# A1 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.378p ps=1.84u w=1.22u l=0.5u
X4 VDD A2 a_692_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X5 a_36_68# A2 ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X6 a_36_68# B1 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X7 ZN B1 a_244_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 VSS VDD C2 C1 B2 B1 A2 A1 ZN VNW VPW
X0 a_291_68# C2 VSS VPW nfet_06v0 ad=98.4f pd=1.06u as=0.361p ps=2.52u w=0.82u l=0.6u
X1 a_1235_68# A2 VSS VPW nfet_06v0 ad=0.172p pd=1.24u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 a_619_484# A1 ZN VNW pfet_06v0 ad=0.51p pd=3.2u as=0.36p ps=1.78u w=1.16u l=0.5u
X3 a_255_484# B1 a_619_484# VNW pfet_06v0 ad=0.302p pd=1.68u as=0.51p ps=3.2u w=1.16u l=0.5u
X4 a_619_484# B2 a_255_484# VNW pfet_06v0 ad=0.302p pd=1.68u as=0.302p ps=1.68u w=1.16u l=0.5u
X5 a_255_484# C2 VDD VNW pfet_06v0 ad=0.302p pd=1.68u as=0.51p ps=3.2u w=1.16u l=0.5u
X6 ZN C1 a_291_68# VPW nfet_06v0 ad=0.338p pd=1.64u as=98.4f ps=1.06u w=0.82u l=0.6u
X7 ZN A1 a_1235_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.172p ps=1.24u w=0.82u l=0.6u
X8 VSS B2 a_744_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.301p ps=1.55u w=0.82u l=0.6u
X9 VDD C1 a_255_484# VNW pfet_06v0 ad=0.51p pd=3.2u as=0.302p ps=1.68u w=1.16u l=0.5u
X10 ZN A2 a_619_484# VNW pfet_06v0 ad=0.36p pd=1.78u as=0.302p ps=1.68u w=1.16u l=0.5u
X11 a_744_68# B1 ZN VPW nfet_06v0 ad=0.301p pd=1.55u as=0.338p ps=1.64u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 B C VDD VSS ZN A1 A2 VNW VPW
X0 VSS B ZN VPW nfet_06v0 ad=0.227p pd=1.91u as=0.134p ps=1.03u w=0.515u l=0.6u
X1 VSS C ZN VPW nfet_06v0 ad=0.134p pd=1.03u as=0.134p ps=1.03u w=0.515u l=0.6u
X2 a_244_68# A2 VSS VPW nfet_06v0 ad=93.6f pd=1.02u as=0.343p ps=2.44u w=0.78u l=0.6u
X3 ZN A1 a_244_68# VPW nfet_06v0 ad=0.203p pd=1.3u as=93.6f ps=1.02u w=0.78u l=0.6u
X4 ZN C VSS VPW nfet_06v0 ad=0.134p pd=1.03u as=0.134p ps=1.03u w=0.515u l=0.6u
X5 VDD C a_1044_488# VNW pfet_06v0 ad=0.353p pd=1.76u as=0.353p ps=1.76u w=1.14u l=0.5u
X6 ZN A1 a_36_488# VNW pfet_06v0 ad=0.296p pd=1.66u as=0.308p ps=1.68u w=1.14u l=0.5u
X7 ZN B VSS VPW nfet_06v0 ad=0.134p pd=1.03u as=0.233p ps=1.48u w=0.515u l=0.6u
X8 ZN A2 a_36_488# VNW pfet_06v0 ad=0.296p pd=1.66u as=0.502p ps=3.16u w=1.14u l=0.5u
X9 a_36_488# A2 ZN VNW pfet_06v0 ad=0.296p pd=1.66u as=0.296p ps=1.66u w=1.14u l=0.5u
X10 a_1044_488# B a_36_488# VNW pfet_06v0 ad=0.353p pd=1.76u as=0.296p ps=1.66u w=1.14u l=0.5u
X11 a_36_488# A1 ZN VNW pfet_06v0 ad=0.308p pd=1.68u as=0.296p ps=1.66u w=1.14u l=0.5u
X12 a_36_488# B a_1492_488# VNW pfet_06v0 ad=0.502p pd=3.16u as=0.353p ps=1.76u w=1.14u l=0.5u
X13 a_636_68# A1 ZN VPW nfet_06v0 ad=93.6f pd=1.02u as=0.203p ps=1.3u w=0.78u l=0.6u
X14 a_1492_488# C VDD VNW pfet_06v0 ad=0.353p pd=1.76u as=0.353p ps=1.76u w=1.14u l=0.5u
X15 VSS A2 a_636_68# VPW nfet_06v0 ad=0.233p pd=1.48u as=93.6f ps=1.02u w=0.78u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A3 VDD VSS ZN A1 A2 VNW VPW
X0 a_672_472# A3 VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 a_36_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X2 ZN A1 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X3 VDD A3 a_1120_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X4 ZN A1 a_1792_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X5 VSS A2 ZN VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X6 VSS A3 ZN VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X7 a_1792_472# A2 a_1568_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X8 VSS A1 ZN VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X9 VDD A3 a_224_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X10 VSS A2 ZN VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X11 a_36_472# A1 ZN VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X12 VSS A3 ZN VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X13 a_1120_472# A2 a_36_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X14 ZN A2 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X15 a_36_472# A2 a_672_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X16 a_36_472# A1 ZN VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X17 a_1568_472# A3 VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X18 ZN A3 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X19 VSS A1 ZN VPW nfet_06v0 ad=0.205p pd=1.81u as=0.121p ps=0.985u w=0.465u l=0.6u
X20 ZN A2 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.205p ps=1.81u w=0.465u l=0.6u
X21 a_224_472# A2 a_36_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
X22 ZN A1 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X23 ZN A3 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 VSS ZN I VDD VNW VPW
X0 ZN I VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 ZN I VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X3 ZN I VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.537p ps=3.32u w=1.22u l=0.5u
X4 VSS I ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X5 VDD I ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_224_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.409p ps=1.89u w=1.22u l=0.5u
X1 VSS A1 ZN VPW nfet_06v0 ad=0.249p pd=2.01u as=0.147p ps=1.09u w=0.565u l=0.6u
X2 a_224_472# A2 VDD VNW pfet_06v0 ad=0.409p pd=1.89u as=0.537p ps=3.32u w=1.22u l=0.5u
X3 ZN A2 VSS VPW nfet_06v0 ad=0.147p pd=1.09u as=0.249p ps=2.01u w=0.565u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D Q VDD VSS CLK VNW VPW
X0 VSS CLK a_36_151# VPW nfet_06v0 ad=0.105p pd=0.925u as=0.178p ps=1.69u w=0.405u l=0.6u
X1 VDD a_2011_527# a_2304_115# VNW pfet_06v0 ad=0.386p pd=1.92u as=0.246p ps=1.46u w=0.945u l=0.5u
X2 a_1004_159# D a_836_159# VPW nfet_06v0 ad=0.207p pd=1.51u as=43.2f ps=0.6u w=0.36u l=0.6u
X3 VSS a_2304_115# Q VPW nfet_06v0 ad=0.359p pd=2.51u as=0.212p ps=1.34u w=0.815u l=0.6u
X4 a_2304_115# a_2011_527# VSS VPW nfet_06v0 ad=0.212p pd=1.34u as=0.233p ps=1.55u w=0.815u l=0.6u
X5 a_1004_159# D a_880_527# VNW pfet_06v0 ad=0.187p pd=1.4u as=54f ps=0.66u w=0.36u l=0.5u
X6 a_2011_527# a_36_151# a_1376_115# VNW pfet_06v0 ad=0.166p pd=1.28u as=0.179p ps=1.36u w=0.36u l=0.5u
X7 a_2296_527# a_448_472# a_2011_527# VNW pfet_06v0 ad=50.4f pd=0.64u as=0.166p ps=1.28u w=0.36u l=0.5u
X8 Q a_2304_115# VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.386p ps=1.92u w=1.22u l=0.5u
X9 VSS a_2304_115# Q VPW nfet_06v0 ad=0.212p pd=1.34u as=0.212p ps=1.34u w=0.815u l=0.6u
X10 a_1376_115# a_1004_159# VDD VNW pfet_06v0 ad=0.179p pd=1.36u as=0.104p ps=0.94u w=0.36u l=0.5u
X11 VDD CLK a_36_151# VNW pfet_06v0 ad=0.225p pd=1.38u as=0.381p ps=2.61u w=0.865u l=0.5u
X12 VDD a_2304_115# Q VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
X13 VSS a_1376_115# a_1328_159# VPW nfet_06v0 ad=0.264p pd=1.82u as=43.2f ps=0.6u w=0.36u l=0.6u
X14 a_2011_527# a_448_472# a_1376_115# VPW nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X15 Q a_2304_115# VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X16 a_448_472# a_36_151# VDD VNW pfet_06v0 ad=0.381p pd=2.61u as=0.225p ps=1.38u w=0.865u l=0.5u
X17 Q a_2304_115# VSS VPW nfet_06v0 ad=0.212p pd=1.34u as=0.212p ps=1.34u w=0.815u l=0.6u
X18 a_1376_115# a_1004_159# VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.264p ps=1.82u w=0.36u l=0.6u
X19 VSS a_2304_115# a_2256_159# VPW nfet_06v0 ad=0.233p pd=1.55u as=43.2f ps=0.6u w=0.36u l=0.6u
X20 Q a_2304_115# VSS VPW nfet_06v0 ad=0.212p pd=1.34u as=0.261p ps=1.45u w=0.815u l=0.6u
X21 a_836_159# a_36_151# VSS VPW nfet_06v0 ad=43.2f pd=0.6u as=0.158p ps=1.6u w=0.36u l=0.6u
X22 a_448_472# a_36_151# VSS VPW nfet_06v0 ad=0.178p pd=1.69u as=0.105p ps=0.925u w=0.405u l=0.6u
X23 a_2256_159# a_36_151# a_2011_527# VPW nfet_06v0 ad=43.2f pd=0.6u as=93.6f ps=0.88u w=0.36u l=0.6u
X24 a_880_527# a_448_472# VDD VNW pfet_06v0 ad=54f pd=0.66u as=0.455p ps=3.25u w=0.36u l=0.5u
X25 a_1348_527# a_36_151# a_1004_159# VNW pfet_06v0 ad=43.2f pd=0.6u as=0.187p ps=1.4u w=0.36u l=0.5u
X26 VDD a_2304_115# Q VNW pfet_06v0 ad=0.537p pd=3.32u as=0.439p ps=1.94u w=1.22u l=0.5u
X27 a_1328_159# a_448_472# a_1004_159# VPW nfet_06v0 ad=43.2f pd=0.6u as=0.207p ps=1.51u w=0.36u l=0.6u
X28 VDD a_1376_115# a_1348_527# VNW pfet_06v0 ad=0.104p pd=0.94u as=43.2f ps=0.6u w=0.36u l=0.5u
X29 VSS a_2011_527# a_2304_115# VPW nfet_06v0 ad=0.261p pd=1.45u as=0.212p ps=1.34u w=0.815u l=0.6u
X30 VDD a_2304_115# a_2296_527# VNW pfet_06v0 ad=0.262p pd=1.68u as=50.4f ps=0.64u w=0.36u l=0.5u
X31 a_2304_115# a_2011_527# VDD VNW pfet_06v0 ad=0.246p pd=1.46u as=0.262p ps=1.68u w=0.945u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A3 B1 B2 VDD VSS ZN A1 A2 VNW VPW
X0 a_468_497# A2 a_244_497# VNW pfet_06v0 ad=0.339p pd=1.71u as=0.339p ps=1.71u w=1.1u l=0.5u
X1 VSS A1 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 VSS A3 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X3 VDD B2 a_2060_497# VNW pfet_06v0 ad=0.482p pd=3.07u as=0.46p ps=1.93u w=1.1u l=0.5u
X4 VDD A3 a_1120_497# VNW pfet_06v0 ad=0.394p pd=1.81u as=0.339p ps=1.71u w=1.1u l=0.5u
X5 a_1588_497# B2 VDD VNW pfet_06v0 ad=0.46p pd=1.93u as=0.394p ps=1.81u w=1.1u l=0.5u
X6 ZN B2 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u
X7 a_244_497# A3 VDD VNW pfet_06v0 ad=0.339p pd=1.71u as=0.482p ps=3.07u w=1.1u l=0.5u
X8 a_36_68# B1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.31p ps=1.68u w=0.82u l=0.6u
X9 ZN A1 a_468_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.339p ps=1.71u w=1.1u l=0.5u
X10 a_1120_497# A2 a_896_497# VNW pfet_06v0 ad=0.339p pd=1.71u as=0.339p ps=1.71u w=1.1u l=0.5u
X11 a_36_68# A3 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X12 a_896_497# A1 ZN VNW pfet_06v0 ad=0.339p pd=1.71u as=0.285p ps=1.62u w=1.1u l=0.5u
X13 ZN B1 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u
X14 a_36_68# A1 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X15 a_36_68# B2 ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.31p ps=1.68u w=0.82u l=0.6u
X16 ZN B1 a_1588_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.46p ps=1.93u w=1.1u l=0.5u
X17 a_36_68# A2 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X18 a_2060_497# B1 ZN VNW pfet_06v0 ad=0.46p pd=1.93u as=0.285p ps=1.62u w=1.1u l=0.5u
X19 VSS A2 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 Z VSS VDD I VNW VPW
X0 VDD I a_36_160# VNW pfet_06v0 ad=0.458p pd=2.02u as=0.449p ps=2.92u w=1.02u l=0.5u
X1 VSS I a_36_160# VPW nfet_06v0 ad=0.151p pd=1.18u as=0.158p ps=1.6u w=0.36u l=0.6u
X2 VDD a_36_160# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X3 Z a_36_160# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.458p ps=2.02u w=1.22u l=0.5u
X4 VSS a_36_160# Z VPW nfet_06v0 ad=0.213p pd=1.85u as=0.126p ps=1u w=0.485u l=0.6u
X5 Z a_36_160# VSS VPW nfet_06v0 ad=0.126p pd=1u as=0.151p ps=1.18u w=0.485u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A2 B1 B2 VDD VSS ZN A1 VNW VPW
X0 a_36_497# B1 VDD VNW pfet_06v0 ad=0.285p pd=1.62u as=0.285p ps=1.62u w=1.1u l=0.5u
X1 a_2356_68# A1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 VDD B1 a_36_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.285p ps=1.62u w=1.1u l=0.5u
X3 a_244_68# B2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
X4 ZN B1 a_244_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X5 a_1468_68# B1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X6 a_36_497# B2 VDD VNW pfet_06v0 ad=0.285p pd=1.62u as=0.285p ps=1.62u w=1.1u l=0.5u
X7 ZN A1 a_2764_68# VPW nfet_06v0 ad=0.416p pd=1.9u as=0.131p ps=1.14u w=0.82u l=0.6u
X8 a_2764_68# A2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X9 VDD B2 a_36_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.285p ps=1.62u w=1.1u l=0.5u
X10 ZN A1 a_36_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.526p ps=2.05u w=1.1u l=0.5u
X11 ZN A1 a_1948_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X12 a_652_68# B1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X13 VSS B2 a_652_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X14 VSS A2 a_3260_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
X15 a_36_497# A2 ZN VNW pfet_06v0 ad=0.482p pd=3.07u as=0.285p ps=1.62u w=1.1u l=0.5u
X16 a_3260_68# A1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.416p ps=1.9u w=0.82u l=0.6u
X17 a_36_497# A1 ZN VNW pfet_06v0 ad=0.285p pd=1.62u as=0.285p ps=1.62u w=1.1u l=0.5u
X18 a_36_497# B1 VDD VNW pfet_06v0 ad=0.285p pd=1.62u as=0.285p ps=1.62u w=1.1u l=0.5u
X19 ZN B1 a_1060_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X20 ZN A1 a_36_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.285p ps=1.62u w=1.1u l=0.5u
X21 a_1948_68# A2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=1.7u w=0.82u l=0.6u
X22 VSS A2 a_2356_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X23 a_1060_68# B2 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X24 VDD B1 a_36_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.285p ps=1.62u w=1.1u l=0.5u
X25 ZN A2 a_36_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.482p ps=1.98u w=1.1u l=0.5u
X26 a_36_497# A2 ZN VNW pfet_06v0 ad=0.285p pd=1.62u as=0.285p ps=1.62u w=1.1u l=0.5u
X27 a_36_497# B2 VDD VNW pfet_06v0 ad=0.482p pd=1.98u as=0.285p ps=1.62u w=1.1u l=0.5u
X28 VSS B2 a_1468_68# VPW nfet_06v0 ad=0.361p pd=1.7u as=0.131p ps=1.14u w=0.82u l=0.6u
X29 ZN A2 a_36_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.285p ps=1.62u w=1.1u l=0.5u
X30 a_36_497# A1 ZN VNW pfet_06v0 ad=0.526p pd=2.05u as=0.285p ps=1.62u w=1.1u l=0.5u
X31 VDD B2 a_36_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.482p ps=3.07u w=1.1u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A2 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.406p pd=1.81u as=0.22p ps=1.37u w=0.845u l=0.5u
X2 ZN A3 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.372p ps=2.57u w=0.845u l=0.5u
X3 a_244_68# A3 a_36_68# VPW nfet_06v0 ad=0.131p pd=1.14u as=0.361p ps=2.52u w=0.82u l=0.6u
X4 VSS A4 a_244_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X5 a_1468_68# A4 VSS VPW nfet_06v0 ad=0.152p pd=1.19u as=0.213p ps=1.34u w=0.82u l=0.6u
X6 VDD A4 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X7 a_1866_68# A2 a_1662_68# VPW nfet_06v0 ad=0.152p pd=1.19u as=0.172p ps=1.24u w=0.82u l=0.6u
X8 ZN A4 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X9 ZN A1 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.406p ps=1.81u w=0.845u l=0.5u
X10 a_3276_68# A1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.416p ps=1.9u w=0.82u l=0.6u
X11 a_652_68# A4 VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X12 a_36_68# A3 a_652_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X13 VDD A2 ZN VNW pfet_06v0 ad=0.372p pd=2.57u as=0.22p ps=1.37u w=0.845u l=0.5u
X14 VDD A3 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X15 VSS A4 a_1060_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X16 ZN A3 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X17 a_2372_68# A1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.416p ps=1.9u w=0.82u l=0.6u
X18 a_36_68# A2 a_2372_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
X19 ZN A1 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.406p ps=1.81u w=0.845u l=0.5u
X20 a_1060_68# A3 a_36_68# VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X21 VDD A2 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X22 VDD A4 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X23 ZN A2 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X24 ZN A1 a_2780_68# VPW nfet_06v0 ad=0.416p pd=1.9u as=0.131p ps=1.14u w=0.82u l=0.6u
X25 a_2780_68# A2 a_36_68# VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X26 ZN A4 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X27 VDD A1 ZN VNW pfet_06v0 ad=0.406p pd=1.81u as=0.22p ps=1.37u w=0.845u l=0.5u
X28 a_36_68# A2 a_3276_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
X29 VDD A3 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X30 a_1662_68# A3 a_1468_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.152p ps=1.19u w=0.82u l=0.6u
X31 ZN A1 a_1866_68# VPW nfet_06v0 ad=0.416p pd=1.9u as=0.152p ps=1.19u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 VDD ZN B A1 A2 VSS A3 VNW VPW
X0 a_468_497# A1 ZN VNW pfet_06v0 ad=0.58p pd=2.15u as=0.401p ps=1.85u w=1.1u l=0.5u
X1 a_244_69# A2 ZN VPW nfet_06v0 ad=0.212p pd=1.34u as=0.414p ps=1.9u w=0.815u l=0.6u
X2 a_780_497# A2 a_468_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.58p ps=2.15u w=1.1u l=0.5u
X3 ZN A1 a_244_69# VPW nfet_06v0 ad=0.414p pd=1.9u as=0.212p ps=1.34u w=0.815u l=0.6u
X4 VDD A3 a_780_497# VNW pfet_06v0 ad=0.591p pd=3.27u as=0.285p ps=1.62u w=1.1u l=0.5u
X5 a_244_69# B VSS VPW nfet_06v0 ad=0.212p pd=1.34u as=0.359p ps=2.51u w=0.815u l=0.6u
X6 ZN B VDD VNW pfet_06v0 ad=0.401p pd=1.85u as=0.497p ps=3.14u w=1.13u l=0.5u
X7 ZN A3 a_244_69# VPW nfet_06v0 ad=0.359p pd=2.51u as=0.212p ps=1.34u w=0.815u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 B C VDD VSS ZN A1 A2 VNW VPW
X0 ZN A2 a_37_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.535p ps=3.31u w=1.22u l=0.5u
X1 VSS B ZN VPW nfet_06v0 ad=0.121p pd=0.985u as=0.212p ps=1.41u w=0.465u l=0.6u
X2 a_37_472# A1 ZN VNW pfet_06v0 ad=0.377p pd=1.83u as=0.316p ps=1.74u w=1.22u l=0.5u
X3 VDD C a_653_472# VNW pfet_06v0 ad=0.535p pd=3.31u as=0.377p ps=1.83u w=1.22u l=0.5u
X4 a_245_90# A2 VSS VPW nfet_06v0 ad=85.2f pd=0.95u as=0.312p ps=2.3u w=0.71u l=0.6u
X5 ZN A1 a_245_90# VPW nfet_06v0 ad=0.212p pd=1.41u as=85.2f ps=0.95u w=0.71u l=0.6u
X6 a_653_472# B a_37_472# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.377p ps=1.83u w=1.22u l=0.5u
X7 ZN C VSS VPW nfet_06v0 ad=0.205p pd=1.81u as=0.121p ps=0.985u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A3 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X1 VDD A1 ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X2 a_1044_68# A2 a_860_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.131p ps=1.14u w=0.82u l=0.6u
X3 a_860_68# A1 ZN VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X4 ZN A2 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X5 VDD A3 ZN VNW pfet_06v0 ad=0.433p pd=2.85u as=0.256p ps=1.5u w=0.985u l=0.5u
X6 VSS A3 a_1044_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.172p ps=1.24u w=0.82u l=0.6u
X7 a_276_68# A3 VSS VPW nfet_06v0 ad=0.115p pd=1.1u as=0.361p ps=2.52u w=0.82u l=0.6u
X8 ZN A3 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.433p ps=2.85u w=0.985u l=0.5u
X9 VDD A2 ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X10 a_452_68# A2 a_276_68# VPW nfet_06v0 ad=0.131p pd=1.14u as=0.115p ps=1.1u w=0.82u l=0.6u
X11 ZN A1 a_452_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.131p ps=1.14u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A2 ZN A1 B C VDD VSS VNW VPW
X0 a_1229_68# B a_36_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.215p ps=1.35u w=0.82u l=0.6u
X1 VDD B ZN VNW pfet_06v0 ad=0.433p pd=2.85u as=0.256p ps=1.5u w=0.985u l=0.5u
X2 ZN A1 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u
X3 a_716_497# A1 ZN VNW pfet_06v0 ad=0.46p pd=1.93u as=0.285p ps=1.62u w=1.1u l=0.5u
X4 a_36_68# B a_1657_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
X5 ZN A2 a_36_68# VPW nfet_06v0 ad=0.312p pd=1.68u as=0.361p ps=2.52u w=0.82u l=0.6u
X6 VDD A2 a_716_497# VNW pfet_06v0 ad=0.379p pd=1.82u as=0.46p ps=1.93u w=1.1u l=0.5u
X7 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.312p ps=1.68u w=0.82u l=0.6u
X8 a_244_497# A2 VDD VNW pfet_06v0 ad=0.46p pd=1.93u as=0.482p ps=3.07u w=1.1u l=0.5u
X9 a_36_68# A2 ZN VPW nfet_06v0 ad=0.215p pd=1.35u as=0.31p ps=1.68u w=0.82u l=0.6u
X10 a_1657_68# C VSS VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X11 ZN B VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.379p ps=1.82u w=0.985u l=0.5u
X12 VDD C ZN VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X13 VSS C a_1229_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.172p ps=1.24u w=0.82u l=0.6u
X14 ZN A1 a_244_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.46p ps=1.93u w=1.1u l=0.5u
X15 ZN C VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 B1 B2 VDD VSS ZN A1 A2 VNW VPW
X0 VDD B1 a_36_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X1 VSS A2 a_1468_69# VPW nfet_06v0 ad=0.359p pd=2.51u as=0.13p ps=1.13u w=0.815u l=0.6u
X2 a_36_472# B2 VDD VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X3 ZN A2 a_36_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X4 a_36_472# A1 ZN VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X5 ZN B1 a_244_69# VPW nfet_06v0 ad=0.226p pd=1.37u as=0.13p ps=1.13u w=0.815u l=0.6u
X6 a_659_69# B1 ZN VPW nfet_06v0 ad=0.116p pd=1.1u as=0.226p ps=1.37u w=0.815u l=0.6u
X7 a_244_69# B2 VSS VPW nfet_06v0 ad=0.13p pd=1.13u as=0.359p ps=2.51u w=0.815u l=0.6u
X8 ZN A1 a_36_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X9 a_1468_69# A1 ZN VPW nfet_06v0 ad=0.13p pd=1.13u as=0.212p ps=1.34u w=0.815u l=0.6u
X10 a_36_472# A2 ZN VNW pfet_06v0 ad=0.535p pd=3.31u as=0.316p ps=1.74u w=1.22u l=0.5u
X11 VSS B2 a_659_69# VPW nfet_06v0 ad=0.212p pd=1.34u as=0.116p ps=1.1u w=0.815u l=0.6u
X12 VDD B2 a_36_472# VNW pfet_06v0 ad=0.316p pd=1.74u as=0.535p ps=3.31u w=1.22u l=0.5u
X13 ZN A1 a_1060_69# VPW nfet_06v0 ad=0.212p pd=1.34u as=0.13p ps=1.13u w=0.815u l=0.6u
X14 a_36_472# B1 VDD VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X15 a_1060_69# A2 VSS VPW nfet_06v0 ad=0.13p pd=1.13u as=0.212p ps=1.34u w=0.815u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 B1 VDD VSS ZN A1 A2 B2 VNW VPW
X0 ZN A1 a_2036_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.46p ps=1.93u w=1.1u l=0.5u
X1 ZN B1 a_244_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.339p ps=1.71u w=1.1u l=0.5u
X2 a_672_497# B1 ZN VNW pfet_06v0 ad=0.394p pd=1.81u as=0.285p ps=1.62u w=1.1u l=0.5u
X3 a_2508_497# A1 ZN VNW pfet_06v0 ad=0.394p pd=1.81u as=0.285p ps=1.62u w=1.1u l=0.5u
X4 VSS B1 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X5 VDD A2 a_2508_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.394p ps=1.81u w=1.1u l=0.5u
X6 VSS B2 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X7 ZN A2 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u
X8 ZN A2 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X9 a_2956_497# A2 VDD VNW pfet_06v0 ad=0.394p pd=1.81u as=0.285p ps=1.62u w=1.1u l=0.5u
X10 VSS B1 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X11 ZN A1 a_2956_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.394p ps=1.81u w=1.1u l=0.5u
X12 ZN A1 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X13 VDD B2 a_1568_497# VNW pfet_06v0 ad=0.394p pd=1.81u as=0.339p ps=1.71u w=1.1u l=0.5u
X14 a_244_497# B2 VDD VNW pfet_06v0 ad=0.339p pd=1.71u as=0.482p ps=3.07u w=1.1u l=0.5u
X15 ZN A1 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u
X16 VDD B2 a_672_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.394p ps=1.81u w=1.1u l=0.5u
X17 a_3404_497# A1 ZN VNW pfet_06v0 ad=0.46p pd=1.93u as=0.285p ps=1.62u w=1.1u l=0.5u
X18 a_36_68# B2 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X19 a_36_68# A2 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X20 a_1120_497# B2 VDD VNW pfet_06v0 ad=0.394p pd=1.81u as=0.285p ps=1.62u w=1.1u l=0.5u
X21 a_36_68# B1 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X22 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.31p ps=1.68u w=0.82u l=0.6u
X23 ZN B1 a_1120_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.394p ps=1.81u w=1.1u l=0.5u
X24 VDD A2 a_3404_497# VNW pfet_06v0 ad=0.482p pd=3.07u as=0.46p ps=1.93u w=1.1u l=0.5u
X25 a_2036_497# A2 VDD VNW pfet_06v0 ad=0.46p pd=1.93u as=0.394p ps=1.81u w=1.1u l=0.5u
X26 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X27 a_36_68# B2 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X28 a_1568_497# B1 ZN VNW pfet_06v0 ad=0.339p pd=1.71u as=0.285p ps=1.62u w=1.1u l=0.5u
X29 a_36_68# B1 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X30 a_36_68# A2 ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.31p ps=1.68u w=0.82u l=0.6u
X31 VSS B2 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A3 B1 B2 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_468_472# VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X1 a_244_68# A1 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 a_244_68# A3 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X3 a_916_472# B1 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
X4 VDD B2 a_916_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X5 ZN B1 a_244_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X6 a_224_472# A3 VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.537p ps=3.32u w=1.22u l=0.5u
X7 VSS A2 a_244_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X8 a_244_68# B2 ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X9 a_468_472# A2 a_224_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A3 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A1 a_448_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X1 ZN A1 VSS VPW nfet_06v0 ad=0.205p pd=1.81u as=0.121p ps=0.985u w=0.465u l=0.6u
X2 a_244_472# A3 VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.537p ps=3.32u w=1.22u l=0.5u
X3 a_448_472# A2 a_244_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.317p ps=1.74u w=1.22u l=0.5u
X4 VSS A2 ZN VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X5 ZN A3 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.205p ps=1.81u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A3 VDD VSS Z A1 A2 VNW VPW
X0 a_224_604# A1 a_36_88# VNW pfet_06v0 ad=0.174p pd=1.18u as=0.246p ps=2u w=0.56u l=0.5u
X1 a_36_88# A2 VSS VPW nfet_06v0 ad=0.14p pd=1.1u as=0.104p ps=0.92u w=0.4u l=0.6u
X2 Z a_36_88# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.389p ps=2.02u w=1.22u l=0.5u
X3 VSS A1 a_36_88# VPW nfet_06v0 ad=0.104p pd=0.92u as=0.176p ps=1.68u w=0.4u l=0.6u
X4 a_448_604# A2 a_224_604# VNW pfet_06v0 ad=0.224p pd=1.36u as=0.174p ps=1.18u w=0.56u l=0.5u
X5 VSS A3 a_36_88# VPW nfet_06v0 ad=0.224p pd=1.52u as=0.14p ps=1.1u w=0.4u l=0.6u
X6 VDD A3 a_448_604# VNW pfet_06v0 ad=0.389p pd=2.02u as=0.224p ps=1.36u w=0.56u l=0.5u
X7 Z a_36_88# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.224p ps=1.52u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 Z VSS VDD I VNW VPW
X0 Z a_224_552# VSS VPW nfet_06v0 ad=0.118p pd=0.975u as=0.118p ps=0.975u w=0.455u l=0.6u
X1 VDD a_224_552# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X2 a_224_552# I VDD VNW pfet_06v0 ad=0.254p pd=1.44u as=0.361p ps=2.52u w=0.82u l=0.5u
X3 a_224_552# I VSS VPW nfet_06v0 ad=0.266p pd=2.09u as=0.266p ps=2.09u w=0.605u l=0.6u
X4 VSS a_224_552# Z VPW nfet_06v0 ad=0.118p pd=0.975u as=0.118p ps=0.975u w=0.455u l=0.6u
X5 VDD a_224_552# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X6 VSS a_224_552# Z VPW nfet_06v0 ad=0.2p pd=1.79u as=0.118p ps=0.975u w=0.455u l=0.6u
X7 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.428p ps=2.02u w=1.22u l=0.5u
X8 Z a_224_552# VSS VPW nfet_06v0 ad=0.118p pd=0.975u as=0.2p ps=1.79u w=0.455u l=0.6u
X9 VDD I a_224_552# VNW pfet_06v0 ad=0.428p pd=2.02u as=0.254p ps=1.44u w=0.82u l=0.5u
X10 Z a_224_552# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 VDD VSS Z A1 A2 VNW VPW
X0 a_728_472# a_56_604# VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.4p ps=2.12u w=1.22u l=0.5u
X1 Z A1 a_728_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X2 VSS A1 a_56_604# VPW nfet_06v0 ad=0.218p pd=1.52u as=93.6f ps=0.88u w=0.36u l=0.6u
X3 a_728_472# A2 Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X4 Z a_56_604# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X5 VSS A2 a_952_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
X6 a_244_604# A2 a_56_604# VNW pfet_06v0 ad=0.146p pd=1.08u as=0.246p ps=2u w=0.56u l=0.5u
X7 a_56_604# A2 VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
X8 a_952_68# A1 Z VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X9 VDD A1 a_244_604# VNW pfet_06v0 ad=0.4p pd=2.12u as=0.146p ps=1.08u w=0.56u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A3 VDD VSS Z A1 A2 VNW VPW
X0 Z a_36_148# VDD VNW pfet_06v0 ad=0.535p pd=3.31u as=0.427p ps=2.17u w=1.22u l=0.5u
X1 a_428_148# A2 a_244_148# VPW nfet_06v0 ad=79.8f pd=0.8u as=60.8f ps=0.7u w=0.38u l=0.6u
X2 Z a_36_148# VSS VPW nfet_06v0 ad=0.341p pd=2.43u as=0.242p ps=1.63u w=0.775u l=0.6u
X3 VSS A3 a_428_148# VPW nfet_06v0 ad=0.242p pd=1.63u as=79.8f ps=0.8u w=0.38u l=0.6u
X4 a_244_148# A1 a_36_148# VPW nfet_06v0 ad=60.8f pd=0.7u as=0.167p ps=1.64u w=0.38u l=0.6u
X5 VDD A1 a_36_148# VNW pfet_06v0 ad=0.139p pd=1.05u as=0.235p ps=1.95u w=0.535u l=0.5u
X6 a_36_148# A2 VDD VNW pfet_06v0 ad=0.139p pd=1.05u as=0.139p ps=1.05u w=0.535u l=0.5u
X7 VDD A3 a_36_148# VNW pfet_06v0 ad=0.427p pd=2.17u as=0.139p ps=1.05u w=0.535u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 B VDD VSS A1 ZN A2 VNW VPW
X0 ZN A1 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X1 a_716_497# A1 ZN VNW pfet_06v0 ad=0.394p pd=1.81u as=0.285p ps=1.62u w=1.1u l=0.5u
X2 VDD B ZN VNW pfet_06v0 ad=0.42p pd=2.79u as=0.248p ps=1.48u w=0.955u l=0.5u
X3 VSS B a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X4 VDD A2 a_716_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.394p ps=1.81u w=1.1u l=0.5u
X5 VSS B a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.307p ps=1.68u w=0.82u l=0.6u
X6 ZN A2 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.361p ps=2.52u w=0.82u l=0.6u
X7 a_36_68# A2 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X8 a_1164_497# A2 VDD VNW pfet_06v0 ad=0.394p pd=1.81u as=0.285p ps=1.62u w=1.1u l=0.5u
X9 VDD A2 a_1612_497# VNW pfet_06v0 ad=0.525p pd=2.13u as=0.339p ps=1.71u w=1.1u l=0.5u
X10 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.31p ps=1.68u w=0.82u l=0.6u
X11 a_36_68# A2 ZN VPW nfet_06v0 ad=0.307p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u
X12 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X13 ZN A1 a_1164_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.394p ps=1.81u w=1.1u l=0.5u
X14 a_1612_497# A1 ZN VNW pfet_06v0 ad=0.339p pd=1.71u as=0.285p ps=1.62u w=1.1u l=0.5u
X15 ZN B VDD VNW pfet_06v0 ad=0.248p pd=1.48u as=0.525p ps=2.13u w=0.955u l=0.5u
X16 a_36_68# B VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X17 ZN A1 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X18 a_36_68# B VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X19 VDD B ZN VNW pfet_06v0 ad=0.248p pd=1.48u as=0.248p ps=1.48u w=0.955u l=0.5u
X20 ZN A2 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X21 a_224_497# A2 VDD VNW pfet_06v0 ad=0.515p pd=2.03u as=0.482p ps=3.07u w=1.1u l=0.5u
X22 ZN B VDD VNW pfet_06v0 ad=0.248p pd=1.48u as=0.248p ps=1.48u w=0.955u l=0.5u
X23 ZN A1 a_224_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.515p ps=2.03u w=1.1u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 VSS A3 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X1 a_1213_472# A2 a_943_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.518p ps=2.07u w=1.22u l=0.5u
X2 VSS A2 ZN VPW nfet_06v0 ad=0.158p pd=1.6u as=93.6f ps=0.88u w=0.36u l=0.6u
X3 a_943_472# A3 a_683_472# VNW pfet_06v0 ad=0.518p pd=2.07u as=0.488p ps=2.02u w=1.22u l=0.5u
X4 VSS A1 ZN VPW nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X5 a_1661_472# A1 ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.409p ps=1.89u w=1.22u l=0.5u
X6 VSS A4 ZN VPW nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X7 a_57_472# A2 a_1661_472# VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X8 ZN A1 VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X9 VDD A4 a_245_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.348p ps=1.79u w=1.22u l=0.5u
X10 ZN A2 VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X11 ZN A4 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=93.6f ps=0.88u w=0.36u l=0.6u
X12 a_245_472# A3 a_57_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.537p ps=3.32u w=1.22u l=0.5u
X13 ZN A3 VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
X14 ZN A1 a_1213_472# VNW pfet_06v0 ad=0.409p pd=1.89u as=0.348p ps=1.79u w=1.22u l=0.5u
X15 a_683_472# A4 VDD VNW pfet_06v0 ad=0.488p pd=2.02u as=0.378p ps=1.84u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 B2 VDD VSS ZN A1 A2 B1 VNW VPW
X0 VDD A2 a_1612_497# VNW pfet_06v0 ad=0.482p pd=3.07u as=0.46p ps=1.93u w=1.1u l=0.5u
X1 ZN B1 a_244_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.339p ps=1.71u w=1.1u l=0.5u
X2 a_672_497# B1 ZN VNW pfet_06v0 ad=0.339p pd=1.71u as=0.285p ps=1.62u w=1.1u l=0.5u
X3 a_1140_497# A2 VDD VNW pfet_06v0 ad=0.46p pd=1.93u as=0.394p ps=1.81u w=1.1u l=0.5u
X4 VSS B1 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X5 VSS B2 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X6 a_36_68# A2 ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.31p ps=1.68u w=0.82u l=0.6u
X7 a_244_497# B2 VDD VNW pfet_06v0 ad=0.339p pd=1.71u as=0.482p ps=3.07u w=1.1u l=0.5u
X8 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.31p ps=1.68u w=0.82u l=0.6u
X9 ZN A1 a_1140_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.46p ps=1.93u w=1.1u l=0.5u
X10 VDD B2 a_672_497# VNW pfet_06v0 ad=0.394p pd=1.81u as=0.339p ps=1.71u w=1.1u l=0.5u
X11 a_1612_497# A1 ZN VNW pfet_06v0 ad=0.46p pd=1.93u as=0.285p ps=1.62u w=1.1u l=0.5u
X12 ZN A1 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u
X13 a_36_68# B2 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X14 a_36_68# B1 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X15 ZN A2 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A3 A4 VDD VSS Z A1 A2 VNW VPW
X0 a_48_148# A1 VDD VNW pfet_06v0 ad=0.156p pd=1.12u as=0.264p ps=2.08u w=0.6u l=0.5u
X1 a_440_148# A2 a_256_148# VPW nfet_06v0 ad=88.2f pd=0.84u as=67.2f ps=0.74u w=0.42u l=0.6u
X2 Z a_48_148# VSS VPW nfet_06v0 ad=0.359p pd=2.51u as=0.226p ps=1.51u w=0.815u l=0.6u
X3 VDD A2 a_48_148# VNW pfet_06v0 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X4 Z a_48_148# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.395p ps=2.02u w=1.22u l=0.5u
X5 a_644_148# A3 a_440_148# VPW nfet_06v0 ad=88.2f pd=0.84u as=88.2f ps=0.84u w=0.42u l=0.6u
X6 a_48_148# A3 VDD VNW pfet_06v0 ad=0.156p pd=1.12u as=0.156p ps=1.12u w=0.6u l=0.5u
X7 VSS A4 a_644_148# VPW nfet_06v0 ad=0.226p pd=1.51u as=88.2f ps=0.84u w=0.42u l=0.6u
X8 VDD A4 a_48_148# VNW pfet_06v0 ad=0.395p pd=2.02u as=0.156p ps=1.12u w=0.6u l=0.5u
X9 a_256_148# A1 a_48_148# VPW nfet_06v0 ad=67.2f pd=0.74u as=0.185p ps=1.72u w=0.42u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A2 B VDD VSS ZN A1 VNW VPW
X0 VDD B a_76_476# VNW pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X1 a_680_68# A1 ZN VPW nfet_06v0 ad=98.4f pd=1.06u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 VDD B a_76_476# VNW pfet_06v0 ad=0.312p pd=1.72u as=0.48p ps=2u w=1.2u l=0.5u
X3 a_76_476# B VDD VNW pfet_06v0 ad=0.528p pd=3.28u as=0.312p ps=1.72u w=1.2u l=0.5u
X4 ZN B VSS VPW nfet_06v0 ad=0.133p pd=1.03u as=0.133p ps=1.03u w=0.51u l=0.6u
X5 ZN A2 a_76_476# VNW pfet_06v0 ad=0.312p pd=1.72u as=0.528p ps=3.28u w=1.2u l=0.5u
X6 a_76_476# A1 ZN VNW pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X7 a_1464_68# A1 ZN VPW nfet_06v0 ad=98.4f pd=1.06u as=0.213p ps=1.34u w=0.82u l=0.6u
X8 ZN A1 a_76_476# VNW pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X9 VSS A2 a_1464_68# VPW nfet_06v0 ad=0.241p pd=1.52u as=98.4f ps=1.06u w=0.82u l=0.6u
X10 a_76_476# A2 ZN VNW pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X11 VSS A2 a_680_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=98.4f ps=1.06u w=0.82u l=0.6u
X12 ZN A2 a_76_476# VNW pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X13 VSS B ZN VPW nfet_06v0 ad=0.133p pd=1.03u as=0.133p ps=1.03u w=0.51u l=0.6u
X14 ZN A1 a_1072_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=98.4f ps=1.06u w=0.82u l=0.6u
X15 a_288_68# A2 VSS VPW nfet_06v0 ad=98.4f pd=1.06u as=0.361p ps=2.52u w=0.82u l=0.6u
X16 a_1072_68# A2 VSS VPW nfet_06v0 ad=98.4f pd=1.06u as=0.213p ps=1.34u w=0.82u l=0.6u
X17 VSS B ZN VPW nfet_06v0 ad=0.224p pd=1.9u as=0.133p ps=1.03u w=0.51u l=0.6u
X18 a_76_476# A1 ZN VNW pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X19 ZN A1 a_288_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=98.4f ps=1.06u w=0.82u l=0.6u
X20 ZN A1 a_76_476# VNW pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X21 a_76_476# A2 ZN VNW pfet_06v0 ad=0.48p pd=2u as=0.312p ps=1.72u w=1.2u l=0.5u
X22 a_76_476# B VDD VNW pfet_06v0 ad=0.312p pd=1.72u as=0.312p ps=1.72u w=1.2u l=0.5u
X23 ZN B VSS VPW nfet_06v0 ad=0.133p pd=1.03u as=0.241p ps=1.52u w=0.51u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 a_1458_68# A3 a_1254_68# VPW nfet_06v0 ad=0.152p pd=1.19u as=0.172p ps=1.24u w=0.82u l=0.6u
X1 a_632_68# A2 a_438_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.152p ps=1.19u w=0.82u l=0.6u
X2 VDD A4 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.372p ps=2.57u w=0.845u l=0.5u
X3 a_244_68# A4 VSS VPW nfet_06v0 ad=0.152p pd=1.19u as=0.361p ps=2.52u w=0.82u l=0.6u
X4 ZN A3 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X5 a_438_68# A3 a_244_68# VPW nfet_06v0 ad=0.152p pd=1.19u as=0.152p ps=1.19u w=0.82u l=0.6u
X6 VDD A2 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X7 ZN A1 a_632_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.172p ps=1.24u w=0.82u l=0.6u
X8 ZN A1 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X9 VDD A1 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X10 a_1060_68# A1 ZN VPW nfet_06v0 ad=0.152p pd=1.19u as=0.213p ps=1.34u w=0.82u l=0.6u
X11 a_1254_68# A2 a_1060_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.152p ps=1.19u w=0.82u l=0.6u
X12 ZN A2 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X13 VSS A4 a_1458_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.152p ps=1.19u w=0.82u l=0.6u
X14 VDD A3 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X15 ZN A4 VDD VNW pfet_06v0 ad=0.372p pd=2.57u as=0.22p ps=1.37u w=0.845u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A2 ZN A1 VSS B VDD VNW VPW
X0 ZN A1 a_692_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.46p ps=1.93u w=1.1u l=0.5u
X1 ZN A2 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 VSS B a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X3 a_36_68# A2 ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.312p ps=1.68u w=0.82u l=0.6u
X4 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.31p ps=1.68u w=0.82u l=0.6u
X5 a_1164_497# A1 ZN VNW pfet_06v0 ad=0.46p pd=1.93u as=0.285p ps=1.62u w=1.1u l=0.5u
X6 ZN B VDD VNW pfet_06v0 ad=0.248p pd=1.48u as=0.42p ps=2.79u w=0.955u l=0.5u
X7 a_692_497# A2 VDD VNW pfet_06v0 ad=0.46p pd=1.93u as=0.372p ps=1.81u w=1.1u l=0.5u
X8 VDD B ZN VNW pfet_06v0 ad=0.372p pd=1.81u as=0.248p ps=1.48u w=0.955u l=0.5u
X9 VDD A2 a_1164_497# VNW pfet_06v0 ad=0.482p pd=3.07u as=0.46p ps=1.93u w=1.1u l=0.5u
X10 a_36_68# B VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X11 ZN A1 a_36_68# VPW nfet_06v0 ad=0.312p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 a_66_473# A3 a_692_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X1 VSS A3 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X2 a_2180_473# A2 a_1920_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X3 a_3220_473# A2 a_66_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X4 a_3740_473# A1 ZN VNW pfet_06v0 ad=0.456p pd=1.96u as=0.486p ps=2.02u w=1.22u l=0.5u
X5 a_1212_473# A3 a_66_473# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.486p ps=2.02u w=1.22u l=0.5u
X6 VSS A3 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X7 a_66_473# A2 a_2700_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X8 a_66_473# A2 a_3740_473# VNW pfet_06v0 ad=0.535p pd=3.31u as=0.456p ps=1.96u w=1.22u l=0.5u
X9 ZN A1 a_2180_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X10 ZN A2 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X11 VDD A4 a_254_473# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.346p ps=1.78u w=1.22u l=0.5u
X12 VSS A4 ZN VPW nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X13 ZN A1 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X14 a_1660_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.02u as=0.377p ps=1.83u w=1.22u l=0.5u
X15 a_2700_473# A1 ZN VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X16 VSS A1 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X17 a_254_473# A3 a_66_473# VNW pfet_06v0 ad=0.346p pd=1.78u as=0.535p ps=3.31u w=1.22u l=0.5u
X18 VSS A4 ZN VPW nfet_06v0 ad=93.6f pd=0.88u as=93.6f ps=0.88u w=0.36u l=0.6u
X19 a_1920_473# A3 a_1660_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X20 VSS A2 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X21 ZN A4 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=93.6f ps=0.88u w=0.36u l=0.6u
X22 ZN A3 VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X23 ZN A4 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=93.6f ps=0.88u w=0.36u l=0.6u
X24 ZN A3 VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
X25 VDD A4 a_1212_473# VNW pfet_06v0 ad=0.377p pd=1.83u as=0.377p ps=1.83u w=1.22u l=0.5u
X26 VSS A1 ZN VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X27 a_692_473# A4 VDD VNW pfet_06v0 ad=0.486p pd=2.02u as=0.377p ps=1.83u w=1.22u l=0.5u
X28 ZN A2 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
X29 VSS A2 ZN VPW nfet_06v0 ad=0.158p pd=1.6u as=0.126p ps=1.06u w=0.36u l=0.6u
X30 ZN A1 a_3220_473# VNW pfet_06v0 ad=0.486p pd=2.02u as=0.486p ps=2.02u w=1.22u l=0.5u
X31 ZN A1 VSS VPW nfet_06v0 ad=0.126p pd=1.06u as=0.126p ps=1.06u w=0.36u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A2 A3 B VDD VSS ZN A1 VNW VPW
X0 VDD A3 a_1612_497# VNW pfet_06v0 ad=0.482p pd=3.07u as=0.46p ps=1.93u w=1.1u l=0.5u
X1 a_960_497# A2 a_692_497# VNW pfet_06v0 ad=0.339p pd=1.71u as=0.46p ps=1.93u w=1.1u l=0.5u
X2 ZN A3 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u
X3 VSS B a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X4 a_36_68# A3 ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.31p ps=1.68u w=0.82u l=0.6u
X5 a_36_68# A2 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.31p ps=1.68u w=0.82u l=0.6u
X6 ZN B VDD VNW pfet_06v0 ad=0.281p pd=1.6u as=0.529p ps=3.14u w=1.08u l=0.5u
X7 a_36_68# A1 ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X8 a_692_497# A3 VDD VNW pfet_06v0 ad=0.46p pd=1.93u as=0.392p ps=1.81u w=1.1u l=0.5u
X9 VDD B ZN VNW pfet_06v0 ad=0.392p pd=1.81u as=0.281p ps=1.6u w=1.08u l=0.5u
X10 a_1612_497# A2 a_1388_497# VNW pfet_06v0 ad=0.46p pd=1.93u as=0.339p ps=1.71u w=1.1u l=0.5u
X11 ZN A2 a_36_68# VPW nfet_06v0 ad=0.31p pd=1.68u as=0.213p ps=1.34u w=0.82u l=0.6u
X12 ZN A1 a_960_497# VNW pfet_06v0 ad=0.285p pd=1.62u as=0.339p ps=1.71u w=1.1u l=0.5u
X13 a_36_68# B VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X14 ZN A1 a_36_68# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X15 a_1388_497# A1 ZN VNW pfet_06v0 ad=0.339p pd=1.71u as=0.285p ps=1.62u w=1.1u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 VDD VSS ZN I VNW VPW
X0 ZN I VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X1 VSS I ZN VPW nfet_06v0 ad=0.211p pd=1.84u as=0.125p ps=1u w=0.48u l=0.6u
X2 ZN I VSS VPW nfet_06v0 ad=0.125p pd=1u as=0.211p ps=1.84u w=0.48u l=0.6u
X3 VDD I ZN VNW pfet_06v0 ad=0.537p pd=3.32u as=0.439p ps=1.94u w=1.22u l=0.5u
X4 ZN I VSS VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
X5 ZN I VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.537p ps=3.32u w=1.22u l=0.5u
X6 VDD I ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
X7 VSS I ZN VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 VSS ZN I VDD VNW VPW
X0 ZN I VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=0.6u
X1 ZN I VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or4_4 A3 A4 VDD VSS Z A1 A2 VNW VPW
X0 VSS a_244_72# Z VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X1 Z a_244_72# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.234p ps=1.52u w=0.82u l=0.6u
X2 a_458_472# A3 a_244_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.348p ps=1.79u w=1.22u l=0.5u
X3 VDD a_244_72# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X4 VSS A4 a_244_72# VPW nfet_06v0 ad=0.234p pd=1.52u as=0.121p ps=0.985u w=0.465u l=0.6u
X5 Z a_244_72# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X6 VSS A2 a_244_72# VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X7 VDD A4 a_1578_472# VNW pfet_06v0 ad=0.518p pd=2.07u as=0.378p ps=1.84u w=1.22u l=0.5u
X8 a_244_472# A4 VDD VNW pfet_06v0 ad=0.348p pd=1.79u as=0.537p ps=3.32u w=1.22u l=0.5u
X9 a_244_72# A1 a_682_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.409p ps=1.89u w=1.22u l=0.5u
X10 VSS A1 a_244_72# VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X11 a_1578_472# A3 a_1364_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.348p ps=1.79u w=1.22u l=0.5u
X12 VDD a_244_72# Z VNW pfet_06v0 ad=0.348p pd=1.79u as=0.348p ps=1.79u w=1.22u l=0.5u
X13 VSS A3 a_244_72# VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X14 a_1120_472# A1 a_244_72# VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X15 a_244_72# A1 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X16 a_1364_472# A2 a_1120_472# VNW pfet_06v0 ad=0.348p pd=1.79u as=0.439p ps=1.94u w=1.22u l=0.5u
X17 Z a_244_72# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.348p ps=1.79u w=1.22u l=0.5u
X18 a_682_472# A2 a_458_472# VNW pfet_06v0 ad=0.409p pd=1.89u as=0.378p ps=1.84u w=1.22u l=0.5u
X19 a_244_72# A2 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
X20 a_244_72# A4 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.205p ps=1.81u w=0.465u l=0.6u
X21 Z a_244_72# VDD VNW pfet_06v0 ad=0.348p pd=1.79u as=0.518p ps=2.07u w=1.22u l=0.5u
X22 VSS a_244_72# Z VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X23 a_244_72# A3 VSS VPW nfet_06v0 ad=0.121p pd=0.985u as=0.121p ps=0.985u w=0.465u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 VDD VSS Z A1 A2 VNW VPW
X0 VSS a_730_497# Z VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X1 a_954_497# A1 a_730_497# VNW pfet_06v0 ad=0.526p pd=2.05u as=0.339p ps=1.71u w=1.1u l=0.5u
X2 a_286_93# A2 a_78_93# VPW nfet_06v0 ad=57.6f pd=0.68u as=0.158p ps=1.6u w=0.36u l=0.6u
X3 Z a_730_497# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X4 a_730_497# a_78_93# VDD VNW pfet_06v0 ad=0.339p pd=1.71u as=0.344p ps=1.89u w=1.1u l=0.5u
X5 Z a_730_497# VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.537p ps=3.32u w=1.22u l=0.5u
X6 a_78_93# A2 VDD VNW pfet_06v0 ad=0.146p pd=1.08u as=0.246p ps=2u w=0.56u l=0.5u
X7 a_730_497# A1 a_730_68# VPW nfet_06v0 ad=0.416p pd=1.9u as=0.213p ps=1.34u w=0.82u l=0.6u
X8 VDD A1 a_78_93# VNW pfet_06v0 ad=0.344p pd=1.89u as=0.146p ps=1.08u w=0.56u l=0.5u
X9 VDD a_730_497# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X10 VSS A1 a_286_93# VPW nfet_06v0 ad=0.218p pd=1.52u as=57.6f ps=0.68u w=0.36u l=0.6u
X11 a_730_68# A2 a_730_497# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.416p ps=1.9u w=0.82u l=0.6u
X12 a_730_68# a_78_93# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X13 VDD A2 a_954_497# VNW pfet_06v0 ad=0.482p pd=3.07u as=0.526p ps=2.05u w=1.1u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A3 A4 VDD VSS ZN A1 A2 VNW VPW
X0 ZN A4 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.372p ps=2.57u w=0.845u l=0.5u
X1 VDD A3 ZN VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X2 ZN A2 VDD VNW pfet_06v0 ad=0.22p pd=1.37u as=0.22p ps=1.37u w=0.845u l=0.5u
X3 VDD A1 ZN VNW pfet_06v0 ad=0.372p pd=2.57u as=0.22p ps=1.37u w=0.845u l=0.5u
X4 a_275_68# A4 VSS VPW nfet_06v0 ad=0.152p pd=1.19u as=0.361p ps=2.52u w=0.82u l=0.6u
X5 a_673_68# A2 a_469_68# VPW nfet_06v0 ad=0.152p pd=1.19u as=0.172p ps=1.24u w=0.82u l=0.6u
X6 a_469_68# A3 a_275_68# VPW nfet_06v0 ad=0.172p pd=1.24u as=0.152p ps=1.19u w=0.82u l=0.6u
X7 ZN A1 a_673_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.152p ps=1.19u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A3 VDD VSS Z A1 A2 VNW VPW
X0 a_952_93# A1 a_728_93# VPW nfet_06v0 ad=57.6f pd=0.68u as=93.6f ps=0.88u w=0.36u l=0.6u
X1 a_728_93# A1 a_718_524# VNW pfet_06v0 ad=0.147p pd=1.09u as=0.161p ps=1.13u w=0.565u l=0.5u
X2 a_1524_472# a_728_93# a_1336_472# VNW pfet_06v0 ad=90.4f pd=0.885u as=0.249p ps=2.01u w=0.565u l=0.5u
X3 a_244_524# A2 a_56_524# VNW pfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.5u
X4 a_718_524# a_56_524# VDD VNW pfet_06v0 ad=0.161p pd=1.13u as=0.194p ps=1.41u w=0.565u l=0.5u
X5 a_718_524# A2 a_728_93# VNW pfet_06v0 ad=0.249p pd=2.01u as=0.147p ps=1.09u w=0.565u l=0.5u
X6 VSS A1 a_56_524# VPW nfet_06v0 ad=0.126p pd=1.06u as=93.6f ps=0.88u w=0.36u l=0.6u
X7 a_1336_472# a_728_93# VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
X8 VDD A1 a_244_524# VNW pfet_06v0 ad=0.194p pd=1.41u as=93.6f ps=0.88u w=0.36u l=0.5u
X9 a_56_524# A2 VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.158p ps=1.6u w=0.36u l=0.6u
X10 VSS A3 a_1336_472# VPW nfet_06v0 ad=0.218p pd=1.52u as=93.6f ps=0.88u w=0.36u l=0.6u
X11 a_2215_68# A3 Z VPW nfet_06v0 ad=0.131p pd=1.14u as=0.213p ps=1.34u w=0.82u l=0.6u
X12 VSS a_728_93# a_2215_68# VPW nfet_06v0 ad=0.361p pd=2.52u as=0.131p ps=1.14u w=0.82u l=0.6u
X13 Z a_1336_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X14 Z A3 a_1936_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.317p ps=1.74u w=1.22u l=0.5u
X15 a_728_93# a_56_524# VSS VPW nfet_06v0 ad=93.6f pd=0.88u as=0.126p ps=1.06u w=0.36u l=0.6u
X16 a_1936_472# a_728_93# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.317p ps=1.74u w=1.22u l=0.5u
X17 VSS A2 a_952_93# VPW nfet_06v0 ad=0.158p pd=1.6u as=57.6f ps=0.68u w=0.36u l=0.6u
X18 VDD A3 a_1524_472# VNW pfet_06v0 ad=0.353p pd=1.96u as=90.4f ps=0.885u w=0.565u l=0.5u
X19 a_1936_472# a_1336_472# VDD VNW pfet_06v0 ad=0.317p pd=1.74u as=0.353p ps=1.96u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 Z I VDD VSS VNW VPW
X0 a_224_472# I VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X1 VDD a_224_472# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X2 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X3 a_224_472# I VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X4 VSS a_224_472# Z VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X5 VSS a_224_472# Z VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X6 VDD I a_224_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X7 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X8 a_224_472# I VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X9 Z a_224_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X10 VSS a_224_472# Z VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X11 VSS a_224_472# Z VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X12 VDD a_224_472# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X13 Z a_224_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X14 Z a_224_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X15 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X16 Z a_224_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X17 VDD I a_224_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X18 VDD a_224_472# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X19 VDD a_224_472# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X20 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X21 Z a_224_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X22 a_224_472# I VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X23 VSS a_224_472# Z VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X24 VDD I a_224_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X25 VSS I a_224_472# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X26 VDD a_224_472# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X27 VSS a_224_472# Z VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X28 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X29 VSS I a_224_472# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X30 a_224_472# I VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
X31 VDD a_224_472# Z VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X32 VSS I a_224_472# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X33 Z a_224_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X34 Z a_224_472# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X35 a_224_472# I VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A3 VDD VSS Z A1 A2 VNW VPW
X0 Z a_47_69# VSS VPW nfet_06v0 ad=0.212p pd=1.34u as=0.212p ps=1.34u w=0.815u l=0.6u
X1 VDD A1 a_47_69# VNW pfet_06v0 ad=0.256p pd=1.5u as=0.433p ps=2.85u w=0.985u l=0.5u
X2 Z a_47_69# VDD VNW pfet_06v0 ad=0.316p pd=1.74u as=0.391p ps=1.91u w=1.22u l=0.5u
X3 a_47_69# A2 VDD VNW pfet_06v0 ad=0.256p pd=1.5u as=0.256p ps=1.5u w=0.985u l=0.5u
X4 VDD a_47_69# Z VNW pfet_06v0 ad=0.535p pd=3.31u as=0.316p ps=1.74u w=1.22u l=0.5u
X5 VSS a_47_69# Z VPW nfet_06v0 ad=0.359p pd=2.51u as=0.212p ps=1.34u w=0.815u l=0.6u
X6 VSS A3 a_439_69# VPW nfet_06v0 ad=0.212p pd=1.34u as=0.171p ps=1.24u w=0.815u l=0.6u
X7 VDD A3 a_47_69# VNW pfet_06v0 ad=0.391p pd=1.91u as=0.256p ps=1.5u w=0.985u l=0.5u
X8 a_255_69# A1 a_47_69# VPW nfet_06v0 ad=0.13p pd=1.13u as=0.359p ps=2.51u w=0.815u l=0.6u
X9 a_439_69# A2 a_255_69# VPW nfet_06v0 ad=0.171p pd=1.24u as=0.13p ps=1.13u w=0.815u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 VDD VSS Z A1 A2 VNW VPW
X0 a_247_68# A1 a_39_68# VPW nfet_06v0 ad=0.13p pd=1.13u as=0.359p ps=2.51u w=0.815u l=0.6u
X1 Z a_39_68# VDD VNW pfet_06v0 ad=0.316p pd=1.74u as=0.428p ps=1.96u w=1.22u l=0.5u
X2 Z a_39_68# VSS VPW nfet_06v0 ad=0.22p pd=1.36u as=0.212p ps=1.34u w=0.815u l=0.6u
X3 VDD a_39_68# Z VNW pfet_06v0 ad=0.535p pd=3.31u as=0.316p ps=1.74u w=1.22u l=0.5u
X4 a_39_68# A1 VDD VNW pfet_06v0 ad=0.278p pd=1.59u as=0.471p ps=3.02u w=1.07u l=0.5u
X5 VSS a_39_68# Z VPW nfet_06v0 ad=0.359p pd=2.51u as=0.22p ps=1.36u w=0.815u l=0.6u
X6 VDD A2 a_39_68# VNW pfet_06v0 ad=0.428p pd=1.96u as=0.278p ps=1.59u w=1.07u l=0.5u
X7 VSS A2 a_247_68# VPW nfet_06v0 ad=0.212p pd=1.34u as=0.13p ps=1.13u w=0.815u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 VDD I VSS Z VNW VPW
X0 a_523_68# a_47_68# VSS VPW nfet_06v0 ad=43.2f pd=0.6u as=93.6f ps=0.88u w=0.36u l=0.6u
X1 a_671_644# a_47_68# a_523_68# VPW nfet_06v0 ad=0.369p pd=2.77u as=43.2f ps=0.6u w=0.36u l=0.6u
X2 a_503_644# a_47_68# VDD VNW pfet_06v0 ad=61.2f pd=0.7u as=0.112p ps=0.98u w=0.36u l=0.5u
X3 VDD a_671_644# a_1127_622# VNW pfet_06v0 ad=0.379p pd=2.37u as=61.2f ps=0.7u w=0.36u l=0.5u
X4 VDD I a_47_68# VNW pfet_06v0 ad=0.112p pd=0.98u as=0.385p ps=2.86u w=0.36u l=0.5u
X5 Z a_895_68# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.283p ps=1.87u w=0.82u l=0.6u
X6 a_1147_68# a_671_644# a_895_68# VPW nfet_06v0 ad=43.8f pd=0.605u as=0.37p ps=2.77u w=0.365u l=0.6u
X7 a_1127_622# a_671_644# a_895_68# VNW pfet_06v0 ad=61.2f pd=0.7u as=0.346p ps=2.64u w=0.36u l=0.5u
X8 VSS a_671_644# a_1147_68# VPW nfet_06v0 ad=0.283p pd=1.87u as=43.8f ps=0.605u w=0.365u l=0.6u
X9 a_671_644# a_47_68# a_503_644# VNW pfet_06v0 ad=0.385p pd=2.86u as=61.2f ps=0.7u w=0.36u l=0.5u
X10 VSS I a_47_68# VPW nfet_06v0 ad=93.6f pd=0.88u as=0.333p ps=2.57u w=0.36u l=0.6u
X11 Z a_895_68# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.379p ps=2.37u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 VDD VSS Z A1 A2 VNW VPW
X0 Z a_56_472# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X1 a_56_472# A1 VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X2 a_244_472# A1 a_56_472# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.537p ps=3.32u w=1.22u l=0.5u
X3 VDD A2 a_244_472# VNW pfet_06v0 ad=0.409p pd=1.89u as=0.317p ps=1.74u w=1.22u l=0.5u
X4 VDD a_56_472# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.348p ps=1.79u w=1.22u l=0.5u
X5 Z a_56_472# VDD VNW pfet_06v0 ad=0.348p pd=1.79u as=0.409p ps=1.89u w=1.22u l=0.5u
X6 VSS a_56_472# Z VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X7 VSS A2 a_56_472# VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 VDD ZN I VSS VNW VPW
X0 ZN I VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.125p pd=1u as=0.211p ps=1.84u w=0.48u l=0.6u
X2 VDD I ZN VNW pfet_06v0 ad=0.378p pd=1.84u as=0.378p ps=1.84u w=1.22u l=0.5u
X3 ZN I VSS VPW nfet_06v0 ad=0.211p pd=1.84u as=0.125p ps=1u w=0.48u l=0.6u
X4 ZN I VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.537p ps=3.32u w=1.22u l=0.5u
X5 VSS I ZN VPW nfet_06v0 ad=0.125p pd=1u as=0.125p ps=1u w=0.48u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A3 VDD VSS Z A1 A2 VNW VPW
X0 VDD A3 a_448_472# VNW pfet_06v0 ad=0.488p pd=2.02u as=0.378p ps=1.84u w=1.22u l=0.5u
X1 VSS A3 a_36_68# VPW nfet_06v0 ad=0.264p pd=1.52u as=0.173p ps=1.18u w=0.665u l=0.6u
X2 Z a_36_68# VDD VNW pfet_06v0 ad=0.378p pd=1.84u as=0.488p ps=2.02u w=1.22u l=0.5u
X3 VSS A1 a_36_68# VPW nfet_06v0 ad=0.173p pd=1.18u as=0.293p ps=2.21u w=0.665u l=0.6u
X4 VSS a_36_68# Z VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X5 a_244_472# A1 a_36_68# VNW pfet_06v0 ad=0.317p pd=1.74u as=0.537p ps=3.32u w=1.22u l=0.5u
X6 a_448_472# A2 a_244_472# VNW pfet_06v0 ad=0.378p pd=1.84u as=0.317p ps=1.74u w=1.22u l=0.5u
X7 Z a_36_68# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.264p ps=1.52u w=0.82u l=0.6u
X8 VDD a_36_68# Z VNW pfet_06v0 ad=0.537p pd=3.32u as=0.378p ps=1.84u w=1.22u l=0.5u
X9 a_36_68# A2 VSS VPW nfet_06v0 ad=0.173p pd=1.18u as=0.173p ps=1.18u w=0.665u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A2 VDD VSS Z A1 VNW VPW
X0 Z a_224_490# VSS VPW nfet_06v0 ad=0.201p pd=1.29u as=0.201p ps=1.29u w=0.775u l=0.6u
X1 VSS a_224_490# Z VPW nfet_06v0 ad=0.341p pd=2.43u as=0.201p ps=1.29u w=0.775u l=0.6u
X2 a_224_490# A1 a_244_69# VPW nfet_06v0 ad=0.215p pd=1.33u as=0.124p ps=1.1u w=0.775u l=0.6u
X3 a_659_69# A1 a_224_490# VPW nfet_06v0 ad=0.11p pd=1.06u as=0.215p ps=1.33u w=0.775u l=0.6u
X4 a_244_69# A2 VSS VPW nfet_06v0 ad=0.124p pd=1.1u as=0.341p ps=2.43u w=0.775u l=0.6u
X5 a_224_490# A2 VDD VNW pfet_06v0 ad=0.292p pd=1.64u as=0.495p ps=3.13u w=1.12u l=0.5u
X6 Z a_224_490# VDD VNW pfet_06v0 ad=0.316p pd=1.74u as=0.412p ps=1.91u w=1.22u l=0.5u
X7 VSS a_224_490# Z VPW nfet_06v0 ad=0.201p pd=1.29u as=0.201p ps=1.29u w=0.775u l=0.6u
X8 VDD A1 a_224_490# VNW pfet_06v0 ad=0.292p pd=1.64u as=0.292p ps=1.64u w=1.12u l=0.5u
X9 VDD a_224_490# Z VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X10 VSS A2 a_659_69# VPW nfet_06v0 ad=0.201p pd=1.29u as=0.11p ps=1.06u w=0.775u l=0.6u
X11 a_224_490# A1 VDD VNW pfet_06v0 ad=0.292p pd=1.64u as=0.292p ps=1.64u w=1.12u l=0.5u
X12 Z a_224_490# VDD VNW pfet_06v0 ad=0.316p pd=1.74u as=0.316p ps=1.74u w=1.22u l=0.5u
X13 VDD A2 a_224_490# VNW pfet_06v0 ad=0.412p pd=1.91u as=0.292p ps=1.64u w=1.12u l=0.5u
X14 VDD a_224_490# Z VNW pfet_06v0 ad=0.535p pd=3.31u as=0.316p ps=1.74u w=1.22u l=0.5u
X15 Z a_224_490# VSS VPW nfet_06v0 ad=0.201p pd=1.29u as=0.201p ps=1.29u w=0.775u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 VDD VSS ZN A1 A2 VNW VPW
X0 ZN a_64_93# VDD VNW pfet_06v0 ad=0.312p pd=1.66u as=0.344p ps=1.89u w=1.1u l=0.5u
X1 a_272_93# A2 a_64_93# VPW nfet_06v0 ad=57.6f pd=0.68u as=0.158p ps=1.6u w=0.36u l=0.6u
X2 VSS A1 a_272_93# VPW nfet_06v0 ad=0.218p pd=1.52u as=57.6f ps=0.68u w=0.36u l=0.6u
X3 a_716_68# a_64_93# VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.218p ps=1.52u w=0.82u l=0.6u
X4 VDD A2 a_930_497# VNW pfet_06v0 ad=0.482p pd=3.07u as=0.553p ps=2.11u w=1.1u l=0.5u
X5 ZN A1 a_716_68# VPW nfet_06v0 ad=0.416p pd=1.9u as=0.213p ps=1.34u w=0.82u l=0.6u
X6 a_64_93# A2 VDD VNW pfet_06v0 ad=0.146p pd=1.08u as=0.246p ps=2u w=0.56u l=0.5u
X7 a_716_68# A2 ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.416p ps=1.9u w=0.82u l=0.6u
X8 VDD A1 a_64_93# VNW pfet_06v0 ad=0.344p pd=1.89u as=0.146p ps=1.08u w=0.56u l=0.5u
X9 a_930_497# A1 ZN VNW pfet_06v0 ad=0.553p pd=2.11u as=0.312p ps=1.66u w=1.1u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS VNW VPW
X0 ZN a_124_24# VSS VPW nfet_06v0 ad=0.361p pd=2.52u as=0.361p ps=2.52u w=0.82u l=0.6u
X1 a_124_24# a_124_24# VDD VNW pfet_06v0 ad=0.537p pd=3.32u as=0.537p ps=3.32u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 VSS ZN I VDD VNW VPW
X0 ZN I VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.317p ps=1.74u w=1.22u l=0.5u
X1 ZN I VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X2 ZN I VSS VPW nfet_06v0 ad=0.213p pd=1.34u as=0.361p ps=2.52u w=0.82u l=0.6u
X3 VDD I ZN VNW pfet_06v0 ad=0.537p pd=3.32u as=0.439p ps=1.94u w=1.22u l=0.5u
X4 VSS I ZN VPW nfet_06v0 ad=0.361p pd=2.52u as=0.213p ps=1.34u w=0.82u l=0.6u
X5 ZN I VDD VNW pfet_06v0 ad=0.439p pd=1.94u as=0.537p ps=3.32u w=1.22u l=0.5u
X6 VSS I ZN VPW nfet_06v0 ad=0.213p pd=1.34u as=0.213p ps=1.34u w=0.82u l=0.6u
X7 VDD I ZN VNW pfet_06v0 ad=0.317p pd=1.74u as=0.439p ps=1.94u w=1.22u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 VSS VDD I2 I1 S0 I3 S1 Z VNW VPW
X0 VDD S1 a_1525_369# VNW pfet_06v0 ad=0.175p pd=1.18u as=0.249p ps=2.01u w=0.565u l=0.5u
X1 a_2929_515# S0 a_1901_156# VNW pfet_06v0 ad=0.203p pd=1.28u as=0.147p ps=1.09u w=0.565u l=0.5u
X2 Z a_1081_112# VSS VPW nfet_06v0 ad=0.167p pd=1.64u as=0.131p ps=1.08u w=0.38u l=0.6u
X3 VSS I3 a_712_156# VPW nfet_06v0 ad=0.131p pd=1.08u as=99.4f ps=0.91u w=0.365u l=0.6u
X4 Z a_1081_112# VDD VNW pfet_06v0 ad=0.343p pd=2.44u as=0.241p ps=1.48u w=0.78u l=0.5u
X5 VSS I0 a_2929_515# VPW nfet_06v0 ad=94.9f pd=0.885u as=94.9f ps=0.885u w=0.365u l=0.6u
X6 VDD I3 a_712_156# VNW pfet_06v0 ad=0.241p pd=1.48u as=0.16p ps=1.13u w=0.565u l=0.5u
X7 a_1901_156# S0 a_2521_156# VPW nfet_06v0 ad=94.9f pd=0.885u as=94.9f ps=0.885u w=0.365u l=0.6u
X8 a_468_156# a_348_112# a_224_515# VPW nfet_06v0 ad=0.113p pd=0.985u as=94.9f ps=0.885u w=0.365u l=0.6u
X9 a_468_156# S0 a_224_515# VNW pfet_06v0 ad=0.186p pd=1.23u as=0.243p ps=1.42u w=0.565u l=0.5u
X10 a_224_515# I2 VDD VNW pfet_06v0 ad=0.243p pd=1.42u as=0.249p ps=2.01u w=0.565u l=0.5u
X11 a_1901_156# S1 a_1081_112# VNW pfet_06v0 ad=0.249p pd=2.01u as=0.249p ps=1.44u w=0.565u l=0.5u
X12 a_712_156# S0 a_468_156# VPW nfet_06v0 ad=99.4f pd=0.91u as=0.113p ps=0.985u w=0.365u l=0.6u
X13 a_348_112# S0 VDD VNW pfet_06v0 ad=0.249p pd=2.01u as=0.175p ps=1.18u w=0.565u l=0.5u
X14 a_1081_112# a_1525_369# a_468_156# VNW pfet_06v0 ad=0.249p pd=1.44u as=0.367p ps=2.43u w=0.565u l=0.5u
X15 a_712_156# a_348_112# a_468_156# VNW pfet_06v0 ad=0.16p pd=1.13u as=0.186p ps=1.23u w=0.565u l=0.5u
X16 a_2521_156# I1 VSS VPW nfet_06v0 ad=94.9f pd=0.885u as=94.9f ps=0.885u w=0.365u l=0.6u
X17 a_224_515# I2 VSS VPW nfet_06v0 ad=94.9f pd=0.885u as=0.161p ps=1.61u w=0.365u l=0.6u
X18 a_348_112# S0 VSS VPW nfet_06v0 ad=0.161p pd=1.61u as=94.9f ps=0.885u w=0.365u l=0.6u
X19 a_2521_156# I1 VDD VNW pfet_06v0 ad=0.147p pd=1.09u as=0.175p ps=1.18u w=0.565u l=0.5u
X20 VSS S1 a_1525_369# VPW nfet_06v0 ad=94.9f pd=0.885u as=0.161p ps=1.61u w=0.365u l=0.6u
X21 VDD I0 a_2929_515# VNW pfet_06v0 ad=0.175p pd=1.18u as=0.203p ps=1.28u w=0.565u l=0.5u
X22 a_2929_515# a_348_112# a_1901_156# VPW nfet_06v0 ad=94.9f pd=0.885u as=94.9f ps=0.885u w=0.365u l=0.6u
X23 a_1081_112# S1 a_468_156# VPW nfet_06v0 ad=0.113p pd=0.985u as=0.265p ps=2.18u w=0.365u l=0.6u
X24 a_1901_156# a_348_112# a_2521_156# VNW pfet_06v0 ad=0.147p pd=1.09u as=0.147p ps=1.09u w=0.565u l=0.5u
X25 a_1901_156# a_1525_369# a_1081_112# VPW nfet_06v0 ad=0.161p pd=1.61u as=0.113p ps=0.985u w=0.365u l=0.6u
.ends

.subckt serv_rf_top clk i_dbus_ack i_dbus_rdt[0] i_dbus_rdt[10] i_dbus_rdt[11] i_dbus_rdt[12]
+ i_dbus_rdt[13] i_dbus_rdt[14] i_dbus_rdt[15] i_dbus_rdt[16] i_dbus_rdt[17] i_dbus_rdt[18]
+ i_dbus_rdt[19] i_dbus_rdt[1] i_dbus_rdt[20] i_dbus_rdt[21] i_dbus_rdt[22] i_dbus_rdt[23]
+ i_dbus_rdt[24] i_dbus_rdt[25] i_dbus_rdt[26] i_dbus_rdt[27] i_dbus_rdt[28] i_dbus_rdt[29]
+ i_dbus_rdt[2] i_dbus_rdt[30] i_dbus_rdt[31] i_dbus_rdt[3] i_dbus_rdt[4] i_dbus_rdt[5]
+ i_dbus_rdt[6] i_dbus_rdt[7] i_dbus_rdt[8] i_dbus_rdt[9] i_ext_rd[0] i_ext_rd[10]
+ i_ext_rd[11] i_ext_rd[12] i_ext_rd[13] i_ext_rd[14] i_ext_rd[15] i_ext_rd[16] i_ext_rd[17]
+ i_ext_rd[18] i_ext_rd[19] i_ext_rd[1] i_ext_rd[20] i_ext_rd[21] i_ext_rd[22] i_ext_rd[23]
+ i_ext_rd[24] i_ext_rd[25] i_ext_rd[26] i_ext_rd[27] i_ext_rd[28] i_ext_rd[29] i_ext_rd[2]
+ i_ext_rd[30] i_ext_rd[31] i_ext_rd[3] i_ext_rd[4] i_ext_rd[5] i_ext_rd[6] i_ext_rd[7]
+ i_ext_rd[8] i_ext_rd[9] i_ext_ready i_ibus_ack i_ibus_rdt[0] i_ibus_rdt[10] i_ibus_rdt[11]
+ i_ibus_rdt[12] i_ibus_rdt[13] i_ibus_rdt[14] i_ibus_rdt[15] i_ibus_rdt[16] i_ibus_rdt[17]
+ i_ibus_rdt[18] i_ibus_rdt[19] i_ibus_rdt[1] i_ibus_rdt[20] i_ibus_rdt[21] i_ibus_rdt[22]
+ i_ibus_rdt[23] i_ibus_rdt[24] i_ibus_rdt[25] i_ibus_rdt[26] i_ibus_rdt[27] i_ibus_rdt[28]
+ i_ibus_rdt[29] i_ibus_rdt[2] i_ibus_rdt[30] i_ibus_rdt[31] i_ibus_rdt[3] i_ibus_rdt[4]
+ i_ibus_rdt[5] i_ibus_rdt[6] i_ibus_rdt[7] i_ibus_rdt[8] i_ibus_rdt[9] i_rst i_timer_irq
+ o_dbus_adr[10] o_dbus_adr[11] o_dbus_adr[12] o_dbus_adr[13] o_dbus_adr[14] o_dbus_adr[15]
+ o_dbus_adr[16] o_dbus_adr[17] o_dbus_adr[18] o_dbus_adr[19] o_dbus_adr[1] o_dbus_adr[20]
+ o_dbus_adr[21] o_dbus_adr[22] o_dbus_adr[23] o_dbus_adr[24] o_dbus_adr[25] o_dbus_adr[26]
+ o_dbus_adr[27] o_dbus_adr[28] o_dbus_adr[29] o_dbus_adr[2] o_dbus_adr[30] o_dbus_adr[31]
+ o_dbus_adr[3] o_dbus_adr[4] o_dbus_adr[5] o_dbus_adr[6] o_dbus_adr[7] o_dbus_adr[8]
+ o_dbus_adr[9] o_dbus_cyc o_dbus_dat[0] o_dbus_dat[10] o_dbus_dat[11] o_dbus_dat[12]
+ o_dbus_dat[13] o_dbus_dat[14] o_dbus_dat[15] o_dbus_dat[16] o_dbus_dat[17] o_dbus_dat[18]
+ o_dbus_dat[19] o_dbus_dat[1] o_dbus_dat[20] o_dbus_dat[21] o_dbus_dat[22] o_dbus_dat[23]
+ o_dbus_dat[24] o_dbus_dat[25] o_dbus_dat[26] o_dbus_dat[27] o_dbus_dat[28] o_dbus_dat[29]
+ o_dbus_dat[2] o_dbus_dat[30] o_dbus_dat[31] o_dbus_dat[3] o_dbus_dat[4] o_dbus_dat[5]
+ o_dbus_dat[6] o_dbus_dat[7] o_dbus_dat[8] o_dbus_dat[9] o_dbus_sel[0] o_dbus_sel[1]
+ o_dbus_sel[2] o_dbus_sel[3] o_dbus_we o_ext_funct3[0] o_ext_funct3[1] o_ext_funct3[2]
+ o_ext_rs1[0] o_ext_rs1[10] o_ext_rs1[11] o_ext_rs1[12] o_ext_rs1[13] o_ext_rs1[14]
+ o_ext_rs1[15] o_ext_rs1[16] o_ext_rs1[17] o_ext_rs1[18] o_ext_rs1[19] o_ext_rs1[1]
+ o_ext_rs1[20] o_ext_rs1[21] o_ext_rs1[22] o_ext_rs1[23] o_ext_rs1[24] o_ext_rs1[25]
+ o_ext_rs1[26] o_ext_rs1[27] o_ext_rs1[28] o_ext_rs1[29] o_ext_rs1[2] o_ext_rs1[30]
+ o_ext_rs1[31] o_ext_rs1[3] o_ext_rs1[4] o_ext_rs1[5] o_ext_rs1[6] o_ext_rs1[7] o_ext_rs1[8]
+ o_ext_rs1[9] o_ext_rs2[0] o_ext_rs2[10] o_ext_rs2[11] o_ext_rs2[12] o_ext_rs2[13]
+ o_ext_rs2[14] o_ext_rs2[15] o_ext_rs2[16] o_ext_rs2[17] o_ext_rs2[18] o_ext_rs2[19]
+ o_ext_rs2[1] o_ext_rs2[20] o_ext_rs2[21] o_ext_rs2[22] o_ext_rs2[23] o_ext_rs2[24]
+ o_ext_rs2[25] o_ext_rs2[26] o_ext_rs2[27] o_ext_rs2[28] o_ext_rs2[29] o_ext_rs2[2]
+ o_ext_rs2[30] o_ext_rs2[31] o_ext_rs2[3] o_ext_rs2[4] o_ext_rs2[5] o_ext_rs2[6]
+ o_ext_rs2[7] o_ext_rs2[8] o_ext_rs2[9] o_ibus_adr[0] o_ibus_adr[10] o_ibus_adr[11]
+ o_ibus_adr[12] o_ibus_adr[13] o_ibus_adr[14] o_ibus_adr[15] o_ibus_adr[16] o_ibus_adr[17]
+ o_ibus_adr[18] o_ibus_adr[19] o_ibus_adr[1] o_ibus_adr[20] o_ibus_adr[21] o_ibus_adr[22]
+ o_ibus_adr[23] o_ibus_adr[24] o_ibus_adr[25] o_ibus_adr[26] o_ibus_adr[27] o_ibus_adr[28]
+ o_ibus_adr[29] o_ibus_adr[2] o_ibus_adr[30] o_ibus_adr[31] o_ibus_adr[3] o_ibus_adr[4]
+ o_ibus_adr[5] o_ibus_adr[6] o_ibus_adr[7] o_ibus_adr[8] o_ibus_adr[9] o_ibus_cyc
+ vdd vss o_mdu_valid o_dbus_adr[0]
X_05903_ rf_ram.memory\[82\]\[0\] _02099_ vss vdd rf_ram.memory\[81\]\[0\] _01715_
+ rf_ram.memory\[83\]\[0\] _01654_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__09523__A2 vss net45 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06337__A2 vss _01755_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09671_ vdd vss _04755_ net1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06883_ vdd vss _02983_ _02750_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__05545__B1 vss _01688_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05834_ vdd vss _02030_ rf_ram.memory\[222\]\[0\] _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08622_ vdd _04086_ _04085_ _00729_ _04058_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08553_ vdd vss _04042_ net249 _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05765_ _01959_ rf_ram.memory\[155\]\[0\] vdd vss _01961_ rf_ram.memory\[154\]\[0\]
+ _01958_ _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07504_ vdd vss _03378_ rf_ram.memory\[363\]\[0\] _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08484_ vdd vss _03996_ rf_ram.memory\[379\]\[0\] _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_61 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11633__I vss net83 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06727__I vss _02819_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_330 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07435_ vdd vss _03335_ rf_ram.memory\[332\]\[0\] _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05696_ rf_ram.memory\[391\]\[0\] _01773_ _01777_ rf_ram.memory\[390\]\[0\] _01892_
+ vss vdd rf_ram.memory\[389\]\[0\] _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_9_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_369 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_706 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_246 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09039__A1 vss _04334_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_739 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_205 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_116_931 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07366_ vdd _03291_ _03290_ _00268_ _03289_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09105_ vdd vss _04386_ rf_ram.memory\[95\]\[1\] _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07297_ vdd _03248_ _03247_ _00242_ _03222_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06317_ _01505_ vdd vss _02512_ rf_ram.memory\[182\]\[1\] _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05787__B vss _01923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06248_ _01928_ vdd vss _02443_ _02440_ _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_116_986 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09036_ vdd vss _04344_ rf_ram.memory\[105\]\[0\] _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_962 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09211__A1 vss _04431_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06179_ _02371_ _02372_ _02373_ _01670_ vdd vss _02374_ _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__09762__A2 vss _04766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09938_ vdd _04928_ _04926_ _01204_ _04921_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1133 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07525__A1 vss _02752_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09869_ vdd _04886_ _04885_ _01177_ _04884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06328__A2 vss _01537_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_998 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10713_ vdd rf_ram.memory\[42\]\[1\] clknet_leaf_131_clk vss _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_823 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10644_ vdd rf_ram.memory\[383\]\[0\] clknet_leaf_107_clk vss _00388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10575_ vdd rf_ram.memory\[324\]\[1\] clknet_leaf_169_clk vss _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_953 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06264__A1 vss _01674_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_567 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_792 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09753__A2 vss _04766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06016__A1 vss _01351_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07764__A1 vss _03521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11127_ vdd rf_ram.memory\[117\]\[1\] clknet_leaf_72_clk vss _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_311_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05716__I vss _01626_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06319__A2 vss _01922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11058_ vdd rf_ram.memory\[139\]\[1\] clknet_leaf_10_clk vss _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10009_ vdd vss _04972_ rf_ram.memory\[277\]\[1\] _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_69 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_326_clk_I vss clknet_5_4__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_444 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09269__A1 vss cpu.genblk3.csr.o_new_irq vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05550_ _01746_ _01563_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_89_1224 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05481_ _01677_ _01633_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_1009 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07220_ vdd _03200_ _03198_ _00213_ _03193_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_333 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_709 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07151_ _03157_ _03013_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_27_586 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06102_ _01625_ rf_ram.memory\[275\]\[1\] vdd vss _02297_ rf_ram.memory\[274\]\[1\]
+ _01623_ _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_89_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_854 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_967 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07082_ vdd vss _03114_ _02781_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_718 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06033_ _01505_ vdd vss _02228_ rf_ram.memory\[574\]\[1\] _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11628__I vss net78 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06231__B vss _01504_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07984_ vdd vss _03676_ _03672_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07507__A1 vss _03360_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06935_ vdd _03019_ _03015_ _00109_ _03018_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09723_ vdd vss _04793_ _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09654_ _04738_ _04740_ vdd vss _04741_ net109 _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06866_ _02972_ vss vdd _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07841__I vss _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05817_ rf_ram.memory\[178\]\[0\] _02013_ vss vdd rf_ram.memory\[177\]\[0\] _01931_
+ rf_ram.memory\[179\]\[0\] _01911_ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_08605_ vdd _04075_ _04074_ _00723_ _04058_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06191__B1 vss _01786_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06797_ vdd vss _02925_ rf_ram.memory\[50\]\[0\] _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09585_ vdd vss _04697_ _04651_ _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05748_ rf_ram.memory\[418\]\[0\] _01944_ vss vdd rf_ram.memory\[417\]\[0\] _01645_
+ rf_ram.memory\[419\]\[0\] _01646_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_78_998 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08536_ vdd vss _04031_ _02865_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08483__A2 vss _03496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_190 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05679_ rf_ram.memory\[450\]\[0\] _01875_ vss vdd rf_ram.memory\[449\]\[0\] _01810_
+ rf_ram.memory\[451\]\[0\] _01646_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_147_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_423 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_199 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08467_ _03983_ vdd vss _03984_ _03981_ _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_174_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07418_ vdd vss _03324_ _02866_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08398_ vdd vss _03935_ rf_ram.memory\[17\]\[1\] _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06494__A1 vss _01371_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_531 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_5_31__f_clk_I vss clknet_3_7_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07349_ vdd vss _03281_ rf_ram.memory\[26\]\[0\] _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_219 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_545 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10360_ vdd rf_ram.memory\[298\]\[0\] clknet_leaf_133_clk vss _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_718 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07994__A1 vss _03672_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09019_ vdd vss _04333_ rf_ram.memory\[108\]\[0\] _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10291_ vdd rf_ram.memory\[525\]\[1\] clknet_leaf_318_clk vss _00035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_1217 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07746__A1 vss _03524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_1112 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_628 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_998 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_661 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09671__A1 vss net1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_300 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_979 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06485__A1 vss rf_ram.memory\[4\]\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05288__A2 vss _01341_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10627_ vdd rf_ram.memory\[406\]\[1\] clknet_leaf_114_clk vss _00371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06237__A1 vss _01768_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1075 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08226__A2 vss _03135_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10558_ vdd rf_ram.memory\[330\]\[0\] clknet_leaf_158_clk vss _00302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10033__A2 vss _02815_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06788__A2 vss _02917_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10489_ vdd rf_ram.memory\[193\]\[1\] clknet_leaf_46_clk vss _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_250_clk_I vss clknet_5_20__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06051__B vss _01629_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05748__B1 vss _01646_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_265_clk_I vss clknet_5_17__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05212__A2 vss _01411_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06720_ vdd vss _02868_ _02797_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06651_ vdd vss _02818_ rf_ram.memory\[346\]\[1\] _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08162__A1 vss net237 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_274 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05602_ rf_ram.memory\[309\]\[0\] _01715_ _01709_ rf_ram.memory\[308\]\[0\] _01798_
+ vss vdd rf_ram.memory\[311\]\[0\] _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__06173__B1 vss _01654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06712__A2 vss _02846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06582_ _02763_ vdd vss _02764_ cpu.immdec.imm11_7\[2\] _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_09370_ _04552_ net208 vdd vss _04557_ net207 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05533_ _01728_ vdd vss _01729_ _01349_ _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_129_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08321_ vdd _03886_ _03885_ _00628_ _03884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08465__A2 vss net1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_694 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05464_ vdd vss _01660_ _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_156_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08252_ vdd vss _03844_ rf_ram.memory\[527\]\[0\] _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07203_ vdd _03189_ _03187_ _00207_ _03161_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_203_clk_I vss clknet_5_24__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09414__A1 vss _04463_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08183_ vdd _03801_ _03799_ _00575_ _03790_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05395_ _01590_ _01564_ vdd vss _01591_ _01587_ _01588_ _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_160_859 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_580 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07134_ vdd vss _03147_ rf_ram.memory\[486\]\[1\] _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07065_ vdd vss _03104_ rf_ram.memory\[375\]\[1\] _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_218_clk_I vss clknet_5_22__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05451__A2 vss _01644_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput231 o_ibus_adr[7] net231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput220 o_ibus_adr[26] net220 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06016_ _02210_ _01569_ vdd vss _02211_ _01351_ _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05356__I vss _01551_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07967_ vdd vss _03665_ _02921_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input36_I vss i_ibus_rdt[11] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06918_ vdd _03006_ _03004_ _00105_ _02975_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09706_ vss _04781_ _04739_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__06951__A2 vss _02829_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07898_ vdd vss _03623_ rf_ram.memory\[461\]\[1\] _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08153__A1 vss _03754_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06849_ vdd vss _02961_ _02958_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07900__A1 vss _02839_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09637_ vdd vss _04727_ _04524_ net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09568_ vdd vss _04684_ _03992_ cpu.immdec.imm30_25\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_176_970 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_149 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08519_ vdd vss _04020_ _02838_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11530_ vdd rf_ram.memory\[30\]\[1\] clknet_leaf_205_clk vss _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_765 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09499_ vss _01059_ _04633_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_851 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_547 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05959__C vss rf_ram.i_raddr\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11461_ vdd rf_ram.memory\[292\]\[0\] clknet_leaf_137_clk vss _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10412_ vdd rf_ram.memory\[494\]\[0\] clknet_leaf_182_clk vss _00156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11392_ _01124_ vdd vss clknet_leaf_225_clk net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10343_ vdd rf_ram.memory\[283\]\[1\] clknet_leaf_178_clk vss _00087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_550 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07967__A1 vss _02921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05978__B1 vss _01655_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07719__A1 vss _03491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10274_ vdd rf_ram.memory\[235\]\[0\] clknet_leaf_276_clk vss _00018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_1223 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08392__A1 vss _03919_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06155__B1 vss _01678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_406 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_812 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09644__A1 vss cpu.mem_bytecnt\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10254__A2 vss _03035_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_275 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_415 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_815 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_517 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11659_ vss net182 net110 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_153_185 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10006__A2 vss _03072_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_25_887 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05180_ vdd vss cpu.decode.opcode\[2\] _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__05885__B vss _01928_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06630__A1 vss _02795_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_1_0_clk clknet_3_1_0_clk vss vdd clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_110_767 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08870_ vdd vss _04241_ rf_ram.memory\[130\]\[1\] _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07821_ vdd vss _03575_ _02761_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_84_clk_I vss clknet_5_10__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07752_ vdd vss _03532_ _02781_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08135__A1 vss _03757_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06146__B1 vss _01725_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07683_ vdd vss _03489_ _02908_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09883__A1 vss _04884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06703_ vdd vss _02857_ rf_ram.memory\[522\]\[0\] _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06634_ vdd _02804_ _02802_ _00023_ _02748_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06697__A1 vss _02781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09422_ vss _01029_ _04586_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_99_clk_I vss clknet_5_14__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_609 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09353_ vdd vss _04547_ _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_clkbuf_leaf_142_clk_I vss clknet_5_27__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_61 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06449__A1 vss _01903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06565_ vdd _02749_ _02748_ _00009_ _02739_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08304_ vdd vss _03876_ rf_ram.memory\[221\]\[0\] _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11641__I vss net120 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09635__A1 vss _04524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05516_ _01602_ vdd vss _01712_ rf_ram.memory\[320\]\[0\] _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06496_ vss _02690_ _01376_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_09284_ vdd vss _04505_ _01485_ _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_366 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_22_clk_I vss clknet_5_3__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05447_ _01643_ vss vdd _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_28_681 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08235_ vdd _03833_ _03831_ _00595_ _03823_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05672__A2 vss _01709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05378_ rf_ram.memory\[555\]\[0\] _01521_ _01532_ rf_ram.memory\[554\]\[0\] _01574_
+ vss vdd rf_ram.memory\[553\]\[0\] _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08166_ vdd vss _03791_ rf_ram.memory\[544\]\[1\] _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_157_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07117_ vdd vss _03137_ rf_ram.memory\[500\]\[0\] _03136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_37_clk_I vss clknet_5_7__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08610__A2 vss _04078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08097_ vdd _03747_ _03745_ _00543_ _03724_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07048_ vdd vss _03093_ rf_ram.memory\[391\]\[1\] _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08374__A1 vss net245 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08999_ vdd _04320_ _04319_ _00872_ _04298_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10181__A1 vss _05049_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08126__A1 vss _02829_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06137__B1 vss _01778_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10961_ vdd rf_ram.memory\[69\]\[1\] clknet_leaf_65_clk vss _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08677__A2 vss _03765_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_151_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_710 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10892_ vdd rf_ram.memory\[214\]\[0\] clknet_leaf_303_clk vss _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_423 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09626__A1 vss _04643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_299 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09021__I vss _04061_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06645__I vss _02812_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11513_ vdd rf_ram.memory\[506\]\[0\] clknet_leaf_197_clk vss _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_355 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_483 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09929__A2 vss _03072_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_859 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05663__A2 vss _01856_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11444_ vdd rf_ram.memory\[5\]\[1\] clknet_leaf_293_clk vss _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08860__I vss _04057_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_1113 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11375_ _01107_ vdd vss clknet_leaf_233_clk net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_61_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_857 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05415__A2 vss _01606_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10326_ vdd rf_ram.memory\[290\]\[0\] clknet_leaf_122_clk vss _00070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10257_ vdd vss _05124_ rf_ram.memory\[9\]\[1\] _05122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08365__A1 vss _03884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10188_ vdd _05082_ _05079_ _01300_ _05081_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06376__B1 vss _01793_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08117__A1 vss _03754_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1118 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09865__A1 vss _04840_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_345 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09617__A1 vss _04637_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05351__A1 vss _01495_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_480 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06350_ _02542_ _02543_ _02544_ _01717_ vdd vss _02545_ _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_29_478 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_415 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_150_clk vdd vss clknet_leaf_150_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_142_601 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06281_ _02475_ vdd vss _02476_ _01951_ _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05301_ _01497_ rf_ram.i_raddr\[1\] vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06851__A1 vss _02927_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08840__A2 vss _04195_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08020_ vdd vss _03700_ _02822_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05232_ vdd vss cpu.immdec.imm24_20\[0\] _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_142_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_133 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05163_ vdd vss _01366_ _01364_ _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09971_ vdd _04948_ _04947_ _01217_ _04918_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06603__A1 vss _01496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08922_ vdd vss _04273_ rf_ram.memory\[389\]\[1\] _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07159__A2 vss _02946_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_784 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_1142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08853_ vdd vss _04230_ rf_ram.memory\[132\]\[1\] _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07804_ vdd vss _03565_ rf_ram.memory\[435\]\[1\] _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08784_ vdd _04187_ _04186_ _00790_ _04167_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05996_ _01528_ vdd vss _02191_ rf_ram.memory\[520\]\[1\] _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07735_ vss _03521_ _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__06119__B1 vss _01668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09856__A1 vss cpu.state.genblk1.misalign_trap_sync_r vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_553 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07666_ vdd vss _03478_ _02866_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_827 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09405_ vdd vss _04575_ _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07597_ vdd _03435_ _03433_ _00355_ _03425_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09608__A1 vss net249 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06617_ vdd _02790_ _02789_ _00020_ _02743_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09459__I1 vss net80 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09336_ vdd vss _04538_ rf_ram.memory\[99\]\[1\] _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06548_ _02733_ _01341_ vdd vss _02734_ _01353_ _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_0_146_984 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09267_ vdd vss cpu.genblk3.csr.mcause31 _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_141_clk vdd vss clknet_leaf_141_clk clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_132_111 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05645__A2 vss _01644_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06479_ _01503_ vdd vss _02674_ rf_ram.memory\[14\]\[1\] _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08218_ _03823_ _03689_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_133_656 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09198_ vdd _04444_ _04442_ _00947_ _04434_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09631__I1 vss net58 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08149_ vdd vss _03780_ rf_ram.memory\[547\]\[1\] _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11160_ vdd rf_ram.memory\[100\]\[0\] clknet_leaf_66_clk vss _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08595__A1 vss _04058_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_676 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11091_ vdd rf_ram.memory\[419\]\[0\] clknet_leaf_98_clk vss _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06070__A2 vss _01677_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10111_ vdd vss _05035_ rf_ram.memory\[392\]\[0\] _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_197 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_max_cap236_I vss _02922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10042_ vdd _04992_ _04990_ _01244_ _04985_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output67_I vss net67 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08898__A2 vss _04257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10154__A1 vss _05046_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06358__B1 vss _01959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_818 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_wire239_I vss _02893_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09847__A1 vss _01382_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10944_ vdd rf_ram.memory\[379\]\[0\] clknet_leaf_103_clk vss _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_164 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_168_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10875_ vdd rf_ram.memory\[203\]\[1\] clknet_leaf_35_clk vss _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05869__C1 vss _01702_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_225 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_1184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10209__A2 vss _03547_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05884__A2 vss _01808_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_729 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_770 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07086__A1 vss _03092_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06833__A1 vss _02930_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_132_clk vdd vss clknet_leaf_132_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09686__I vss _04766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_5 vss _01804_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11427_ vdd rf_ram.memory\[249\]\[0\] clknet_leaf_212_clk vss _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05719__I vss _01536_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11358_ vdd rf_ram.memory\[72\]\[0\] clknet_leaf_22_clk vss _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08586__A1 vss _04062_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10309_ vdd rf_ram.memory\[516\]\[1\] clknet_leaf_271_clk vss _00053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08338__A1 vss _03884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11289_ _01024_ vdd vss clknet_leaf_249_clk net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xclkbuf_leaf_199_clk vdd vss clknet_leaf_199_clk clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06349__B1 vss _01811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05850_ _02033_ _02045_ _01362_ vdd vss _02046_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__07561__A2 vss _02917_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05454__I vss _01601_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07520_ vdd _03387_ _03386_ _00326_ _03356_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_64 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05781_ rf_ram.memory\[131\]\[0\] _01608_ _01606_ rf_ram.memory\[130\]\[0\] _01977_
+ vss vdd rf_ram.memory\[129\]\[0\] _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07451_ vdd _03344_ _03343_ _00300_ _03323_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_1165 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07382_ vdd _03301_ _03300_ _00274_ _03289_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06402_ _01707_ vdd vss _02597_ rf_ram.memory\[86\]\[1\] _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_85_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07077__A1 vss _02788_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_370 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06333_ vdd vss _02528_ rf_ram.memory\[217\]\[1\] _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09121_ vdd _04395_ _04393_ _00919_ _04367_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_781 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_123_clk vdd vss clknet_leaf_123_clk clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06824__A1 vss _02927_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06264_ _02447_ _02458_ _01569_ vdd vss _02459_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__05627__A2 vss _01687_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09052_ vdd _04353_ _04352_ _00892_ _04331_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06195_ _02389_ vdd vss _02390_ _01769_ _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08003_ vdd _03688_ _03687_ _00508_ _03686_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05215_ _01414_ vdd vss _01415_ cpu.immdec.imm11_7\[0\] cpu.immdec.imm24_20\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_124_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05146_ _01349_ _01348_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08577__A1 vss _04026_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_473 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xmax_cap241 net241 _02882_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06052__A2 vss _01631_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09954_ vdd vss _04938_ _04911_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08329__A1 vss _03887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08905_ vdd vss _04262_ rf_ram.memory\[126\]\[1\] _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10136__A1 vss _05049_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_80 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09885_ vdd _04895_ _04893_ _01184_ _04887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09264__C vss _02713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08836_ vdd vss _04220_ rf_ram.memory\[469\]\[0\] _04219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07001__A1 vss _03053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_339 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05979_ _01525_ vdd vss _02175_ rf_ram.memory\[10\]\[0\] _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09829__A1 vss _04837_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08767_ vdd vss _04177_ _02945_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07718_ vdd vss _03511_ rf_ram.memory\[380\]\[1\] _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08698_ vdd _04133_ _04131_ _00758_ _04129_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09280__B vss cpu.genblk3.csr.o_new_irq vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1243 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07649_ vdd vss _03468_ rf_ram.memory\[405\]\[1\] _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_726 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output105_I vss net105 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10660_ vdd rf_ram.memory\[37\]\[0\] clknet_leaf_129_clk vss _00404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05866__A2 vss _01989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_578 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_189 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_893 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09319_ cpu.immdec.imm11_7\[4\] _04521_ net35 _04526_ _04528_ vss vdd cpu.immdec.imm11_7\[3\]
+ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_10591_ vdd rf_ram.memory\[320\]\[1\] clknet_leaf_165_clk vss _00335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_114_clk vdd vss clknet_leaf_114_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_152_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05539__I vss _01536_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11212_ vdd rf_ram.memory\[70\]\[0\] clknet_leaf_65_clk vss _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09765__B1 vss _04760_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08568__A1 vss net247 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07240__A1 vss _03193_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11143_ vdd rf_ram.memory\[10\]\[1\] clknet_leaf_35_clk vss _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput75 o_dbus_adr[18] net75 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11074_ vdd rf_ram.memory\[469\]\[1\] clknet_leaf_54_clk vss _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10127__A1 vss _05014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput86 o_dbus_adr[29] net86 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput97 o_dbus_cyc net97 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10025_ vdd _04981_ _04979_ _01238_ _04953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06200__C1 vss _01726_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08740__A1 vss _04157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_648 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05554__A1 vss _01603_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10927_ vdd rf_ram.memory\[174\]\[1\] clknet_leaf_8_clk vss _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06319__B vss _01923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07059__A1 vss _03092_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10858_ vdd rf_ram.memory\[527\]\[0\] clknet_leaf_315_clk vss _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_105_clk vdd vss clknet_leaf_105_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10789_ vdd rf_ram.memory\[562\]\[1\] clknet_leaf_323_clk vss _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_147_1039 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05877__C vss _01569_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_17__f_clk vdd vss clknet_5_17__leaf_clk clknet_3_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_1114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_998 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05449__I vss _01609_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09756__B1 vss _04760_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_8__f_clk_I vss clknet_3_2_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07231__A1 vss _02829_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06034__A2 vss _01538_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06951_ vdd vss _03029_ _02766_ _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05902_ _01602_ vdd vss _02098_ rf_ram.memory\[80\]\[0\] _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09670_ _04753_ _04739_ vdd vss _04754_ net124 _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_158_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06882_ vdd _02982_ _02980_ _00093_ _02975_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_89 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08621_ vdd vss _04086_ rf_ram.memory\[529\]\[0\] _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05833_ _01928_ vdd vss _02029_ _02026_ _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_1099 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08552_ vdd _04041_ _04039_ _00704_ _04026_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_462 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05764_ vdd vss _01960_ rf_ram.memory\[153\]\[0\] _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07503_ vdd vss _03377_ _02781_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08483_ vdd vss _03995_ net244 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_832 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_821 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07434_ vdd vss _03334_ _02788_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05695_ vdd vss _01891_ rf_ram.memory\[388\]\[0\] _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1065 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_126 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_329 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_175_898 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_770 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07365_ vdd vss _03291_ rf_ram.memory\[251\]\[0\] _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09104_ vdd _04385_ _04384_ _00912_ _04364_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07296_ vdd vss _03248_ rf_ram.memory\[25\]\[0\] _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06316_ _02509_ _02510_ vdd vss _02511_ _02507_ _02508_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__08798__A1 vss _02787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06247_ _01719_ _01925_ rf_ram.memory\[443\]\[1\] _02441_ vdd vss _02442_ rf_ram.memory\[442\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_09035_ vdd vss _04343_ net249 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_1247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_557 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06273__A2 vss _01958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input66_I vss i_timer_irq vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05359__I vss _01516_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06178_ rf_ram.memory\[498\]\[1\] _02373_ vss vdd rf_ram.memory\[497\]\[1\] _01668_
+ rf_ram.memory\[499\]\[1\] _01763_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_13_484 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06025__A2 vss _01544_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05129_ vdd vss _01332_ cpu.decode.op21 _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09937_ vdd vss _04928_ rf_ram.memory\[340\]\[1\] _04926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10109__A1 vss _05017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08970__A1 vss _04301_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06430__C1 vss _01696_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05295__S vss _01491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07525__A2 vss _03390_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09868_ vdd vss _04886_ rf_ram.memory\[60\]\[0\] _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09799_ vdd _04843_ _04842_ _01149_ _04837_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08819_ vdd _04209_ _04207_ _00803_ _04205_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_169_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07289__A1 vss _03225_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_692 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10712_ vdd rf_ram.memory\[42\]\[0\] clknet_leaf_134_clk vss _00456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05839__A2 vss _01649_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_331 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10643_ vdd rf_ram.memory\[402\]\[1\] clknet_leaf_96_clk vss _00387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10574_ vdd rf_ram.memory\[324\]\[0\] clknet_leaf_169_clk vss _00318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_965 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1235 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08789__A1 vss _04167_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06653__I vss _02742_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07461__A1 vss _03323_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_524 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07213__A1 vss _03190_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06421__C1 vss _01786_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11126_ vdd rf_ram.memory\[117\]\[0\] clknet_leaf_72_clk vss _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08961__A1 vss _04266_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06321__C vss _01978_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11057_ vdd rf_ram.memory\[139\]\[0\] clknet_leaf_10_clk vss _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08713__A1 vss _04129_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10008_ vdd _04971_ _04970_ _01231_ _04950_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06828__I vss _02945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_478 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05732__I vss _01563_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_326_clk vdd vss clknet_leaf_326_clk clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_819 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_854 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05480_ vdd vss _01676_ rf_ram.memory\[350\]\[0\] _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_638 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07150_ vdd _03156_ _03154_ _00187_ _03126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06563__I vss _02747_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06255__A2 vss _01808_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06101_ vdd vss _02296_ rf_ram.memory\[273\]\[1\] _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07081_ vdd _03113_ _03111_ _00161_ _03092_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_180_890 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06032_ _02225_ _02226_ vdd vss _02227_ _02223_ _02224_ _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_26_1275 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06007__A2 vss _01511_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1128 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07983_ vdd _03675_ _03673_ _00501_ _03654_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09722_ _04791_ _04792_ vdd vss _04793_ net105 _04790_ net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06934_ vdd vss _03019_ rf_ram.memory\[297\]\[1\] _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08704__A1 vss _02991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09653_ vss _04740_ _04739_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06865_ vdd vss _02971_ _02773_ _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_145_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05816_ _01923_ vdd vss _02012_ rf_ram.memory\[176\]\[0\] _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_1095 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09584_ vdd vss _04696_ _04477_ cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08604_ vdd vss _04075_ rf_ram.memory\[164\]\[0\] _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_467 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_618 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08535_ vdd _04030_ _04028_ _00698_ _04026_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06796_ vdd vss _02924_ _02921_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05747_ _01756_ vdd vss _01943_ rf_ram.memory\[416\]\[0\] _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_317_clk vdd vss clknet_leaf_317_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05678_ _01756_ vdd vss _01874_ rf_ram.memory\[448\]\[0\] _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08466_ _02709_ vdd vss _03983_ cpu.state.init_done _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07691__A1 vss _03488_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07417_ _03323_ _03013_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08397_ vdd _03934_ _03933_ _00656_ _03919_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_107_228 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07348_ vdd vss _03280_ _02813_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06246__A2 vss _01918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06406__C vss _01670_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07279_ vdd _03237_ _03235_ _00235_ _03225_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_143_570 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07443__A1 vss _03326_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_412 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_765 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output172_I vss net172 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07994__A2 vss _02923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09018_ vdd vss _04332_ _02787_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10290_ vdd rf_ram.memory\[525\]\[0\] clknet_leaf_314_clk vss _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09196__A1 vss _04431_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08943__A1 vss _04269_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06403__C1 vss _01763_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1217 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_308_clk vdd vss clknet_leaf_308_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_84_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06485__A2 vss _01643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10626_ vdd rf_ram.memory\[406\]\[0\] clknet_leaf_114_clk vss _00370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05693__B1 vss _01786_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_740 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_362 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06316__C vss _01860_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07434__A1 vss _02788_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10557_ vdd rf_ram.memory\[368\]\[1\] clknet_leaf_148_clk vss _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10488_ vdd rf_ram.memory\[193\]\[0\] clknet_leaf_45_clk vss _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08934__A1 vss _02953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05727__I vss _01550_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06332__B vss _01551_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11109_ vdd rf_ram.memory\[124\]\[1\] clknet_leaf_85_clk vss _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_75_58 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06650_ vdd _02817_ _02816_ _00026_ _02743_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08162__A2 vss _03765_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05601_ _01707_ vdd vss _01797_ rf_ram.memory\[310\]\[0\] _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05462__I vss _01563_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_229 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_1208 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05920__A1 vss _01909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09111__A1 vss _04367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05381__C1 vss _01540_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06581_ vdd vss _02763_ _02732_ _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05532_ _01723_ _01727_ vdd vss _01728_ _01720_ _01722_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_129_331 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08320_ vdd vss _03886_ rf_ram.memory\[242\]\[0\] _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05463_ _01658_ vdd vss _01659_ _01651_ _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_145_824 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06476__A2 vss _01633_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08251_ vdd vss _03843_ _02845_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07202_ vdd vss _03189_ rf_ram.memory\[273\]\[1\] _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08182_ vdd vss _03801_ rf_ram.memory\[541\]\[1\] _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05394_ rf_ram.memory\[571\]\[0\] _01540_ _01544_ rf_ram.memory\[570\]\[0\] _01590_
+ vss vdd rf_ram.memory\[569\]\[0\] _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__06228__A2 vss _01755_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1229 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07133_ vdd _03146_ _03145_ _00180_ _03123_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07064_ vdd _03103_ _03102_ _00154_ _03087_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_765 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05987__A1 vss _01348_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput210 o_ibus_adr[17] net210 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_30_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09178__A1 vss _03134_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11639__I vss net98 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput232 o_ibus_adr[8] net232 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput221 o_ibus_adr[27] net221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06015_ vdd _01351_ _02209_ _02210_ _02204_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_57_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_763 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07966_ vdd _03664_ _03662_ _00495_ _03654_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06400__A2 vss _01801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06917_ vdd vss _03006_ rf_ram.memory\[298\]\[1\] _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09705_ vdd vss _04780_ _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input29_I vss i_dbus_rdt[5] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_94_clk vdd vss clknet_leaf_94_clk clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07897_ vss _03622_ _03359_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09636_ vdd _04726_ _01433_ _01103_ _04524_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07900__A2 vss _03547_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_229 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06848_ _02960_ vss vdd _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06779_ _02911_ vss vdd _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_09567_ vss _01077_ _04683_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09102__A1 vss _02908_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_796 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09498_ _01491_ vdd vss _04633_ cpu.alu.cmp_r _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08518_ vdd _04019_ _04017_ _00692_ _03956_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_1043 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1009 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06467__A2 vss _01682_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_310_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08449_ _03967_ net34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_163_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_777 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11460_ vdd rf_ram.memory\[345\]\[1\] clknet_leaf_167_clk vss _01192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07416__A1 vss _03292_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06219__A2 vss _01785_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10411_ vdd rf_ram.memory\[375\]\[1\] clknet_leaf_111_clk vss _00155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11391_ _01123_ vdd vss clknet_leaf_228_clk net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10342_ vdd rf_ram.memory\[283\]\[0\] clknet_leaf_178_clk vss _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07967__A2 vss _02954_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_325_clk_I vss clknet_5_4__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_398 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09169__A1 vss _04397_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_798 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05978__B2 vss rf_ram.memory\[13\]\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10273_ vdd rf_ram.memory\[234\]\[1\] clknet_leaf_261_clk vss _00017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05991__B vss _02186_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_85_clk vdd vss clknet_leaf_85_clk clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_185_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05363__C1 vss _01554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1170 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_413 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_616 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_971 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_470 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07655__A1 vss _03458_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06458__A2 vss _01508_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09644__A2 vss _01376_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_643 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_120 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_462 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_154_676 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11658_ vss net180 net108 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_83_298 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_438 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_693 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10609_ vdd rf_ram.memory\[355\]\[1\] clknet_leaf_156_clk vss _00353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11589_ vdd rf_ram.memory\[213\]\[0\] clknet_leaf_302_clk vss _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08080__A1 vss _03721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06062__B vss _01504_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08907__A1 vss _02959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06630__A2 vss _02801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05457__I vss _01518_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07820_ vdd _03574_ _03572_ _00439_ _03557_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09580__A1 vss _01391_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07751_ vdd _03531_ _03529_ _00413_ _03524_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06394__A1 vss _01972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09332__A1 vss _04466_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_76_clk vdd vss clknet_leaf_76_clk clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06702_ vdd vss _02856_ _02775_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07682_ _03488_ _03355_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06633_ vdd vss _02804_ rf_ram.memory\[293\]\[1\] _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07894__A1 vss _02836_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_240 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06697__A2 vss _02846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09421_ _02707_ vdd vss _04586_ net91 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06564_ vdd vss _02749_ rf_ram.memory\[200\]\[1\] _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09352_ _04540_ net231 vdd vss _04547_ net230 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07646__A1 vss _03071_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05515_ _01711_ _01613_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08303_ vdd vss _03875_ _03230_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09635__A2 vss net60 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06237__B vss _02431_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05657__B1 vss _01778_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06495_ _02235_ _02462_ _02689_ vdd vss _00001_ _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_16_800 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09283_ vdd vss _04504_ _01393_ _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05446_ vdd vss _01642_ rf_ram.memory\[382\]\[0\] _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_665 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_345 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08234_ vdd vss _03833_ rf_ram.memory\[531\]\[1\] _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05141__B vss cpu.state.genblk1.misalign_trap_sync_r vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_624 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08165_ vss _03790_ _03689_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_05377_ _01528_ vdd vss _01573_ rf_ram.memory\[552\]\[0\] _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_160_646 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07116_ vdd vss _03136_ _02915_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_825 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08096_ vdd vss _03747_ rf_ram.memory\[557\]\[1\] _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07047_ _03092_ _03017_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05367__I vss _01562_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_571 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08374__A2 vss _03903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08998_ vdd vss _04320_ rf_ram.memory\[112\]\[0\] _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_103_1092 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07949_ _03654_ _03359_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09323__A1 vss net243 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_67_clk vdd vss clknet_leaf_67_clk clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_825 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output135_I vss net135 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08126__A2 vss _03765_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10960_ vdd rf_ram.memory\[69\]\[0\] clknet_leaf_65_clk vss _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07885__A1 vss _03587_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10891_ vdd rf_ram.memory\[240\]\[1\] clknet_leaf_215_clk vss _00635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05345__C1 vss _01540_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09619_ vdd _04705_ _01333_ _01093_ _04643_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09874__A2 vss _01418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1029 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_289 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_407 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05360__A2 vss _01501_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06147__B vss _01650_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11512_ vdd rf_ram.memory\[305\]\[1\] clknet_leaf_144_clk vss _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_120 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_150_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11443_ vdd rf_ram.memory\[5\]\[0\] clknet_leaf_293_clk vss _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_264_clk_I vss clknet_5_17__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_123 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06661__I vss _02825_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_685 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08062__A1 vss net242 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11374_ vdd rf_ram.memory\[78\]\[1\] clknet_leaf_61_clk vss _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10325_ vdd rf_ram.memory\[291\]\[1\] clknet_leaf_123_clk vss _00069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_1289 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10256_ vdd _05123_ _05122_ _01327_ _02819_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_279_clk_I vss clknet_5_17__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_202_clk_I vss clknet_5_25__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10172__A2 vss _03134_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10187_ vdd vss _05082_ rf_ram.memory\[190\]\[1\] _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_58_clk vdd vss clknet_leaf_58_clk clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09314__A1 vss _04524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09314__B2 vss cpu.immdec.imm11_7\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_217_clk_I vss clknet_5_22__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_413 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07628__A1 vss _03425_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_468 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_665 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05300_ _01496_ vss vdd rf_ram.i_raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06280_ vss vdd rf_ram.memory\[149\]\[1\] _01968_ rf_ram.memory\[151\]\[1\] _01959_
+ _01940_ rf_ram.memory\[150\]\[1\] _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_182_793 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05231_ _01405_ cpu.branch_op vdd vss _01431_ cpu.bufreg.i_sh_signed net134 vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_188_36 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05162_ vdd vss _01365_ cpu.genblk3.csr.o_new_irq _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07800__A1 vss _03557_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09970_ vdd vss _04948_ rf_ram.memory\[464\]\[0\] _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_510 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08921_ vdd _04272_ _04271_ _00842_ _04266_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08852_ vdd _04229_ _04228_ _00816_ _04202_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07803_ vdd _03564_ _03563_ _00432_ _03554_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_49_clk vdd vss clknet_leaf_49_clk clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08783_ vdd vss _04187_ rf_ram.memory\[141\]\[0\] _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05995_ vss vdd rf_ram.memory\[527\]\[1\] _01521_ rf_ram.memory\[525\]\[1\] _01517_
+ _01511_ rf_ram.memory\[524\]\[1\] _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_07734_ vdd _03520_ _03518_ _00407_ _03491_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09305__A1 vss _04463_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07665_ vdd _03477_ _03475_ _00381_ _03458_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07867__A1 vss _03590_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09856__A2 vss _01413_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06616_ vdd vss _02790_ rf_ram.memory\[236\]\[0\] _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09404_ _04539_ net226 vdd vss _04575_ net225 _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07596_ vdd vss _03435_ rf_ram.memory\[315\]\[1\] _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05650__I vss _01536_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09122__I vss _02742_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09608__A2 vss _04507_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07619__A1 vss _02904_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09335_ vdd _04537_ _04536_ _00991_ _04463_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06547_ vdd vss _02733_ _01352_ cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08292__A1 vss _03855_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06478_ _02669_ _02672_ vdd vss _02673_ _02661_ _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09266_ vdd _04491_ _04481_ _00968_ _04480_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05429_ vdd vss _01625_ _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_28_490 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08217_ vdd _03822_ _03821_ _00588_ _03820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09197_ vdd vss _04444_ rf_ram.memory\[82\]\[1\] _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_419 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08148_ vdd _03779_ _03778_ _00562_ _03754_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08044__A1 vss _03690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08079_ vdd vss _03737_ rf_ram.memory\[560\]\[0\] _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10110_ vdd vss _05034_ net250 _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11090_ vdd rf_ram.memory\[128\]\[1\] clknet_leaf_26_clk vss _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05802__B1 vss _01520_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10041_ vdd vss _04992_ rf_ram.memory\[305\]\[1\] _04990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09544__A1 vss _04478_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07858__A1 vss _02728_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10943_ vdd cpu.state.ibus_cyc clknet_leaf_255_clk vss _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05869__B1 vss _01625_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05560__I vss _01601_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10874_ vdd rf_ram.memory\[203\]\[0\] clknet_leaf_35_clk vss _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_3_0_0_clk clknet_3_0_0_clk vss vdd clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__05333__A2 vss _01524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1200 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06656__I vss _02821_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_1209 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_232 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08283__A1 vss _03230_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1244 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_793 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10090__A1 vss _03445_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_164 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_83_clk_I vss clknet_5_11__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_955 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11426_ vdd rf_ram.memory\[259\]\[1\] clknet_leaf_201_clk vss _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08035__A1 vss _02991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_931 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06046__B1 vss _01608_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11357_ vdd rf_ram.memory\[73\]\[1\] clknet_leaf_22_clk vss _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_688 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1075 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_98_clk_I vss clknet_5_14__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10308_ vdd rf_ram.memory\[516\]\[0\] clknet_leaf_271_clk vss _00052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11288_ vdd net225 clknet_leaf_248_clk vss _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_141_clk_I vss clknet_5_27__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05735__I vss _01626_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ vdd vss _05113_ _02737_ _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05557__C1 vss _01636_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_21_clk_I vss clknet_5_3__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05780_ _01923_ vdd vss _01976_ rf_ram.memory\[128\]\[0\] _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_156_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1014 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_1144 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07450_ vdd vss _03344_ rf_ram.memory\[368\]\[0\] _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05470__I vss _01643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1095 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_36_clk_I vss clknet_5_6__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07381_ vdd vss _03301_ rf_ram.memory\[266\]\[0\] _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06401_ _01746_ vdd vss _02596_ _02594_ _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_17_405 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07077__A2 vss _02911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06332_ _01551_ vdd vss _02527_ rf_ram.memory\[216\]\[1\] _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_427 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_298 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09120_ vdd vss _04395_ rf_ram.memory\[575\]\[1\] _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10081__A1 vss _05014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09051_ vdd vss _04353_ rf_ram.memory\[102\]\[0\] _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_235 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06263_ _02457_ vdd vss _02458_ _01350_ _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08002_ vdd vss _03688_ rf_ram.memory\[465\]\[0\] _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_600 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06194_ rf_ram.memory\[477\]\[1\] _01848_ _01863_ rf_ram.memory\[476\]\[1\] _02389_
+ vss vdd rf_ram.memory\[479\]\[1\] _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_130_616 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_605 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1165 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05214_ vdd vss _01414_ net134 _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09774__A1 vss _04637_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmax_cap253 net253 _01568_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05145_ _01347_ vdd vss _01348_ cpu.csr_imm _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xmax_cap242 net242 _02865_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_109_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09953_ vdd _04937_ _04935_ _01210_ _04921_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11647__I vss net128 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09526__A1 vss _03967_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05260__A1 vss _01436_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08904_ vdd _04261_ _04260_ _00836_ _04234_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_395 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09884_ vdd vss _04895_ rf_ram.memory\[229\]\[1\] _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08835_ vdd vss _04219_ _03672_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08766_ vdd _04176_ _04174_ _00783_ _04170_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07717_ vdd _03510_ _03509_ _00400_ _03488_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_5_25__f_clk_I vss clknet_3_6_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input11_I vss i_dbus_rdt[18] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05978_ rf_ram.memory\[12\]\[0\] _02174_ vss vdd rf_ram.memory\[15\]\[0\] _01653_
+ rf_ram.memory\[13\]\[0\] _01655_ _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_178_852 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_614 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_80 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08697_ vdd vss _04133_ rf_ram.memory\[153\]\[1\] _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09280__C vss _01391_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07648_ vdd _03467_ _03466_ _00374_ _03455_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07579_ vdd _03424_ _03423_ _00348_ _03422_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08691__I vss _04061_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08265__A1 vss _03823_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09318_ vdd vss _04527_ _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10590_ vdd rf_ram.memory\[320\]\[0\] clknet_leaf_165_clk vss _00334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10072__A1 vss _04985_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_533 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05618__A3 vss _01813_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_635 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09249_ vss _04478_ _04477_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__08017__A1 vss _03686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06144__C vss _01717_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11211_ vdd rf_ram.memory\[82\]\[1\] clknet_leaf_47_clk vss _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08568__A2 vss _03949_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11142_ vdd rf_ram.memory\[10\]\[0\] clknet_leaf_35_clk vss _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_373 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09517__A1 vss _04643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput76 o_dbus_adr[19] net76 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_179_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11073_ vdd rf_ram.memory\[469\]\[0\] clknet_leaf_54_clk vss _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06160__B vss _01746_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput87 o_dbus_adr[2] net87 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput98 o_dbus_dat[0] net98 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10024_ vdd vss _04981_ rf_ram.memory\[246\]\[1\] _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06200__B1 vss _01725_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_920 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05504__B vss _01620_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10926_ vdd rf_ram.memory\[174\]\[0\] clknet_leaf_8_clk vss _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10857_ vdd rf_ram.memory\[528\]\[1\] clknet_leaf_309_clk vss _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10063__A1 vss _03445_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_235 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10788_ vdd rf_ram.memory\[562\]\[0\] clknet_leaf_323_clk vss _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_758 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08256__A1 vss _02845_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06335__B vss _01928_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08008__A1 vss _02730_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11409_ vdd rf_ram.memory\[77\]\[0\] clknet_leaf_20_clk vss _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09756__B2 vss net118 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07945__I vss _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07231__A2 vss _03040_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05778__C1 vss _01925_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06950_ vdd _03028_ _03026_ _00115_ _03018_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_182_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input3_I vss i_dbus_rdt[10] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06881_ vdd vss _02982_ rf_ram.memory\[301\]\[1\] _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05901_ rf_ram.memory\[84\]\[0\] _02097_ vss vdd rf_ram.memory\[87\]\[0\] _01763_
+ rf_ram.memory\[85\]\[0\] _01656_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__05465__I vss _01499_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06990__A1 vss _03053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05832_ _01959_ rf_ram.memory\[219\]\[0\] vdd vss _02028_ rf_ram.memory\[218\]\[0\]
+ _01940_ _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08620_ vdd vss _04085_ _02760_ _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05545__A2 vss _01623_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06742__A1 vss _02881_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08551_ vdd vss _04041_ rf_ram.memory\[119\]\[1\] _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05950__C1 vss _01635_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05763_ _01959_ vss vdd _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08495__A1 vss _03953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07502_ vdd _03376_ _03374_ _00319_ _03360_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05694_ _01790_ vdd vss _01890_ _01887_ _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_89_485 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08482_ vdd _03994_ _03993_ _00681_ _03991_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07433_ vdd _03333_ _03331_ _00293_ _03326_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_1180 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09103_ vdd vss _04385_ rf_ram.memory\[95\]\[0\] _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07364_ vdd vss _03290_ _03055_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_398 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09995__A1 vss _04953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07295_ vdd vss _03247_ _02984_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06315_ rf_ram.memory\[184\]\[1\] _02510_ vss vdd rf_ram.memory\[187\]\[1\] _01773_
+ rf_ram.memory\[185\]\[1\] _01848_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__08798__A2 vss _04195_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06246_ vdd vss _02441_ rf_ram.memory\[441\]\[1\] _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06245__B vss _01923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09034_ vdd _04342_ _04340_ _00885_ _04334_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_796 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09747__B2 vss net115 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09747__A1 vss net114 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_696 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06177_ _01526_ vdd vss _02372_ rf_ram.memory\[496\]\[1\] _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_7_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05128_ vdd vss cpu.decode.op26 _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input59_I vss i_ibus_rdt[4] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09936_ vdd _04927_ _04926_ _01203_ _04918_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06430__B1 vss _01848_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_280_clk vdd vss clknet_leaf_280_clk clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06981__A1 vss _03014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05784__A2 vss _01770_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09867_ vdd vss _04885_ _02838_ _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06194__C1 vss _01696_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09798_ vdd vss _04843_ rf_ram.memory\[58\]\[0\] _04842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08818_ vdd vss _04209_ rf_ram.memory\[137\]\[1\] _04207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06733__A1 vss _02876_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_23__f_clk vdd vss clknet_5_23__leaf_clk clknet_3_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08749_ vdd _04165_ _04164_ _00777_ _04126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_184_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10711_ vdd rf_ram.memory\[40\]\[1\] clknet_leaf_134_clk vss _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_1063 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1074 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_803 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_371 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10642_ vdd rf_ram.memory\[402\]\[0\] clknet_leaf_96_clk vss _00386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_579 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08238__A1 vss _03820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10573_ vdd rf_ram.memory\[364\]\[1\] clknet_leaf_162_clk vss _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10045__A1 vss _04982_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09986__A1 vss _02915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_588 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_465 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_1062 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_958 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05994__B vss _01506_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08410__A1 vss _02761_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06421__B1 vss _01772_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11125_ vdd rf_ram.memory\[118\]\[1\] clknet_leaf_73_clk vss _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_271_clk vdd vss clknet_leaf_271_clk clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_43_1067 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11056_ vdd rf_ram.memory\[149\]\[1\] clknet_leaf_1_clk vss _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09910__A1 vss _04887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10007_ vdd vss _04971_ rf_ram.memory\[277\]\[0\] _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05527__A2 vss _01706_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06724__A1 vss _02820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_647 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08477__A1 vss _01491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_682 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_568 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10909_ vdd rf_ram.memory\[189\]\[1\] clknet_leaf_26_clk vss _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_516 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1248 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_853 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_393 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09977__A1 vss _04950_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_763 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06100_ _01615_ vdd vss _02295_ rf_ram.memory\[272\]\[1\] _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07080_ vdd vss _03113_ rf_ram.memory\[492\]\[1\] _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_54_374 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06031_ rf_ram.memory\[562\]\[1\] _02226_ vss vdd rf_ram.memory\[561\]\[1\] _01555_
+ rf_ram.memory\[563\]\[1\] _01554_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_160_1026 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_777 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07982_ vdd vss _03675_ rf_ram.memory\[478\]\[1\] _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_466 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_262_clk vdd vss clknet_leaf_262_clk clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09721_ vdd vss _04792_ _04781_ net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06933_ _03018_ vss vdd _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09901__A1 vss _03319_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06864_ _02970_ _02819_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06176__C1 vss _01519_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09652_ vss _04739_ net1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XANTENNA__08704__A2 vss _04078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05923__C1 vss _01625_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05815_ rf_ram.memory\[181\]\[0\] _01772_ _01799_ rf_ram.memory\[180\]\[0\] _02011_
+ vss vdd rf_ram.memory\[183\]\[0\] _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08603_ vdd vss _04074_ net241 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09583_ vdd vss _04695_ _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06795_ _02923_ _02922_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_05746_ rf_ram.memory\[420\]\[0\] _01942_ vss vdd rf_ram.memory\[423\]\[0\] _01646_
+ rf_ram.memory\[421\]\[0\] _01810_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_179_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06191__A2 vss _01856_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08534_ vdd vss _04030_ rf_ram.memory\[69\]\[1\] _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_400 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_811 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05677_ rf_ram.memory\[453\]\[0\] _01810_ _01666_ rf_ram.memory\[452\]\[0\] _01873_
+ vss vdd rf_ram.memory\[455\]\[0\] _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__07140__A1 vss _03126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_477 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08465_ vdd vss _03982_ _01381_ net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_161_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07416_ vdd _03322_ _03320_ _00287_ _03292_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08396_ vdd vss _03934_ rf_ram.memory\[17\]\[0\] _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_858 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10027__A1 vss _04911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09968__A1 vss _04921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07347_ vdd _03279_ _03277_ _00261_ _03260_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_812 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_385 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07278_ vdd vss _03237_ rf_ram.memory\[417\]\[1\] _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09017_ vss _04331_ _04057_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06229_ rf_ram.memory\[411\]\[1\] _01726_ _01801_ rf_ram.memory\[410\]\[1\] _02424_
+ vss vdd rf_ram.memory\[409\]\[1\] _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09440__I0 vss net70 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06403__B1 vss _01656_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_253_clk vdd vss clknet_leaf_253_clk clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09919_ vdd _04916_ _04915_ _01197_ _04884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06706__A1 vss _02826_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06182__A2 vss _01846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_945 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_438 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08459__A1 vss net120 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07131__A1 vss _02806_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_414 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_308 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_458 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10625_ vdd rf_ram.memory\[388\]\[1\] clknet_leaf_95_clk vss _00369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09959__A1 vss _04911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10018__A1 vss _04950_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10186__I vss _02747_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1210 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07434__A2 vss _02815_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10556_ vdd rf_ram.memory\[368\]\[0\] clknet_leaf_148_clk vss _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_1254 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10487_ vdd rf_ram.memory\[196\]\[1\] clknet_leaf_42_clk vss _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_254 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05996__A2 vss _01524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08934__A2 vss _03559_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1010 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07198__A1 vss _03161_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_244_clk vdd vss clknet_leaf_244_clk clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_764 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05748__A2 vss _01662_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11108_ vdd rf_ram.memory\[124\]\[0\] clknet_leaf_85_clk vss _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06945__A1 vss _03018_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08698__A1 vss _04129_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11039_ _00776_ rf_ram.i_raddr\[3\] vdd vss clknet_leaf_275_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_177_928 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07370__A1 vss _02781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05600_ _01791_ _01795_ vdd vss _01796_ _01775_ _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06173__A2 vss _01652_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_455 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1080 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05381__B1 vss _01539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06580_ vdd vss _02734_ _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_05531_ rf_ram.memory\[328\]\[0\] _01727_ vss vdd rf_ram.memory\[331\]\[0\] _01726_
+ rf_ram.memory\[329\]\[0\] _01725_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_157_652 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05899__B vss _01746_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05462_ _01658_ _01563_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_117_505 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08250_ vdd _03842_ _03840_ _00601_ _03823_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07201_ vdd _03188_ _03187_ _00206_ _03157_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08181_ vdd _03800_ _03799_ _00574_ _03787_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_508 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07132_ vdd vss _03146_ rf_ram.memory\[486\]\[0\] _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_491 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05393_ _01528_ vdd vss _01589_ rf_ram.memory\[568\]\[0\] _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08622__A1 vss _04058_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07063_ vdd vss _03103_ rf_ram.memory\[375\]\[0\] _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput200 o_ext_rs2[8] net200 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09178__A2 vss _04418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput211 o_ibus_adr[18] net211 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput233 o_ibus_adr[9] net233 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput222 o_ibus_adr[28] net222 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06014_ _02207_ _02208_ vdd vss _02209_ _02205_ _02206_ _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07189__A1 vss _02836_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_235_clk vdd vss clknet_leaf_235_clk clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05739__A2 vss _01804_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06397__C1 vss _01773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06936__A1 vss _02766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07965_ vdd vss _03664_ rf_ram.memory\[470\]\[1\] _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11655__I vss net105 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06916_ vdd _03005_ _03004_ _00104_ _02970_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09704_ _04768_ _04779_ vdd vss _04780_ net100 _04767_ net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__06749__I vss _02888_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07896_ vdd _03621_ _03620_ _00468_ _03619_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09350__A2 vss _03991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09635_ vdd vss _04726_ _04524_ net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06847_ vdd vss _02959_ _02750_ _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_179_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05911__A2 vss _01787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06778_ vdd vss _02910_ _02764_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08964__I vss _04057_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_764 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09566_ _04678_ vdd vss _04683_ cpu.immdec.imm30_25\[1\] _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10248__A1 vss _02825_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09102__A2 vss _04005_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07113__A1 vss _03126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05729_ _01925_ vss vdd _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09497_ _04630_ _04631_ _01440_ vdd vss _04632_ _04628_ _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_08517_ vdd vss _04019_ rf_ram.memory\[172\]\[1\] _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08861__A1 vss _02983_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08448_ vdd _03966_ _03964_ _00675_ _03956_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_184_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_817 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10410_ vdd rf_ram.memory\[375\]\[0\] clknet_leaf_111_clk vss _00154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_869 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08379_ vdd _03923_ _03920_ _00649_ _03922_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11390_ _01122_ vdd vss clknet_leaf_228_clk net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10341_ vdd rf_ram.memory\[284\]\[1\] clknet_leaf_173_clk vss _00085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05978__A2 vss _01643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10272_ vdd rf_ram.memory\[234\]\[0\] clknet_leaf_261_clk vss _00016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_226_clk vdd vss clknet_leaf_226_clk clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05991__C vss _01373_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06155__A2 vss _01677_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07352__A1 vss _03260_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_725 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05902__A2 vss _01863_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_230 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05363__B1 vss _01555_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_909 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_572 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07104__A1 vss _02915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10239__A1 vss _02737_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05512__B vss _01707_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_745 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08852__A1 vss _04202_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11657_ net179 vss vdd net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_36_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10608_ vdd rf_ram.memory\[355\]\[0\] clknet_leaf_156_clk vss _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11588_ vdd rf_ram.memory\[208\]\[1\] clknet_leaf_32_clk vss _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_193 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10539_ vdd rf_ram.memory\[247\]\[1\] clknet_leaf_213_clk vss _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_714 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05969__A2 vss _01682_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06343__B vss _01916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_217_clk vdd vss clknet_leaf_217_clk clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_561 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08907__A2 vss _04038_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06918__A1 vss _02975_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07750_ vdd vss _03531_ rf_ram.memory\[377\]\[1\] _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06701_ vdd _02855_ _02853_ _00039_ _02826_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06146__A2 vss _01724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07681_ vdd _03487_ _03485_ _00387_ _03458_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07343__A1 vss _03055_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06632_ vdd _02803_ _02802_ _00022_ _02743_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07894__A2 vss _02844_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09420_ vss _01028_ _04585_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09096__A1 vss _04367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09351_ vdd vss _04546_ _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06563_ _02748_ _02747_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05514_ rf_ram.memory\[324\]\[0\] _01710_ vss vdd rf_ram.memory\[327\]\[0\] _01654_
+ rf_ram.memory\[325\]\[0\] _01656_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_08302_ vdd _03874_ _03872_ _00621_ _03855_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09282_ _04503_ vdd vss _00972_ _04497_ _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_173_953 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07646__A2 vss _03089_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_994 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06237__C vss net254 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06494_ vdd vss _02689_ _01371_ _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08233_ vdd _03832_ _03831_ _00594_ _03820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05445_ _01641_ vss vdd _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__05141__C vss cpu.genblk3.csr.o_new_irq vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05376_ rf_ram.memory\[557\]\[0\] _01517_ _01511_ rf_ram.memory\[556\]\[0\] _01572_
+ vss vdd rf_ram.memory\[559\]\[0\] _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08164_ vdd _03789_ _03788_ _00568_ _03787_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_193 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_995 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07115_ _03135_ vss vdd _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08095_ vdd _03746_ _03745_ _00542_ _03721_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06253__B vss _01805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06082__A1 vss _01603_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_360 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07046_ vdd _03091_ _03090_ _00148_ _03087_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_185 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_208_clk vdd vss clknet_leaf_208_clk clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09020__A1 vss _04331_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_257 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06909__A1 vss _02822_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1060 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input41_I vss i_ibus_rdt[16] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07582__A1 vss _03425_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08997_ vdd vss _04319_ _02945_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06385__A2 vss _01918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05593__B1 vss _01786_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07948_ vdd _03653_ _03652_ _00488_ _03651_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06137__A2 vss _01777_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07879_ vdd vss _03611_ rf_ram.memory\[446\]\[0\] _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output128_I vss net128 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09323__A2 vss _04037_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10890_ vdd rf_ram.memory\[240\]\[0\] clknet_leaf_214_clk vss _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05345__B1 vss _01539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09618_ vdd _04707_ _01460_ _01092_ _04643_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_1106 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05896__A1 vss _01769_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09549_ vdd vss _04669_ _01447_ _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_1139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09087__A1 vss _02983_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_520 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_633 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08834__A1 vss _04205_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11511_ vdd rf_ram.memory\[305\]\[0\] clknet_leaf_150_clk vss _01243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_327 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_379 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05986__C vss _01493_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11442_ _01174_ vdd vss clknet_leaf_239_clk cpu.state.genblk1.misalign_trap_sync_r
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11373_ vdd rf_ram.memory\[78\]\[0\] clknet_leaf_60_clk vss _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10324_ vdd rf_ram.memory\[291\]\[0\] clknet_leaf_135_clk vss _00068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08062__A2 vss _03693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_360 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09011__A1 vss _04301_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10255_ vdd vss _05123_ rf_ram.memory\[9\]\[0\] _05122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05820__A1 vss _01768_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_881 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_1000 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10186_ _05081_ _02747_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07573__A1 vss _03389_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06376__A2 vss _01863_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05584__B1 vss _01778_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06128__A2 vss _01692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07325__A1 vss _03257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09314__A2 vss net63 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07628__A2 vss _03452_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_920 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05639__A1 vss _01527_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08825__A1 vss _02828_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06300__A2 vss _01846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_485 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_759 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_236 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05230_ vdd vss _01429_ _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_181_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_461 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_686 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05161_ vdd vss cpu.state.genblk1.misalign_trap_sync_r _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__05468__I vss _01514_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09250__A1 vss _04478_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08920_ vdd vss _04272_ rf_ram.memory\[389\]\[0\] _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09002__A1 vss _02953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08851_ vdd vss _04229_ rf_ram.memory\[132\]\[0\] _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_1032 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07802_ vdd vss _03564_ rf_ram.memory\[435\]\[0\] _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08782_ vdd vss _04186_ net243 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05994_ _01506_ vdd vss _02189_ rf_ram.memory\[526\]\[1\] _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07733_ vdd vss _03520_ rf_ram.memory\[397\]\[1\] _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06119__A2 vss _01509_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_4__f_clk vdd vss clknet_5_4__leaf_clk clknet_3_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07664_ vdd vss _03477_ rf_ram.memory\[385\]\[1\] _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_324_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1080 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_369 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_509 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05878__A1 vss _01368_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06615_ vdd vss _02789_ _02766_ _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09403_ vdd vss _04574_ _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07595_ vdd _03434_ _03433_ _00354_ _03422_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_149_268 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06248__B vss _01928_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09069__A1 vss _04334_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07619__A2 vss _03390_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09334_ vdd vss _04537_ rf_ram.memory\[99\]\[0\] _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06546_ rf_ram_if.wen0_r rf_ram_if.wen1_r _01347_ vdd vss _02732_ rf_ram_if.rtrig1
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_146_964 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_121 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06477_ _02671_ vdd vss _02672_ _01903_ _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_339_clk_I vss clknet_5_0__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09265_ vdd vss _04491_ cpu.genblk3.csr.mstatus_mpie _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09196_ vdd _04443_ _04442_ _00946_ _04431_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05428_ _01624_ vss vdd _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_69_1246 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08216_ vdd vss _03822_ rf_ram.memory\[534\]\[0\] _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_198 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08147_ vdd vss _03779_ rf_ram.memory\[547\]\[0\] _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05359_ _01555_ vss vdd _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09241__A1 vss _01418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_155 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08078_ vdd vss _03736_ _02945_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07029_ vdd vss _03079_ _02738_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10040_ vdd _04991_ _04990_ _01243_ _04982_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09544__A2 vss net42 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07555__A1 vss _03393_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06358__A2 vss _01940_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_601 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_98_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10942_ vdd rf_ram_if.rdata1 clknet_leaf_280_clk vss _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07858__A2 vss _02869_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09313__I vss _03992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10873_ vdd rf_ram.memory\[192\]\[1\] clknet_leaf_46_clk vss _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08807__A1 vss _04170_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08283__A2 vss _02788_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10090__A2 vss _03009_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_986 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1060 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_135 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09232__A1 vss _04463_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_989 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11425_ vdd rf_ram.memory\[259\]\[0\] clknet_leaf_201_clk vss _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08035__A2 vss _03693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_954 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11356_ vdd rf_ram.memory\[73\]\[0\] clknet_leaf_20_clk vss _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07794__A1 vss _03557_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10307_ vdd rf_ram.memory\[517\]\[1\] clknet_leaf_273_clk vss _00051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11287_ vdd net223 clknet_leaf_243_clk vss _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07546__A1 vss _02921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06349__A2 vss _01801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10238_ vdd _05112_ _05110_ _01320_ _02825_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10169_ vdd _05070_ _05069_ _01293_ _05046_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05557__B1 vss _01645_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_1074 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_1204 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06400_ rf_ram.memory\[91\]\[1\] _01646_ _01801_ rf_ram.memory\[90\]\[1\] _02595_
+ vss vdd rf_ram.memory\[89\]\[1\] _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07380_ vdd vss _03300_ _02775_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_512 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06331_ _01978_ vdd vss _02526_ _02523_ _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06262_ _02454_ _02455_ _02456_ _01717_ vdd vss _02457_ _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_143_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09050_ vdd vss _04352_ _02805_ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06285__A1 vss _01972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_940 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_753 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08001_ vdd vss _03687_ _02761_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_4_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05213_ _01385_ cpu.state.o_cnt\[2\] vdd vss _01413_ cpu.state.cnt_r\[3\] cpu.mem_bytecnt\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__09223__A1 vss _04434_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06193_ vdd vss _02388_ rf_ram.memory\[478\]\[1\] _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05144_ _01347_ vss vdd rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07785__A1 vss _03521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09952_ vdd vss _04937_ rf_ram.memory\[337\]\[1\] _04935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1029 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08903_ vdd vss _04261_ rf_ram.memory\[126\]\[0\] _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05260__A2 vss _01437_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09883_ vdd _04894_ _04893_ _01183_ _04884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08834_ vdd _04218_ _04216_ _00809_ _04205_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_139_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_263_clk_I vss clknet_5_17__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08765_ vdd vss _04176_ rf_ram.memory\[145\]\[1\] _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07716_ vdd vss _03510_ rf_ram.memory\[380\]\[0\] _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05977_ _01503_ vdd vss _02173_ rf_ram.memory\[14\]\[0\] _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_79_133 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11663__I vss net114 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_1114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05661__I vss _01695_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08696_ vdd _04132_ _04131_ _00757_ _04126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07647_ vdd vss _03467_ rf_ram.memory\[405\]\[0\] _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06512__A2 vss cpu.decode.opcode\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07578_ vdd vss _03424_ rf_ram.memory\[356\]\[0\] _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_278_clk_I vss clknet_5_17__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11368__CLK vss clknet_5_20__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_238 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06529_ vdd vss net234 _02714_ _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09317_ cpu.immdec.imm11_7\[3\] _04521_ net64 _04526_ _04527_ vss vdd cpu.immdec.imm11_7\[2\]
+ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__05610__B vss _01805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1043 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_661 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_951 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_201_clk_I vss clknet_5_25__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_887 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output195_I vss net195 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_258 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09248_ vss _04477_ net34 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__05484__C1 vss _01679_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09179_ vdd vss _04433_ rf_ram.memory\[84\]\[0\] _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09214__A1 vss net240 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_217 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11210_ vdd rf_ram.memory\[82\]\[0\] clknet_leaf_47_clk vss _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09765__A2 vss _04766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_976 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07776__A1 vss _03524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11141_ vdd rf_ram.memory\[110\]\[1\] clknet_leaf_69_clk vss _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_998 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_max_cap241_I vss _02882_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_216_clk_I vss clknet_5_22__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output72_I vss net72 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11072_ vdd rf_ram.memory\[459\]\[1\] clknet_leaf_52_clk vss _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput99 o_dbus_dat[10] net99 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput88 o_dbus_adr[30] net88 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput77 o_dbus_adr[20] net77 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10023_ vdd _04980_ _04979_ _01237_ _04950_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07700__A1 vss _02945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_659 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10925_ vdd rf_ram.memory\[59\]\[1\] clknet_leaf_296_clk vss _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06503__A2 vss cpu.genblk3.csr.o_new_irq vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1070 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_158 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1165 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10856_ vdd rf_ram.memory\[528\]\[0\] clknet_leaf_309_clk vss _00600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_867 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_238 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06267__A1 vss _01373_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10787_ vdd rf_ram.memory\[563\]\[1\] clknet_leaf_332_clk vss _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08256__A2 vss _02972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10063__A2 vss _02866_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_397 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11408_ vdd rf_ram.memory\[269\]\[1\] clknet_5_28__leaf_clk vss _01140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09756__A2 vss _04766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07767__A1 vss _02752_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06351__B vss _01350_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05778__B1 vss _01912_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11339_ vdd cpu.immdec.imm19_12_20\[5\] clknet_leaf_215_clk vss _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06880_ vdd _02981_ _02980_ _00092_ _02970_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05900_ _01707_ vdd vss _02096_ rf_ram.memory\[86\]\[0\] _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_175_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_1114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05831_ vdd vss _02027_ rf_ram.memory\[217\]\[0\] _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06742__A2 vss _02883_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08550_ vdd _04040_ _04039_ _00703_ _04023_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_453 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05481__I vss _01633_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05950__B1 vss _01609_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05762_ _01958_ vss vdd _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07501_ vdd vss _03376_ rf_ram.memory\[324\]\[1\] _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05693_ _01786_ rf_ram.memory\[387\]\[0\] vdd vss _01889_ rf_ram.memory\[386\]\[0\]
+ _01856_ _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_134_53 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08481_ vdd vss _03994_ cpu.state.ibus_cyc _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_186_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07432_ vdd vss _03333_ rf_ram.memory\[370\]\[1\] _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_158 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09692__B2 vss net128 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_322 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_309 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09102_ vdd vss _04384_ _02908_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07363_ _03289_ _03013_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07294_ vdd _03246_ _03244_ _00241_ _03225_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06314_ _01916_ vdd vss _02509_ rf_ram.memory\[186\]\[1\] _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_1205 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06245_ _01923_ vdd vss _02440_ rf_ram.memory\[440\]\[1\] _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09033_ vdd vss _04342_ rf_ram.memory\[106\]\[1\] _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_770 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_285 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06176_ rf_ram.memory\[500\]\[1\] _02371_ vss vdd rf_ram.memory\[503\]\[1\] _01519_
+ rf_ram.memory\[501\]\[1\] _01668_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_130_469 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_475 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1093 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_661 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05769__B1 vss _01953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09935_ vdd vss _04927_ rf_ram.memory\[340\]\[0\] _04926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_1174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09866_ _04884_ _04396_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_102_1147 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08817_ vdd _04208_ _04207_ _00802_ _04202_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08183__A1 vss _03790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_82_clk_I vss clknet_5_11__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06194__B1 vss _01848_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07930__A1 vss _02991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09797_ vdd vss _04842_ net245 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_913 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08748_ vdd vss _04165_ rf_ram.memory\[147\]\[0\] _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09683__A1 vss net1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08679_ vdd _04121_ _04120_ _00751_ _04094_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10710_ vdd rf_ram.memory\[40\]\[0\] clknet_leaf_134_clk vss _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_467 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_97_clk_I vss clknet_5_14__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10641_ vdd rf_ram.memory\[384\]\[1\] clknet_leaf_92_clk vss _00385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_140_clk_I vss clknet_5_27__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10572_ vdd rf_ram.memory\[364\]\[0\] clknet_leaf_162_clk vss _00316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_945 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09986__A2 vss _03083_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_992 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_20_clk_I vss clknet_5_3__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_155_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07749__A1 vss _03521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_935 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08410__A2 vss _03903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_35_clk_I vss clknet_5_6__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11124_ vdd rf_ram.memory\[118\]\[0\] clknet_leaf_76_clk vss _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11055_ vdd rf_ram.memory\[149\]\[0\] clknet_leaf_1_clk vss _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10006_ vdd vss _04970_ _02940_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_157_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_261 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1078 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10908_ vdd rf_ram.memory\[189\]\[0\] clknet_leaf_13_clk vss _00652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08477__A2 vss _03989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05696__C1 vss _01848_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_670 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_169 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_309 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_108_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_377 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06346__B vss _01805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10839_ vdd rf_ram.memory\[537\]\[1\] clknet_leaf_314_clk vss _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09977__A2 vss _04951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_578 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07988__A1 vss _03654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06030_ _01552_ vdd vss _02225_ rf_ram.memory\[560\]\[1\] _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1146 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07981_ vdd _03674_ _03673_ _00500_ _03651_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06932_ _03017_ _02747_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09720_ _04791_ vss vdd _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09901__A2 vss _02984_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06863_ vdd _02969_ _02967_ _00087_ _02930_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07912__A1 vss _03619_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06176__B1 vss _01668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09651_ vdd vss _04738_ net98 _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05425__B vss _01620_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05923__B1 vss _01702_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_913 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05814_ _01505_ vdd vss _02010_ rf_ram.memory\[182\]\[0\] _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08602_ vdd _04073_ _04071_ _00722_ _04062_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09582_ vdd _04694_ _04678_ _04695_ cpu.immdec.imm30_25\[5\] vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06794_ vdd vss _02922_ _02773_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05745_ _01805_ vdd vss _01941_ rf_ram.memory\[422\]\[0\] _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08533_ vdd _04029_ _04028_ _00697_ _04023_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_272 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_1231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_642 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05676_ _01805_ vdd vss _01872_ rf_ram.memory\[454\]\[0\] _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08464_ vdd _03981_ _01399_ _01442_ _01447_ vss _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_07415_ vdd vss _03322_ rf_ram.memory\[334\]\[1\] _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08395_ vdd vss _03933_ _02761_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10027__A2 vss _02829_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_731 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07346_ vdd vss _03279_ rf_ram.memory\[253\]\[1\] _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_550 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07979__A1 vss _03672_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_846 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_323 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07277_ vdd _03236_ _03235_ _00234_ _03222_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_252 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09016_ vdd _04330_ _04328_ _00879_ _04301_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06228_ _01615_ vdd vss _02423_ rf_ram.memory\[408\]\[1\] _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06770__I vss _02903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_570 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06159_ _01688_ rf_ram.memory\[491\]\[1\] vdd vss _02354_ rf_ram.memory\[490\]\[1\]
+ _01687_ _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09440__I1 vss net71 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05611__C1 vss _01726_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09918_ vdd vss _04916_ rf_ram.memory\[343\]\[0\] _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output158_I vss net158 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08156__A1 vss net238 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1029 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09849_ vdd vss _01169_ _02713_ _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_1137 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_1218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07131__A2 vss _02911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_889 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10624_ vdd rf_ram.memory\[388\]\[0\] clknet_leaf_94_clk vss _00368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09959__A2 vss _02954_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05693__A2 vss _01856_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06890__A1 vss _02788_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_640 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_824 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10555_ vdd rf_ram.memory\[331\]\[1\] clknet_leaf_151_clk vss _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_561 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_559 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09477__B vss _03989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_745 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10486_ vdd rf_ram.memory\[196\]\[0\] clknet_leaf_43_clk vss _00230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_1168 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06642__A1 vss _02756_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_581 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08395__A1 vss _02761_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09431__I1 vss net67 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05602__C1 vss _01713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11107_ vdd rf_ram.memory\[389\]\[1\] clknet_leaf_116_clk vss _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09895__A1 vss _04887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11038_ _00775_ vdd vss clknet_leaf_285_clk rf_ram.i_raddr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07370__A2 vss _03253_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05530_ _01726_ _01635_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_115_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_77 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05461_ rf_ram.memory\[378\]\[0\] _01657_ vss vdd rf_ram.memory\[377\]\[0\] _01656_
+ rf_ram.memory\[379\]\[0\] _01654_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xclkbuf_leaf_180_clk vdd vss clknet_leaf_180_clk clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_138_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_908 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06330__B1 vss _02019_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05684__A2 vss _01770_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06076__B vss _01684_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07200_ vdd vss _03188_ rf_ram.memory\[273\]\[0\] _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_1068 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_331 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08180_ vdd vss _03800_ rf_ram.memory\[541\]\[0\] _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05392_ rf_ram.memory\[573\]\[0\] _01555_ _01538_ rf_ram.memory\[572\]\[0\] _01588_
+ vss vdd rf_ram.memory\[575\]\[0\] _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07131_ vdd vss _03145_ _02806_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07686__I vss _03359_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05436__A2 vss _01631_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07062_ vdd vss _03102_ _03082_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput201 o_ext_rs2[9] net201 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_3_965 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput223 o_ibus_adr[29] net223 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput212 o_ibus_adr[19] net212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput234 o_ibus_cyc net234 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06013_ rf_ram.memory\[538\]\[1\] _02208_ vss vdd rf_ram.memory\[537\]\[1\] _01539_
+ rf_ram.memory\[539\]\[1\] _01540_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__07189__A2 vss _02984_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06397__B1 vss _01772_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1253 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10193__A1 vss _05081_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06936__A2 vss _02883_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07964_ vdd _03663_ _03662_ _00494_ _03651_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08138__A1 vss _03754_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07895_ vdd vss _03621_ rf_ram.memory\[461\]\[0\] _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06915_ vdd vss _03005_ rf_ram.memory\[298\]\[0\] _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09703_ vdd vss _04779_ _04740_ net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09886__A1 vss _03892_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06846_ _02958_ _02940_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09634_ vdd _04725_ _01380_ _01102_ _04524_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05372__A1 vss _01347_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09638__A1 vss _04524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06777_ _02909_ vss vdd _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11671__I vss cpu.ctrl.pc vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09565_ vdd _04681_ _04680_ _04682_ _03992_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05728_ _01923_ vdd vss _01924_ rf_ram.memory\[440\]\[0\] _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08310__A1 vss _03852_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09496_ vdd _04630_ _01388_ _04631_ cpu.alu.cmp_r vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08516_ vdd _04018_ _04017_ _00691_ _03953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_171_clk vdd vss clknet_leaf_171_clk clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05659_ _01783_ vdd vss _01855_ rf_ram.memory\[472\]\[0\] _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08447_ vdd vss _03966_ rf_ram.memory\[176\]\[1\] _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08861__A2 vss _03559_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06872__A1 vss _02975_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08378_ vdd vss _03923_ rf_ram.memory\[186\]\[1\] _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_306 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07329_ vdd vss _03269_ rf_ram.memory\[271\]\[0\] _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06085__C1 vss _01654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10340_ vdd rf_ram.memory\[284\]\[0\] clknet_leaf_173_clk vss _00084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06624__A1 vss cpu.immdec.imm11_7\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06433__C vss _01978_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10271_ vdd rf_ram.memory\[233\]\[1\] clknet_leaf_277_clk vss _00015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_1141 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09316__I vss _03992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09629__A1 vss _04524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1168 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10239__A2 vss _03071_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07104__A2 vss _03072_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_162_clk vdd vss clknet_leaf_162_clk clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_167_995 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_494 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06863__A1 vss _02930_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05666__A2 vss _01543_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11656_ net178 vss vdd net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10607_ vdd rf_ram.memory\[316\]\[1\] clknet_leaf_154_clk vss _00351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09801__A1 vss _04840_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11587_ vdd rf_ram.memory\[208\]\[0\] clknet_leaf_300_clk vss _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_380 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10538_ vdd rf_ram.memory\[247\]\[0\] clknet_leaf_208_clk vss _00282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06615__A1 vss _02766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06091__A2 vss _01706_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10469_ vdd rf_ram.memory\[260\]\[1\] clknet_leaf_195_clk vss _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08368__A1 vss _02983_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_946 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09654__C vss _04740_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07040__A1 vss _03053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09317__C2 vss cpu.immdec.imm11_7\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06700_ vdd vss _02855_ rf_ram.memory\[523\]\[1\] _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07680_ vdd vss _03487_ rf_ram.memory\[402\]\[1\] _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07343__A2 vss _02960_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08540__A1 vss _04026_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06000__C1 vss _01540_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06631_ vdd vss _02803_ rf_ram.memory\[293\]\[0\] _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_540 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_759 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09350_ _04540_ net230 vdd vss _04546_ net229 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06562_ _02747_ vss vdd _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_48_916 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05513_ _01709_ _01508_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08301_ vdd vss _03874_ rf_ram.memory\[244\]\[1\] _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09281_ vdd vss _04503_ cpu.genblk3.csr.mcause3_0\[2\] _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_47_426 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_153_clk vdd vss clknet_leaf_153_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06854__A1 vss _02839_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_53 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05657__A2 vss _01785_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06493_ _02687_ _01373_ vdd vss _02688_ _02519_ _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08232_ vdd vss _03832_ rf_ram.memory\[531\]\[0\] _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_976 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_196 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05444_ _01640_ _01499_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_28_673 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_155 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05375_ _01506_ vdd vss _01571_ rf_ram.memory\[558\]\[0\] _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08163_ vdd vss _03789_ rf_ram.memory\[544\]\[0\] _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08094_ vdd vss _03746_ rf_ram.memory\[557\]\[0\] _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07114_ vdd vss _03134_ _02716_ _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__06606__A1 vss _02766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_164 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06534__B vss _01347_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07045_ vdd vss _03091_ rf_ram.memory\[391\]\[0\] _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1027 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10166__A1 vss _05049_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06909__A2 vss _02997_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_19__f_clk_I vss clknet_3_4_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08996_ vdd _04318_ _04316_ _00871_ _04301_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07031__A1 vss _03050_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07947_ vdd vss _03653_ rf_ram.memory\[456\]\[0\] _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05664__I vss _01563_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input34_I vss i_ibus_ack vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07878_ vdd vss _03610_ _02916_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08531__A1 vss _02794_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06829_ vdd vss _02947_ _02935_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09617_ vdd _04719_ _04717_ _01091_ _04637_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05613__B vss _01650_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09548_ _04668_ vdd vss _01073_ _04667_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06428__C vss _01860_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07098__A1 vss _02921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09087__A2 vss _03765_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_144_clk vdd vss clknet_leaf_144_clk clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11510_ vdd rf_ram.memory\[326\]\[1\] clknet_leaf_143_clk vss _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_325 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09479_ _03989_ vdd vss _04617_ cpu.bufreg.i_sh_signed net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_163_442 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06845__A1 vss _02930_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_347 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_155 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11441_ vdd cpu.mem_if.signbit clknet_leaf_233_clk vss _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_199 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11372_ _01104_ vdd vss clknet_leaf_235_clk cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08598__A1 vss _02794_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06073__A2 vss _01626_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10323_ vdd rf_ram.memory\[50\]\[1\] clknet_leaf_288_clk vss _00067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05805__C1 vss _01953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10157__A1 vss _02787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10254_ vdd vss _05122_ net249 _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10185_ vdd _05080_ _05079_ _01299_ _05078_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05574__I vss _01530_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05887__A2 vss _01918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07089__A1 vss _03087_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_135_clk vdd vss clknet_leaf_135_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08825__A2 vss _04195_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1073 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06836__A1 vss _02927_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_155 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_259 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11639_ net170 vss vdd net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_125 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08125__I vss _03692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08589__A1 vss _04058_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05160_ vdd vss _01363_ _01334_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__06064__A2 vss _01666_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09250__A2 vss cpu.bufreg.i_sh_signed vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09002__A2 vss _04303_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05811__A2 vss _01641_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1201 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08850_ vdd vss _04228_ net241 _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07801_ vdd vss _03563_ _02866_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_174_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08781_ vdd _04185_ _04183_ _00789_ _04170_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05993_ _01594_ _01950_ _02188_ vdd vss _00000_ _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_07732_ vdd _03519_ _03518_ _00406_ _03488_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07663_ vdd _03476_ _03475_ _00380_ _03455_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09561__I0 vss cpu.immdec.imm30_25\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_225 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_819 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05878__A2 vss _02046_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09402_ _04564_ net225 vdd vss _04574_ net223 _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06614_ _02788_ _02787_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_07594_ vdd vss _03434_ rf_ram.memory\[315\]\[0\] _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09333_ vdd vss _04536_ net240 _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07204__I vss _03013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_61 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_126_clk vdd vss clknet_leaf_126_clk clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06545_ _02730_ vdd vss _02731_ cpu.immdec.imm11_7\[3\] _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_47_245 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06476_ vss vdd rf_ram.memory\[31\]\[1\] _01607_ rf_ram.memory\[29\]\[1\] _01609_
+ _01633_ rf_ram.memory\[28\]\[1\] _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_29_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1037 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06827__A1 vss _02716_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09264_ _04490_ _02713_ vdd vss _00967_ _04486_ _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09195_ vdd vss _04443_ rf_ram.memory\[82\]\[0\] _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05427_ _01623_ _01605_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08215_ vdd vss _03821_ _03798_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06264__B vss _02458_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_648 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08146_ vdd vss _03778_ _02888_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_30_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05358_ _01554_ vss vdd _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09241__A2 vss _03989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05289_ vdd vss _01431_ _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08077_ vdd _03735_ _03733_ _00535_ _03724_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_1172 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_1025 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10139__A1 vss _05046_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06460__C1 vss _01655_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07028_ vdd _03078_ _03076_ _00143_ _03053_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05802__A2 vss _01989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_91 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07004__A1 vss _03050_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08979_ vdd _04308_ _04307_ _00864_ _04298_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08504__A1 vss _03956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10941_ vdd rf_ram_if.rdata0\[1\] clknet_leaf_280_clk vss _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06439__B vss _01601_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05869__A2 vss _01606_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10872_ vdd rf_ram.memory\[192\]\[0\] clknet_leaf_46_clk vss _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_217 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_1176 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_117_clk vdd vss clknet_leaf_117_clk clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_93_340 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06818__A1 vss _02930_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_965 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_659 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06174__B vss _01629_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11424_ vdd rf_ram.memory\[7\]\[1\] clknet_leaf_293_clk vss _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09768__B1 vss _04760_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_478 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07243__A1 vss _03190_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06046__A2 vss _01606_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11355_ _01087_ vdd vss clknet_leaf_259_clk cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08991__A1 vss _04301_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11286_ vdd net222 clknet_leaf_242_clk vss _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10306_ vdd rf_ram.memory\[517\]\[0\] clknet_leaf_270_clk vss _00050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10237_ vdd vss _05112_ rf_ram.memory\[208\]\[1\] _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06203__C1 vss _01811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07546__A2 vss _02889_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10168_ vdd vss _05070_ rf_ram.memory\[447\]\[0\] _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_1021 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10099_ vdd _05027_ _05025_ _01266_ _05017_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_1042 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_832 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05253__B vss cpu.mem_bytecnt\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06068__C vss net253 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_690 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09440__S vss _04593_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_108_clk vdd vss clknet_leaf_108_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_130_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06330_ _02019_ rf_ram.memory\[211\]\[1\] vdd vss _02525_ rf_ram.memory\[210\]\[1\]
+ _01804_ _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07482__A1 vss _03360_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06261_ rf_ram.memory\[418\]\[1\] _02456_ vss vdd rf_ram.memory\[417\]\[1\] _01645_
+ rf_ram.memory\[419\]\[1\] _01646_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_120_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06084__B vss _01707_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_637 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05479__I vss _01602_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09759__B1 vss _04760_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08000_ _03686_ _03685_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05212_ vdd vss _01412_ _01375_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06192_ _01860_ vdd vss _02387_ _02384_ _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_484 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1009 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1106 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05143_ _01341_ _01345_ vdd vss _01346_ _01332_ _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XANTENNA__07694__I vss _03100_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09951_ vdd _04936_ _04935_ _01209_ _04918_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08982__A1 vss net242 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08902_ vdd vss _04260_ _02916_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08734__A1 vss _04129_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09882_ vdd vss _04894_ rf_ram.memory\[229\]\[0\] _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08833_ vdd vss _04218_ rf_ram.memory\[459\]\[1\] _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05976_ _02168_ _02171_ vdd vss _02172_ _02160_ _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08764_ vdd _04175_ _04174_ _00782_ _04167_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07715_ vdd vss _03509_ _02839_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08695_ vdd vss _04132_ rf_ram.memory\[153\]\[0\] _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07646_ vdd vss _03466_ _03071_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_1126 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07577_ vdd vss _03423_ _02882_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06528_ vdd vss cpu.state.ibus_cyc _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09316_ _04526_ _03992_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07473__A1 vss _03356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_401 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09247_ vdd vss _04476_ _03967_ net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06276__A2 vss _01664_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_261 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05484__B1 vss _01678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06459_ _01525_ vdd vss _02654_ rf_ram.memory\[48\]\[1\] _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_185_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output188_I vss net188 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09178_ vdd vss _04432_ _03134_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09214__A2 vss _04418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07225__A1 vss _03193_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_264 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08129_ vdd vss _03768_ rf_ram.memory\[551\]\[1\] _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_955 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06028__A2 vss _01532_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11140_ vdd rf_ram.memory\[110\]\[0\] clknet_leaf_69_clk vss _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_865 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput67 o_dbus_adr[10] net67 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_179_1032 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11071_ vdd rf_ram.memory\[459\]\[0\] clknet_leaf_52_clk vss _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput78 o_dbus_adr[21] net78 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput89 o_dbus_adr[31] net89 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10022_ vdd vss _04980_ rf_ram.memory\[246\]\[0\] _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06200__A2 vss _01724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_810 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09150__A1 vss _04401_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_338_clk vdd vss clknet_leaf_338_clk clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_85_104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10924_ vdd rf_ram.memory\[59\]\[0\] clknet_leaf_296_clk vss _00668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10855_ vdd rf_ram.memory\[52\]\[1\] clknet_leaf_297_clk vss _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07464__A1 vss _02921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_9_clk_I vss clknet_5_0__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10786_ vdd rf_ram.memory\[563\]\[0\] clknet_leaf_329_clk vss _00530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05299__I vss _01494_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_927 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_133_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11407_ vdd rf_ram.memory\[269\]\[0\] clknet_leaf_191_clk vss _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07216__A1 vss _02883_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06019__A2 vss _01524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11338_ vdd cpu.csr_imm clknet_leaf_216_clk vss _01070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_605 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_323_clk_I vss clknet_5_4__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06351__C vss _02545_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11269_ vdd net204 clknet_leaf_246_clk vss _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08716__A1 vss _04126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_338_clk_I vss clknet_5_0__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05830_ _01551_ vdd vss _02026_ rf_ram.memory\[216\]\[0\] _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_168_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_118_99 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05762__I vss _01640_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07500_ vdd _03375_ _03374_ _00318_ _03356_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06079__B vss _01620_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09141__A1 vss net245 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_329_clk vdd vss clknet_leaf_329_clk clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05761_ _01956_ vdd vss _01957_ rf_ram.memory\[152\]\[0\] _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05692_ vdd vss _01888_ rf_ram.memory\[385\]\[0\] _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08480_ _01418_ vdd vss _03993_ _02713_ _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_07431_ vdd _03332_ _03331_ _00292_ _03323_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_3_7_0_clk_I vss clknet_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05711__B vss _01660_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_537 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07362_ vdd _03288_ _03286_ _00267_ _03260_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_169_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09101_ vdd _04383_ _04381_ _00911_ _04367_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06313_ rf_ram.memory\[189\]\[1\] _01793_ _01677_ rf_ram.memory\[188\]\[1\] _02508_
+ vss vdd rf_ram.memory\[191\]\[1\] _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__06258__A2 vss _01940_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_710 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07293_ vdd vss _03246_ rf_ram.memory\[468\]\[1\] _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06244_ _01790_ vdd vss _02439_ _02436_ _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09032_ vdd _04341_ _04340_ _00884_ _04331_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07207__A1 vss _03190_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06175_ _01504_ vdd vss _02370_ rf_ram.memory\[502\]\[1\] _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_60_549 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1061 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_240 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_284 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09934_ vdd vss _04926_ _04911_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_695 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06430__A2 vss _01863_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09865_ vdd _04883_ _04881_ _01176_ _04840_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08816_ vdd vss _04208_ rf_ram.memory\[137\]\[0\] _04207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_1060 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07930__A2 vss _03547_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09796_ vdd _04841_ _04838_ _01148_ _04840_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05959_ _02153_ _02154_ vdd vss _02155_ _02151_ _02152_ rf_ram.i_raddr\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08747_ vdd vss _04164_ net242 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08678_ vdd vss _04121_ rf_ram.memory\[559\]\[0\] _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_684 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07629_ _03455_ vss vdd _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output103_I vss net103 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06497__A2 vss _01375_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10640_ vdd rf_ram.memory\[384\]\[0\] clknet_leaf_92_clk vss _00384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_740 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_874 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_356 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07446__A1 vss _03323_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10571_ vdd rf_ram.memory\[325\]\[1\] clknet_leaf_171_clk vss _00315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06249__A2 vss _01531_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_754 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_434 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_445 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_793 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09199__A1 vss _02805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08946__A1 vss _04266_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1172 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06421__A2 vss _01799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11123_ vdd rf_ram.memory\[11\]\[1\] clknet_leaf_37_clk vss _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11054_ vdd rf_ram.memory\[141\]\[1\] clknet_leaf_9_clk vss _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1312 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10005_ vdd _04969_ _04967_ _01230_ _04953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05582__I vss _01695_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05932__A1 vss _01350_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_58_115 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07685__A1 vss _03488_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_835 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_295 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10907_ vdd rf_ram.memory\[180\]\[1\] clknet_leaf_19_clk vss _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05696__B1 vss _01773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_129 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10838_ vdd rf_ram.memory\[537\]\[0\] clknet_leaf_312_clk vss _00582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10769_ vdd rf_ram.memory\[572\]\[1\] clknet_leaf_304_clk vss _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_584 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_262_clk_I vss clknet_5_17__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_590 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_1148 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05757__I vss _01695_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_763 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06412__A2 vss _01915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07980_ vdd vss _03674_ rf_ram.memory\[478\]\[0\] _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06931_ vdd _03016_ _03015_ _00108_ _03014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_277_clk_I vss clknet_5_16__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09650_ _04737_ vss vdd _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06862_ vdd vss _02969_ rf_ram.memory\[283\]\[1\] _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1181 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05492__I vss _01624_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08601_ vdd vss _04073_ rf_ram.memory\[165\]\[1\] _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06793_ vss _02921_ _02868_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_leaf_200_clk_I vss clknet_5_25__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05813_ _02008_ _01860_ vdd vss _02009_ _02005_ _02006_ _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_59_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09581_ _04678_ _04476_ vdd vss _04694_ _03992_ _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09114__A1 vss _04364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08532_ vdd vss _04029_ rf_ram.memory\[69\]\[0\] _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05744_ _01940_ vss vdd _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07676__A1 vss _03458_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06479__A2 vss _01640_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08463_ vdd vss _03980_ _03971_ _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07414_ vdd _03321_ _03320_ _00286_ _03289_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05675_ _01869_ _01870_ vdd vss _01871_ _01867_ _01868_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA_clkbuf_leaf_215_clk_I vss clknet_5_19__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08394_ vdd _03932_ _03930_ _00655_ _03922_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07428__A1 vss _03326_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07345_ vdd _03278_ _03277_ _00260_ _03257_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_652 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07276_ vdd vss _03236_ rf_ram.memory\[417\]\[0\] _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07979__A2 vss _02917_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_220 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_30_clk vdd vss clknet_leaf_30_clk clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_941 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06227_ _02421_ vdd vss _02422_ _01603_ _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_143_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09015_ vdd vss _04330_ rf_ram.memory\[10\]\[1\] _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_195 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08928__A1 vss _04269_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_223 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05667__I vss _01633_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input64_I vss i_ibus_rdt[9] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06158_ vdd vss _02353_ rf_ram.memory\[489\]\[1\] _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07600__A1 vss _03422_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06089_ _01707_ vdd vss _02284_ rf_ram.memory\[334\]\[1\] _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06403__A2 vss _01509_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05611__B1 vss _01725_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09917_ vdd vss _04915_ _04911_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_1092 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_97_clk vdd vss clknet_leaf_97_clk clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08156__A2 vss _03765_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06167__A1 vss _01603_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09848_ _04870_ _04872_ vdd vss _04873_ cpu.ctrl.i_jump _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09779_ vdd _04830_ _04828_ _01142_ _04637_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_1029 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_470 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_180_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10623_ vdd rf_ram.memory\[407\]\[1\] clknet_leaf_102_clk vss _00367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06890__A2 vss _02801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_581 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_187_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10554_ vdd rf_ram.memory\[331\]\[0\] clknet_leaf_152_clk vss _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_21_clk vdd vss clknet_leaf_21_clk clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_load_slew254_I vss _01361_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08092__A1 vss _03724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_860 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10485_ vdd rf_ram.memory\[418\]\[1\] clknet_leaf_98_clk vss _00229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08919__A1 vss _02794_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05577__I vss _01695_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1278 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_711 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08395__A2 vss _02997_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07792__I vss _03359_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05602__B1 vss _01715_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11106_ vdd rf_ram.memory\[389\]\[0\] clknet_leaf_118_clk vss _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_88_clk vdd vss clknet_leaf_88_clk clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09344__A1 vss net224 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09344__B2 vss net227 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1175 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11037_ vdd rf_ram.i_raddr\[1\] clknet_leaf_275_clk vss _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_571 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05381__A2 vss _01538_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07658__A1 vss _03455_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05460_ vdd vss _01656_ _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_74_438 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05391_ _01506_ vdd vss _01587_ rf_ram.memory\[574\]\[0\] _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_131_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07130_ vdd _03144_ _03142_ _00179_ _03126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_12_clk vdd vss clknet_leaf_12_clk clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08083__A1 vss _03668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_549 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07830__A1 vss _03557_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07061_ vss _03101_ _03100_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_clkbuf_leaf_81_clk_I vss clknet_5_11__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05487__I vss _01682_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_699 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput224 o_ibus_adr[2] net224 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput213 o_ibus_adr[1] net213 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput202 o_ibus_adr[0] net202 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06012_ _01552_ vdd vss _02207_ rf_ram.memory\[536\]\[1\] _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_96_clk_I vss clknet_5_14__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_79_clk vdd vss clknet_leaf_79_clk clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09335__A1 vss _04463_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07963_ vdd vss _03663_ rf_ram.memory\[470\]\[0\] _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07894_ vdd vss _03620_ _02836_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06914_ vdd vss _03004_ _02775_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09702_ vdd vss _04778_ _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_179_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06845_ vdd _02957_ _02955_ _00081_ _02930_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09886__A2 vss _02822_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09633_ vdd vss _04725_ _04524_ net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09564_ vdd vss _04681_ _03992_ net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_154_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08515_ vdd vss _04018_ rf_ram.memory\[172\]\[0\] _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09638__A2 vss _01391_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_1__f_clk_I vss clknet_3_0_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06776_ vdd vss _02908_ _02779_ _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05727_ vss _01923_ _01550_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09495_ vdd vss _04630_ _01442_ _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_1035 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_654 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05658_ _01790_ vdd vss _01854_ _01851_ _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_34_clk_I vss clknet_5_6__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08446_ vdd _03965_ _03964_ _00674_ _03953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_484 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08377_ _03922_ _03689_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_169_clk_I vss clknet_5_30__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07328_ vdd vss _03268_ _02958_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05589_ _01785_ vss vdd _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_972 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06085__B1 vss _01656_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07259_ vdd _03224_ _03223_ _00228_ _03222_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07821__A1 vss _02761_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_49_clk_I vss clknet_5_12__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_757 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06624__A2 vss _02730_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05832__B1 vss _01959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output170_I vss net170 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10270_ vdd rf_ram.memory\[233\]\[0\] clknet_leaf_277_clk vss _00014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_1067 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_107_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05346__B vss _01528_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07888__A1 vss _02959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05363__A2 vss _01538_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06560__A1 vss _01369_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09629__A2 vss net55 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06177__B vss _01526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_65_961 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11655_ vss net177 net105 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05520__C1 vss _01715_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10606_ vdd rf_ram.memory\[316\]\[0\] clknet_leaf_154_clk vss _00350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11586_ vdd rf_ram.memory\[237\]\[1\] clknet_leaf_284_clk vss _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_58 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10537_ vdd rf_ram.memory\[248\]\[1\] clknet_leaf_212_clk vss _00281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06615__A2 vss _02788_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10468_ vdd rf_ram.memory\[260\]\[0\] clknet_leaf_195_clk vss _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08368__A2 vss _03903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09565__A1 vss _03992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06379__A1 vss _01768_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10399_ vdd rf_ram.memory\[218\]\[1\] clknet_leaf_302_clk vss _00143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_1_clk vdd vss clknet_leaf_1_clk clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09317__B2 vss cpu.immdec.imm11_7\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09317__A1 vss _04526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06630_ vdd vss _02802_ _02795_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06000__B1 vss _01539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06551__A1 vss _02731_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1079 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06866__I vss _02971_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_749 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06561_ vdd _02745_ rf_ram_if.wdata1_r\[1\] _02746_ _01353_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05512_ _01707_ vdd vss _01708_ rf_ram.memory\[326\]\[0\] _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06492_ _02630_ _02687_ _02603_ _01372_ _02686_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_08300_ vdd _03873_ _03872_ _00620_ _03852_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09280_ cpu.genblk3.csr.o_new_irq _01391_ vdd vss _04502_ cpu.genblk3.csr.mcause3_0\[3\]
+ _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_185_793 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05443_ _01630_ _01638_ vdd vss _01639_ _01612_ _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_144_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_524 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08231_ vdd vss _03831_ _03798_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06854__A2 vss _02941_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_657 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_460 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_96 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_999 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08162_ vdd vss _03788_ net237 _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08056__A1 vss _03134_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05374_ _01566_ _01569_ vdd vss _01570_ _01351_ _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_160_638 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07803__A1 vss _03554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07113_ vdd _03133_ _03131_ _00173_ _03126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_1153 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08093_ vdd vss _03745_ _02843_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_817 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06606__A2 vss _02781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07044_ vdd vss _03090_ _02829_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05290__A1 vss _01434_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_349 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08995_ vdd vss _04318_ rf_ram.memory\[113\]\[1\] _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05578__C1 vss _01773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07946_ vdd vss _03652_ _02728_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05593__A2 vss _01785_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06790__A1 vss _02873_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input27_I vss i_dbus_rdt[3] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07877_ vdd _03609_ _03607_ _00461_ _03590_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_817 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08531__A2 vss _04005_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08477__B vss net65 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09616_ vdd vss _04719_ rf_ram.memory\[72\]\[1\] _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05345__A2 vss _01538_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06828_ _02946_ vss vdd _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_149_941 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09547_ net43 _04650_ cpu.immdec.imm19_12_20\[7\] vdd vss _04668_ _04478_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06759_ vdd _02896_ _02895_ _00056_ _02873_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_164_900 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08295__A1 vss _03852_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07098__A2 vss _02946_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_624 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_257 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09478_ vdd _04615_ _02705_ _04616_ _02703_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_657 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_780 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08429_ vdd vss _03955_ rf_ram.memory\[59\]\[0\] _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_164_988 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_1077 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08047__A1 vss _03686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11440_ _01172_ cpu.mem_bytecnt\[1\] vdd vss clknet_leaf_241_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_132_841 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08598__A2 vss _04067_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11371_ _01103_ net134 vdd vss clknet_leaf_236_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
X_10322_ vdd rf_ram.memory\[50\]\[0\] clknet_leaf_288_clk vss _00066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_485 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05805__B1 vss _01516_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09547__A1 vss _04478_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_29__f_clk vdd vss clknet_5_29__leaf_clk clknet_3_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10157__A2 vss _02921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10253_ vdd _05121_ _05119_ _01326_ _02825_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_861 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10184_ vdd vss _05080_ rf_ram.memory\[190\]\[0\] _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05584__A2 vss _01777_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_817 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05590__I vss _01695_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06686__I vss _02845_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_513 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_500 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_785 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11638_ vss net162 net89 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_126_189 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11569_ vdd rf_ram.memory\[238\]\[0\] clknet_leaf_285_clk vss _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_485 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09438__S vss _04593_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09538__A1 vss _04526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09665__C vss _04740_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05272__A1 vss cpu.ctrl.pc vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06370__B vss _01684_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1170 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1181 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07800_ vdd _03562_ _03560_ _00431_ _03557_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08780_ vdd vss _04185_ rf_ram.memory\[142\]\[1\] _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07731_ vdd vss _03519_ rf_ram.memory\[397\]\[0\] _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05575__A2 vss _01770_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05992_ vdd vss _02188_ _01371_ _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05980__C1 vss _01653_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07662_ vdd vss _03476_ rf_ram.memory\[385\]\[0\] _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09710__A1 vss _04781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07593_ vdd vss _03433_ _02935_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09401_ vdd vss _04573_ _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06613_ vdd vss _02787_ _02716_ _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_09332_ vdd _04535_ _04533_ _00990_ _04466_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08277__A1 vss _03855_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06544_ vdd vss _02730_ _01347_ _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__10084__A1 vss _05017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_613 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06475_ vdd vss _02670_ rf_ram.memory\[30\]\[1\] _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09263_ vdd vss _04490_ _01484_ _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05426_ _01615_ vdd vss _01622_ rf_ram.memory\[360\]\[0\] _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_161_903 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09194_ vdd vss _04442_ net236 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08214_ _03820_ _03685_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_8_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08029__A1 vss _03690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_295 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06264__C vss _01569_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09777__A1 vss _04634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08145_ vdd _03777_ _03775_ _00561_ _03757_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05357_ _01552_ vdd vss _01553_ rf_ram.memory\[528\]\[0\] _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_688 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_293 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08076_ vdd vss _03735_ rf_ram.memory\[561\]\[1\] _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05288_ vdd _01485_ _01341_ cpu.o_wdata1 _01389_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_1161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06460__B1 vss _01518_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07027_ vdd vss _03078_ rf_ram.memory\[218\]\[1\] _03076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08201__A1 vss _03787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08978_ vdd vss _04308_ rf_ram.memory\[116\]\[0\] _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05566__A2 vss _01644_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07929_ vdd _03641_ _03639_ _00481_ _03622_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output133_I vss net133 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_658 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_124 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09701__A1 vss net99 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06515__A1 vss cpu.alu.i_rs1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10940_ vdd rf_ram_if.rgnt clknet_leaf_256_clk vss _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_1074 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_557 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_831 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10871_ vdd rf_ram.memory\[204\]\[1\] clknet_leaf_34_clk vss _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10075__A1 vss _04982_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_1236 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_925 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_156 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_920 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_189 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11423_ vdd rf_ram.memory\[7\]\[0\] clknet_leaf_294_clk vss _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_953 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11354_ vdd cpu.immdec.imm24_20\[4\] clknet_leaf_280_clk vss _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10305_ vdd rf_ram.memory\[518\]\[1\] clknet_leaf_268_clk vss _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11285_ vdd net221 clknet_leaf_242_clk vss _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10236_ vdd _05111_ _05110_ _01319_ _02819_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06203__B1 vss _01725_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10167_ vdd vss _05069_ _02908_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05557__A2 vss _01644_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06754__A1 vss _02876_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10098_ vdd vss _05027_ rf_ram.memory\[351\]\[1\] _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_1077 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_1055 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_1039 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_1038 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_174_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_29_224 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06260_ _01756_ vdd vss _02455_ rf_ram.memory\[416\]\[1\] _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_72_536 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09759__A1 vss net118 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05211_ _01404_ vdd vss _01411_ _01401_ _01403_ _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_0_5_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_777 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06191_ _01786_ rf_ram.memory\[475\]\[1\] vdd vss _02386_ rf_ram.memory\[474\]\[1\]
+ _01856_ _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09759__B2 vss net119 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_794 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_636 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_41_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05142_ _01337_ _01345_ _01334_ _01344_ cpu.immdec.imm24_20\[0\] vdd vss vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_09950_ vdd vss _04936_ rf_ram.memory\[337\]\[0\] _04935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08982__A2 vss _04303_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_321 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_292_clk vdd vss clknet_leaf_292_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08901_ vdd _04259_ _04257_ _00835_ _04237_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_3_3_0_clk_I vss clknet_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05796__A2 vss _01846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09931__A1 vss _04918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_12__f_clk vdd vss clknet_5_12__leaf_clk clknet_3_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_110_376 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09881_ vdd vss _04893_ _03309_ _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05548__A2 vss _01697_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08832_ vdd _04217_ _04216_ _00808_ _04202_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_1242 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05975_ _02170_ vdd vss _02171_ _01903_ _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05953__C1 vss _01655_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08763_ vdd vss _04175_ rf_ram.memory\[145\]\[0\] _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07714_ vdd _03508_ _03506_ _00399_ _03491_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08498__A1 vss _02736_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09631__S vss _04526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08694_ vdd vss _04131_ _02983_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1214 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07645_ vdd _03465_ _03463_ _00373_ _03458_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07576_ vss _03422_ _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__09998__A1 vss _04950_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10057__A1 vss _04985_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_886 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06527_ vss _02714_ _02713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09315_ vdd vss _04525_ _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06458_ rf_ram.memory\[53\]\[1\] _01655_ _01508_ rf_ram.memory\[52\]\[1\] _02653_
+ vss vdd rf_ram.memory\[55\]\[1\] _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_09246_ vdd vss _00964_ _02714_ _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06275__B vss _01956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_413 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05409_ _01605_ vss vdd _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_17_975 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09177_ _04431_ _04396_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06389_ vdd vss _02584_ rf_ram.memory\[65\]\[1\] _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_102_811 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08422__A1 vss net243 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08128_ vdd _03767_ _03766_ _00554_ _03754_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_283_clk vdd vss clknet_leaf_283_clk clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08059_ vss _03724_ _03689_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_179_1000 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11070_ vdd rf_ram.memory\[135\]\[1\] clknet_leaf_15_clk vss _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05787__A2 vss _01922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10021_ vdd vss _04979_ _03309_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput68 o_dbus_adr[11] net68 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput79 o_dbus_adr[22] net79 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06736__A1 vss _02873_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_444 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07161__A1 vss _03157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10923_ vdd rf_ram.memory\[173\]\[1\] clknet_leaf_4_clk vss _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10854_ vdd rf_ram.memory\[52\]\[0\] clknet_leaf_297_clk vss _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10048__A1 vss _03445_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_410 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_717 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06185__B vss _01693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_322 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_547 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10785_ vdd rf_ram.memory\[564\]\[1\] clknet_leaf_326_clk vss _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06121__C1 vss _01668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07464__A2 vss _02904_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_344 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08661__A1 vss _04097_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07795__I vss _03088_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07216__A2 vss _02941_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11406_ _01138_ vdd vss clknet_leaf_233_clk net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09461__I0 vss net80 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11337_ vdd cpu.immdec.imm19_12_20\[3\] clknet_leaf_217_clk vss _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_274_clk vdd vss clknet_leaf_274_clk clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05778__A2 vss _01649_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11268_ vdd net203 clknet_leaf_248_clk vss _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11199_ vdd rf_ram.memory\[87\]\[1\] clknet_leaf_49_clk vss _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10219_ vdd vss _05101_ _02996_ _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_118_45 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05935__C1 vss _01607_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_411 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05760_ vss _01956_ _01526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_178_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09141__A2 vss _04005_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05950__A2 vss _01633_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07035__I vss net235 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05691_ _01783_ vdd vss _01887_ rf_ram.memory\[384\]\[0\] _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05702__A2 vss _01614_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07430_ vdd vss _03332_ rf_ram.memory\[370\]\[0\] _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_1003 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_696 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07361_ vdd vss _03288_ rf_ram.memory\[268\]\[1\] _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_812 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_368 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09100_ vdd vss _04383_ rf_ram.memory\[96\]\[1\] _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06312_ _02004_ vdd vss _02507_ rf_ram.memory\[190\]\[1\] _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_72_322 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_210 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07292_ vdd _03245_ _03244_ _00240_ _03222_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_127_273 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09031_ vdd vss _04341_ rf_ram.memory\[106\]\[0\] _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08652__A1 vss net237 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06243_ _01857_ rf_ram.memory\[435\]\[1\] vdd vss _02438_ rf_ram.memory\[434\]\[1\]
+ _01856_ _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_26_794 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06174_ _01629_ vdd vss _02369_ _02367_ _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08404__A1 vss _03922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09452__I0 vss net76 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1040 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10211__A1 vss _05078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_978 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_265_clk vdd vss clknet_leaf_265_clk clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06966__A1 vss _03018_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05769__A2 vss _01958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09933_ vdd _04925_ _04923_ _01202_ _04921_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09864_ vdd vss _04883_ rf_ram.memory\[5\]\[1\] _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08815_ vdd vss _04207_ net249 _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06194__A2 vss _01863_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09795_ vdd vss _04841_ rf_ram.memory\[80\]\[1\] _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05941__A2 vss _01682_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05958_ rf_ram.memory\[51\]\[0\] _01653_ _01499_ rf_ram.memory\[50\]\[0\] _02154_
+ vss vdd rf_ram.memory\[49\]\[0\] _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08746_ vdd vss _00776_ _04157_ _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05889_ _01978_ vdd vss _02085_ _02082_ _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07143__A1 vss _03123_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08677_ vdd vss _04120_ _02953_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07628_ vdd _03454_ _03452_ _00367_ _03425_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08891__A1 vss _04237_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05902__B vss _01602_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1055 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07559_ vdd vss _03412_ rf_ram.memory\[358\]\[1\] _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_322 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10570_ vdd rf_ram.memory\[325\]\[0\] clknet_leaf_163_clk vss _00314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_867 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_232 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09229_ _04463_ _04396_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_17_761 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09199__A2 vss _04418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_731 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_630 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_256_clk vdd vss clknet_leaf_256_clk clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11122_ vdd rf_ram.memory\[11\]\[0\] clknet_leaf_37_clk vss _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11053_ vdd rf_ram.memory\[141\]\[0\] clknet_leaf_9_clk vss _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06709__A1 vss _02820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10004_ vdd vss _04969_ rf_ram.memory\[504\]\[1\] _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07382__A1 vss _03289_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06185__A2 vss _01782_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08882__A1 vss net240 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10906_ vdd rf_ram.memory\[180\]\[0\] clknet_leaf_19_clk vss _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09070__I vss _04057_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_508 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10837_ vdd rf_ram.memory\[538\]\[1\] clknet_leaf_314_clk vss _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08634__A1 vss _04062_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10768_ vdd rf_ram.memory\[572\]\[0\] clknet_leaf_327_clk vss _00512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_163 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10699_ vdd rf_ram.memory\[412\]\[1\] clknet_leaf_91_clk vss _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_563 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_703 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05999__A2 vss _01502_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_247_clk vdd vss clknet_leaf_247_clk clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06948__A1 vss _03014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09446__S vss _04593_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05620__A1 vss net252 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06930_ vdd vss _03016_ rf_ram.memory\[297\]\[0\] _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_180_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input1_I vss i_dbus_ack vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06861_ vdd _02968_ _02967_ _00086_ _02927_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05908__C1 vss _01931_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06176__A2 vss _01509_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08600_ vdd _04072_ _04071_ _00721_ _04058_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05923__A2 vss _01677_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05812_ rf_ram.memory\[185\]\[0\] _01848_ _01711_ rf_ram.memory\[184\]\[0\] _02008_
+ vss vdd rf_ram.memory\[187\]\[0\] _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_06792_ vdd _02920_ _02918_ _00065_ _02876_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09580_ cpu.immdec.imm7 _04691_ _04692_ vdd vss _04693_ _01391_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_0_175_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05743_ _01937_ _01938_ vdd vss _01939_ _01935_ _01936_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08531_ vdd vss _04028_ _02794_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07125__A1 vss _03126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05674_ rf_ram.memory\[457\]\[0\] _01725_ _01724_ rf_ram.memory\[456\]\[0\] _01870_
+ vss vdd rf_ram.memory\[459\]\[0\] _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08462_ vdd vss _03979_ _03972_ _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07413_ vdd vss _03321_ rf_ram.memory\[334\]\[0\] _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08393_ vdd vss _03932_ rf_ram.memory\[199\]\[1\] _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_439 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07344_ vdd vss _03278_ rf_ram.memory\[253\]\[0\] _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_804 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08625__A1 vss _02821_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07275_ vdd vss _03235_ _02899_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06226_ rf_ram.memory\[412\]\[1\] _02421_ vss vdd rf_ram.memory\[415\]\[1\] _01608_
+ rf_ram.memory\[413\]\[1\] _01702_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__06100__A2 vss _01614_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09014_ vdd _04329_ _04328_ _00878_ _04298_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_287 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_238_clk vdd vss clknet_leaf_238_clk clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09050__A1 vss _02805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06157_ _01684_ vdd vss _02352_ rf_ram.memory\[488\]\[1\] _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06088_ _02281_ _02282_ vdd vss _02283_ _02279_ _02280_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_112_983 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_90 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input57_I vss i_ibus_rdt[31] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09916_ vdd _04914_ _04912_ _01196_ _04887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_8_clk_I vss clknet_5_0__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07364__A1 vss _03055_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09847_ _01391_ vdd vss _04872_ _01382_ _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05914__A2 vss _01915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09778_ vdd vss _04830_ rf_ram.memory\[77\]\[1\] _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07116__A1 vss _02915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08729_ vss _04152_ _04077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA_output213_I vss net213 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_972 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05632__B vss _01620_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_222 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_322_clk_I vss clknet_5_4__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11671_ vss net202 cpu.ctrl.pc vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_160 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_614 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10622_ vdd rf_ram.memory\[407\]\[0\] clknet_leaf_102_clk vss _00366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_316 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_519 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_193 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10553_ vdd rf_ram.memory\[36\]\[1\] clknet_leaf_130_clk vss _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_1273 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_337_clk_I vss clknet_5_0__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1148 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10484_ vdd rf_ram.memory\[418\]\[0\] clknet_leaf_98_clk vss _00228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_229_clk vdd vss clknet_leaf_229_clk clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08919__A2 vss _03559_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_909 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05850__A1 vss _01674_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11105_ vdd rf_ram.memory\[439\]\[1\] clknet_leaf_79_clk vss _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09344__A2 vss _03991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06158__A2 vss _01626_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07355__A1 vss _03257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1154 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11036_ vdd rf_ram_if.rtrig0 clknet_leaf_278_clk vss _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05669__A1 vss _01769_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06315__C1 vss _01773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08855__A1 vss net240 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1026 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06330__A2 vss _01804_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08607__A1 vss _04062_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05390_ _01584_ _01585_ vdd vss _01586_ _01582_ _01583_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_166_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_153_850 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_461 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_450 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06094__A1 vss _01349_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_360 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07060_ vdd vss _03100_ _02764_ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_82_483 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06373__B vss _02004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08083__A2 vss _03083_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06011_ rf_ram.memory\[541\]\[1\] _01555_ _01538_ rf_ram.memory\[540\]\[1\] _02206_
+ vss vdd rf_ram.memory\[543\]\[1\] _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09032__A1 vss _04331_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput214 o_ibus_adr[20] net214 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput203 o_ibus_adr[10] net203 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput225 o_ibus_adr[30] net225 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06397__A2 vss _01711_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07962_ vdd vss _03662_ _02836_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09701_ _04768_ _04777_ vdd vss _04778_ net99 _04767_ net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_07893_ vss _03619_ _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06913_ vdd _03003_ _03001_ _00103_ _02975_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06844_ vdd vss _02957_ rf_ram.memory\[303\]\[1\] _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09632_ vss _01101_ _04724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09099__A1 vss _04364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_701 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09563_ vdd vss cpu.immdec.imm30_25\[2\] _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08514_ vdd vss _04017_ _02787_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06775_ vdd _02907_ _02905_ _00061_ _02876_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05726_ vss _01922_ _01536_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_72_1074 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09494_ _04627_ vdd vss _04629_ _01439_ _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05657_ rf_ram.memory\[467\]\[0\] _01852_ vdd vss _01853_ rf_ram.memory\[466\]\[0\]
+ _01785_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_92_214 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_1096 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08445_ vdd vss _03965_ rf_ram.memory\[176\]\[0\] _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05588_ _01783_ vdd vss _01784_ rf_ram.memory\[288\]\[0\] _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08376_ vdd _03921_ _03920_ _00648_ _03919_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_198 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07327_ vdd _03267_ _03265_ _00253_ _03260_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_563 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_541 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09271__A1 vss _01364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07258_ vdd vss _03224_ rf_ram.memory\[418\]\[0\] _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07821__A2 vss _03234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_224 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09023__A1 vss _04334_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06209_ _02403_ vdd vss _02404_ _01368_ _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07189_ vdd vss _03181_ _02836_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_881 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_1290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07893__I vss _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07585__A1 vss _03422_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06388__A2 vss _01922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_997 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_964 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07337__A1 vss _03260_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07888__A2 vss _03234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_531 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1130 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_261_clk_I vss clknet_5_17__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08837__A1 vss _04202_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05362__B vss _01505_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05520__B1 vss _01713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_828 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11654_ net176 vss vdd net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__06312__A2 vss _01641_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_276_clk_I vss clknet_5_16__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10605_ vdd rf_ram.memory\[356\]\[1\] clknet_leaf_157_clk vss _00349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_826 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_163 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_861 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_552 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11585_ vdd rf_ram.memory\[237\]\[0\] clknet_leaf_284_clk vss _01317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09262__A1 vss _01461_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10536_ vdd rf_ram.memory\[248\]\[0\] clknet_leaf_212_clk vss _00280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_1043 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10467_ vdd rf_ram.memory\[261\]\[1\] clknet_leaf_195_clk vss _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09014__A1 vss _04298_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10398_ vdd rf_ram.memory\[218\]\[0\] clknet_leaf_302_clk vss _00142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_214_clk_I vss clknet_5_19__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07328__A1 vss _02958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09317__A2 vss net64 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11019_ vdd rf_ram.memory\[154\]\[1\] clknet_leaf_330_clk vss _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_229_clk_I vss clknet_5_23__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06368__B vss _02004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06551__A2 vss _02736_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07043__I vss _03088_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06560_ vdd vss _02745_ _01369_ rf_ram_if.wdata0_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_143_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05511_ _01707_ _01503_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06491_ _02685_ vdd vss _02686_ net252 _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_173_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05442_ _01637_ vdd vss _01638_ _01527_ _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07500__A1 vss _03356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_940 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08230_ vdd _03830_ _03828_ _00593_ _03823_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_126_861 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_280 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05373_ _01569_ _01568_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08161_ vss _03787_ _03685_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__09253__A1 vss _01366_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08056__A2 vss _03693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1019 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07112_ vdd vss _03133_ rf_ram.memory\[488\]\[1\] _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08092_ vdd _03744_ _03742_ _00541_ _03724_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07043_ vss _03089_ _03088_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_141_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08994_ vdd _04317_ _04316_ _00870_ _04298_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05578__B1 vss _01772_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07945_ _03651_ _03355_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_48_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_177_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1115 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07876_ vdd vss _03609_ rf_ram.memory\[463\]\[1\] _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09615_ vdd _04718_ _04717_ _01090_ _04634_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_1136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06827_ vdd vss _02945_ _02716_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__06278__B vss _01494_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_28__f_clk_I vss clknet_3_7_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08819__A1 vss _04205_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09546_ vdd vss cpu.immdec.imm19_12_20\[8\] _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06758_ vdd vss _02896_ rf_ram.memory\[514\]\[0\] _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05709_ rf_ram.memory\[402\]\[0\] _01905_ vss vdd rf_ram.memory\[401\]\[0\] _01656_
+ rf_ram.memory\[403\]\[0\] _01763_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_65_203 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09477_ _03989_ vdd vss _04615_ _02703_ _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_164_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05910__B vss _01916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08428_ vdd vss _03954_ _02822_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_225 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06689_ vdd _02848_ _02847_ _00034_ _02820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_642 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_1260 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_175_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_135 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08359_ vdd vss _03911_ rf_ram.memory\[183\]\[0\] _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_184_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06058__A1 vss _01527_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11370_ _01102_ vdd vss clknet_leaf_235_clk cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10321_ vdd rf_ram.memory\[510\]\[1\] clknet_leaf_221_clk vss _00065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05281__A2 vss _01478_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09547__A2 vss net43 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output88_I vss net88 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07558__A1 vss _03389_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10252_ vdd vss _05121_ rf_ram.memory\[28\]\[1\] _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10183_ vdd vss _05079_ _02916_ _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05357__B vss _01552_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07730__A1 vss _02844_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_80_clk_I vss clknet_5_11__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06188__B vss _01790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1029 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_463 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_940 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_731 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_95_clk_I vss clknet_5_14__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_967 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_636 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09235__A1 vss _04466_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_228 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11637_ vss net161 net88 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11568_ vdd rf_ram.memory\[190\]\[1\] clknet_leaf_25_clk vss _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_965 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10519_ vdd rf_ram.memory\[26\]\[1\] clknet_leaf_209_clk vss _00263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11499_ vdd rf_ram.memory\[277\]\[0\] clknet_leaf_178_clk vss _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_153_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09538__A2 vss net39 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_33_clk_I vss clknet_5_6__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09454__S vss _04593_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07730_ vdd vss _03518_ _02844_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05991_ _02186_ _01373_ vdd vss _02187_ _02017_ _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_168_clk_I vss clknet_5_30__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05980__B1 vss _01714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07661_ vdd vss _03475_ net238 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_48_clk_I vss clknet_5_12__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09710__A2 vss net6 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06524__A2 vss _02709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07592_ vdd _03432_ _03430_ _00353_ _03425_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_1072 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09400_ _04564_ net223 vdd vss _04573_ net222 _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06612_ vdd vss _02786_ _02785_ _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09331_ vdd vss _04535_ rf_ram.memory\[309\]\[1\] _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06543_ vdd vss cpu.immdec.imm11_7\[4\] _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_1_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1089 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1164 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06474_ _01563_ vdd vss _02669_ _02666_ _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09262_ _04488_ vdd vss _04489_ _01461_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_106_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05425_ _01620_ vdd vss _01621_ _01616_ _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_172_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09226__A1 vss _04431_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09193_ vdd _04441_ _04439_ _00945_ _04434_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08213_ vdd _03819_ _03817_ _00587_ _03790_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_921 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_559 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08144_ vdd vss _03777_ rf_ram.memory\[548\]\[1\] _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05356_ vss _01552_ _01551_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_105_1103 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08075_ vdd _03734_ _03733_ _00534_ _03721_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05287_ vdd vss _01485_ _01341_ _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07026_ vdd _03077_ _03076_ _00142_ _03050_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05263__A2 vss _01460_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08201__A2 vss _03811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06212__A1 vss _01769_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08977_ vdd vss _04307_ _03134_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07928_ vdd vss _03641_ rf_ram.memory\[458\]\[1\] _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05905__B vss _01660_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05971__B1 vss _01624_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06787__I vss _02916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07859_ vdd vss _03599_ rf_ram.memory\[40\]\[0\] _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output126_I vss net126 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1112 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07712__A1 vss _03488_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_158 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10870_ vdd rf_ram.memory\[204\]\[0\] clknet_leaf_34_clk vss _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09529_ vdd vss _04656_ cpu.immdec.imm19_12_20\[2\] _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07411__I vss _02814_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05640__B vss _01756_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1073 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_1090 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_786 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11422_ vdd rf_ram.memory\[74\]\[1\] clknet_leaf_35_clk vss _01154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09768__A2 vss _04766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06471__B vss _01550_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11353_ _01085_ vdd vss clknet_leaf_216_clk cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_21_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_659 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10304_ vdd rf_ram.memory\[518\]\[0\] clknet_leaf_269_clk vss _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11284_ vdd net220 clknet_leaf_243_clk vss _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10235_ vdd vss _05111_ rf_ram.memory\[208\]\[0\] _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_1219 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10166_ vdd _05068_ _05066_ _01292_ _05049_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07951__A1 vss _03654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10097_ vdd _05026_ _05025_ _01265_ _05014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05534__C vss _01361_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1006 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10999_ vdd rf_ram.memory\[162\]\[1\] clknet_leaf_334_clk vss _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_556 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09208__A1 vss _04434_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_910 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_797 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05493__A2 vss _01626_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06190_ vdd vss _02385_ rf_ram.memory\[473\]\[1\] _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09759__A2 vss _04766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05210_ vdd vss _01410_ _01408_ _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05141_ _01336_ cpu.state.genblk1.misalign_trap_sync_r cpu.genblk3.csr.o_new_irq
+ vdd vss _01344_ _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__05776__I vss _01615_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_434 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xmax_cap235 net235 _03082_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09248__I vss net34 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap246 net246 _02780_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08900_ vdd vss _04259_ rf_ram.memory\[429\]\[1\] _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09880_ vdd _04892_ _04890_ _01182_ _04887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08831_ vdd vss _04217_ rf_ram.memory\[459\]\[0\] _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09392__B1 vss _04564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07942__A1 vss _03619_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05725__B vss _01790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05974_ vss vdd rf_ram.memory\[31\]\[0\] _01607_ rf_ram.memory\[29\]\[0\] _01617_
+ _01633_ rf_ram.memory\[28\]\[0\] _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__05953__B1 vss _01653_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08762_ vdd vss _04174_ _02760_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07713_ vdd vss _03508_ rf_ram.memory\[3\]\[1\] _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08498__A2 vss _02867_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_125 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09695__A1 vss net128 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08693_ vdd _04130_ _04127_ _00756_ _04129_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07644_ vdd vss _03465_ rf_ram.memory\[387\]\[1\] _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09695__B2 vss net129 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1106 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07575_ vdd _03421_ _03419_ _00347_ _03393_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_901 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06526_ _02713_ vss vdd net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_09314_ vss vdd cpu.immdec.imm11_7\[1\] _04522_ cpu.immdec.imm11_7\[2\] _04521_ net63
+ _04524_ _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__05469__C1 vss _01519_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06130__B1 vss _01778_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06457_ _01503_ vdd vss _02652_ rf_ram.memory\[54\]\[1\] _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_17_921 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_781 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09245_ _04473_ _04474_ vdd vss _04475_ cpu.genblk3.csr.o_new_irq _01413_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05408_ vdd vss _01604_ rf_ram.memory\[356\]\[0\] _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05484__A2 vss _01677_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_105 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_1035 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_233 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09176_ vdd _04430_ _04428_ _00939_ _04401_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06388_ _01551_ vdd vss _02583_ rf_ram.memory\[64\]\[1\] _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08422__A2 vss _03949_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05339_ _01506_ vdd vss _01535_ rf_ram.memory\[518\]\[0\] _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08127_ vdd vss _03767_ rf_ram.memory\[551\]\[0\] _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05619__C vss net253 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08058_ vdd _03723_ _03722_ _00528_ _03721_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05641__C1 vss _01715_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07009_ vdd _03066_ _03065_ _00136_ _03050_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10020_ vdd _04978_ _04976_ _01236_ _04953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput69 o_dbus_adr[12] net69 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08186__A1 vss _03787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_957 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10922_ vdd rf_ram.memory\[173\]\[0\] clknet_leaf_5_clk vss _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_117 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_309 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_854 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05172__A1 vss _01351_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10853_ vdd rf_ram.memory\[530\]\[1\] clknet_leaf_309_clk vss _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10048__A2 vss _02923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1095 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_887 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10784_ vdd rf_ram.memory\[564\]\[0\] clknet_leaf_325_clk vss _00528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05370__B vss _01351_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1113 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_898 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_572 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06121__B1 vss _01519_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1135 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05880__C1 vss _02019_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09610__A1 vss _04634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11405_ vdd net121 clknet_leaf_230_clk vss _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09461__I1 vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11336_ vdd cpu.immdec.imm19_12_20\[2\] clknet_leaf_218_clk vss _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_787 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11267_ _01002_ vdd vss clknet_leaf_248_clk net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08177__A1 vss _03790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07924__A1 vss _03622_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11198_ vdd rf_ram.memory\[87\]\[0\] clknet_leaf_49_clk vss _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10218_ vdd _05100_ _05098_ _01312_ _05081_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10149_ vdd _05058_ _05057_ _01285_ _05046_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05935__B1 vss _01609_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_445 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05690_ _01746_ vdd vss _01886_ _01883_ _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05163__A1 vss _01364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07360_ vdd _03287_ _03286_ _00266_ _03257_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_1101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1112 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06095__C vss _01361_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06311_ _02502_ _02505_ vdd vss _02506_ _02494_ _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_07291_ vdd vss _03245_ rf_ram.memory\[468\]\[0\] _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09030_ vdd vss _04340_ net247 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08652__A2 vss _04067_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06242_ vdd vss _02437_ rf_ram.memory\[433\]\[1\] _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__06663__A1 vss _02826_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_378 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_762 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_406 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06173_ rf_ram.memory\[507\]\[1\] _01654_ _01652_ rf_ram.memory\[506\]\[1\] _02368_
+ vss vdd rf_ram.memory\[505\]\[1\] _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09452__I1 vss net77 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09932_ vdd vss _04925_ rf_ram.memory\[341\]\[1\] _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_653 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05623__C1 vss _01679_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08168__A1 vss _02881_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07915__A1 vss _02844_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09863_ vdd _04882_ _04881_ _01175_ _04837_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05455__B vss _01650_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09794_ _04840_ _04400_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08814_ vdd _04206_ _04203_ _00801_ _04205_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08745_ vdd vss _04163_ _01495_ _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05957_ _01525_ vdd vss _02153_ rf_ram.memory\[48\]\[0\] _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09668__A1 vss net120 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05888_ rf_ram.memory\[67\]\[0\] _02083_ vdd vss _02084_ rf_ram.memory\[66\]\[0\]
+ _01804_ _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_95_415 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08340__A1 vss _03887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08676_ vdd _04119_ _04117_ _00750_ _04097_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07627_ vdd vss _03454_ rf_ram.memory\[407\]\[1\] _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05154__A1 vss _01347_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07558_ vdd _03411_ _03410_ _00340_ _03389_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06286__B vss _01923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06509_ _02696_ vdd vss _00006_ _02697_ _02698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_180_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07489_ vdd vss _03369_ rf_ram.memory\[325\]\[0\] _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_857 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_559 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09228_ vdd _04462_ _04460_ _00959_ _04434_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output193_I vss net193 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1044 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09159_ vdd _04420_ _04419_ _00932_ _04397_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_776 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11121_ vdd rf_ram.memory\[120\]\[1\] clknet_leaf_85_clk vss _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output70_I vss net70 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11052_ vdd rf_ram.memory\[142\]\[1\] clknet_leaf_6_clk vss _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10003_ vdd _04968_ _04967_ _01229_ _04950_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_1124 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09659__A1 vss net120 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1146 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_776 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08331__A1 vss _03892_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1243 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_192_clk vdd vss clknet_leaf_192_clk clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_129_506 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10905_ vdd rf_ram.memory\[186\]\[1\] clknet_leaf_19_clk vss _00649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_303 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08882__A2 vss _03547_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05696__A2 vss _01777_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10836_ vdd rf_ram.memory\[538\]\[0\] clknet_leaf_270_clk vss _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_678 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09831__A1 vss _04840_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10767_ vdd rf_ram.memory\[573\]\[1\] clknet_leaf_327_clk vss _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10698_ vdd rf_ram.memory\[412\]\[0\] clknet_leaf_91_clk vss _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_531 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1242 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_551 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11319_ _01052_ vdd vss clknet_leaf_263_clk net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09898__A1 vss _04884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06860_ vdd vss _02968_ rf_ram.memory\[283\]\[0\] _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05908__B1 vss _01911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05811_ _01916_ vdd vss _02007_ rf_ram.memory\[186\]\[0\] _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08570__A1 vss _04023_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06791_ vdd vss _02920_ rf_ram.memory\[510\]\[1\] _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05742_ rf_ram.memory\[424\]\[0\] _01938_ vss vdd rf_ram.memory\[427\]\[0\] _01811_
+ rf_ram.memory\[425\]\[0\] _01810_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_145_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08530_ vdd _04027_ _04024_ _00696_ _04026_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05673_ _01650_ vdd vss _01869_ rf_ram.memory\[458\]\[0\] _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08461_ vdd vss _03978_ cpu.bufreg2.o_sh_done_r _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_159_174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07412_ vdd vss _03320_ _03319_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05687__A2 vss _01782_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_183_clk vdd vss clknet_leaf_183_clk clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08392_ vdd _03931_ _03930_ _00654_ _03919_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_174_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09822__A1 vss _03309_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07343_ vdd vss _03277_ _03055_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08625__A2 vss _02881_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07274_ vss _03234_ _03039_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_45_356 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06225_ vdd vss _02420_ rf_ram.memory\[414\]\[1\] _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09013_ vdd vss _04329_ rf_ram.memory\[10\]\[0\] _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_570 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_50 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08389__A1 vss _03922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09425__I1 vss net94 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_951 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06156_ _02350_ vdd vss _02351_ _01675_ _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__09050__A2 vss _04339_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10196__A1 vss _05078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06087_ rf_ram.memory\[322\]\[1\] _02282_ vss vdd rf_ram.memory\[321\]\[1\] _01715_
+ rf_ram.memory\[323\]\[1\] _01654_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__05611__A2 vss _01724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09915_ vdd vss _04914_ rf_ram.memory\[344\]\[1\] _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09846_ vdd vss _04871_ _01452_ _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07364__A2 vss _02822_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09777_ vdd _04829_ _04828_ _01141_ _04634_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06989_ vdd vss _03054_ rf_ram.memory\[227\]\[1\] _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05913__B vss _01790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08728_ vdd _04151_ _04149_ _00770_ _04129_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06795__I vss _02922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_815 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07116__A2 vss _03135_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08313__A1 vss _03230_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08659_ vdd _04109_ _04108_ _00743_ _04094_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_174_clk vdd vss clknet_leaf_174_clk clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05678__A2 vss _01649_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10120__A1 vss _03008_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06875__A1 vss _02970_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11670_ net194 vss vdd net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_824 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10621_ vdd rf_ram.memory\[352\]\[1\] clknet_leaf_157_clk vss _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_941 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_846 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_339 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_222 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10552_ vdd rf_ram.memory\[36\]\[0\] clknet_leaf_205_clk vss _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_553 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_704 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06463__C vss _01568_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05835__C1 vss _02019_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10483_ vdd rf_ram.memory\[41\]\[1\] clknet_leaf_132_clk vss _00227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07052__A1 vss _03087_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05602__A2 vss _01709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11104_ vdd rf_ram.memory\[439\]\[0\] clknet_leaf_79_clk vss _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11035_ vdd rf_ram.memory\[148\]\[1\] clknet_leaf_0_clk vss _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08552__A1 vss _04026_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1207 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_165_clk vdd vss clknet_leaf_165_clk clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_157_612 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06315__B1 vss _01848_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_234 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08855__A2 vss _04195_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_976 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_645 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_678 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_306 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09804__A1 vss _04837_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10819_ vdd rf_ram.memory\[547\]\[1\] clknet_leaf_317_clk vss _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_171_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09280__A2 vss _01341_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09457__S vss _04604_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06010_ _01505_ vdd vss _02205_ rf_ram.memory\[542\]\[1\] _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05841__A2 vss _01915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput226 o_ibus_adr[31] net226 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput215 o_ibus_adr[21] net215 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput204 o_ibus_adr[11] net204 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_51_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07961_ vdd _03661_ _03659_ _00493_ _03654_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09256__I vss _01356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08791__A1 vss _04170_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06912_ vdd vss _03003_ rf_ram.memory\[27\]\[1\] _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09700_ vdd vss _04777_ _04740_ net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07892_ vdd _03618_ _03616_ _00467_ _03590_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08543__A1 vss _04023_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06843_ vdd _02956_ _02955_ _00080_ _02927_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09631_ _04526_ vdd vss _04724_ cpu.decode.opcode\[1\] net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_136_1010 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05733__B vss _01928_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06774_ vdd vss _02907_ rf_ram.memory\[512\]\[1\] _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09562_ vss _01076_ _04679_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05725_ _01790_ vdd vss _01921_ _01917_ _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08513_ vdd _04016_ _04015_ _00690_ _04009_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06548__C vss _01341_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_156_clk vdd vss clknet_leaf_156_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10102__A1 vss _05014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09493_ _04627_ vdd vss _04628_ _01439_ _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06306__B1 vss _01520_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05656_ vdd vss _01852_ rf_ram.memory\[465\]\[0\] _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08444_ vdd vss _03964_ _02945_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05587_ _01783_ vss vdd _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08375_ vdd vss _03921_ rf_ram.memory\[186\]\[0\] _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07326_ vdd vss _03267_ rf_ram.memory\[255\]\[1\] _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_131 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06085__A2 vss _01709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07282__A1 vss _03222_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05817__C1 vss _01931_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_484 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07257_ vdd vss _03223_ _02894_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1036 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10169__A1 vss _05046_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06208_ _02402_ net254 vdd vss _02403_ _01674_ _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_07188_ vdd _03180_ _03178_ _00201_ _03161_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05832__A2 vss _01940_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_573 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06139_ _02330_ _02333_ vdd vss _02334_ _02322_ _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07034__A1 vss _02779_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_781 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08782__A1 vss net243 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output156_I vss net156 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1199 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09829_ vdd _04861_ _04860_ _01161_ _04837_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05643__B vss _01504_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1007 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_147_clk vdd vss clknet_leaf_147_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_83_204 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11653_ net175 vss vdd net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10604_ vdd rf_ram.memory\[356\]\[0\] clknet_leaf_152_clk vss _00348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06474__B vss _01563_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_478 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11584_ vdd rf_ram.memory\[212\]\[1\] clknet_leaf_30_clk vss _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10535_ vdd rf_ram.memory\[265\]\[1\] clknet_leaf_140_clk vss _00279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06076__A2 vss _01692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_586 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07273__A1 vss _03225_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_134 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10466_ vdd rf_ram.memory\[261\]\[0\] clknet_leaf_138_clk vss _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_589 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_729 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10397_ vdd rf_ram.memory\[245\]\[1\] clknet_leaf_214_clk vss _00141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07328__A2 vss _02954_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08525__A1 vss net248 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11018_ vdd rf_ram.memory\[154\]\[0\] clknet_leaf_329_clk vss _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06000__A2 vss _01538_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_910 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_138_clk vdd vss clknet_leaf_138_clk clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05510_ _01706_ vss vdd _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06490_ _02684_ net254 vdd vss _02685_ _01349_ _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06839__A1 vss _02779_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05441_ vss vdd rf_ram.memory\[367\]\[0\] _01636_ rf_ram.memory\[365\]\[0\] _01610_
+ _01634_ rf_ram.memory\[364\]\[0\] _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_158_976 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_173_968 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06384__B vss _01551_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08160_ vdd _03786_ _03784_ _00567_ _03757_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_172_445 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07111_ vdd _03132_ _03131_ _00172_ _03123_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05372_ _01567_ vdd vss _01347_ _01568_ cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XANTENNA_clkbuf_leaf_7_clk_I vss clknet_5_0__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09253__A2 vss _01418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08091_ vdd vss _03744_ rf_ram.memory\[558\]\[1\] _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_310_clk vdd vss clknet_leaf_310_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07042_ vdd vss _03088_ _02830_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__05814__A2 vss _01631_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1199 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_307 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_156 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05728__B vss _01923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07016__A1 vss _03053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_321_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08764__A1 vss _04167_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08993_ vdd vss _04317_ rf_ram.memory\[113\]\[0\] _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07944_ vdd _03650_ _03648_ _00487_ _03622_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_1007 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07875_ vdd _03608_ _03607_ _00460_ _03587_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08516__A1 vss _03953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05463__B vss _01658_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06826_ vdd _02944_ _02942_ _00075_ _02930_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09614_ vdd vss _04718_ rf_ram.memory\[72\]\[0\] _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_336_clk_I vss clknet_5_0__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_228 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05750__A1 vss _01350_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_921 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_129_clk vdd vss clknet_leaf_129_clk clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_532 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09545_ _04666_ vdd vss _01072_ _01595_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06757_ vdd vss _02895_ _02881_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05708_ _01903_ vdd vss _01904_ rf_ram.memory\[400\]\[0\] _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_148_442 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06688_ vdd vss _02848_ rf_ram.memory\[525\]\[0\] _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09476_ vss _01055_ _04614_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_784 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_998 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05639_ _01834_ vdd vss _01835_ _01527_ _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08427_ _03953_ vss vdd _03685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_108_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06294__B vss _01928_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_467 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_618 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08358_ vdd vss _03910_ net235 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07309_ vdd vss _03256_ rf_ram.memory\[257\]\[1\] _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07255__A1 vss _03193_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08289_ vdd vss _03867_ rf_ram.memory\[192\]\[0\] _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_301_clk vdd vss clknet_leaf_301_clk clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10320_ vdd rf_ram.memory\[510\]\[0\] clknet_leaf_211_clk vss _00064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05805__A2 vss _01692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_679 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10251_ vdd _05120_ _05119_ _01325_ _02819_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07007__A1 vss _02738_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08755__A1 vss _04167_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10182_ _05078_ _02742_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_156_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09180__A1 vss _04431_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_587 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_261 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_535 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06297__A2 vss _01523_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05820__C vss _01569_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_765 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11636_ vss net159 net86 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06049__A2 vss _01617_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07246__A1 vss _02882_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_938 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11567_ vdd rf_ram.memory\[190\]\[0\] clknet_leaf_24_clk vss _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08994__A1 vss _04298_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10518_ vdd rf_ram.memory\[26\]\[0\] clknet_leaf_211_clk vss _00262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_898 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11498_ vdd rf_ram.memory\[504\]\[1\] clknet_leaf_185_clk vss _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10449_ vdd rf_ram.memory\[483\]\[1\] clknet_leaf_186_clk vss _00193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08746__A1 vss _04157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06221__A2 vss _01846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05990_ _02129_ _02186_ _02102_ _01372_ _02185_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__09171__A1 vss _04401_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06379__B vss _02573_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07660_ vdd _03474_ _03472_ _00379_ _03458_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07591_ vdd vss _03432_ rf_ram.memory\[355\]\[1\] _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_172_1040 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_217 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06611_ vdd vss _02785_ _02717_ _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09330_ vdd _04534_ _04533_ _00989_ _04463_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_153_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_53 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06542_ _02728_ _02727_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07485__A1 vss _03356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1007 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09261_ cpu.decode.co_ebreak _01460_ vdd vss _04488_ cpu.mem_bytecnt\[1\] _01385_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_06473_ _01624_ rf_ram.memory\[27\]\[1\] vdd vss _02668_ rf_ram.memory\[26\]\[1\]
+ _01686_ _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_30_1029 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08212_ vdd vss _03819_ rf_ram.memory\[535\]\[1\] _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09192_ vdd vss _04441_ rf_ram.memory\[83\]\[1\] _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05424_ _01620_ _01493_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_56_793 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05355_ _01551_ _01550_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08143_ vdd _03776_ _03775_ _00560_ _03754_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_240 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08074_ vdd vss _03734_ rf_ram.memory\[561\]\[0\] _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05286_ _01480_ vdd vss _01484_ _01468_ _01481_ _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_07025_ vdd vss _03077_ rf_ram.memory\[218\]\[0\] _03076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_260_clk_I vss clknet_5_17__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1006 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06460__A2 vss _01499_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08737__A1 vss _01369_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_194 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1196 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1147 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08976_ vdd _04306_ _04304_ _00863_ _04301_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input32_I vss i_dbus_rdt[8] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_275_clk_I vss clknet_5_16__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07927_ vdd _03640_ _03639_ _00480_ _03619_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09162__A1 vss net235 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07858_ vdd vss _03598_ _02728_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_78_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_515 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07789_ vdd vss _03555_ _03039_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06809_ vdd vss _02933_ rf_ram.memory\[290\]\[0\] _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_1211 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output119_I vss net119 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09528_ _04651_ _04655_ vdd vss _01066_ _04646_ _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_213_clk_I vss clknet_5_19__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09459_ _04604_ vdd vss _04606_ net79 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06279__A2 vss _01523_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07228__A1 vss _03190_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_106 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11421_ vdd rf_ram.memory\[74\]\[0\] clknet_leaf_24_clk vss _01153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08976__A1 vss _04301_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11352_ vdd cpu.immdec.imm24_20\[2\] clknet_leaf_280_clk vss _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_228_clk_I vss clknet_5_23__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10303_ vdd rf_ram.memory\[51\]\[1\] clknet_leaf_286_clk vss _00047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06451__A2 vss _01530_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11283_ vdd net219 clknet_leaf_243_clk vss _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08728__A1 vss _04129_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10234_ vdd vss _05110_ _02737_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10165_ vdd vss _05068_ rf_ram.memory\[448\]\[1\] _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06203__A2 vss _01724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07400__A1 vss _03292_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10096_ vdd vss _05026_ rf_ram.memory\[351\]\[0\] _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06199__B vss _01650_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09153__A1 vss _04397_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1080 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1091 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_504 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10998_ vdd rf_ram.memory\[162\]\[0\] clknet_leaf_334_clk vss _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_793 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_264 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11619_ vss net141 net69 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_167_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08967__A1 vss _04298_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06427__C1 vss _01679_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1103 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05140_ _01342_ vdd vss _01343_ cpu.decode.co_mem_word cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_52_251 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_616 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_476 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_695 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap247 net247 _02774_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_40_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xmax_cap236 net236 _02922_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_110_345 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08719__A1 vss _02983_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09465__S vss _04604_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08830_ vdd vss _04216_ net246 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05973_ vdd vss _02169_ rf_ram.memory\[30\]\[0\] _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08761_ vdd _04173_ _04009_ _00781_ _04172_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_174_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07712_ vdd _03507_ _03506_ _00398_ _03488_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08692_ vdd vss _04130_ rf_ram.memory\[154\]\[1\] _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07643_ vdd _03464_ _03463_ _00372_ _03455_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05741__B vss _01756_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07574_ vdd vss _03421_ rf_ram.memory\[317\]\[1\] _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09313_ _04524_ vss vdd _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__07458__A1 vss _03326_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06525_ vss net97 _02712_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05469__B1 vss _01664_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_60_clk vdd vss clknet_leaf_60_clk clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06456_ _01562_ vdd vss _02651_ _02649_ _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09244_ vdd vss cpu.genblk3.csr.timer_irq_r _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05407_ _01603_ vss vdd _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_145_275 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09175_ vdd vss _04430_ rf_ram.memory\[85\]\[1\] _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08958__A1 vss _04269_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06387_ _01928_ vdd vss _02582_ _02579_ _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_465 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08126_ vdd vss _03766_ _02829_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05338_ _01529_ _01533_ vdd vss _01534_ _01507_ _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_273 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07630__A1 vss _02882_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1258 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08057_ vdd vss _03723_ rf_ram.memory\[564\]\[0\] _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05269_ _01459_ _01463_ cpu.genblk3.csr.mstatus_mie _01467_ vdd vss _01468_ _01363_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__05641__B1 vss _01654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_334 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07008_ vdd vss _03066_ rf_ram.memory\[223\]\[0\] _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_94_clk_I vss clknet_5_14__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08959_ vdd vss _04295_ net246 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_1007 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09135__A1 vss _04401_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_802 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07697__A1 vss _03488_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10921_ vdd rf_ram.memory\[29\]\[1\] clknet_leaf_206_clk vss _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_1041 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_12__f_clk_I vss clknet_3_3_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05172__A2 vss _01362_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10852_ vdd rf_ram.memory\[530\]\[0\] clknet_leaf_308_clk vss _00596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_152_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07449__A1 vss _02946_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1182 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10783_ vdd rf_ram.memory\[565\]\[1\] clknet_leaf_326_clk vss _00527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_186_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_164_540 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_51_clk vdd vss clknet_leaf_51_clk clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_32_clk_I vss clknet_5_6__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_167_clk_I vss clknet_5_30__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08949__A1 vss _02983_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05880__B1 vss _01912_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11404_ _01136_ vdd vss clknet_leaf_231_clk net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_23_958 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07621__A1 vss _03422_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06424__A2 vss _01641_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_47_clk_I vss clknet_5_12__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11335_ vdd cpu.immdec.imm19_12_20\[1\] clknet_leaf_217_clk vss _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11266_ _01001_ vdd vss clknet_leaf_247_clk net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10217_ vdd vss _05100_ rf_ram.memory\[207\]\[1\] _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11197_ vdd rf_ram.memory\[88\]\[1\] clknet_leaf_58_clk vss _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05826__B vss _01551_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10148_ vdd vss _05058_ rf_ram.memory\[451\]\[0\] _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_105_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10079_ vdd vss _05015_ _02814_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09126__A1 vss _04397_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07688__A1 vss _03491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_356 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_345 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05561__B vss _01756_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07290_ vdd vss _03244_ _02836_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_1049 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_220 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_42_clk vdd vss clknet_leaf_42_clk clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06310_ _02504_ vdd vss _02505_ _01552_ _02503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_143_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06241_ _01916_ vdd vss _02436_ rf_ram.memory\[432\]\[1\] _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_84_195 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07860__A1 vss _03587_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06172_ _01756_ vdd vss _02367_ rf_ram.memory\[504\]\[1\] _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07612__A1 vss _03425_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09931_ vdd _04924_ _04923_ _01201_ _04918_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05623__B1 vss _01793_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_874 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08168__A2 vss _02909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09862_ vdd vss _04882_ rf_ram.memory\[5\]\[0\] _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07915__A2 vss _02869_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09793_ vdd _04839_ _04838_ _01147_ _04837_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08813_ vdd vss _04206_ rf_ram.memory\[138\]\[1\] _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05387__C1 vss _01554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05956_ rf_ram.memory\[52\]\[0\] _02152_ vss vdd rf_ram.memory\[55\]\[0\] _01518_
+ rf_ram.memory\[53\]\[0\] _01655_ _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_08744_ vdd vss _00775_ _04157_ _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09117__A1 vss _02908_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07679__A1 vss _03455_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05887_ vdd vss _02083_ rf_ram.memory\[65\]\[0\] _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08675_ vdd vss _04119_ rf_ram.memory\[156\]\[1\] _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07626_ vdd _03453_ _03452_ _00366_ _03422_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05471__B vss _01526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05154__A2 vss _01356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07557_ vdd vss _03411_ rf_ram.memory\[358\]\[0\] _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_518 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_33_clk vdd vss clknet_leaf_33_clk clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_36_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06508_ _01423_ _01398_ vdd vss _02698_ _01412_ _01383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_48_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_365 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07488_ vdd vss _03368_ _02795_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09227_ vdd vss _04462_ rf_ram.memory\[339\]\[1\] _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06439_ _01601_ vdd vss _02634_ rf_ram.memory\[40\]\[1\] _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_91_677 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output186_I vss net186 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09158_ vdd vss _04420_ rf_ram.memory\[88\]\[0\] _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07603__A1 vss _02935_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1078 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08109_ vdd vss _03755_ net247 _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09089_ vdd _04376_ _04375_ _00906_ _04364_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11120_ vdd rf_ram.memory\[120\]\[0\] clknet_leaf_86_clk vss _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_1218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11051_ vdd rf_ram.memory\[142\]\[0\] clknet_leaf_7_clk vss _00788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10002_ vdd vss _04968_ rf_ram.memory\[504\]\[0\] _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07417__I vss _03013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05378__C1 vss _01517_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05393__A2 vss _01524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06590__A1 vss _02752_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1173 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10904_ vdd rf_ram.memory\[186\]\[0\] clknet_leaf_20_clk vss _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06342__A1 vss _01972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08331__A2 vss _02984_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10835_ vdd rf_ram.memory\[53\]\[1\] clknet_leaf_285_clk vss _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_1179 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_220 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_24_clk vdd vss clknet_leaf_24_clk clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_140 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08095__A1 vss _03721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_869 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_549 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10766_ vdd rf_ram.memory\[573\]\[0\] clknet_leaf_327_clk vss _00510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07842__A1 vss _02953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10697_ vdd rf_ram.memory\[433\]\[1\] clknet_leaf_82_clk vss _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_275 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_1129 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_289 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_928 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11318_ _01051_ vdd vss clknet_leaf_263_clk net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_26_1259 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11249_ _00985_ cpu.immdec.imm11_7\[3\] vdd vss clknet_leaf_279_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_98_1095 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05810_ rf_ram.memory\[189\]\[0\] _01793_ _01677_ rf_ram.memory\[188\]\[0\] _02006_
+ vss vdd rf_ram.memory\[191\]\[0\] _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_59_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06790_ vdd _02919_ _02918_ _00064_ _02873_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05741_ _01756_ vdd vss _01937_ rf_ram.memory\[426\]\[0\] _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_171_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06387__B vss _01928_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05672_ rf_ram.memory\[461\]\[0\] _01721_ _01709_ rf_ram.memory\[460\]\[0\] _01868_
+ vss vdd rf_ram.memory\[463\]\[0\] _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_89_287 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08460_ vdd vss _03977_ net124 _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_187_484 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07411_ vss _03319_ _02814_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_08391_ vdd vss _03931_ rf_ram.memory\[199\]\[0\] _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05541__C1 vss _01678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07342_ vdd _03276_ _03274_ _00259_ _03260_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_15_clk vdd vss clknet_leaf_15_clk clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_169_1045 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09822__A2 vss _02984_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_86 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07833__A1 vss _03554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07273_ vdd _03233_ _03231_ _00233_ _03225_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_305 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_955 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06224_ _02415_ _02418_ vdd vss _02419_ _02407_ _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_09012_ vdd vss _04328_ _02774_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_896 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06155_ rf_ram.memory\[493\]\[1\] _01678_ _01677_ rf_ram.memory\[492\]\[1\] _02350_
+ vss vdd rf_ram.memory\[495\]\[1\] _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09586__A1 vss net134 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_999 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05310__I vss _01505_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_799 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06086_ _01602_ vdd vss _02281_ rf_ram.memory\[320\]\[1\] _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09914_ vdd _04913_ _04912_ _01195_ _04884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09338__A1 vss net65 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1061 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_1102 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09845_ vdd vss _04870_ _01413_ _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08010__A1 vss _02959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09776_ vdd vss _04829_ rf_ram.memory\[77\]\[0\] _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06988_ _03053_ _03017_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05375__A2 vss _01502_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05939_ rf_ram.memory\[43\]\[0\] _02134_ vdd vss _02135_ rf_ram.memory\[42\]\[0\]
+ _01605_ _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08727_ vdd vss _04151_ rf_ram.memory\[14\]\[1\] _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_405 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08658_ vdd vss _04109_ rf_ram.memory\[15\]\[0\] _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08313__A2 vss _02839_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06324__A1 vss net251 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07609_ vdd vss _03443_ rf_ram.memory\[353\]\[0\] _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10120__A2 vss _03547_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output101_I vss net101 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08589_ vdd _04065_ _04064_ _00717_ _04058_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10620_ vdd rf_ram.memory\[352\]\[0\] clknet_leaf_158_clk vss _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08077__A1 vss _03724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10551_ vdd rf_ram.memory\[332\]\[1\] clknet_leaf_165_clk vss _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06627__A2 vss cpu.immdec.imm11_7\[4\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10482_ vdd rf_ram.memory\[41\]\[0\] clknet_leaf_132_clk vss _00226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05835__B1 vss _01968_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11103_ vdd rf_ram.memory\[125\]\[1\] clknet_leaf_83_clk vss _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08001__A1 vss _02761_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11034_ vdd rf_ram.memory\[148\]\[0\] clknet_leaf_0_clk vss _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_1219 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09501__A1 vss _03445_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_224 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_443 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10818_ vdd rf_ram.memory\[547\]\[0\] clknet_leaf_317_clk vss _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08068__A1 vss net236 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07815__A1 vss _03557_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_510 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10749_ vdd rf_ram.memory\[480\]\[1\] clknet_leaf_186_clk vss _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_828 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_165 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09568__A1 vss _03992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput205 o_ibus_adr[12] net205 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput216 o_ibus_adr[22] net216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_26_1023 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput227 o_ibus_adr[3] net227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_26_1034 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08240__A1 vss _03823_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07960_ vdd vss _03661_ rf_ram.memory\[480\]\[1\] _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06911_ vdd _03002_ _03001_ _00102_ _02970_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_4_clk vdd vss clknet_leaf_4_clk clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09473__S vss _04604_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07891_ vdd vss _03618_ rf_ram.memory\[445\]\[1\] _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06842_ vdd vss _02956_ rf_ram.memory\[303\]\[0\] _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06554__A1 vss _01369_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05357__A2 vss _01511_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06896__I vss _02991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09630_ vdd _04723_ _01382_ _01100_ _04643_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06773_ vdd _02906_ _02905_ _00060_ _02873_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09561_ _04678_ vdd vss _04679_ cpu.immdec.imm30_25\[0\] _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05724_ _01911_ rf_ram.memory\[435\]\[0\] vdd vss _01920_ rf_ram.memory\[434\]\[0\]
+ _01856_ _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_136_1044 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08512_ vdd vss _04016_ _01353_ rf_ram_if.wen0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_246 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05305__I vss _01500_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09492_ vdd vss _04627_ _01490_ _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__05514__C1 vss _01654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05655_ _01693_ vdd vss _01851_ rf_ram.memory\[464\]\[0\] _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08443_ vdd _03963_ _03961_ _00673_ _03956_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_476 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05586_ _01782_ _01682_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_92_238 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08374_ vdd vss _03920_ net245 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07806__A1 vss _02916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07325_ vdd _03266_ _03265_ _00252_ _03257_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_964 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_18__f_clk vdd vss clknet_5_18__leaf_clk clknet_3_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07256_ _03222_ _03013_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05817__B1 vss _01911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_614 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06207_ _02401_ vdd vss _02402_ _01350_ _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09559__A1 vss _01491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1015 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07187_ vdd vss _03180_ rf_ram.memory\[198\]\[1\] _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_861 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06138_ _02332_ vdd vss _02333_ _01675_ _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_input62_I vss i_ibus_rdt[7] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08231__A1 vss _03798_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06069_ vdd vss _02264_ rf_ram.memory\[350\]\[1\] _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08782__A2 vss _04152_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05596__A2 vss _01735_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05924__B vss _01783_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09828_ vdd vss _04861_ rf_ram.memory\[62\]\[0\] _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06545__A1 vss cpu.immdec.imm11_7\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_1242 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09759_ _04760_ _04817_ vdd vss _04818_ net118 _04766_ net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__08298__A1 vss _03309_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_955 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05520__A2 vss _01652_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11652_ vss net174 net102 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_182_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10603_ vdd rf_ram.memory\[317\]\[1\] clknet_leaf_154_clk vss _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_143 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11583_ vdd rf_ram.memory\[212\]\[0\] clknet_leaf_30_clk vss _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10534_ vdd rf_ram.memory\[265\]\[0\] clknet_leaf_140_clk vss _00278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_1202 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_513 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10465_ vdd rf_ram.memory\[262\]\[1\] clknet_leaf_196_clk vss _00209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10396_ vdd rf_ram.memory\[245\]\[0\] clknet_leaf_214_clk vss _00140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05818__C vss _01978_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06784__A1 vss _02876_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09722__A1 vss net105 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08525__A2 vss _02869_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05339__A2 vss _01502_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11017_ vdd rf_ram.memory\[155\]\[1\] clknet_leaf_332_clk vss _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_224 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_785 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05440_ _01636_ _01635_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_172_424 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09789__A1 vss _04637_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05371_ vdd vss _01567_ _01355_ _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_51_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_88 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1026 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07110_ vdd vss _03132_ rf_ram.memory\[488\]\[0\] _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_55_496 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_176 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_885 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08090_ vdd _03743_ _03742_ _00540_ _03721_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07041_ _03087_ _03013_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_23_360 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08213__A1 vss _03790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09961__A1 vss _04918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10020__A1 vss _04953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08992_ vdd vss _04316_ net248 _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05578__A2 vss _01711_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1043 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06775__A1 vss _02876_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07943_ vdd vss _03650_ rf_ram.memory\[43\]\[1\] _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05983__C1 vss _01635_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_85 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07874_ vdd vss _03608_ rf_ram.memory\[463\]\[0\] _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09713__A1 vss _04781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06825_ vdd vss _02944_ rf_ram.memory\[287\]\[1\] _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09613_ vdd vss _04717_ net250 _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_1247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09544_ net42 _04650_ cpu.immdec.imm19_12_20\[6\] vdd vss _04666_ _04478_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06756_ _02894_ vss vdd _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10087__A1 vss _05014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05707_ _01903_ _01525_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06687_ vdd vss _02847_ _02844_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09475_ _04604_ vdd vss _04614_ net88 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_136_616 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_1161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05638_ rf_ram.memory\[509\]\[0\] _01610_ _01644_ rf_ram.memory\[508\]\[0\] _01834_
+ vss vdd rf_ram.memory\[511\]\[0\] _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08426_ vdd _03952_ _03950_ _00667_ _03922_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05502__A2 vss _01697_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_649 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_441 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_90 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05569_ _01762_ _01764_ vdd vss _01765_ _01760_ _01761_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_110_1069 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08357_ vdd _03909_ _03907_ _00641_ _03887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_150_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_800 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07308_ vdd _03255_ _03254_ _00246_ _03222_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08288_ vdd vss _03866_ _03230_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_1199 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08452__A1 vss _01369_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07239_ vdd vss _03212_ rf_ram.memory\[422\]\[1\] _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_833 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_395 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_179 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05266__A1 vss _01409_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10250_ vdd vss _05120_ rf_ram.memory\[28\]\[0\] _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07007__A2 vss _02909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08204__A1 vss _03798_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06215__B1 vss _01778_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10011__A1 vss _04911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_398 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10181_ vdd _05077_ _05075_ _01298_ _05049_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06766__A1 vss _02873_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05974__C1 vss _01607_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09704__B2 vss net101 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07191__A1 vss _03157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05741__A2 vss _01808_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_897 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_763 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11635_ vss net158 net85 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_181_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07246__A2 vss _03040_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11566_ vdd rf_ram.memory\[202\]\[1\] clknet_leaf_36_clk vss _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08443__A1 vss _03956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1010 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_855 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10517_ vdd rf_ram.memory\[253\]\[1\] clknet_leaf_218_clk vss _00261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05829__B vss _01978_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_477 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11497_ vdd rf_ram.memory\[504\]\[0\] clknet_leaf_186_clk vss _01229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_376 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10448_ vdd rf_ram.memory\[483\]\[0\] clknet_leaf_197_clk vss _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10379_ vdd rf_ram.memory\[428\]\[1\] clknet_leaf_99_clk vss _00123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09943__A1 vss _04921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06757__A1 vss _02881_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05564__B vss _01504_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05980__A2 vss _01643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06379__C vss _01569_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05717__C1 vss _01912_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07590_ vdd _03431_ _03430_ _00352_ _03422_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_853 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06610_ vdd _02784_ _02782_ _00019_ _02748_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_730 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06541_ vdd vss _02727_ _02716_ _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_06472_ vdd vss _02667_ rf_ram.memory\[25\]\[1\] _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09260_ vdd vss _04487_ cpu.state.cnt_r\[3\] cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05423_ _01608_ rf_ram.memory\[355\]\[0\] vdd vss _01619_ rf_ram.memory\[354\]\[0\]
+ _01606_ _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_146_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08211_ vdd _03818_ _03817_ _00586_ _03787_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08682__A1 vss _02821_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_975 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_435 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09191_ vdd _04440_ _04439_ _00944_ _04431_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_517 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_260 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_474 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_411 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_788 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05354_ _01550_ _01525_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08434__A1 vss _02971_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08142_ vdd vss _03776_ rf_ram.memory\[548\]\[0\] _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05739__B vss _01805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06445__B1 vss _01607_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_295_clk vdd vss clknet_leaf_295_clk clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05285_ vdd vss _01483_ _01405_ _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10241__A1 vss _02819_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08073_ vdd vss _03733_ _02761_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_285 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07024_ vdd vss _03076_ _02738_ _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06996__A1 vss _03053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05263__A4 vss _01461_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09934__A1 vss _04911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06748__A1 vss _02779_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08737__A2 vss _04157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08975_ vdd vss _04306_ rf_ram.memory\[117\]\[1\] _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05956__C1 vss _01518_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07926_ vdd vss _03640_ rf_ram.memory\[458\]\[0\] _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input25_I vss i_dbus_rdt[30] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09162__A2 vss _04418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05971__A2 vss _01686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07857_ vdd _03597_ _03595_ _00453_ _03590_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07173__A1 vss _03161_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_617 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07788_ _03554_ vss vdd _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__05723__A2 vss _01918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06808_ vdd vss _02932_ _02801_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06920__A1 vss _02773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05921__C vss _01660_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09527_ vdd vss _04655_ cpu.immdec.imm19_12_20\[1\] _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06739_ vss _02881_ _02845_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_38_216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09458_ vss _01046_ _04605_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_901 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1032 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08409_ vdd _03941_ _03939_ _00661_ _03922_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09389_ vdd vss _04567_ _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_35_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_660 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11420_ vdd rf_ram.memory\[75\]\[1\] clknet_leaf_24_clk vss _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_693 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05239__A1 vss _01434_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_286_clk vdd vss clknet_leaf_286_clk clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_50_915 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11351_ vdd cpu.immdec.imm24_20\[1\] clknet_leaf_258_clk vss _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10302_ vdd rf_ram.memory\[51\]\[0\] clknet_leaf_286_clk vss _00046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06987__A1 vss _03050_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11282_ vdd net218 clknet_leaf_244_clk vss _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09925__A1 vss _04918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10233_ vdd _05109_ _05107_ _01318_ _05081_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_683 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10164_ vdd _05067_ _05066_ _01291_ _05046_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10095_ vdd vss _05025_ _02814_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05962__A2 vss _01536_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_6_clk_I vss clknet_5_2__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__S vss _03967_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07164__A1 vss _02889_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08900__A2 vss _04257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_210_clk vdd vss clknet_leaf_210_clk clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05714__A2 vss _01510_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_650 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06911__A1 vss _02970_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_300 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10997_ vdd rf_ram.memory\[549\]\[1\] clknet_leaf_308_clk vss _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_193 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_320_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08664__A1 vss _04094_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_761 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08416__A1 vss _02959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11618_ vss net140 net68 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06427__B1 vss _01793_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10223__A1 vss _05081_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_277_clk vdd vss clknet_leaf_277_clk clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06978__A1 vss _03018_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11549_ vdd rf_ram.memory\[453\]\[0\] clknet_leaf_122_clk vss _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_994 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_674 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1148 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05278__C vss _01366_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmax_cap237 net237 _02903_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xmax_cap248 net248 _02760_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09916__A1 vss _04887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08719__A2 vss _04005_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05402__A1 vss _01347_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05972_ _01563_ vdd vss _02168_ _02165_ _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05953__A2 vss _01661_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09481__S vss _01411_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08760_ vdd vss _04173_ _01353_ rf_ram_if.wen1_r vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07155__A1 vss _03157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07711_ vdd vss _03507_ rf_ram.memory\[3\]\[0\] _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08691_ _04129_ _04061_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07642_ vdd vss _03464_ rf_ram.memory\[387\]\[0\] _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_201_clk vdd vss clknet_leaf_201_clk clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_75_1266 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05705__A2 vss _01623_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06902__A1 vss _02867_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07573_ vdd _03420_ _03419_ _00346_ _03389_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_368 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_508 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09312_ _02721_ _04523_ vdd vss _00982_ _04520_ _04521_ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__05313__I vss _01508_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06524_ _02710_ _02711_ vdd vss _02712_ cpu.state.init_done _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__06130__A2 vss _01777_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_958 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06455_ rf_ram.memory\[59\]\[1\] _01653_ _01661_ rf_ram.memory\[58\]\[1\] _02650_
+ vss vdd rf_ram.memory\[57\]\[1\] _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_17_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09243_ vdd vss _04473_ _04471_ _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09174_ vdd _04429_ _04428_ _00938_ _04397_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05406_ _01602_ _01601_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08407__A1 vss _03919_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06386_ _01925_ rf_ram.memory\[75\]\[1\] vdd vss _02581_ rf_ram.memory\[74\]\[1\]
+ _01808_ _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_17_967 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06418__B1 vss _01911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10214__A1 vss _03892_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05337_ rf_ram.memory\[523\]\[0\] _01521_ _01532_ rf_ram.memory\[522\]\[0\] _01533_
+ vss vdd rf_ram.memory\[521\]\[0\] _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
Xclkbuf_leaf_268_clk vdd vss clknet_leaf_268_clk clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08125_ _03765_ _03692_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_43_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06969__A1 vss _02788_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_414 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07630__A2 vss _03089_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05268_ vdd vss _01467_ _01465_ _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08056_ vdd vss _03722_ _03134_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07007_ vdd vss _03065_ _02738_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05199_ _01399_ cpu.decode.opcode\[2\] vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_12_683 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_661 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07394__A1 vss _03292_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06197__A2 vss _01719_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08958_ vdd _04294_ _04292_ _00857_ _04269_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_904 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08889_ vdd _04252_ _04251_ _00830_ _04234_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07909_ vdd _03629_ _03627_ _00473_ _03622_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07146__A1 vss _02761_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10920_ vdd rf_ram.memory\[29\]\[0\] clknet_leaf_207_clk vss _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_1080 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08894__A1 vss _04234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06354__C1 vss _01959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_834 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_514 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10851_ vdd rf_ram.memory\[531\]\[1\] clknet_leaf_310_clk vss _00595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07449__A2 vss _03101_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_711 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08646__A1 vss _04097_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10782_ vdd rf_ram.memory\[565\]\[0\] clknet_leaf_326_clk vss _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06121__A2 vss _01500_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_859 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_539 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08949__A2 vss _04038_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11403_ _01135_ vdd vss clknet_leaf_231_clk net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09446__I0 vss net73 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_259_clk vdd vss clknet_leaf_259_clk clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09071__A1 vss net248 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_696 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11334_ vdd cpu.immdec.imm19_12_20\[0\] clknet_leaf_216_clk vss _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09566__S vss _04678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11265_ vdd net231 clknet_leaf_247_clk vss _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10216_ vdd _05099_ _05098_ _01311_ _05078_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11196_ vdd rf_ram.memory\[88\]\[0\] clknet_leaf_58_clk vss _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07385__A1 vss _02992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10147_ vdd vss _05057_ _03672_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05935__A2 vss _01633_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10078_ _05014_ _04396_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_89_403 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07613__I vss _02800_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_806 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06360__A2 vss _01846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_85_664 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_0_clk vdd vss clknet_0_clk clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_155_574 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06240_ _02434_ vdd vss _02435_ _01909_ _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__06112__A2 vss _01631_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_939 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_274_clk_I vss clknet_5_16__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_438 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09062__A1 vss _04331_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06171_ _02365_ vdd vss _02366_ _01527_ _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_180_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09930_ vdd vss _04924_ rf_ram.memory\[341\]\[0\] _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_289_clk_I vss clknet_5_18__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09861_ vdd vss _04881_ _02794_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09792_ vdd vss _04839_ rf_ram.memory\[80\]\[0\] _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_212_clk_I vss clknet_5_19__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08812_ _04205_ _04061_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05387__B1 vss _01555_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1020 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05308__I vss _01503_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05955_ _01503_ vdd vss _02151_ rf_ram.memory\[54\]\[0\] _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08743_ vdd vss _04162_ _04160_ _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09117__A2 vss _03692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07128__A1 vss _03123_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07523__I vss _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05886_ _01551_ vdd vss _02082_ rf_ram.memory\[64\]\[0\] _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08876__A1 vss _04237_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_227_clk_I vss clknet_5_23__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08674_ vdd _04118_ _04117_ _00749_ _04094_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07625_ vdd vss _03453_ rf_ram.memory\[407\]\[0\] _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_812 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07556_ vdd vss _03410_ _02806_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_5_4__f_clk_I vss clknet_3_1_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06507_ vdd vss _02697_ cpu.ctrl.pc_plus_offset_cy_r _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07487_ vdd _03367_ _03365_ _00313_ _03360_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09226_ vdd _04461_ _04460_ _00958_ _04431_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07300__A1 vss net239 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_314 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1034 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06438_ _02632_ vdd vss _02633_ _01903_ _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_91_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09157_ vdd vss _04419_ _02991_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06369_ rf_ram.memory\[245\]\[1\] _01610_ _01634_ rf_ram.memory\[244\]\[1\] _02564_
+ vss vdd rf_ram.memory\[247\]\[1\] _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_32_723 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07603__A2 vss _02813_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08800__A1 vss _04167_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08108_ vss _03754_ _03685_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09088_ vdd vss _04376_ rf_ram.memory\[569\]\[0\] _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output179_I vss net179 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08039_ vdd _03711_ _03709_ _00521_ _03690_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05927__B vss _02004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11050_ vdd rf_ram.memory\[143\]\[1\] clknet_leaf_10_clk vss _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10001_ vdd vss _04967_ _02910_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05378__B1 vss _01521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1115 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_222 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06590__A2 vss _02766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08867__A1 vss net239 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10903_ vdd rf_ram.memory\[185\]\[1\] clknet_leaf_17_clk vss _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10834_ vdd rf_ram.memory\[53\]\[0\] clknet_leaf_286_clk vss _00578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08619__A1 vss _04062_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_322 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10765_ vdd rf_ram.memory\[465\]\[1\] clknet_leaf_127_clk vss _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09292__A1 vss _04466_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06493__B vss _02687_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07842__A2 vss _03234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10696_ vdd rf_ram.memory\[433\]\[0\] clknet_leaf_82_clk vss _00440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09419__I0 vss net90 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09044__A1 vss _04334_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05853__A1 vss _01951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_583 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_1243 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_520 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_942 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11317_ _01050_ vdd vss clknet_leaf_262_clk net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_26_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_463 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07358__A1 vss _02788_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11248_ _00984_ vdd vss clknet_leaf_280_clk cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11179_ vdd rf_ram.memory\[94\]\[1\] clknet_leaf_55_clk vss _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05908__A2 vss _01706_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_920 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05740_ rf_ram.memory\[429\]\[0\] _01725_ _01724_ rf_ram.memory\[428\]\[0\] _01936_
+ vss vdd rf_ram.memory\[431\]\[0\] _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__06318__C1 vss _01773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_929 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07530__A1 vss _03393_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05671_ _01707_ vdd vss _01867_ rf_ram.memory\[462\]\[0\] _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06333__A2 vss _01515_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07410_ vdd _03318_ _03316_ _00285_ _03292_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05541__B1 vss _01679_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08390_ vdd vss _03930_ _03892_ _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_198 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07341_ vdd vss _03276_ rf_ram.memory\[270\]\[1\] _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_308 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_831 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_371 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_93_clk_I vss clknet_5_14__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_522 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_574 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07272_ vdd vss _03233_ rf_ram.memory\[193\]\[1\] _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_171_864 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06223_ _02417_ vdd vss _02418_ _01675_ _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09011_ vdd _04327_ _04325_ _00877_ _04301_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09035__A1 vss net249 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_188 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_712 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_967 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_268 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06154_ vdd vss _02349_ rf_ram.memory\[494\]\[1\] _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07597__A1 vss _03425_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05747__B vss _01756_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06085_ rf_ram.memory\[324\]\[1\] _02280_ vss vdd rf_ram.memory\[327\]\[1\] _01654_
+ rf_ram.memory\[325\]\[1\] _01656_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_106_1063 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_151_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09913_ vdd vss _04913_ rf_ram.memory\[344\]\[0\] _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09844_ vdd vss _01168_ _02714_ _04869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08010__A2 vss _03693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_80 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_31_clk_I vss clknet_5_6__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09775_ vdd vss _04828_ net243 _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06987_ vdd _03052_ _03051_ _00128_ _03050_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05938_ vdd vss _02134_ rf_ram.memory\[41\]\[0\] _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08849__A1 vss _04205_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08726_ vdd _04150_ _04149_ _00769_ _04126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06309__C1 vss _01953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_46_clk_I vss clknet_5_12__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08657_ vdd vss _04108_ _02953_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05869_ rf_ram.memory\[242\]\[0\] _02065_ vss vdd rf_ram.memory\[241\]\[0\] _01702_
+ rf_ram.memory\[243\]\[0\] _01625_ _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_68_439 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07608_ vdd vss _03442_ _02898_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_76_461 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08588_ vdd vss _04065_ rf_ram.memory\[167\]\[0\] _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07539_ vdd vss _03400_ rf_ram.memory\[360\]\[1\] _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10550_ vdd rf_ram.memory\[332\]\[0\] clknet_leaf_165_clk vss _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_146_371 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05501__I vss _01514_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06627__A3 vss _02730_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_104_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10481_ vdd rf_ram.memory\[420\]\[1\] clknet_leaf_104_clk vss _00225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09026__A1 vss _04331_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09209_ vdd vss _04451_ net241 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_1238 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_121_216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08812__I vss _04061_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07588__A1 vss _02889_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11102_ vdd rf_ram.memory\[125\]\[0\] clknet_leaf_83_clk vss _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_119_clk_I vss clknet_5_12__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_120_1049 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08001__A2 vss _02832_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11033_ vdd rf_ram.memory\[14\]\[1\] clknet_leaf_294_clk vss _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09501__A2 vss _02899_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07512__A1 vss _03360_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06315__A2 vss _01711_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_951 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_850 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1156 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10817_ vdd rf_ram.memory\[548\]\[1\] clknet_leaf_319_clk vss _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08068__A2 vss _03729_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_639 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_691 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10748_ vdd rf_ram.memory\[480\]\[0\] clknet_leaf_197_clk vss _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05411__I vss _01518_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_965 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_442 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_544 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10679_ vdd rf_ram.memory\[374\]\[1\] clknet_leaf_110_clk vss _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07579__A1 vss _03422_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput217 o_ibus_adr[23] net217 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput206 o_ibus_adr[13] net206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput228 o_ibus_adr[4] net228 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06251__A1 vss _01909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_293 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06910_ vdd vss _03002_ rf_ram.memory\[27\]\[0\] _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07890_ vdd _03617_ _03616_ _00466_ _03587_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07751__A1 vss _03524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06841_ vdd vss _02955_ _02935_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09740__A2 vss net16 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06772_ vdd vss _02906_ rf_ram.memory\[512\]\[0\] _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09560_ vdd vss _04678_ _04477_ _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_188_750 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05723_ vdd vss _01919_ rf_ram.memory\[433\]\[0\] _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_136_1056 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09491_ vdd vss _04626_ cpu.alu.i_rs1 _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08511_ _01366_ vdd vss _04015_ _03989_ _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07503__A1 vss _02781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1066 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08442_ vdd vss _03963_ rf_ram.memory\[175\]\[1\] _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06306__A2 vss _01989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05514__B1 vss _01656_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05654_ _01849_ vdd vss _01850_ _01769_ _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_65_409 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_461 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_466 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05585_ _01746_ vdd vss _01781_ _01776_ _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_850 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08373_ _03919_ _03685_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_19_859 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07806__A2 vss _03559_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_511 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07324_ vdd vss _03266_ rf_ram.memory\[255\]\[0\] _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07255_ vdd _03221_ _03219_ _00227_ _03193_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_731 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05321__I vss _01516_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06206_ _02399_ _02400_ vdd vss _02401_ _02397_ _02398_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06490__A1 vss _01349_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_171_694 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07186_ vdd _03179_ _03178_ _00200_ _03157_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_182_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05477__B vss _01672_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06137_ vss vdd rf_ram.memory\[293\]\[1\] _01793_ rf_ram.memory\[295\]\[1\] _01778_
+ _01777_ rf_ram.memory\[294\]\[1\] _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_14_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08231__A2 vss _02866_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06068_ _02262_ net253 vdd vss _02263_ _01600_ _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA_input55_I vss i_ibus_rdt[2] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07742__A1 vss _02788_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09827_ vdd vss _04860_ _03668_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09758_ vdd vss _04817_ _04804_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08709_ vdd vss _04140_ net235 _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09689_ _04768_ _04769_ vdd vss _04770_ net126 _04767_ net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__08298__A2 vss _03135_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05940__B vss _01563_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_450 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11651_ net173 vss vdd net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09247__A1 vss _03967_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10602_ vdd rf_ram.memory\[317\]\[0\] clknet_leaf_154_clk vss _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_500 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11582_ vdd rf_ram.memory\[23\]\[1\] clknet_leaf_290_clk vss _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_818 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10533_ vdd rf_ram.memory\[24\]\[1\] clknet_leaf_209_clk vss _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_load_slew245_I vss _02812_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1035 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10464_ vdd rf_ram.memory\[262\]\[0\] clknet_leaf_196_clk vss _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06490__C vss net254 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06481__A1 vss rf_ram.memory\[10\]\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10395_ vdd rf_ram.memory\[222\]\[1\] clknet_leaf_295_clk vss _00139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_1208 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09574__S vss _03967_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05441__C1 vss _01636_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07981__A1 vss _03651_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11016_ vdd rf_ram.memory\[155\]\[0\] clknet_leaf_332_clk vss _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_5_24__f_clk vdd vss clknet_5_24__leaf_clk clknet_3_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05406__I vss _01601_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1099 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_556 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09486__A1 vss _01375_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_731 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09238__A1 vss _04463_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_617 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_135 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1005 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_762 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_431 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_28_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05370_ vdd _01351_ _01565_ _01566_ _01557_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_396 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07040_ vdd _03086_ _03084_ _00147_ _03053_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_545 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08991_ vdd _04315_ _04313_ _00869_ _04301_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_167_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07942_ vdd _03649_ _03648_ _00486_ _03619_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05983__B1 vss _01714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07873_ vdd vss _03607_ _02836_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09713__A2 vss net7 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1220 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06824_ vdd _02943_ _02942_ _00074_ _02927_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07724__A1 vss _03491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09612_ vdd _04716_ _04714_ _01089_ _04637_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09543_ _04665_ vdd vss _01071_ _01732_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05316__I vss _01496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09477__A1 vss _02703_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06755_ vdd vss _02893_ _02773_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_188_580 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05706_ rf_ram.memory\[404\]\[0\] _01902_ vss vdd rf_ram.memory\[407\]\[0\] _01763_
+ rf_ram.memory\[405\]\[0\] _01656_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_149_934 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_411 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_556 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_718 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09474_ vss _01054_ _04613_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06686_ _02846_ vss vdd _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_05637_ vdd vss _01833_ rf_ram.memory\[510\]\[0\] _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08425_ vdd vss _03952_ rf_ram.memory\[173\]\[1\] _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08356_ vdd vss _03909_ rf_ram.memory\[182\]\[1\] _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_127 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_691 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07307_ vdd vss _03255_ rf_ram.memory\[257\]\[0\] _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05568_ rf_ram.memory\[259\]\[0\] _01763_ _01500_ rf_ram.memory\[258\]\[0\] _01764_
+ vss vdd rf_ram.memory\[257\]\[0\] _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_80_209 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_144_661 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08287_ vdd _03865_ _03863_ _00615_ _03855_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05499_ _01695_ _01518_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_33_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08452__A2 vss _01496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07238_ vdd _03211_ _03210_ _00220_ _03190_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06463__A1 vss _01599_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_478 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07169_ vdd vss _03169_ _02915_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08204__A2 vss _02992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10011__A2 vss _02839_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10180_ vdd vss _05077_ rf_ram.memory\[202\]\[1\] _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05974__B1 vss _01617_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09407__B vss _01344_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08507__A3 vss cpu.immdec.imm11_7\[4\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07715__A1 vss _02839_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_854 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_606 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08140__A1 vss _03757_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_932 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_723 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_285 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_902 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11634_ vss net157 net84 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_604 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_469 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11565_ vdd rf_ram.memory\[202\]\[0\] clknet_leaf_36_clk vss _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_648 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11496_ vdd rf_ram.memory\[276\]\[1\] clknet_leaf_189_clk vss _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10516_ vdd rf_ram.memory\[253\]\[0\] clknet_leaf_219_clk vss _00260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10447_ vdd rf_ram.memory\[496\]\[1\] clknet_leaf_198_clk vss _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10378_ vdd rf_ram.memory\[428\]\[0\] clknet_leaf_99_clk vss _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07954__A1 vss _03651_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06757__A2 vss _02894_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1217 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05717__B1 vss _01911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06390__B1 vss _02019_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05580__B vss _01693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06540_ vdd vss _02726_ _02719_ _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_158_775 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06471_ _01550_ vdd vss _02666_ rf_ram.memory\[24\]\[1\] _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_87_375 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_1183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08131__A1 vss _02805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05422_ vdd vss _01618_ rf_ram.memory\[353\]\[0\] _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08210_ vdd vss _03818_ rf_ram.memory\[535\]\[0\] _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08682__A2 vss _04078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09190_ vdd vss _04440_ rf_ram.memory\[83\]\[0\] _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08434__A2 vss _03949_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_659 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08141_ vdd vss _03775_ net241 _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05353_ rf_ram.memory\[532\]\[0\] _01549_ vss vdd rf_ram.memory\[535\]\[0\] _01520_
+ rf_ram.memory\[533\]\[0\] _01516_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_05284_ vdd vss _01482_ _01442_ cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08072_ vdd _03732_ _03730_ _00533_ _03724_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05653__C1 vss _01848_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07023_ vdd _03075_ _03073_ _00141_ _03053_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08198__A1 vss _03790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09934__A2 vss _03135_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08974_ vdd _04305_ _04304_ _00862_ _04298_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05956__B1 vss _01655_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05420__A2 vss _01614_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07925_ vdd vss _03639_ _02774_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09698__A1 vss net129 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09698__B2 vss net99 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07856_ vdd vss _03597_ rf_ram.memory\[430\]\[1\] _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08370__A1 vss _03884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07787_ vdd _03553_ _03551_ _00427_ _03524_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06807_ vdd _02931_ _02928_ _00069_ _02930_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input18_I vss i_dbus_rdt[24] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09526_ vdd vss _04654_ _03967_ _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_06738_ vdd _02880_ _02878_ _00051_ _02876_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08122__A1 vss _03754_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09457_ _04604_ vdd vss _04605_ net78 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_583 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06669_ vdd vss _02833_ _02829_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08408_ vdd vss _03941_ rf_ram.memory\[178\]\[1\] _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09388_ _04564_ net217 vdd vss _04567_ net216 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08339_ vdd vss _03898_ rf_ram.memory\[240\]\[1\] _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09473__I1 vss net88 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_439 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_119 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11350_ _01082_ vdd vss clknet_leaf_216_clk cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06605__I vss _02780_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05649__C vss net253 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05644__C1 vss _01519_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10301_ vdd rf_ram.memory\[520\]\[1\] clknet_leaf_316_clk vss _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_675 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08189__A1 vss _03668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_692 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11281_ vdd net217 clknet_leaf_244_clk vss _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09386__B1 vss _04564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10232_ vdd vss _05109_ rf_ram.memory\[237\]\[1\] _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10163_ vdd vss _05067_ rf_ram.memory\[448\]\[0\] _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05665__B vss _01860_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10094_ vdd _05024_ _05022_ _01264_ _05017_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09689__A1 vss net126 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05384__C vss _01495_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07164__A2 vss _03158_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_804 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_1058 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05175__A1 vss _01375_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_550 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10996_ vdd rf_ram.memory\[549\]\[0\] clknet_leaf_324_clk vss _00733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_915 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09861__A1 vss _02794_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_548 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_378 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_924 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08416__A2 vss _03945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09613__A1 vss net250 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11617_ vss net139 net67 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_957 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11548_ vdd rf_ram.memory\[454\]\[1\] clknet_leaf_121_clk vss _01280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11479_ vdd rf_ram.memory\[336\]\[0\] clknet_leaf_177_clk vss _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_512 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_640 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap238 net238 _02898_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_21_651 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07927__A1 vss _03619_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_695 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06060__C1 vss _01656_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1025 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05402__A2 vss _01478_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07710_ vdd vss _03506_ net240 _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05971_ _01624_ rf_ram.memory\[27\]\[0\] vdd vss _02167_ rf_ram.memory\[26\]\[0\]
+ _01686_ _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__08352__A1 vss _03887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08690_ vdd _04128_ _04127_ _00755_ _04126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_815 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07641_ vdd vss _03463_ _02889_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07572_ vdd vss _03420_ rf_ram.memory\[317\]\[0\] _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06902__A2 vss _02939_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_695 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09311_ vdd vss _04523_ _04477_ net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06523_ vdd vss _02711_ _01399_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_150_1170 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09852__A1 vss _01385_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05469__A2 vss _01509_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06454_ _01601_ vdd vss _02649_ rf_ram.memory\[56\]\[1\] _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06666__A1 vss cpu.immdec.imm11_7\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09242_ net66 vdd vss _04472_ cpu.genblk3.csr.mie_mtie cpu.genblk3.csr.mstatus_mie
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09173_ vdd vss _04429_ rf_ram.memory\[85\]\[0\] _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06385_ vdd vss _02580_ rf_ram.memory\[73\]\[1\] _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05874__C1 vss _01696_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05405_ _01601_ rf_ram.i_raddr\[2\] vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_8_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09604__A1 vss _04478_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_225 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10214__A2 vss _02954_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08124_ vdd _03764_ _03762_ _00553_ _03757_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05336_ _01532_ _01531_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06969__A2 vss _03040_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07091__A1 vss _03092_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_95 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08055_ _03721_ _03685_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05267_ _01386_ cpu.genblk3.csr.mcause3_0\[0\] vdd vss _01466_ cpu.genblk3.csr.mcause31
+ _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_141_483 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05641__A2 vss _01652_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07006_ vdd _03064_ _03062_ _00135_ _03053_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05198_ vdd vss _01398_ cpu.ctrl.pc_plus_offset_cy_r _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07256__I vss _03013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08591__A1 vss _04062_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08957_ vdd vss _04294_ rf_ram.memory\[120\]\[1\] _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08888_ vdd vss _04252_ rf_ram.memory\[479\]\[0\] _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07908_ vdd vss _03629_ rf_ram.memory\[460\]\[1\] _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07839_ vdd vss _03586_ rf_ram.memory\[411\]\[1\] _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07146__A2 vss _02911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08343__A1 vss _03884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06354__B1 vss _01968_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10850_ vdd rf_ram.memory\[531\]\[0\] clknet_leaf_306_clk vss _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06106__B1 vss _01679_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09509_ vdd _04640_ _04639_ _01062_ _04634_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_846 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10781_ vdd rf_ram.memory\[566\]\[1\] clknet_leaf_325_clk vss _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06657__A1 vss _02815_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1105 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_827 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11402_ _01134_ vdd vss clknet_leaf_230_clk net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09446__I1 vss net74 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09071__A2 vss _04005_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05880__A2 vss _01755_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_264 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07082__A1 vss _02781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11333_ vdd cpu.immdec.imm31 clknet_leaf_236_clk vss _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_21__f_clk_I vss clknet_3_5_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06290__C1 vss _01857_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11264_ vdd net230 clknet_leaf_247_clk vss _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07909__A1 vss _03622_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10215_ vdd vss _05099_ rf_ram.memory\[207\]\[0\] _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06042__C1 vss _01610_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07385__A2 vss _02997_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11195_ vdd rf_ram.memory\[159\]\[1\] clknet_leaf_5_clk vss _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08582__A1 vss _04058_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10146_ vdd _05056_ _05054_ _01284_ _05049_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_391 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06003__C vss _01495_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10077_ vdd _05013_ _05011_ _01258_ _04985_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10141__A1 vss _05049_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08885__A2 vss _04248_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05699__A2 vss _01543_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_195_clk vdd vss clknet_leaf_195_clk clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_173_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_1165 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05414__I vss _01609_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09834__A1 vss _04837_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10979_ vdd rf_ram.memory\[168\]\[1\] clknet_leaf_1_clk vss _00716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06648__A1 vss _02813_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_258 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06170_ rf_ram.memory\[509\]\[1\] _01645_ _01644_ rf_ram.memory\[508\]\[1\] _02365_
+ vss vdd rf_ram.memory\[511\]\[1\] _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__05871__A2 vss _01641_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1071 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_275 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_269 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_450 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06820__A1 vss _02799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_623 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05623__A2 vss _01677_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_342 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09860_ _02714_ vdd vss _01174_ _04877_ _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08573__A1 vss _02945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09791_ vdd vss _04838_ _02945_ _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08811_ vdd _04204_ _04203_ _00800_ _04202_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05954_ _01562_ vdd vss _02150_ _02148_ _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08742_ vdd _01506_ _04158_ _04161_ _01498_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_1076 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08325__A1 vss _03035_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08673_ vdd vss _04118_ rf_ram.memory\[156\]\[0\] _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07624_ vdd vss _03452_ _03082_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06887__A1 vss _02970_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_186_clk vdd vss clknet_leaf_186_clk clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05885_ _01928_ vdd vss _02081_ _02078_ _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_166_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05324__I vss _01519_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07555_ vdd _03409_ _03407_ _00339_ _03393_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07486_ vdd vss _03367_ rf_ram.memory\[365\]\[1\] _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06639__A1 vss _02743_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_211 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08635__I vss _04057_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1160 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06506_ _02696_ vdd vss _00005_ _02692_ _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09225_ vdd vss _04461_ rf_ram.memory\[339\]\[0\] _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07300__A2 vss _02941_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06437_ rf_ram.memory\[45\]\[1\] _01609_ _01633_ rf_ram.memory\[44\]\[1\] _02632_
+ vss vdd rf_ram.memory\[47\]\[1\] _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__05847__C1 vss _01725_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09156_ vss _04418_ _04004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06368_ _02004_ vdd vss _02563_ rf_ram.memory\[246\]\[1\] _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10199__A1 vss _02908_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_5_clk_I vss clknet_5_1__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05862__A2 vss _01523_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_110_clk vdd vss clknet_leaf_110_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07064__A1 vss _03087_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_91 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05319_ _01515_ _01514_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08107_ vdd _03753_ _03751_ _00547_ _03724_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06299_ _02493_ vdd vss _02494_ _01552_ _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09087_ vdd vss _04375_ _02983_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1068 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08038_ vdd vss _03711_ rf_ram.memory\[568\]\[1\] _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_987 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06104__B vss _01684_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10000_ vdd _04966_ _04964_ _01228_ _04953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09989_ vdd vss _04960_ rf_ram.memory\[503\]\[1\] _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_5__f_clk vdd vss clknet_5_5__leaf_clk clknet_3_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_177_clk vdd vss clknet_leaf_177_clk clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08867__A2 vss _04195_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_334_clk_I vss clknet_5_0__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06878__A1 vss _02935_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10902_ vdd rf_ram.memory\[185\]\[0\] clknet_leaf_17_clk vss _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09816__A1 vss _04840_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10833_ vdd rf_ram.memory\[540\]\[1\] clknet_leaf_273_clk vss _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10764_ vdd rf_ram.memory\[465\]\[0\] clknet_leaf_126_clk vss _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_974 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06493__C vss _01373_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_884 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_361 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10695_ vdd rf_ram.memory\[413\]\[1\] clknet_leaf_83_clk vss _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_819 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_713 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_101_clk vdd vss clknet_leaf_101_clk clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07055__A1 vss _02806_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_543 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06802__A1 vss _02801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11316_ _01049_ vdd vss clknet_leaf_262_clk net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07358__A2 vss _03253_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08555__A1 vss _04023_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05409__I vss _01499_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11247_ vdd cpu.immdec.imm11_7\[1\] clknet_leaf_279_clk vss _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11178_ vdd rf_ram.memory\[94\]\[0\] clknet_leaf_57_clk vss _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10129_ vdd _05045_ _05043_ _01278_ _05017_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06030__A2 vss _01511_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08307__A1 vss _03855_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_168_clk vdd vss clknet_leaf_168_clk clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_136_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10114__A1 vss _05017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06318__B1 vss _01772_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_954 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06869__A1 vss _02970_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05670_ _01861_ _01865_ vdd vss _01866_ _01850_ _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09807__A1 vss _02774_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1003 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07340_ vdd _03275_ _03274_ _00258_ _03257_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_654 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07294__A1 vss _03225_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06097__A2 vss _01735_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09010_ vdd vss _04327_ rf_ram.memory\[110\]\[1\] _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07271_ vdd _03232_ _03231_ _00232_ _03222_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06222_ rf_ram.memory\[391\]\[1\] _01778_ _01777_ rf_ram.memory\[390\]\[1\] _02417_
+ vss vdd rf_ram.memory\[389\]\[1\] _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09035__A2 vss _04339_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05844__A2 vss _01808_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07046__A1 vss _03087_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06153_ _02347_ vdd vss _02348_ _01597_ _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_13_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06254__C1 vss _01726_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08794__A1 vss _04167_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06084_ _01707_ vdd vss _02279_ rf_ram.memory\[326\]\[1\] _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09912_ vdd vss _04912_ _04911_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08546__A1 vss _02764_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05319__I vss _01514_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_172 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09843_ vdd vss cpu.state.cnt_r\[2\] _04869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06006__C1 vss _01520_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09774_ vdd _04827_ _04825_ _01140_ _04637_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06986_ vdd vss _03052_ rf_ram.memory\[227\]\[0\] _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_159_clk vdd vss clknet_leaf_159_clk clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10105__A1 vss _02800_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05937_ _01601_ vdd vss _02133_ rf_ram.memory\[40\]\[0\] _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08725_ vdd vss _04150_ rf_ram.memory\[14\]\[0\] _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06309__B1 vss _01516_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05868_ _01684_ vdd vss _02064_ rf_ram.memory\[240\]\[0\] _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08656_ vdd _04107_ _04105_ _00742_ _04097_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07607_ vdd _03441_ _03439_ _00359_ _03425_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08587_ vdd vss _04064_ _02828_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07538_ vdd _03399_ _03398_ _00332_ _03389_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_165_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05532__B2 vss _01727_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05799_ _01494_ vdd vss _01995_ _01992_ _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_119_542 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07285__A1 vss _02836_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07469_ _03355_ vss vdd _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_331_clk vdd vss clknet_leaf_331_clk clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10480_ vdd rf_ram.memory\[420\]\[0\] clknet_leaf_103_clk vss _00224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09208_ vdd _04450_ _04448_ _00951_ _04434_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05835__A2 vss _01755_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09139_ vdd vss _04408_ rf_ram.memory\[169\]\[1\] _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_543 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_392 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07588__A2 vss _03390_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_885 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11101_ vdd rf_ram.memory\[126\]\[1\] clknet_leaf_78_clk vss _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05599__A1 vss _01675_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06260__A2 vss _01755_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_1250 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11032_ vdd rf_ram.memory\[14\]\[0\] clknet_leaf_294_clk vss _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05673__B vss _01650_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06012__A2 vss _01511_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06488__C vss rf_ram.i_raddr\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_273_clk_I vss clknet_5_16__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_407 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1008 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157_637 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_288_clk_I vss clknet_5_18__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_484 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10816_ vdd rf_ram.memory\[548\]\[0\] clknet_leaf_319_clk vss _00560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_361 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10747_ vdd rf_ram.memory\[481\]\[1\] clknet_leaf_187_clk vss _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_211_clk_I vss clknet_5_28__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_322_clk vdd vss clknet_leaf_322_clk clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10678_ vdd rf_ram.memory\[374\]\[0\] clknet_leaf_110_clk vss _00422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05826__A2 vss _01537_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07028__A1 vss _03053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08776__A1 vss _04170_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput207 o_ibus_adr[14] net207 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_leaf_226_clk_I vss clknet_5_23__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_727 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput229 o_ibus_adr[5] net229 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput218 o_ibus_adr[24] net218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_142_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_1237 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06840_ _02954_ vss vdd _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_171_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_88 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06771_ vdd vss _02905_ _02881_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05722_ _01918_ vss vdd _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_09490_ vdd _01442_ _01342_ _04625_ cpu.bne_or_bge vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08510_ _04013_ vdd vss _04014_ _04010_ _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_188_784 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07503__A2 vss _03101_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_401 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05653_ vss vdd rf_ram.memory\[469\]\[0\] _01848_ rf_ram.memory\[471\]\[0\] _01786_
+ _01785_ rf_ram.memory\[470\]\[0\] _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_08441_ vdd _03962_ _03961_ _00672_ _03953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_50 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05584_ _01778_ rf_ram.memory\[299\]\[0\] vdd vss _01780_ rf_ram.memory\[298\]\[0\]
+ _01777_ _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08372_ vdd _03918_ _03916_ _00647_ _03887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07267__A1 vss _03225_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07323_ vdd vss _03265_ _03055_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_313_clk vdd vss clknet_leaf_313_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_45_123 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07254_ vdd vss _03221_ rf_ram.memory\[41\]\[1\] _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05817__A2 vss _01856_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06205_ rf_ram.memory\[451\]\[1\] _01811_ _01801_ rf_ram.memory\[450\]\[1\] _02400_
+ vss vdd rf_ram.memory\[449\]\[1\] _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__07019__A1 vss _03055_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1028 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07185_ vdd vss _03179_ rf_ram.memory\[198\]\[0\] _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_565 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08767__A1 vss _02945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05477__C vss net253 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06136_ vdd vss _02331_ rf_ram.memory\[292\]\[1\] _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06067_ _02256_ _01599_ _02261_ vdd vss _02262_ _02253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__06242__A2 vss _01787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_979 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08519__A1 vss _02838_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input48_I vss i_ibus_rdt[23] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09826_ vdd _04859_ _04857_ _01160_ _04840_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06969_ vdd vss _03041_ _02788_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05753__A1 vss _01372_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09757_ vdd vss _04816_ _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06545__A3 vss _02730_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_1135 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08708_ vdd _04139_ _04137_ _00762_ _04129_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09688_ vdd vss _04769_ _04740_ net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08639_ _04097_ _04061_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_11650_ net172 vss vdd net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09247__A2 vss net56 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_473 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10601_ vdd rf_ram.memory\[357\]\[1\] clknet_leaf_155_clk vss _00345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11581_ vdd rf_ram.memory\[23\]\[0\] clknet_leaf_207_clk vss _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_304_clk vdd vss clknet_leaf_304_clk clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_153_128 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10532_ vdd rf_ram.memory\[24\]\[0\] clknet_leaf_209_clk vss _00276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_925 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_860 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_578 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_835 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10463_ vdd rf_ram.memory\[273\]\[1\] clknet_leaf_188_clk vss _00207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06481__A2 vss _01686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08758__A1 vss _04170_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10394_ vdd rf_ram.memory\[222\]\[0\] clknet_leaf_300_clk vss _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_502 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_885 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06233__A2 vss _01634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05441__B1 vss _01610_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09183__A1 vss _04434_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05992__A1 vss _01371_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11015_ vdd rf_ram.memory\[559\]\[1\] clknet_leaf_323_clk vss _00752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_92_clk_I vss clknet_5_11__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06536__A3 vss _01341_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07497__A1 vss _03360_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05850__C vss _01362_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_905 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_968 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06518__I vss _01411_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_150_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08997__A1 vss _02945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_30_clk_I vss clknet_5_6__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_476 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_454 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_165_clk_I vss clknet_5_27__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_835 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06472__A2 vss _01514_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08749__A1 vss _04126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_45_clk_I vss clknet_5_12__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05432__B1 vss _01625_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08990_ vdd vss _04315_ rf_ram.memory\[114\]\[1\] _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07941_ vdd vss _03649_ rf_ram.memory\[43\]\[0\] _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09174__A1 vss _04397_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05983__A1 vss rf_ram.memory\[4\]\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07872_ vdd _03606_ _03604_ _00459_ _03590_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06202__B vss _01805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06823_ vdd vss _02943_ rf_ram.memory\[287\]\[0\] _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08921__A1 vss _04266_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09611_ vdd vss _04716_ rf_ram.memory\[73\]\[1\] _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_103_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09542_ net41 _04650_ cpu.immdec.imm19_12_20\[5\] vdd vss _04665_ _04478_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06754_ vdd _02892_ _02890_ _00055_ _02876_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05705_ _01504_ vdd vss _01901_ rf_ram.memory\[406\]\[0\] _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_92_97 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_90_clk vdd vss clknet_leaf_90_clk clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07488__A1 vss _02795_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09473_ _04604_ vdd vss _04613_ net86 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06685_ _02734_ vdd vss _02845_ _02730_ _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_176_776 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_118_clk_I vss clknet_5_12__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05636_ _01824_ _01828_ _01831_ vdd vss _01832_ _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_08424_ vdd _03951_ _03950_ _00666_ _03919_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_624 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05332__I vss _01527_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_798 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_404 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05567_ vdd vss _01763_ _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_08355_ vdd _03908_ _03907_ _00640_ _03884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07306_ vdd vss _03254_ _02899_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06448__C1 vss _01609_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_774 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_605 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05498_ _01693_ vdd vss _01694_ rf_ram.memory\[336\]\[0\] _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08286_ vdd vss _03865_ rf_ram.memory\[204\]\[1\] _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07237_ vdd vss _03211_ rf_ram.memory\[422\]\[0\] _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07660__A1 vss _03458_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_375 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07168_ vdd _03168_ _03166_ _00193_ _03161_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_5_30__f_clk vdd vss clknet_5_30__leaf_clk clknet_3_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07412__A1 vss _03319_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06215__A2 vss _01777_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06119_ rf_ram.memory\[261\]\[1\] _01668_ _01509_ rf_ram.memory\[260\]\[1\] _02314_
+ vss vdd rf_ram.memory\[263\]\[1\] _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_100_710 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05423__B1 vss _01608_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07099_ vdd vss _03125_ rf_ram.memory\[48\]\[0\] _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output154_I vss net154 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07715__A2 vss _03496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09809_ vdd _04849_ _04848_ _01153_ _04837_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_1218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_81_clk vdd vss clknet_leaf_81_clk clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06151__A1 vss _01768_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11633_ vss net156 net83 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_270 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_757 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08979__A1 vss _04298_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11564_ vdd rf_ram.memory\[20\]\[1\] clknet_leaf_292_clk vss _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07651__A1 vss net239 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11495_ vdd rf_ram.memory\[276\]\[0\] clknet_leaf_189_clk vss _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10515_ vdd rf_ram.memory\[270\]\[1\] clknet_leaf_191_clk vss _00259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06454__A2 vss _01613_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10446_ vdd rf_ram.memory\[496\]\[0\] clknet_leaf_198_clk vss _00190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07403__A1 vss _03289_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_716 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10377_ vdd rf_ram.memory\[22\]\[1\] clknet_leaf_209_clk vss _00121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06801__I vss _02819_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05417__I vss _01508_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06022__B vss _01506_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05861__B vss _01494_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_72_clk vdd vss clknet_leaf_72_clk clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06470_ _01493_ vdd vss _02665_ _02662_ _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08131__A2 vss _03765_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_253 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05421_ _01617_ vss vdd _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07890__A1 vss _03587_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08140_ vdd _03774_ _03772_ _00559_ _03757_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_638 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05352_ _01505_ vdd vss _01548_ rf_ram.memory\[534\]\[0\] _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_125_150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06445__A2 vss _01605_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05283_ _01452_ vdd vss _01481_ _01442_ _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08071_ vdd vss _03732_ rf_ram.memory\[562\]\[1\] _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05653__B1 vss _01786_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07022_ vdd vss _03075_ rf_ram.memory\[245\]\[1\] _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_140_164 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08973_ vdd vss _04305_ rf_ram.memory\[117\]\[0\] _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_80_1188 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07924_ vdd _03638_ _03636_ _00479_ _03622_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05327__I vss _01509_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07855_ vdd _03596_ _03595_ _00452_ _03587_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07786_ vdd vss _03553_ rf_ram.memory\[416\]\[1\] _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06806_ vdd vss _02931_ rf_ram.memory\[291\]\[1\] _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09525_ vdd vss _04653_ _01491_ _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06737_ vdd vss _02880_ rf_ram.memory\[517\]\[1\] _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_754 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06668_ vss _02832_ _02831_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xclkbuf_leaf_63_clk vdd vss clknet_leaf_63_clk clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09456_ _04604_ _01411_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05619_ _01814_ net253 vdd vss _01815_ _01768_ _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08407_ vdd _03940_ _03939_ _00660_ _03919_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_163_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09387_ vdd vss _04566_ _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06599_ vdd vss _02777_ rf_ram.memory\[234\]\[0\] _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08338_ vdd _03897_ _03896_ _00634_ _03884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_621 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06436__A2 vss _01530_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08269_ vdd _03854_ _03853_ _00608_ _03852_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_952 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06107__B vss _01746_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05644__B1 vss _01668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11280_ _01015_ vdd vss clknet_leaf_245_clk net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10300_ vdd rf_ram.memory\[520\]\[0\] clknet_leaf_316_clk vss _00044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_378 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08189__A2 vss _03072_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10231_ vdd _05108_ _05107_ _01317_ _05078_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09386__B2 vss net216 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_max_cap248_I vss _02760_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10162_ vdd vss _05066_ _02831_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05947__A1 vss _01903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output79_I vss net79 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10093_ vdd vss _05024_ rf_ram.memory\[310\]\[1\] _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09138__A1 vss _04397_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1072 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_816 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_1026 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05175__A2 vss _01376_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_54_clk vdd vss clknet_leaf_54_clk clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10995_ vdd rf_ram.memory\[539\]\[1\] clknet_leaf_313_clk vss _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09310__A1 vss _01491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06124__A1 vss _01674_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09861__A2 vss _03035_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_335 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07872__A1 vss _03590_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09613__A2 vss _04507_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11616_ vss net169 net96 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_413 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07624__A1 vss _03082_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11547_ vdd rf_ram.memory\[454\]\[0\] clknet_leaf_121_clk vss _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06427__A2 vss _01677_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_952 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_440 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06017__B vss _01506_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_928 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11478_ vdd rf_ram.memory\[337\]\[1\] clknet_leaf_175_clk vss _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_337 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10429_ vdd rf_ram.memory\[488\]\[1\] clknet_leaf_222_clk vss _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_546 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06060__B1 vss _01763_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05970_ vdd vss _02166_ rf_ram.memory\[25\]\[0\] _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05147__I vss _01349_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07640_ vdd _03462_ _03460_ _00371_ _03458_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07571_ vdd vss _03419_ _02935_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_45_clk vdd vss clknet_leaf_45_clk clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06522_ _01405_ _01375_ vdd vss _02710_ _01442_ _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_48_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09310_ _04013_ _03967_ vdd vss _04522_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_119_916 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07863__A1 vss _02774_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06453_ _02647_ vdd vss _02648_ _01526_ _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06666__A2 vss cpu.immdec.imm11_7\[4\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_763 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09241_ vdd vss _04471_ _01418_ _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_576 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09172_ vdd vss _04428_ _03071_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06384_ _01551_ vdd vss _02579_ rf_ram.memory\[72\]\[1\] _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_84_891 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05874__B1 vss _01793_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05404_ _01600_ _01599_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_185_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06418__A2 vss _01706_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05335_ _01531_ _01530_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08123_ vdd vss _03764_ rf_ram.memory\[552\]\[1\] _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_43_232 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09604__A2 vss cpu.immdec.imm30_25\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1217 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08054_ vdd _03720_ _03718_ _00527_ _03690_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_827 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05266_ vdd vss _01465_ _01409_ _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07005_ vdd vss _03064_ rf_ram.memory\[224\]\[1\] _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_652 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05766__B vss _01564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05197_ vdd vss _01397_ _01389_ _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08040__A1 vss net235 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ vdd _04293_ _04292_ _00856_ _04266_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input30_I vss i_dbus_rdt[6] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08887_ vdd vss _04251_ _03672_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07907_ vdd _03628_ _03627_ _00472_ _03619_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07838_ vdd _03585_ _03584_ _00446_ _03554_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09540__A1 vss _04478_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1033 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07769_ vdd _03542_ _03541_ _00420_ _03521_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05562__C1 vss _01715_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09508_ vdd vss _04640_ rf_ram.memory\[279\]\[0\] _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_36_clk vdd vss clknet_leaf_36_clk clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_79_674 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_1010 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_335 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10780_ vdd rf_ram.memory\[566\]\[0\] clknet_leaf_325_clk vss _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_549 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06657__A2 vss _02822_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_735 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1038 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09439_ vss _01037_ _04595_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_152_705 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_749 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06409__A2 vss _01510_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11401_ _01133_ vdd vss clknet_leaf_227_clk net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_105_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_690 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07082__A2 vss _02911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11332_ vdd cpu.genblk3.csr.timer_irq_r clknet_leaf_240_clk vss _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05676__B vss _01805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06290__B1 vss _01931_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09359__A1 vss net233 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11263_ vdd net229 clknet_leaf_251_clk vss _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10214_ vdd vss _05098_ _03892_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11194_ vdd rf_ram.memory\[159\]\[0\] clknet_leaf_4_clk vss _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_1281 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05395__C vss _01564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06042__B1 vss _01608_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10145_ vdd vss _05056_ rf_ram.memory\[452\]\[1\] _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_882 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09662__I vss net120 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10076_ vdd vss _05013_ rf_ram.memory\[308\]\[1\] _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09531__A1 vss _04526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06300__B vss _01956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_337 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05553__C1 vss _01625_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_27_clk vdd vss clknet_leaf_27_clk clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08098__A1 vss _02787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10978_ vdd rf_ram.memory\[168\]\[0\] clknet_leaf_1_clk vss _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06648__A2 vss _02815_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_724 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06526__I vss net65 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05856__B1 vss _01959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05430__I vss _01514_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09598__A1 vss _04478_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_917 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1202 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_298 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_1115 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06820__A2 vss _02939_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_679 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_77 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08022__A1 vss _03686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09770__A1 vss net243 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08573__A2 vss _03945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08810_ vdd vss _04204_ rf_ram.memory\[138\]\[0\] _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_376 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09790_ _04837_ _04396_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05387__A2 vss _01538_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05953_ vss vdd rf_ram.memory\[57\]\[0\] _01655_ rf_ram.memory\[59\]\[0\] _01653_
+ _01661_ rf_ram.memory\[58\]\[0\] _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_08741_ vdd vss _04160_ _02718_ _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_108_61 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05884_ rf_ram.memory\[75\]\[0\] _02079_ vdd vss _02080_ rf_ram.memory\[74\]\[0\]
+ _01808_ _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08325__A2 vss _03072_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08672_ vdd vss _04117_ _02838_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07623_ vdd _03451_ _03449_ _00365_ _03425_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05605__I vss _01661_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1065 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_18_clk vdd vss clknet_leaf_18_clk clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_75_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_860 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07554_ vdd vss _03409_ rf_ram.memory\[31\]\[1\] _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08916__I vss _04061_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07485_ vdd _03366_ _03365_ _00312_ _03356_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07836__A1 vss _02822_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_370 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06505_ vdd vss _02696_ _01409_ _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_48_379 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09224_ vdd vss _04460_ _03319_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06436_ vdd vss _02631_ rf_ram.memory\[46\]\[1\] _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05847__B1 vss _01811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_880 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_418 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05340__I vss _01508_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09589__A1 vss _03967_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05311__A2 vss _01502_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_360 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10199__A2 vss _03902_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09155_ vdd _04417_ _04415_ _00931_ _04401_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06367_ _02558_ _02561_ vdd vss _02562_ _02550_ _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_130_911 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09086_ vdd _04374_ _04372_ _00905_ _04367_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_1036 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08261__A1 vss _03230_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05318_ _01514_ _01513_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08106_ vdd vss _03753_ rf_ram.memory\[555\]\[1\] _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06298_ rf_ram.memory\[166\]\[1\] _02493_ vss vdd rf_ram.memory\[165\]\[1\] _01516_
+ rf_ram.memory\[167\]\[1\] _01520_ _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_130_955 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_101_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05249_ _01446_ _01448_ vdd vss _01449_ _01428_ _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_08037_ vdd _03710_ _03709_ _00520_ _03686_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_134 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_482 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09988_ vdd _04959_ _04958_ _01223_ _04950_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05378__A2 vss _01532_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06575__A1 vss _01562_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157_1100 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08939_ vdd vss _04283_ net245 _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output234_I vss net234 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06120__B vss _01526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_235 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05515__I vss _01613_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10901_ vdd rf_ram.memory\[184\]\[1\] clknet_leaf_20_clk vss _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06327__A1 vss _01951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06878__A2 vss _02844_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_279 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_605 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_819 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10832_ vdd rf_ram.memory\[540\]\[0\] clknet_leaf_273_clk vss _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_638 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_690 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10763_ vdd rf_ram.memory\[466\]\[1\] clknet_leaf_125_clk vss _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10694_ vdd rf_ram.memory\[413\]\[0\] clknet_leaf_91_clk vss _00438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_513 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_502 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_215 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_963 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07055__A2 vss _02869_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06802__A2 vss _02889_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1109 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11315_ _01048_ vdd vss clknet_leaf_267_clk net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06014__C vss _01564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11246_ vdd cpu.immdec.imm11_7\[0\] clknet_leaf_258_clk vss _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11177_ vdd rf_ram.memory\[95\]\[1\] clknet_leaf_62_clk vss _00913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06566__A1 vss _01496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08510__B vss _04013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10128_ vdd vss _05045_ rf_ram.memory\[475\]\[1\] _05043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1165 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_1206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10059_ vdd vss _05003_ rf_ram.memory\[507\]\[0\] _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06030__B vss _01552_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05526__C1 vss _01713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_988 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05541__A2 vss _01687_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_791 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07818__A1 vss _03554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09807__A2 vss _04004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1037 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07270_ vdd vss _03232_ rf_ram.memory\[193\]\[0\] _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_636 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06221_ vdd vss _02416_ rf_ram.memory\[388\]\[1\] _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_115_237 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06152_ _02346_ vdd vss _02347_ net252 _02319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08243__A1 vss _03820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06254__B1 vss _01725_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10050__A1 vss _04982_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06083_ _02274_ _02277_ vdd vss _02278_ _02266_ _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__09991__A1 vss _02727_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_65 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09911_ _04911_ vss vdd _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xclkbuf_leaf_7_clk vdd vss clknet_leaf_7_clk clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1_696 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06006__B1 vss _01516_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08546__A2 vss _02867_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09842_ vdd vss _01167_ _02714_ _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09773_ vdd vss _04827_ rf_ram.memory\[269\]\[1\] _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08724_ vdd vss _04149_ _02971_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06985_ vdd vss _03051_ _02766_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10105__A2 vss _02992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05936_ _02131_ vdd vss _02132_ _01903_ _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__05335__I vss _01530_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05780__A2 vss _01915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05867_ rf_ram.memory\[245\]\[0\] _01610_ _01634_ rf_ram.memory\[244\]\[0\] _02063_
+ vss vdd rf_ram.memory\[247\]\[0\] _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08655_ vdd vss _04107_ rf_ram.memory\[160\]\[1\] _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07606_ vdd vss _03441_ rf_ram.memory\[314\]\[1\] _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_238 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08586_ vdd _04063_ _04059_ _00716_ _04062_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07537_ vdd vss _03399_ rf_ram.memory\[360\]\[0\] _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05798_ _01520_ rf_ram.memory\[163\]\[0\] vdd vss _01994_ rf_ram.memory\[162\]\[0\]
+ _01958_ _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_91_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07285__A2 vss _03083_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07468_ vdd _03354_ _03352_ _00307_ _03326_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_1234 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08482__A1 vss _03991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06419_ _01928_ vdd vss _02614_ _02611_ _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09207_ vdd vss _04450_ rf_ram.memory\[6\]\[1\] _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07399_ vdd vss _03312_ rf_ram.memory\[248\]\[1\] _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output184_I vss net184 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09138_ vdd _04407_ _04406_ _00924_ _04397_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_894 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11100_ vdd rf_ram.memory\[126\]\[0\] clknet_leaf_78_clk vss _00836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06115__B vss _01756_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09069_ vdd _04363_ _04361_ _00899_ _04334_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06796__A1 vss _02921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1240 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11031_ vdd rf_ram.memory\[89\]\[1\] clknet_leaf_59_clk vss _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05954__B vss _01562_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06548__A1 vss _01353_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05771__A2 vss _01523_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_903 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_435 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06720__A1 vss _02797_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10815_ vdd rf_ram.memory\[54\]\[1\] clknet_leaf_297_clk vss _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_885 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10746_ vdd rf_ram.memory\[481\]\[0\] clknet_leaf_197_clk vss _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05287__A1 vss _01341_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10677_ vdd rf_ram.memory\[393\]\[1\] clknet_leaf_116_clk vss _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06009__C vss _01494_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_360 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08225__A1 vss _03823_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10032__A1 vss _04985_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09973__A1 vss _04921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_771 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05848__C vss _01717_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput208 o_ibus_adr[15] net208 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_142_1210 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput219 o_ibus_adr[25] net219 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_103_1205 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05995__C1 vss _01521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09725__B2 vss net107 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11229_ vdd cpu.bufreg.i_sh_signed clknet_leaf_257_clk vss _00965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06539__A1 vss _02723_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_175_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_175_1041 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06770_ _02904_ vss vdd _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_164_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05721_ _01916_ vdd vss _01917_ rf_ram.memory\[432\]\[0\] _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_136_1036 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10099__A1 vss _05017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_4_clk_I vss clknet_5_1__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05652_ _01848_ _01617_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_76_1193 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08440_ vdd vss _03962_ rf_ram.memory\[175\]\[0\] _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05514__A2 vss _01709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_77 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06711__A1 vss _02826_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05583_ vdd vss _01779_ rf_ram.memory\[297\]\[0\] _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_105_62 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08371_ vdd vss _03918_ rf_ram.memory\[185\]\[1\] _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07322_ vdd _03264_ _03262_ _00251_ _03260_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_293 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09498__S vss _01491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_349 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07253_ vdd _03220_ _03219_ _00226_ _03190_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06204_ _01756_ vdd vss _02399_ rf_ram.memory\[448\]\[1\] _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_121_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07184_ vdd vss _03178_ _02738_ _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07019__A2 vss _03072_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_533 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11620__I vss net70 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1007 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09964__A1 vss _03445_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06135_ _01790_ vdd vss _02330_ _02327_ _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10023__A1 vss _04950_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_333_clk_I vss clknet_5_4__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08767__A2 vss _04152_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06778__A1 vss _02764_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06066_ _02258_ _02259_ _02260_ _01670_ vdd vss _02261_ _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_69_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09716__A1 vss _04781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08519__A2 vss _03949_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09825_ vdd vss _04859_ rf_ram.memory\[249\]\[1\] _04857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06968_ _03040_ vss vdd _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_154_1103 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09756_ _04760_ _04815_ vdd vss _04816_ net117 _04766_ net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__06950__A1 vss _03018_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05919_ rf_ram.memory\[124\]\[0\] _02115_ vss vdd rf_ram.memory\[127\]\[0\] _01786_
+ rf_ram.memory\[125\]\[0\] _01931_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09687_ _04768_ vss vdd _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08707_ vdd vss _04139_ rf_ram.memory\[152\]\[1\] _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06899_ vdd _02994_ _02993_ _00098_ _02970_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_1146 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1233 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08638_ vdd _04096_ _04095_ _00735_ _04094_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05505__A2 vss _01537_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06702__A1 vss _02775_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08569_ vdd vss _04052_ rf_ram.memory\[170\]\[0\] _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10600_ vdd rf_ram.memory\[357\]\[0\] clknet_leaf_155_clk vss _00344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11580_ vdd rf_ram.memory\[207\]\[1\] clknet_leaf_34_clk vss _01312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_293 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_438 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10531_ vdd rf_ram.memory\[266\]\[1\] clknet_leaf_192_clk vss _00275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05269__A1 vss _01363_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_505 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10462_ vdd rf_ram.memory\[273\]\[0\] clknet_leaf_189_clk vss _00206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09404__B1 vss _04539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10393_ vdd rf_ram.memory\[223\]\[1\] clknet_leaf_33_clk vss _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06769__A1 vss _02716_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09707__A1 vss _04781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11014_ vdd rf_ram.memory\[559\]\[0\] clknet_leaf_323_clk vss _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07194__A1 vss _02813_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_330 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06941__A1 vss _02738_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_240_clk vdd vss clknet_leaf_240_clk clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_750 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08694__A1 vss _02983_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05901__C1 vss _01763_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08446__A1 vss _03953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08997__A2 vss _04303_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10729_ vdd rf_ram.memory\[460\]\[1\] clknet_leaf_51_clk vss _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10253__A1 vss _02825_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_959 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10005__A1 vss _04953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09946__A1 vss _04918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07940_ vdd vss _03648_ _02781_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05983__A2 vss _01643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07871_ vdd vss _03606_ rf_ram.memory\[408\]\[1\] _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06822_ vdd vss _02942_ _02909_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06393__C1 vss _01912_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09610_ vdd _04715_ _04714_ _01088_ _04634_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_1255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_231_clk vdd vss clknet_leaf_231_clk clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09541_ _04664_ vdd vss _01070_ _01354_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06753_ vdd vss _02892_ rf_ram.memory\[515\]\[1\] _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05704_ _01629_ vdd vss _01900_ _01898_ _01899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__07488__A2 vss _02815_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09472_ vss _01053_ _04612_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06684_ _02844_ _02843_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_05635_ _01830_ vdd vss _01831_ _01603_ _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08423_ vdd vss _03951_ rf_ram.memory\[173\]\[0\] _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_928 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05566_ _01526_ vdd vss _01762_ rf_ram.memory\[256\]\[0\] _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08354_ vdd vss _03908_ rf_ram.memory\[182\]\[0\] _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_293 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10244__A1 vss _02727_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07305_ vss _03253_ _02940_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__06448__B1 vss _01607_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_298_clk vdd vss clknet_leaf_298_clk clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05497_ _01693_ vss vdd _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08285_ vdd _03864_ _03863_ _00614_ _03852_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_414 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06999__A1 vss _03050_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07236_ vdd vss _03210_ _02806_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_272_clk_I vss clknet_5_16__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07167_ vdd vss _03168_ rf_ram.memory\[483\]\[1\] _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07412__A2 vss _02972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06118_ _01504_ vdd vss _02313_ rf_ram.memory\[262\]\[1\] _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input60_I vss i_ibus_rdt[5] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_1102 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07098_ vdd vss _03124_ _02921_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_287_clk_I vss clknet_5_18__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06049_ vdd vss _02244_ rf_ram.memory\[361\]\[1\] _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05974__A2 vss _01633_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1008 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07176__A1 vss _03157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_210_clk_I vss clknet_5_25__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_222_clk vdd vss clknet_leaf_222_clk clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09808_ vdd vss _04849_ rf_ram.memory\[74\]\[0\] _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09739_ _04804_ vss vdd _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05523__I vss _01686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08676__A1 vss _04097_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_225_clk_I vss clknet_5_23__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_15__f_clk_I vss clknet_3_3_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08428__A1 vss _02822_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11632_ vss net155 net82 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_289_clk vdd vss clknet_leaf_289_clk clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_108_866 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11563_ vdd rf_ram.memory\[20\]\[0\] clknet_leaf_292_clk vss _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_745 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07100__A1 vss _03123_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_296 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07651__A2 vss _03089_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11494_ vdd rf_ram.memory\[296\]\[1\] clknet_leaf_137_clk vss _01226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_1002 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10514_ vdd rf_ram.memory\[270\]\[0\] clknet_leaf_190_clk vss _00258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_650 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09928__A1 vss _04921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_633 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10445_ vdd rf_ram.memory\[484\]\[1\] clknet_leaf_185_clk vss _00189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_672 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_368 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1154 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08600__A1 vss _04058_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10376_ vdd rf_ram.memory\[22\]\[0\] clknet_leaf_209_clk vss _00120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05965__A2 vss _01682_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06303__B vss _01494_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_213_clk vdd vss clknet_leaf_213_clk clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05717__A2 vss _01706_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06914__A1 vss _02775_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06390__A2 vss _01808_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_722 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05433__I vss _01563_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08667__A1 vss _02959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1103 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_232 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05420_ _01615_ vdd vss _01616_ rf_ram.memory\[352\]\[0\] _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06142__A2 vss _01799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_427 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10226__A1 vss _05078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05351_ _01546_ vdd vss _01547_ _01495_ _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09467__I0 vss net83 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_967 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09092__A1 vss net238 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_279 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_482 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05248__A4 vss _01388_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05282_ cpu.alu.i_rs1 _01480_ _01342_ vss _01479_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_08070_ vdd _03731_ _03730_ _00532_ _03721_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09919__A1 vss _04884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07021_ vdd _03074_ _03073_ _00140_ _03050_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_70_299 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06213__B vss _01693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08972_ vdd vss _04304_ _03071_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05608__I vss _01640_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05956__A2 vss _01508_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07923_ vdd vss _03638_ rf_ram.memory\[441\]\[1\] _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07158__A1 vss _03161_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07854_ vdd vss _03596_ rf_ram.memory\[430\]\[0\] _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_204_clk vdd vss clknet_leaf_204_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05169__B1 vss _01367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05708__A2 vss _01634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06805_ _02930_ _02825_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07785_ vdd _03552_ _03551_ _00426_ _03521_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06381__A2 vss _01531_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_834 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09524_ vdd vss _04652_ _01419_ _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05343__I vss _01516_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06736_ vdd _02879_ _02878_ _00050_ _02873_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06667_ vdd vss _02831_ _02736_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_94_815 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09455_ vss _01045_ _04603_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05618_ _01813_ vdd vss _01814_ _01600_ _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_137_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06133__A2 vss _01787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07330__A1 vss _03257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08406_ vdd vss _03940_ rf_ram.memory\[178\]\[0\] _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05892__A1 vss _01972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09386_ _04564_ net216 vdd vss _04566_ net215 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06598_ vdd vss _02776_ _02766_ _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_268 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05549_ rf_ram.memory\[283\]\[0\] _01744_ vdd vss _01745_ rf_ram.memory\[282\]\[0\]
+ _01687_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08337_ vdd vss _03897_ rf_ram.memory\[240\]\[0\] _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_403 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_91_clk_I vss clknet_5_11__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08830__A1 vss net246 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08268_ vdd vss _03854_ rf_ram.memory\[197\]\[0\] _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07219_ vdd vss _03200_ rf_ram.memory\[260\]\[1\] _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10230_ vdd vss _05108_ rf_ram.memory\[237\]\[0\] _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08199_ vdd vss _03811_ _03798_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_14_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06123__B vss _01349_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10161_ vdd _05065_ _05063_ _01290_ _05049_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10092_ vdd _05023_ _05022_ _01263_ _05014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05518__I vss _01513_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08897__A1 vss net243 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1103 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_164_clk_I vss clknet_5_27__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06109__C1 vss _01625_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10994_ vdd rf_ram.memory\[539\]\[0\] clknet_leaf_313_clk vss _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08649__A1 vss _04094_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_44_clk_I vss clknet_5_12__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09310__A2 vss _04013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06124__A2 vss _02306_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_325 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_179_clk_I vss clknet_5_29__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10208__A1 vss _05081_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_904 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11615_ vss net168 net95 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_170_728 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07624__A2 vss _03089_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_994 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11546_ vdd rf_ram.memory\[475\]\[1\] clknet_leaf_44_clk vss _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_59_clk_I vss clknet_5_9__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_102_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05635__A1 vss _01603_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11477_ vdd rf_ram.memory\[337\]\[0\] clknet_leaf_168_clk vss _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_666 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_992 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10428_ vdd rf_ram.memory\[488\]\[0\] clknet_leaf_184_clk vss _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10359_ vdd rf_ram.memory\[27\]\[1\] clknet_leaf_210_clk vss _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06033__B vss _01505_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_117_clk_I vss clknet_5_14__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05938__A2 vss _01513_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05428__I vss _01518_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07560__A1 vss _03393_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07570_ vdd _03418_ _03416_ _00345_ _03393_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_163 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06521_ cpu.state.cnt_r\[3\] cpu.state.cnt_r\[2\] vdd vss _02709_ cpu.state.cnt_r\[1\]
+ cpu.state.cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_09240_ vdd _04470_ _04468_ _00963_ _04466_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06115__A2 vss _01755_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07312__A1 vss _02904_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_859 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_325 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07863__A2 vss _02869_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06452_ rf_ram.memory\[61\]\[1\] _01609_ _01633_ rf_ram.memory\[60\]\[1\] _02647_
+ vss vdd rf_ram.memory\[63\]\[1\] _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__06666__A3 vss _02730_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_904 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_961 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09171_ vdd _04427_ _04425_ _00937_ _04401_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06383_ _02577_ vdd vss _02578_ _01972_ _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09065__A1 vss net237 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05403_ _01346_ _01598_ vdd vss _01599_ _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_17_937 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_797 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07615__A2 vss _03446_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05334_ _01530_ _01499_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08122_ vdd _03763_ _03762_ _00552_ _03754_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_406 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08053_ vdd vss _03720_ rf_ram.memory\[565\]\[1\] _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05265_ _01337_ vdd vss _01464_ _01333_ cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_07004_ vdd _03063_ _03062_ _00134_ _03050_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_1085 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07379__A1 vss _03292_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05196_ _01394_ _01395_ vdd vss _01396_ cpu.decode.opcode\[0\] cpu.decode.opcode\[1\]
+ _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08040__A2 vss _03693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08955_ vdd vss _04293_ rf_ram.memory\[120\]\[0\] _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05929__A2 vss _01922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07906_ vdd vss _03628_ rf_ram.memory\[460\]\[0\] _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08886_ vdd _04250_ _04248_ _00829_ _04237_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input23_I vss i_dbus_rdt[29] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08879__A1 vss _04234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07837_ vdd vss _03585_ rf_ram.memory\[411\]\[0\] _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07551__A1 vss _02909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09540__A2 vss net40 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06354__A2 vss _01614_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1072 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07768_ vdd vss _03542_ rf_ram.memory\[393\]\[0\] _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05562__B1 vss _01654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09507_ vdd vss _04639_ _02958_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_826 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06719_ _02730_ vdd vss _02867_ _02798_ _02729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_07699_ vdd _03499_ _03497_ _00393_ _03491_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06106__A2 vss _01687_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1078 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1044 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1033 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09438_ _04593_ vdd vss _04595_ net69 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_81_306 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09369_ vdd vss _04556_ _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_164_588 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_279 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06118__B vss _01504_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_471 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11400_ _01132_ vdd vss clknet_leaf_227_clk net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08803__A1 vss net243 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_531 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11331_ vdd rf_ram.memory\[279\]\[1\] clknet_leaf_191_clk vss _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05957__B vss _01525_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1140 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11262_ vdd net228 clknet_leaf_251_clk vss _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10213_ vdd _05097_ _05095_ _01310_ _05081_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11193_ vdd rf_ram.memory\[8\]\[1\] clknet_leaf_39_clk vss _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10144_ vdd _05055_ _05054_ _01283_ _05046_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10075_ vdd _05012_ _05011_ _01257_ _04982_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09531__A2 vss net37 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_30__f_clk_I vss clknet_3_7_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_940 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05553__B1 vss _01678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1100 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09295__A1 vss _04463_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10977_ vdd rf_ram.memory\[16\]\[1\] clknet_leaf_289_clk vss _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_196 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08098__A2 vss _03729_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_831 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_566 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09047__A1 vss _04331_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06028__B vss _01505_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_862 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11529_ vdd rf_ram.memory\[30\]\[0\] clknet_leaf_205_clk vss _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1024 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_496 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06281__A1 vss _01951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06542__I vss _02727_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09770__A2 vss _03253_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xload_slew254 net254 _01361_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xload_slew243 net243 vss vdd _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05952_ _01601_ vdd vss _02148_ rf_ram.memory\[56\]\[0\] _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08740_ vdd vss _00774_ _04157_ _04159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05883_ vdd vss _02079_ rf_ram.memory\[73\]\[0\] _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08671_ vdd _04116_ _04114_ _00748_ _04097_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07622_ vdd vss _03451_ rf_ram.memory\[352\]\[1\] _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07533__A1 vss _03389_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_95 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06336__A2 vss _01531_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_647 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_1039 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07553_ vdd _03408_ _03407_ _00338_ _03389_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_645 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11623__I vss net73 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07484_ vdd vss _03366_ rf_ram.memory\[365\]\[0\] _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07836__A2 vss _03559_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_511 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_76_656 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06504_ vdd vss _02695_ _01408_ _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09223_ vdd _04459_ _04457_ _00957_ _04434_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06435_ _02618_ _02629_ net251 vdd vss _02630_ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_133_216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_99_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09154_ vdd vss _04417_ rf_ram.memory\[159\]\[1\] _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08105_ vdd _03752_ _03751_ _00546_ _03721_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06366_ _02560_ vdd vss _02561_ _01951_ _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09085_ vdd vss _04374_ rf_ram.memory\[98\]\[1\] _04372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_114_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08261__A2 vss _02844_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05317_ vdd vss _01513_ _01512_ _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_4_661 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06297_ vdd vss _02492_ rf_ram.memory\[164\]\[1\] _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_141_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05248_ cpu.alu.cmp_r _01388_ vdd vss _01448_ _01442_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_08036_ vdd vss _03710_ rf_ram.memory\[568\]\[0\] _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05179_ vdd vss _00002_ _01377_ _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07772__A1 vss _03008_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09987_ vdd vss _04959_ rf_ram.memory\[503\]\[0\] _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09761__A2 vss net23 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08938_ vdd _04282_ _04280_ _00849_ _04269_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06401__B vss _01746_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08869_ vdd _04240_ _04239_ _00822_ _04234_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output227_I vss net227 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10900_ vdd rf_ram.memory\[184\]\[0\] clknet_leaf_18_clk vss _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_100 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10831_ vdd rf_ram.memory\[541\]\[1\] clknet_leaf_312_clk vss _00575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_314 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_382 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10762_ vdd rf_ram.memory\[466\]\[0\] clknet_leaf_124_clk vss _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_998 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10693_ vdd rf_ram.memory\[434\]\[1\] clknet_leaf_80_clk vss _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_547 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05687__B vss _01693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06263__A1 vss _01350_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11314_ _01047_ vdd vss clknet_leaf_267_clk net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_22_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11245_ vdd rf_ram.memory\[63\]\[1\] clknet_leaf_292_clk vss _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09201__A1 vss _04431_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11176_ vdd rf_ram.memory\[95\]\[0\] clknet_leaf_56_clk vss _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09752__A2 vss net20 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10127_ vdd _05044_ _05043_ _01277_ _05014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10058_ vdd vss _05002_ _02821_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07515__A1 vss _03356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06318__A2 vss _01711_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05526__B1 vss _01721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09268__A1 vss _01418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_976 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06220_ _01790_ vdd vss _02415_ _02412_ _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_182_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08752__I vss _04057_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06151_ _02345_ net253 vdd vss _02346_ _01768_ _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_06082_ _02276_ vdd vss _02277_ _01603_ _02275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09991__A2 vss _02801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09910_ vdd _04910_ _04908_ _01194_ _04887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07754__A1 vss _03521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09841_ vdd vss _01166_ _02714_ _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09772_ vdd _04826_ _04825_ _01139_ _04634_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06984_ _03050_ _03013_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05765__B1 vss _01959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05935_ rf_ram.memory\[45\]\[0\] _01609_ _01633_ rf_ram.memory\[44\]\[0\] _02131_
+ vss vdd rf_ram.memory\[47\]\[0\] _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08723_ vdd _04148_ _04146_ _00768_ _04129_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06309__A2 vss _01683_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05866_ _02004_ vdd vss _02062_ rf_ram.memory\[246\]\[0\] _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08654_ vdd _04106_ _04105_ _00741_ _04094_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07605_ vdd _03440_ _03439_ _00358_ _03422_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05797_ vdd vss _01993_ rf_ram.memory\[161\]\[0\] _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08585_ vdd vss _04063_ rf_ram.memory\[168\]\[1\] _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07536_ vdd vss _03398_ _02728_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_166_628 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1075 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_864 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_147_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_935 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07467_ vdd vss _03354_ rf_ram.memory\[32\]\[1\] _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09206_ vdd _04449_ _04448_ _00950_ _04431_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_8_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_199 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06418_ _01706_ _01911_ rf_ram.memory\[123\]\[1\] _02612_ vdd vss _02613_ rf_ram.memory\[122\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_106_238 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07398_ vdd _03311_ _03310_ _00280_ _03289_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06493__A1 vss _02519_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06349_ rf_ram.memory\[194\]\[1\] _02544_ vss vdd rf_ram.memory\[193\]\[1\] _01725_
+ rf_ram.memory\[195\]\[1\] _01811_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09137_ vdd vss _04407_ rf_ram.memory\[169\]\[0\] _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09068_ vdd vss _04363_ rf_ram.memory\[0\]\[1\] _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07993__A1 vss _03654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_956 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06796__A2 vss _02923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_589 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08019_ vdd _03699_ _03697_ _00513_ _03690_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_5_13__f_clk vdd vss clknet_5_13__leaf_clk clknet_3_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11030_ vdd rf_ram.memory\[89\]\[0\] clknet_leaf_48_clk vss _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06131__B vss _01746_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05220__A2 vss _01418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08170__A1 vss _03787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06720__A2 vss _02867_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10814_ vdd rf_ram.memory\[54\]\[0\] clknet_leaf_297_clk vss _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1148 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_935 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10745_ vdd rf_ram.memory\[456\]\[1\] clknet_leaf_50_clk vss _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_164_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10676_ vdd rf_ram.memory\[393\]\[0\] clknet_leaf_116_clk vss _00420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05287__A2 vss _01484_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_681 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_512 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_821 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_539 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07984__A1 vss _03672_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput209 o_ibus_adr[16] net209 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05995__B1 vss _01517_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11228_ _00964_ cpu.genblk3.csr.o_new_irq vdd vss clknet_leaf_240_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_177_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07736__A1 vss _02813_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11159_ vdd rf_ram.memory\[101\]\[1\] clknet_leaf_66_clk vss _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09489__A1 vss _02690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05720_ vss _01916_ _01550_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_76_1161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05651_ vdd vss _01847_ rf_ram.memory\[468\]\[0\] _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_81_34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08370_ vdd _03917_ _03916_ _00646_ _03884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07321_ vdd vss _03264_ rf_ram.memory\[272\]\[1\] _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05582_ _01778_ _01695_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_18_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07252_ vdd vss _03220_ rf_ram.memory\[41\]\[0\] _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_350 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_653 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_344 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06203_ rf_ram.memory\[453\]\[1\] _01725_ _01724_ rf_ram.memory\[452\]\[1\] _02398_
+ vss vdd rf_ram.memory\[455\]\[1\] _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07183_ vdd _03177_ _03175_ _00199_ _03161_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_895 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06227__A1 vss _01603_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06216__B vss _01746_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06134_ _01786_ rf_ram.memory\[291\]\[1\] vdd vss _02329_ rf_ram.memory\[290\]\[1\]
+ _01785_ _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_60_139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09964__A2 vss _02829_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07975__A1 vss _03651_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06778__A2 vss _02830_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06065_ rf_ram.memory\[370\]\[1\] _02260_ vss vdd rf_ram.memory\[369\]\[1\] _01664_
+ rf_ram.memory\[371\]\[1\] _01519_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_44_1149 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07727__A1 vss _03488_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09824_ vdd _04858_ _04857_ _01159_ _04837_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06967_ vdd vss _03039_ _02797_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_09755_ vdd vss _04815_ _04804_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05918_ vdd vss _02114_ rf_ram.memory\[126\]\[0\] _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06898_ vdd vss _02994_ rf_ram.memory\[280\]\[0\] _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05753__A3 vss _01948_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09686_ _04767_ vss vdd _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08706_ vdd _04138_ _04137_ _00761_ _04126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_764 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1283 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05849_ _02039_ _01350_ _02044_ vdd vss _02045_ _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_08637_ vdd vss _04096_ rf_ram.memory\[162\]\[0\] _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06163__B1 vss _01696_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06702__A2 vss _02846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08568_ vdd vss _04051_ net247 _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_182_929 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07519_ vdd vss _03387_ rf_ram.memory\[322\]\[0\] _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_661 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08499_ vss _04005_ _04004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_10530_ vdd rf_ram.memory\[266\]\[0\] clknet_leaf_192_clk vss _00274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_536 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06466__A1 vss _01903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_333 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05674__C1 vss _01726_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10461_ vdd rf_ram.memory\[474\]\[1\] clknet_leaf_43_clk vss _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_286 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_815 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07966__A1 vss _03654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10392_ vdd rf_ram.memory\[223\]\[0\] clknet_leaf_33_clk vss _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_1216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05965__B vss _01601_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05441__A2 vss _01634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09707__A2 vss net5 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_1015 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11013_ vdd rf_ram.memory\[156\]\[1\] clknet_leaf_3_clk vss _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07194__A2 vss _02832_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1283 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_504 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06941__A2 vss _02972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08143__A1 vss _03754_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_414 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09891__A1 vss _02922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08694__A2 vss _04078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05901__B1 vss _01656_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09643__A1 vss _04637_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_272 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10728_ vdd rf_ram.memory\[460\]\[0\] clknet_leaf_119_clk vss _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_158 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10659_ vdd rf_ram.memory\[398\]\[1\] clknet_leaf_117_clk vss _00403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06209__A1 vss _01368_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07957__A1 vss _02903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05432__A2 vss _01623_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06090__C1 vss _01713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1074 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07709__A1 vss _03491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07870_ vdd _03605_ _03604_ _00458_ _03587_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08382__A1 vss _03919_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05166__I vss _01347_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06821_ vss _02941_ _02940_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__06393__B1 vss _01925_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09540_ net40 _04650_ cpu.csr_imm vdd vss _04664_ _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06752_ vdd _02891_ _02890_ _00054_ _02873_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05703_ rf_ram.memory\[410\]\[0\] _01899_ vss vdd rf_ram.memory\[409\]\[0\] _01721_
+ rf_ram.memory\[411\]\[0\] _01726_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09471_ _04604_ vdd vss _04612_ net85 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_148_403 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_548 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08422_ vdd vss _03950_ net243 _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06683_ vdd vss _02843_ _02750_ _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_153_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05634_ rf_ram.memory\[486\]\[0\] _01830_ vss vdd rf_ram.memory\[485\]\[0\] _01678_
+ rf_ram.memory\[487\]\[0\] _01688_ _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_19_615 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06696__A1 vss _02826_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05565_ rf_ram.memory\[261\]\[0\] _01668_ _01509_ rf_ram.memory\[260\]\[0\] _01761_
+ vss vdd rf_ram.memory\[263\]\[0\] _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08353_ vdd vss _03907_ _03008_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09634__A1 vss _04524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10244__A2 vss _02958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07304_ vdd _03252_ _03250_ _00245_ _03225_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08284_ vdd vss _03864_ rf_ram.memory\[204\]\[0\] _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11631__I vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07235_ vdd _03209_ _03207_ _00219_ _03193_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05496_ _01692_ vss vdd _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_171_472 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_81_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09398__B1 vss _04564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05671__A2 vss _01808_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07166_ vdd _03167_ _03166_ _00192_ _03157_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06117_ _01629_ vdd vss _02312_ _02310_ _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07948__A1 vss _03651_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07097_ vss _03123_ _03013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__05423__A2 vss _01606_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06048_ _01615_ vdd vss _02243_ rf_ram.memory\[360\]\[1\] _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06081__C1 vss _01702_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input53_I vss i_ibus_rdt[28] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06620__A1 vss _02723_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09807_ vdd vss _04848_ _02774_ _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07999_ _03685_ _02742_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09738_ vdd vss _04803_ _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_119_1043 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_403 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09669_ _04752_ vdd vss _04753_ _04737_ _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09873__A1 vss _02713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_209 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06687__A1 vss _02844_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05895__C1 vss _01773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09625__A1 vss _04637_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_581 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_570 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08428__A2 vss _02869_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11631_ vss net154 net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_166_277 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11562_ vdd rf_ram.memory\[447\]\[1\] clknet_leaf_79_clk vss _01294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_856 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10513_ vdd rf_ram.memory\[254\]\[1\] clknet_leaf_217_clk vss _00257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_681 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_1041 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11493_ vdd rf_ram.memory\[296\]\[0\] clknet_leaf_137_clk vss _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_826 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_load_slew243_I vss _02843_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_656 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_196 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1025 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05662__A2 vss _01787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10444_ vdd rf_ram.memory\[484\]\[0\] clknet_leaf_186_clk vss _00188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_3_clk_I vss clknet_5_1__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07939__A1 vss _03622_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10375_ vdd rf_ram.memory\[230\]\[1\] clknet_leaf_279_clk vss _00119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_1057 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10171__A1 vss _05049_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05178__A1 vss _01369_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06914__A2 vss _02801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_846 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08667__A2 vss _04078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_332_clk_I vss clknet_5_4__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06678__A1 vss _02836_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_902 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157_299 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05350_ _01542_ _01545_ vdd vss _01546_ _01535_ _01541_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09467__I1 vss net84 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09092__A2 vss _04339_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05638__C1 vss _01636_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_995 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_697 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05281_ vdd vss _01479_ _01342_ _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_656 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05653__A2 vss _01785_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07020_ vdd vss _03074_ rf_ram.memory\[245\]\[0\] _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_689 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_556 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06063__C1 vss _01519_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06602__A1 vss _02748_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08971_ _04303_ vss vdd _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_07922_ vdd _03637_ _03636_ _00478_ _03619_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05810__C1 vss _01679_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07853_ vdd vss _03595_ _02971_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08355__A1 vss _03884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05169__A1 vss _01353_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06804_ vdd _02929_ _02928_ _00068_ _02927_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11626__I vss net76 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1004 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07784_ vdd vss _03552_ rf_ram.memory\[416\]\[0\] _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08107__A1 vss _03724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_78_334 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06735_ vdd vss _02879_ rf_ram.memory\[517\]\[0\] _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09855__A1 vss _02713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09523_ vdd vss _04651_ _03992_ net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_531 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06669__A1 vss _02829_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_367 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06666_ _02730_ vdd vss _02830_ cpu.immdec.imm11_7\[3\] cpu.immdec.imm11_7\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_09454_ _04593_ vdd vss _04603_ net77 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05617_ _01807_ _01809_ _01812_ _01658_ vdd vss _01813_ _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_137_929 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08405_ vdd vss _03939_ net236 _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09385_ vdd vss _04565_ _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_176_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08336_ vdd vss _03896_ _03309_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_5_7__f_clk_I vss clknet_3_1_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06597_ _02775_ net247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09607__A1 vss _04643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05548_ vdd vss _01744_ rf_ram.memory\[281\]\[0\] _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_140_clk vdd vss clknet_leaf_140_clk clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08830__A2 vss _02832_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05479_ _01675_ _01602_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07094__A1 vss _03087_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08267_ vdd vss _03853_ _03230_ _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06841__A1 vss _02935_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07218_ vdd _03199_ _03198_ _00212_ _03190_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_859 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05644__A2 vss _01509_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08198_ vdd _03810_ _03808_ _00581_ _03790_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07149_ vdd vss _03156_ rf_ram.memory\[497\]\[1\] _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06404__B vss _01602_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10160_ vdd vss _05065_ rf_ram.memory\[44\]\[1\] _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10091_ vdd vss _05023_ rf_ram.memory\[310\]\[0\] _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08346__A1 vss _02731_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_1029 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08897__A2 vss _03547_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1126 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06109__B1 vss _01678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10993_ vdd rf_ram.memory\[529\]\[1\] clknet_leaf_308_clk vss _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_962 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05883__A2 vss _01918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11614_ vss net167 net94 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_409 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_131_clk vdd vss clknet_leaf_131_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11545_ vdd rf_ram.memory\[475\]\[0\] clknet_leaf_44_clk vss _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11476_ vdd rf_ram.memory\[338\]\[1\] clknet_leaf_175_clk vss _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06293__C1 vss _01610_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1119 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_407 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10427_ vdd rf_ram.memory\[501\]\[1\] clknet_leaf_220_clk vss _00171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_870 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06314__B vss _01916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10358_ vdd rf_ram.memory\[27\]\[0\] clknet_leaf_210_clk vss _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_687 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06060__A2 vss _01500_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10289_ vdd rf_ram.memory\[476\]\[1\] clknet_leaf_121_clk vss _00033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_1141 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10144__A1 vss _05046_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_198_clk vdd vss clknet_leaf_198_clk clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_178_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06899__A1 vss _02970_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_109 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05444__I vss _01499_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_271_clk_I vss clknet_5_16__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05571__A1 vss _01674_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09837__A1 vss cpu.mem_bytecnt\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_687 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_153 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06520_ _02708_ vdd vss _00004_ _02700_ _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_518 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07312__A2 vss _03253_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06451_ vdd vss _02646_ rf_ram.memory\[62\]\[1\] _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_710 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10937__D vss cpu.o_wdata0 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1162 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05402_ vdd vss _01598_ _01347_ _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_286_clk_I vss clknet_5_18__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09170_ vdd vss _04427_ rf_ram.memory\[86\]\[1\] _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06382_ rf_ram.memory\[77\]\[1\] _01912_ _01649_ rf_ram.memory\[76\]\[1\] _02577_
+ vss vdd rf_ram.memory\[79\]\[1\] _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09065__A2 vss _03945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05874__A2 vss _01863_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_122_clk vdd vss clknet_leaf_122_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06208__C vss net254 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07076__A1 vss _03092_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05333_ _01528_ vdd vss _01529_ rf_ram.memory\[520\]\[0\] _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08121_ vdd vss _03763_ rf_ram.memory\[552\]\[0\] _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_154_781 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05626__A2 vss _01626_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06284__C1 vss _01911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08052_ vdd _03719_ _03718_ _00526_ _03686_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05264_ vdd vss _01462_ _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07003_ vdd vss _03063_ rf_ram.memory\[224\]\[0\] _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06036__C1 vss _01539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05195_ cpu.decode.opcode\[1\] vdd vss _01395_ cpu.decode.opcode\[2\] cpu.decode.opcode\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_clkbuf_leaf_224_clk_I vss clknet_5_22__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_1085 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08954_ vdd vss _04292_ _02991_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07905_ vdd vss _03627_ _02787_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08885_ vdd vss _04250_ rf_ram.memory\[419\]\[1\] _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_189_clk vdd vss clknet_leaf_189_clk clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07836_ vdd vss _03584_ _02822_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05354__I vss _01525_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_239_clk_I vss clknet_5_21__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07767_ vdd vss _03541_ _02752_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input16_I vss i_dbus_rdt[22] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07551__A2 vss _02997_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1095 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09506_ vdd _04638_ _04635_ _01061_ _04637_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06718_ _02866_ _02865_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_07698_ vdd vss _03499_ rf_ram.memory\[382\]\[1\] _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08500__A1 vss _02953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06649_ vdd vss _02817_ rf_ram.memory\[346\]\[0\] _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09437_ vss _01036_ _04594_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09368_ _04552_ net207 vdd vss _04556_ net206 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_113_clk vdd vss clknet_leaf_113_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_118_995 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09299_ vdd vss _04515_ rf_ram.memory\[66\]\[0\] _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07067__A1 vss _02915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08319_ vdd vss _03885_ _03309_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_144_280 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06814__A1 vss _02935_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11330_ vdd rf_ram.memory\[279\]\[0\] clknet_leaf_191_clk vss _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08803__A2 vss _03945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05529__I vss _01714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08567__A1 vss _04026_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_max_cap253_I vss _01568_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06290__A2 vss _01799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11261_ _00996_ vdd vss clknet_leaf_250_clk net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_output84_I vss net84 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1197 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_659 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10212_ vdd vss _05097_ rf_ram.memory\[442\]\[1\] _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11192_ vdd rf_ram.memory\[8\]\[0\] clknet_leaf_39_clk vss _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06042__A2 vss _01606_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10143_ vdd vss _05055_ rf_ram.memory\[452\]\[0\] _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08319__A1 vss _03309_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10074_ vdd vss _05012_ rf_ram.memory\[308\]\[0\] _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09819__A1 vss _04837_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10976_ vdd rf_ram.memory\[16\]\[0\] clknet_leaf_289_clk vss _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_156 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05856__A2 vss _01940_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_104_clk vdd vss clknet_leaf_104_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_25_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11528_ vdd rf_ram.memory\[350\]\[1\] clknet_leaf_168_clk vss _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06044__B vss _01615_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11459_ vdd rf_ram.memory\[345\]\[0\] clknet_leaf_167_clk vss _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08558__A1 vss _02865_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05439__I vss _01518_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06018__C1 vss _01521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07230__A1 vss _03193_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06033__A2 vss _01502_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input8_I vss i_dbus_rdt[15] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xload_slew244 net244 _02821_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10117__A1 vss _05014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05951_ _02146_ vdd vss _02147_ _01526_ _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05882_ _01551_ vdd vss _02078_ rf_ram.memory\[72\]\[0\] _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08670_ vdd vss _04116_ rf_ram.memory\[157\]\[1\] _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07621_ vdd _03450_ _03449_ _00364_ _03422_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_90_clk_I vss clknet_5_11__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_1007 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08730__A1 vss _03134_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_637 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07552_ vdd vss _03408_ rf_ram.memory\[31\]\[0\] _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06503_ vdd vss _02694_ cpu.state.init_done cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07483_ vdd vss _03365_ _02844_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07297__A1 vss _03222_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_134 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_342 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09222_ vdd vss _04459_ rf_ram.memory\[349\]\[1\] _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_748 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06434_ _02628_ vdd vss _02629_ _01350_ _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__05847__A2 vss _01801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1152 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07049__A1 vss _03092_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09153_ vdd _04416_ _04415_ _00930_ _04397_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_510 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06365_ rf_ram.memory\[231\]\[1\] _01959_ _01940_ rf_ram.memory\[230\]\[1\] _02560_
+ vss vdd rf_ram.memory\[229\]\[1\] _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_146_1028 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05316_ vdd vss _01512_ _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
X_08104_ vdd vss _03752_ rf_ram.memory\[555\]\[0\] _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_565 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09084_ vdd _04373_ _04372_ _00904_ _04364_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06296_ _02490_ _01362_ vdd vss _02491_ _01674_ _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA_clkbuf_leaf_163_clk_I vss clknet_5_30__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05247_ vdd vss _01342_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__06272__A2 vss _01515_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08035_ vdd vss _03709_ _02991_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05178_ _01378_ vdd vss _01379_ _01369_ rf_ram.rdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_13_996 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07221__A1 vss _02752_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_43_clk_I vss clknet_5_13__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06024__A2 vss _01524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07772__A2 vss _03496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09986_ vdd vss _04958_ _02915_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10108__A1 vss rf_ram.memory\[312\]\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08937_ vdd vss _04282_ rf_ram.memory\[399\]\[1\] _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_178_clk_I vss clknet_5_31__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08868_ vdd vss _04240_ rf_ram.memory\[130\]\[0\] _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07819_ vdd vss _03574_ rf_ram.memory\[413\]\[1\] _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_58_clk_I vss clknet_5_9__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08721__A1 vss _04126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1205 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_101_clk_I vss clknet_5_14__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05535__A1 vss _01368_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08799_ vdd vss _04197_ rf_ram.memory\[140\]\[0\] _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10830_ vdd rf_ram.memory\[541\]\[0\] clknet_leaf_274_clk vss _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10761_ vdd rf_ram.memory\[477\]\[1\] clknet_leaf_120_clk vss _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_334_clk vdd vss clknet_leaf_334_clk clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_164_331 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10692_ vdd rf_ram.memory\[434\]\[0\] clknet_leaf_81_clk vss _00436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_116_clk_I vss clknet_5_14__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05838__A2 vss _01531_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_156 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_578 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_329 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07739__I vss _03359_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05968__B vss _01493_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11313_ _01046_ vdd vss clknet_leaf_263_clk net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11244_ vdd rf_ram.memory\[63\]\[0\] clknet_leaf_292_clk vss _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07474__I vss _02747_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11175_ vdd rf_ram.memory\[96\]\[1\] clknet_leaf_63_clk vss _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10126_ vdd vss _05044_ rf_ram.memory\[475\]\[0\] _05043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05774__A1 vss _01951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10057_ vdd _05001_ _04999_ _01250_ _04985_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_410 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05722__I vss _01514_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07279__A1 vss _03225_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10959_ vdd rf_ram.memory\[49\]\[1\] clknet_leaf_297_clk vss _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_325_clk vdd vss clknet_leaf_325_clk clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06487__C1 vss _01714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_167 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_116_707 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06239__C1 vss _01931_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08779__A1 vss _04167_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05878__B vss _01597_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06150_ _02344_ vdd vss _02345_ _01600_ _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_102_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06254__A2 vss _01724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07451__A1 vss _03323_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06081_ vss vdd rf_ram.memory\[341\]\[1\] _01702_ rf_ram.memory\[343\]\[1\] _01688_
+ _01623_ rf_ram.memory\[342\]\[1\] _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_0_1082 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_760 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07203__A1 vss _03161_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_782 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1180 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06006__A2 vss _01523_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09840_ _02714_ vdd vss _01165_ _04867_ _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06983_ vdd _03049_ _03047_ _00127_ _03018_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08951__A1 vss _04266_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09771_ vdd vss _04826_ rf_ram.memory\[269\]\[0\] _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05934_ vdd vss _02130_ rf_ram.memory\[46\]\[0\] _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08722_ vdd vss _04148_ rf_ram.memory\[89\]\[1\] _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08703__A1 vss _04129_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_935 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11634__I vss net84 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08653_ vdd vss _04106_ rf_ram.memory\[160\]\[0\] _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05865_ _02057_ _02060_ vdd vss _02061_ _02049_ _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07604_ vdd vss _03440_ rf_ram.memory\[314\]\[0\] _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08584_ _04062_ _04061_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05796_ _01956_ vdd vss _01992_ rf_ram.memory\[160\]\[0\] _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07535_ vdd _03397_ _03395_ _00331_ _03393_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_316_clk vdd vss clknet_leaf_316_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_123 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07466_ vdd _03353_ _03352_ _00306_ _03323_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06417_ vdd vss _02612_ rf_ram.memory\[121\]\[1\] _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_92_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09205_ vdd vss _04449_ rf_ram.memory\[6\]\[0\] _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07397_ vdd vss _03311_ rf_ram.memory\[248\]\[0\] _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06348_ _01650_ vdd vss _02543_ rf_ram.memory\[192\]\[1\] _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09136_ vdd vss _04406_ net249 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06245__A2 vss _01922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09067_ vdd _04362_ _04361_ _00898_ _04331_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_535 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06279_ vdd vss _02474_ rf_ram.memory\[148\]\[1\] _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08018_ vdd vss _03699_ rf_ram.memory\[572\]\[1\] _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06412__B vss _01916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09969_ vdd vss _04947_ _03672_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05508__A1 vss _01603_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_579 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06181__A1 vss _01600_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10813_ vdd rf_ram.memory\[550\]\[1\] clknet_leaf_318_clk vss _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_307_clk vdd vss clknet_leaf_307_clk clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_94_240 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_476 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10744_ vdd rf_ram.memory\[456\]\[0\] clknet_leaf_49_clk vss _00488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_180_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07681__A1 vss _03458_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_301 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10675_ vdd rf_ram.memory\[394\]\[1\] clknet_leaf_113_clk vss _00419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06484__A2 vss _01640_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1034 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07469__I vss _02742_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07433__A1 vss _03326_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_518 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_570 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1089 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_181 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07984__A2 vss _02866_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_719 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09186__A1 vss _04431_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11227_ vdd rf_ram.memory\[319\]\[1\] clknet_leaf_153_clk vss _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07736__A2 vss _03496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08933__A1 vss _04269_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11158_ vdd rf_ram.memory\[101\]\[0\] clknet_leaf_66_clk vss _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10109_ vdd _05033_ _05031_ _01270_ _05017_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11089_ vdd rf_ram.memory\[128\]\[0\] clknet_leaf_25_clk vss _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05650_ _01846_ vss vdd _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05581_ _01777_ _01686_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_169_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07320_ vdd _03263_ _03262_ _00250_ _03257_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_85_251 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_470 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_684 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07672__A1 vss _02904_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07251_ vdd vss _03219_ _02752_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_1071 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06475__A2 vss _01530_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06202_ _01805_ vdd vss _02397_ rf_ram.memory\[454\]\[1\] _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07182_ vdd vss _03177_ rf_ram.memory\[1\]\[1\] _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_1100 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07424__A1 vss _03319_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06133_ vdd vss _02328_ rf_ram.memory\[289\]\[1\] _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_131_529 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_941 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06064_ _01526_ vdd vss _02259_ rf_ram.memory\[368\]\[1\] _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__11629__I vss net79 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_286 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08924__A1 vss _02838_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09823_ vdd vss _04858_ rf_ram.memory\[249\]\[0\] _04857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06966_ vdd _03038_ _03036_ _00121_ _03018_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09754_ vdd vss _04814_ _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05917_ _01928_ vdd vss _02113_ _02110_ _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06897_ vdd vss _02993_ _02958_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05790__C vss _01349_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09685_ _04733_ vdd vss _04766_ _04739_ _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_20_1194 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08705_ vdd vss _04138_ rf_ram.memory\[152\]\[0\] _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_93_clk vdd vss clknet_leaf_93_clk clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05848_ _02041_ _02042_ _02043_ _01717_ vdd vss _02044_ _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_90_1115 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08636_ vdd vss _04095_ _02893_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09101__A1 vss _04367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08567_ vdd _04050_ _04048_ _00710_ _04026_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05779_ _01974_ vdd vss _01975_ _01972_ _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07518_ vdd vss _03386_ _03319_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08498_ vdd vss _04004_ _02736_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_175_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07663__A1 vss _03455_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07449_ vdd vss _03343_ _02946_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05674__B1 vss _01725_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10460_ vdd rf_ram.memory\[474\]\[0\] clknet_leaf_43_clk vss _00204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06407__B vss _01660_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_788 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_1077 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05311__B vss _01506_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_885 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06218__A2 vss _01787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09119_ vdd _04394_ _04393_ _00918_ _04364_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_220 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10391_ vdd rf_ram.memory\[224\]\[1\] clknet_leaf_275_clk vss _00135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_754 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06921__I vss _03008_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06142__B vss _01602_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08915__A1 vss _04266_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11012_ vdd rf_ram.memory\[156\]\[0\] clknet_leaf_29_clk vss _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_84_clk vdd vss clknet_leaf_84_clk clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09340__B2 vss net213 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09340__A1 vss cpu.ctrl.pc vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09891__A2 vss _03035_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08583__I vss _02747_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_481 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10727_ vdd rf_ram.memory\[444\]\[1\] clknet_leaf_54_clk vss _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06457__A2 vss _01661_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06317__B vss _01505_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07406__A1 vss _03100_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10658_ vdd rf_ram.memory\[398\]\[0\] clknet_leaf_117_clk vss _00402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06209__A2 vss _02376_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10589_ vdd rf_ram.memory\[360\]\[1\] clknet_leaf_159_clk vss _00333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07957__A2 vss _03158_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05875__C vss _01860_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06090__B1 vss _01715_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09159__A1 vss _04397_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_177_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08906__A1 vss _04237_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05447__I vss _01508_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06820_ vdd vss _02940_ _02799_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__05196__A2 vss cpu.decode.opcode\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_45 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06751_ vdd vss _02891_ rf_ram.memory\[515\]\[0\] _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05702_ _01615_ vdd vss _01898_ rf_ram.memory\[408\]\[0\] _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_75_clk vdd vss clknet_leaf_75_clk clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06682_ vdd _02842_ _02840_ _00033_ _02826_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_516 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09470_ vss _01052_ _04611_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08421_ _03949_ vss vdd _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_25_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_175_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_426 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05633_ vdd vss _01829_ rf_ram.memory\[484\]\[0\] _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05353__C1 vss _01520_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_640 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05564_ _01504_ vdd vss _01760_ rf_ram.memory\[262\]\[0\] _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08352_ vdd _03906_ _03904_ _00639_ _03887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07645__A1 vss _03458_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05495_ _01629_ vdd vss _01691_ _01685_ _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07303_ vdd vss _03252_ rf_ram.memory\[258\]\[1\] _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06448__A2 vss _01661_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08283_ vdd vss _03863_ _03230_ _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07234_ vdd vss _03209_ rf_ram.memory\[423\]\[1\] _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_788 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05131__B vss cpu.decode.co_ebreak vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_490 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07165_ vdd vss _03167_ rf_ram.memory\[483\]\[0\] _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06116_ rf_ram.memory\[267\]\[1\] _01654_ _01652_ rf_ram.memory\[266\]\[1\] _02311_
+ vss vdd rf_ram.memory\[265\]\[1\] _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07096_ vdd _03122_ _03120_ _00167_ _03092_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08070__A1 vss _03721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06741__I vss net241 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06047_ _01620_ vdd vss _02242_ _02239_ _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06081__B1 vss _01688_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_893 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_112_584 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_869 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input46_I vss i_ibus_rdt[21] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07998_ vdd _03684_ _03682_ _00507_ _03654_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09806_ vdd _04847_ _04845_ _01152_ _04840_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09737_ _04791_ _04802_ vdd vss _04803_ net111 _04790_ net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06949_ vdd vss _03028_ rf_ram.memory\[232\]\[1\] _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_66_clk vdd vss clknet_leaf_66_clk clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_1106 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09668_ vdd net123 _03975_ _04752_ net120 vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09873__A2 vss _01413_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_508 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09599_ _04707_ _04708_ vdd vss _01084_ _04700_ _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__06687__A2 vss _02846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output202_I vss net202 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1049 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08619_ vdd _04084_ _04082_ _00728_ _04062_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05895__B1 vss _01772_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11630_ vss net153 net80 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07636__A1 vss _03008_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11561_ vdd rf_ram.memory\[447\]\[0\] clknet_leaf_53_clk vss _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06439__A2 vss _01613_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10512_ vdd rf_ram.memory\[254\]\[0\] clknet_leaf_220_clk vss _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11492_ vdd rf_ram.memory\[503\]\[1\] clknet_leaf_220_clk vss _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_438 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10443_ vdd rf_ram.memory\[497\]\[1\] clknet_leaf_221_clk vss _00187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_1059 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_696 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08061__A1 vss _03724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10374_ vdd rf_ram.memory\[230\]\[0\] clknet_leaf_278_clk vss _00118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_24__f_clk_I vss clknet_3_6_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08578__I vss _02742_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_57_clk vdd vss clknet_leaf_57_clk clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06127__A1 vss _01769_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_869 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1154 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06678__A2 vss _02839_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07875__A1 vss _03587_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06047__B vss _01620_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05638__B1 vss _01610_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_70_224 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05280_ vdd vss cpu.csr_imm _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_125_175 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05886__B vss _01551_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08052__A1 vss _03686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06063__B1 vss _01664_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08970_ vdd _04302_ _04299_ _00861_ _04301_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05810__B1 vss _01793_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07921_ vdd vss _03637_ rf_ram.memory\[441\]\[0\] _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07852_ vdd _03594_ _03592_ _00451_ _03590_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09552__A1 vss _04478_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06366__A1 vss _01951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10162__A2 vss _02904_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06803_ vdd vss _02929_ rf_ram.memory\[291\]\[0\] _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1043 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput1 vss net1 i_dbus_ack vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_07783_ vdd vss _03551_ net237 _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_48_clk vdd vss clknet_leaf_48_clk clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09522_ vdd vss _04649_ _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_06734_ vdd vss _02878_ _02795_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09855__A2 vss _01418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06669__A2 vss _02832_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05326__C1 vss _01521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09453_ vss _01044_ _04602_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06665_ _02829_ _02828_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_05616_ rf_ram.memory\[312\]\[0\] _01812_ vss vdd rf_ram.memory\[315\]\[0\] _01811_
+ rf_ram.memory\[313\]\[0\] _01810_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_143_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08404_ vdd _03938_ _03936_ _00659_ _03922_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09384_ _04564_ net215 vdd vss _04565_ net214 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07618__A1 vss _03425_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08335_ vdd _03895_ _03893_ _00633_ _03887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06596_ vdd vss _02774_ _02773_ _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05547_ _01684_ vdd vss _01743_ rf_ram.memory\[280\]\[0\] _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_34_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05478_ _01674_ _01349_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08266_ _03852_ _03685_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06841__A2 vss _02954_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07217_ vdd vss _03199_ rf_ram.memory\[260\]\[0\] _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08197_ vdd vss _03810_ rf_ram.memory\[538\]\[1\] _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09268__B vss _01366_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05796__B vss _01956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07148_ vdd _03155_ _03154_ _00186_ _03123_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09791__A1 vss _02945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07079_ vdd _03112_ _03111_ _00160_ _03087_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10090_ vdd vss _05022_ _03445_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08346__A2 vss _02797_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05565__C1 vss _01519_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_39_clk vdd vss clknet_leaf_39_clk clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05580__A2 vss _01692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10992_ vdd rf_ram.memory\[529\]\[0\] clknet_leaf_307_clk vss _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07857__A1 vss _03590_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_215 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05550__I vss _01563_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11613_ vss net166 net93 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_0_clk_I vss clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11544_ vdd rf_ram.memory\[438\]\[1\] clknet_leaf_117_clk vss _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08282__A1 vss _03855_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_224 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11475_ vdd rf_ram.memory\[338\]\[0\] clknet_leaf_175_clk vss _01207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05635__A3 vss _01830_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06293__B1 vss _01608_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10426_ vdd rf_ram.memory\[501\]\[0\] clknet_leaf_220_clk vss _00170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08034__A1 vss _03690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_498 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09782__A1 vss _04634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10357_ vdd rf_ram.memory\[2\]\[1\] clknet_leaf_292_clk vss _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06596__A1 vss _02773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10288_ vdd rf_ram.memory\[476\]\[0\] clknet_leaf_123_clk vss _00032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09534__A1 vss _04526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1197 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05571__A2 vss _01751_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09837__A2 vss _01385_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07848__A1 vss _02813_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_1103 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06450_ _02641_ _02644_ vdd vss _02645_ _02633_ _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_132_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05460__I vss _01655_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_850 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05401_ _01596_ vdd vss _01369_ _01597_ _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_06381_ vdd vss _02576_ rf_ram.memory\[78\]\[1\] _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08273__A1 vss _03230_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_382 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08120_ vdd vss _03762_ _02728_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_1288 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05332_ _01528_ vss vdd _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_43_224 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_1070 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06284__B1 vss _01912_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_909 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08051_ vdd vss _03719_ rf_ram.memory\[565\]\[0\] _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05263_ _01386_ _01461_ vdd vss _01462_ cpu.state.cnt_r\[3\] _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_4_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07002_ vdd vss _03062_ _03055_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08025__A1 vss _02813_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_644 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06036__B1 vss _01540_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05194_ vdd cpu.branch_op _01393_ _01394_ _01380_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06587__A1 vss _02743_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08953_ vdd _04291_ _04289_ _00855_ _04269_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07904_ vdd _03626_ _03624_ _00471_ _03622_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09525__A1 vss _01491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11637__I vss net88 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08884_ vdd _04249_ _04248_ _00828_ _04234_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_83 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07835_ vdd _03583_ _03581_ _00445_ _03557_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07766_ vdd _03540_ _03538_ _00419_ _03524_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05562__A2 vss _01652_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09505_ vdd vss _04638_ rf_ram.memory\[289\]\[1\] _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06717_ vdd vss _02865_ _02779_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_clkbuf_leaf_2_clk_I vss clknet_5_1__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07697_ vdd _03498_ _03497_ _00392_ _03488_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_1058 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08500__A2 vss _04005_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09436_ _04593_ vdd vss _04594_ net68 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06648_ vdd vss _02816_ _02813_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_727 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_146 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06511__A1 vss cpu.alu.i_rs1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09367_ vdd vss _04555_ _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06579_ _02761_ _02760_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_118_963 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09298_ vdd vss _04514_ net239 _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07067__A2 vss _02972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08318_ _03884_ _03685_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_19_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06814__A2 vss _02904_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08249_ vdd vss _03842_ rf_ram.memory\[528\]\[1\] _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06415__B vss _01790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11260_ _00995_ vdd vss clknet_leaf_250_clk net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_clkbuf_leaf_331_clk_I vss clknet_5_1__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1078 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10211_ vdd _05096_ _05095_ _01309_ _05078_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11191_ vdd rf_ram.memory\[90\]\[1\] clknet_leaf_57_clk vss _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_max_cap246_I vss _02780_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06578__A1 vss _02750_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10142_ vdd vss _05054_ _03672_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output77_I vss net77 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10073_ vdd vss _05011_ _03445_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xoutput190 o_ext_rs2[28] net190 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_98_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08319__A2 vss _02923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09516__A1 vss _04524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09017__I vss _04057_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_wire249_I vss _02751_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05553__A2 vss _01634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06750__A1 vss _02881_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10975_ vdd rf_ram.memory\[170\]\[1\] clknet_leaf_8_clk vss _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_124 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_5_0__f_clk vdd vss clknet_5_0__leaf_clk clknet_3_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09687__I vss _04760_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_393 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08255__A1 vss _03823_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11527_ vdd rf_ram.memory\[350\]\[0\] clknet_leaf_168_clk vss _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10062__A1 vss _04985_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_909 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_785 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11458_ vdd rf_ram.memory\[263\]\[1\] clknet_leaf_138_clk vss _01190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_476 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08007__A1 vss _03690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06018__B1 vss _01517_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10409_ vdd rf_ram.memory\[38\]\[1\] clknet_leaf_129_clk vss _00153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08558__A2 vss _03158_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06569__A1 vss _02738_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11389_ _01121_ vdd vss clknet_leaf_225_clk net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_68_69 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09507__A1 vss _02958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05241__A1 vss _01343_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xload_slew245 net245 _02812_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05950_ rf_ram.memory\[61\]\[0\] _01609_ _01633_ rf_ram.memory\[60\]\[0\] _02146_
+ vss vdd rf_ram.memory\[63\]\[0\] _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__05792__A2 vss _01523_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1036 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_53 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05881_ _02076_ vdd vss _02077_ _01972_ _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07620_ vdd vss _03450_ rf_ram.memory\[352\]\[0\] _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1057 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08730__A2 vss _04152_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05544__A2 vss _01626_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07551_ vdd vss _03407_ _02909_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06502_ _01471_ vdd vss _02693_ cpu.state.cnt_r\[2\] _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07482_ vdd _03364_ _03362_ _00311_ _03360_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09221_ vdd _04458_ _04457_ _00956_ _04431_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06433_ _02626_ _02627_ vdd vss _02628_ _02624_ _02625_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_57_872 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_173_365 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_760 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09152_ vdd vss _04416_ rf_ram.memory\[159\]\[0\] _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08246__A1 vss _03798_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06364_ vdd vss _02559_ rf_ram.memory\[228\]\[1\] _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08103_ vdd vss _03751_ _02780_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05315_ _01511_ _01510_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_163_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_590 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09083_ vdd vss _04373_ rf_ram.memory\[98\]\[0\] _04372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06295_ _02483_ _02486_ _02489_ _01349_ vdd vss _02490_ _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_25_780 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08034_ vdd _03708_ _03706_ _00519_ _03690_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05246_ vdd _01445_ _01443_ _01446_ _01442_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_953 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_1148 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05177_ vdd vss rf_ram.regzero _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__07221__A2 vss _03040_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07845__I vss _03359_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08450__B vss _03967_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09985_ vdd _04957_ _04955_ _01222_ _04953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08936_ vdd _04281_ _04280_ _00848_ _04266_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08867_ vdd vss _04239_ net239 _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07818_ vdd _03573_ _03572_ _00438_ _03554_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_1255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07580__I vss _03359_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08798_ vdd vss _04196_ _02787_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07749_ vdd _03530_ _03529_ _00412_ _03521_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output115_I vss net115 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_614 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08485__A1 vss _03953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10760_ vdd rf_ram.memory\[477\]\[0\] clknet_leaf_120_clk vss _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10691_ vdd rf_ram.memory\[414\]\[1\] clknet_leaf_91_clk vss _00435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09419_ _02707_ vdd vss _04585_ net90 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_168_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_866 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_259 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_680 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09985__A1 vss _04953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_875 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_566 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_869 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06145__B vss _01805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_955 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11312_ _01045_ vdd vss clknet_leaf_265_clk net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA_clkbuf_leaf_270_clk_I vss clknet_5_16__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11243_ vdd rf_ram.memory\[66\]\[1\] clknet_leaf_60_clk vss _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05984__B vss _01525_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11174_ vdd rf_ram.memory\[96\]\[0\] clknet_leaf_62_clk vss _00910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_285_clk_I vss clknet_5_18__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06971__A1 vss _03014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10125_ vdd vss _05043_ net244 _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xclkbuf_leaf_270_clk vdd vss clknet_leaf_270_clk clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10056_ vdd vss _05001_ rf_ram.memory\[34\]\[1\] _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_1306 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05526__A2 vss _01709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_468 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10958_ vdd rf_ram.memory\[49\]\[0\] clknet_leaf_296_clk vss _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_1041 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_535 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_223_clk_I vss clknet_5_29__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06487__B1 vss _01635_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06039__C vss _01362_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10889_ vdd rf_ram.memory\[217\]\[1\] clknet_leaf_301_clk vss _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08228__A1 vss _03820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10035__A1 vss _04982_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_538 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06239__B1 vss _01911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_238_clk_I vss clknet_5_21__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_368 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06080_ vdd vss _02275_ rf_ram.memory\[340\]\[1\] _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_402 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09728__A1 vss net107 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_98 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08400__A1 vss _03892_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05214__A1 vss net134 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06982_ vdd vss _03049_ rf_ram.memory\[426\]\[1\] _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09770_ vdd vss _04825_ net243 _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_3_6_0_clk_I vss clknet_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06962__A1 vss _03035_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05765__A2 vss _01958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_261_clk vdd vss clknet_leaf_261_clk clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05933_ _02117_ _02128_ net251 vdd vss _02129_ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_08721_ vdd _04147_ _04146_ _00767_ _04126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09900__A1 vss _04887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08652_ vdd vss _04105_ net237 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07603_ vdd vss _03439_ _02935_ _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06714__A1 vss _02820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05864_ _02059_ vdd vss _02060_ _01951_ _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_178_446 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06190__A2 vss _01787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_934 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08583_ _04061_ _02747_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05795_ _01990_ vdd vss _01991_ _01552_ _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07534_ vdd vss _03397_ rf_ram.memory\[321\]\[1\] _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07465_ vdd vss _03353_ rf_ram.memory\[32\]\[0\] _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_308 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_168 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06416_ _01916_ vdd vss _02611_ rf_ram.memory\[120\]\[1\] _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09204_ vdd vss _04448_ _02805_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_360 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07396_ vdd vss _03310_ _03309_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09135_ vdd _04405_ _04403_ _00923_ _04401_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06347_ rf_ram.memory\[196\]\[1\] _02542_ vss vdd rf_ram.memory\[199\]\[1\] _01713_
+ rf_ram.memory\[197\]\[1\] _01721_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_72_683 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09066_ vdd vss _04362_ rf_ram.memory\[0\]\[0\] _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06278_ _01494_ vdd vss _02473_ _02470_ _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05229_ vdd vss _01429_ cpu.alu.i_rs1 cpu.alu.add_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08017_ vdd _03698_ _03697_ _00512_ _03686_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_788 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1232 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1145 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09968_ vdd _04946_ _04944_ _01216_ _04921_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05756__A2 vss _01501_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_252_clk vdd vss clknet_leaf_252_clk clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08919_ vdd vss _04271_ _02794_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output232_I vss net232 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06953__A1 vss _03014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09899_ vdd vss _04904_ rf_ram.memory\[263\]\[1\] _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06166__C1 vss _01702_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05823__I vss _01695_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10812_ vdd rf_ram.memory\[550\]\[0\] clknet_leaf_318_clk vss _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10743_ vdd rf_ram.memory\[43\]\[1\] clknet_leaf_128_clk vss _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05979__B vss _01525_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_403 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06469__B1 vss _01624_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07130__A1 vss _03126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10674_ vdd rf_ram.memory\[394\]\[0\] clknet_leaf_116_clk vss _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06654__I vss _02819_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09958__A1 vss _04921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_741 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_661 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1057 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_763 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08630__A1 vss _02794_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05995__A2 vss _01511_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11226_ vdd rf_ram.memory\[319\]\[0\] clknet_leaf_153_clk vss _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11157_ vdd rf_ram.memory\[102\]\[1\] clknet_leaf_63_clk vss _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_243_clk vdd vss clknet_leaf_243_clk clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05747__A2 vss _01755_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10108_ vdd vss _05033_ rf_ram.memory\[312\]\[1\] _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11088_ vdd rf_ram.memory\[12\]\[1\] clknet_leaf_295_clk vss _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10039_ vdd vss _04991_ rf_ram.memory\[305\]\[0\] _04990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06172__A2 vss _01755_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1027 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1147 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_162_clk_I vss clknet_5_30__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_939 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05580_ _01693_ vdd vss _01776_ rf_ram.memory\[296\]\[0\] _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_98_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10256__A1 vss _02819_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_42_clk_I vss clknet_5_13__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05889__B vss _01978_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07121__A1 vss _02829_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07250_ vdd _03218_ _03216_ _00225_ _03193_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_365 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_190 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09949__A1 vss net248 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_335 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_177_clk_I vss clknet_5_31__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10008__A1 vss _04950_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06201_ _02394_ _02395_ vdd vss _02396_ _02392_ _02393_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__05683__A1 vss _01368_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07181_ vdd _03176_ _03175_ _00198_ _03157_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_823 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07424__A2 vss _02844_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06132_ _01783_ vdd vss _02327_ rf_ram.memory\[288\]\[1\] _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_57_clk_I vss clknet_5_9__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1243 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_100_clk_I vss clknet_5_14__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06063_ rf_ram.memory\[372\]\[1\] _02258_ vss vdd rf_ram.memory\[375\]\[1\] _01519_
+ rf_ram.memory\[373\]\[1\] _01664_ _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__07188__A1 vss _03161_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08924__A2 vss _04038_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09822_ vdd vss _04857_ _03309_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_115_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06935__A1 vss _03018_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09753_ _04760_ _04813_ vdd vss _04814_ net116 _04766_ net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06965_ vdd vss _03038_ rf_ram.memory\[22\]\[1\] _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11645__I vss net126 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08704_ vdd vss _04137_ _02991_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06148__C1 vss _01811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05916_ _01706_ _01911_ rf_ram.memory\[123\]\[0\] _02111_ vdd vss _02112_ rf_ram.memory\[122\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_09684_ _04764_ _04765_ vdd vss _01112_ _04763_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06739__I vss _02845_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08688__A1 vss _02812_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06896_ _02992_ vss vdd _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_167_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05847_ rf_ram.memory\[194\]\[0\] _02043_ vss vdd rf_ram.memory\[193\]\[0\] _01725_
+ rf_ram.memory\[195\]\[0\] _01811_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_08635_ _04094_ _04057_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_167_917 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07360__A1 vss _03257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06163__A2 vss _01687_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_539 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08566_ vdd vss _04050_ rf_ram.memory\[509\]\[1\] _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07517_ vdd _03385_ _03383_ _00325_ _03360_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05910__A2 vss _01915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05778_ rf_ram.memory\[133\]\[0\] _01912_ _01649_ rf_ram.memory\[132\]\[0\] _01974_
+ vss vdd rf_ram.memory\[135\]\[0\] _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_65_904 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08497_ vdd _04003_ _04001_ _00687_ _03956_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_200 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05799__B vss _01494_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07448_ vdd _03342_ _03340_ _00299_ _03326_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_696 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1172 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_376 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06320__C1 vss _01931_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07379_ vdd _03299_ _03297_ _00273_ _03292_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_368 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09118_ vdd vss _04394_ rf_ram.memory\[575\]\[0\] _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08612__A1 vss _04058_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10390_ vdd rf_ram.memory\[224\]\[0\] clknet_leaf_275_clk vss _00134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09049_ vdd _04351_ _04349_ _00891_ _04334_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05977__A2 vss _01640_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_377 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07179__A1 vss _02899_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_225_clk vdd vss clknet_leaf_225_clk clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11011_ vdd rf_ram.memory\[157\]\[1\] clknet_leaf_3_clk vss _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06926__A1 vss _02975_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_1038 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05981__C vss _01562_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08679__A1 vss _04094_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09340__A2 vss _03991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06154__A2 vss _01543_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08864__I vss _04061_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_438 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05901__A2 vss _01709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10238__A1 vss _02825_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07103__A1 vss _03126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_786 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_414 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10726_ vdd rf_ram.memory\[444\]\[0\] clknet_leaf_78_clk vss _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10657_ vdd rf_ram.memory\[380\]\[1\] clknet_leaf_106_clk vss _00401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_869 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_688 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_496 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10588_ vdd rf_ram.memory\[360\]\[0\] clknet_leaf_159_clk vss _00332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07406__A2 vss _03135_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06209__A3 vss _02403_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_344 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08603__A1 vss net241 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_552 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_185 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_1043 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1027 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11209_ vdd rf_ram.memory\[83\]\[1\] clknet_leaf_47_clk vss _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_216_clk vdd vss clknet_leaf_216_clk clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07590__A1 vss _03422_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06393__A2 vss _01719_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06750_ vdd vss _02890_ _02881_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05701_ _01896_ vdd vss _01897_ _01603_ _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06681_ vdd vss _02842_ rf_ram.memory\[476\]\[1\] _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06145__A2 vss _01804_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07342__A1 vss _03260_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05632_ _01620_ vdd vss _01828_ _01825_ _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08420_ vdd _03948_ _03946_ _00665_ _03922_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_148_449 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05353__B1 vss _01516_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05563_ _01629_ vdd vss _01759_ _01757_ _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08351_ vdd vss _03906_ rf_ram.memory\[181\]\[1\] _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_172_920 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05494_ _01688_ rf_ram.memory\[347\]\[0\] vdd vss _01690_ rf_ram.memory\[346\]\[0\]
+ _01687_ _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07302_ vdd _03251_ _03250_ _00244_ _03222_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08282_ vdd _03862_ _03860_ _00613_ _03855_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08842__A1 vss _04202_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07233_ vdd _03208_ _03207_ _00218_ _03190_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07164_ vdd vss _03166_ _02889_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06115_ _01756_ vdd vss _02310_ rf_ram.memory\[264\]\[1\] _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07095_ vdd vss _03122_ rf_ram.memory\[502\]\[1\] _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06046_ _01608_ rf_ram.memory\[355\]\[1\] vdd vss _02241_ rf_ram.memory\[354\]\[1\]
+ _01606_ _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_67_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_207_clk vdd vss clknet_leaf_207_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06908__A1 vss _02975_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06369__C1 vss _01636_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_1246 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07997_ vdd vss _03684_ rf_ram.memory\[466\]\[1\] _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06384__A2 vss _01922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ vdd vss _04847_ rf_ram.memory\[75\]\[1\] _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input39_I vss i_ibus_rdt[14] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09570__A2 vss _04678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09736_ vdd vss _04802_ _04781_ net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06948_ vdd _03027_ _03026_ _00114_ _03014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05373__I vss _01568_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09667_ _04750_ _04751_ vdd vss _01109_ _04747_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06136__A2 vss _01735_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06879_ vdd vss _02981_ rf_ram.memory\[301\]\[0\] _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07333__A1 vss _03055_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1044 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1006 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08618_ vdd vss _04084_ rf_ram.memory\[163\]\[1\] _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09873__A3 vss _03989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_747 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09598_ _04700_ vdd vss _04708_ _04478_ cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_49_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08549_ vdd vss _04040_ rf_ram.memory\[119\]\[0\] _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09086__A1 vss _04367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07636__A2 vss _03089_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11560_ vdd rf_ram.memory\[448\]\[1\] clknet_leaf_112_clk vss _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10511_ vdd rf_ram.memory\[271\]\[1\] clknet_leaf_194_clk vss _00255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_975 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11491_ vdd rf_ram.memory\[503\]\[0\] clknet_leaf_221_clk vss _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06932__I vss _02747_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10442_ vdd rf_ram.memory\[497\]\[0\] clknet_leaf_221_clk vss _00186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_1173 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10373_ vdd rf_ram.memory\[231\]\[1\] clknet_leaf_276_clk vss _00117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_371 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_185 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06375__A2 vss _01989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_38_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09077__A1 vss _03668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07627__A2 vss _03452_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08824__A1 vss _04205_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06328__B vss _01551_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10709_ vdd rf_ram.memory\[430\]\[1\] clknet_leaf_97_clk vss _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_931 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_614 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_951 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_51_483 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05458__I vss _01653_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07920_ vdd vss _03636_ _02983_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09001__A1 vss _04301_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07851_ vdd vss _03594_ rf_ram.memory\[410\]\[1\] _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09552__A2 vss net44 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07563__A1 vss _03389_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07782_ vdd _03550_ _03548_ _00425_ _03524_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06802_ vdd vss _02928_ _02801_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput2 vss net2 i_dbus_rdt[0] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_826 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09521_ vdd vss _04649_ _03967_ _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06733_ vdd _02877_ _02874_ _00049_ _02876_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05193__I vss cpu.decode.co_ebreak vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06118__A2 vss _01662_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05326__B1 vss _01517_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09452_ _04593_ vdd vss _04602_ net76 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06664_ vdd vss _02828_ _02779_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05615_ _01811_ _01635_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_93_306 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09068__A1 vss rf_ram.memory\[0\]\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05877__A1 vss _01768_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08403_ vdd vss _03938_ rf_ram.memory\[209\]\[1\] _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09383_ vss _04564_ _04539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_19_403 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06595_ vdd vss _02773_ _01512_ _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__07618__A2 vss _03446_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05546_ _01620_ vdd vss _01742_ _01739_ _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08334_ vdd vss _03895_ rf_ram.memory\[217\]\[1\] _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08009__I vss _03692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05142__B vss _01344_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_644 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_564 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08815__A1 vss net249 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05477_ _01672_ net253 vdd vss _01673_ _01600_ _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_85_1004 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08265_ vdd _03851_ _03849_ _00607_ _03823_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07216_ vdd vss _03198_ _02883_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08196_ vdd _03809_ _03808_ _00580_ _03787_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09240__A1 vss _04466_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07147_ vdd vss _03155_ rf_ram.memory\[497\]\[0\] _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06054__A1 vss _01527_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_872 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05368__I vss _01563_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1060 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07078_ vdd vss _03112_ rf_ram.memory\[492\]\[0\] _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09791__A2 vss _04507_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06029_ rf_ram.memory\[565\]\[1\] _01555_ _01538_ rf_ram.memory\[564\]\[1\] _02224_
+ vss vdd rf_ram.memory\[567\]\[1\] _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_96_1100 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06357__A2 vss _01515_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05565__B1 vss _01668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_303 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06109__A2 vss _01634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07306__A1 vss _02899_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09719_ _04790_ vss vdd _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_10991_ vdd rf_ram.memory\[163\]\[1\] clknet_leaf_338_clk vss _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06927__I vss _02742_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09059__A1 vss _04334_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11612_ vss net165 net92 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_182_547 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08806__A1 vss rf_ram.memory\[13\]\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_19__f_clk vdd vss clknet_5_19__leaf_clk clknet_3_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_65_575 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11543_ vdd rf_ram.memory\[438\]\[0\] clknet_leaf_53_clk vss _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1213 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11474_ vdd rf_ram.memory\[33\]\[1\] clknet_leaf_202_clk vss _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10425_ vdd rf_ram.memory\[48\]\[1\] clknet_leaf_208_clk vss _00169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10356_ vdd rf_ram.memory\[2\]\[0\] clknet_leaf_206_clk vss _00100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10287_ vdd rf_ram.memory\[455\]\[1\] clknet_leaf_122_clk vss _00031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09534__A2 vss net38 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1165 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07545__A1 vss _03393_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06348__A2 vss _01649_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09298__A1 vss net239 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07848__A2 vss _03559_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_864 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_185_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_717 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05400_ vdd vss _01596_ cpu.immdec.imm24_20\[3\] _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06380_ vdd _02575_ _01597_ _01368_ _02547_ vss _02574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_12_1245 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05897__B vss _01684_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08273__A2 vss _02889_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05331_ _01527_ vss vdd _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_56_586 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05262_ vdd vss _01461_ cpu.decode.op26 _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08050_ vdd vss _03718_ _03071_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_45 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07001_ vdd _03061_ _03059_ _00133_ _03053_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05193_ vss _01393_ cpu.decode.co_ebreak vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08025__A2 vss _03693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08952_ vdd vss _04291_ rf_ram.memory\[121\]\[1\] _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08499__I vss _04004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08883_ vdd vss _04249_ rf_ram.memory\[419\]\[0\] _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07903_ vdd vss _03626_ rf_ram.memory\[444\]\[1\] _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07536__A1 vss _02728_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07834_ vdd vss _03583_ rf_ram.memory\[432\]\[1\] _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_1042 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07765_ vdd vss _03540_ rf_ram.memory\[394\]\[1\] _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11653__I vss net103 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_612 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07696_ vdd vss _03498_ rf_ram.memory\[382\]\[0\] _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09504_ _04637_ _04400_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_56_1150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06716_ vdd _02864_ _02862_ _00045_ _02826_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_853 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06647_ vss _02815_ _02814_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09435_ _04593_ _01411_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_59_391 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09366_ _04552_ net206 vdd vss _04555_ net205 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06578_ vdd vss _02760_ _02750_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05529_ vdd vss _01725_ _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_09297_ vdd _04513_ _04511_ _00977_ _04466_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08317_ vdd _03883_ _03881_ _00627_ _03855_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_133_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_625 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08248_ vdd _03841_ _03840_ _00600_ _03820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_921 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10210_ vdd vss _05096_ rf_ram.memory\[442\]\[0\] _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09213__A1 vss _04434_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06027__A1 vss _01495_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08179_ vdd vss _03799_ _03798_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_11190_ vdd rf_ram.memory\[90\]\[0\] clknet_leaf_57_clk vss _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_820 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09764__A2 vss net25 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10141_ vdd _05053_ _05051_ _01282_ _05049_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06431__B vss _01923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput180 o_ext_rs2[19] net180 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10072_ vdd _05010_ _05008_ _01256_ _04985_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput191 o_ext_rs2[29] net191 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09516__A2 vss net57 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05250__A2 vss _01382_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07527__A1 vss _03389_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06750__A2 vss _02889_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10974_ vdd rf_ram.memory\[170\]\[0\] clknet_leaf_336_clk vss _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_823 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_975 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11526_ vdd rf_ram.memory\[308\]\[1\] clknet_leaf_144_clk vss _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06266__A1 vss _01372_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_854 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_753 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwire252 net252 _01734_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_11457_ vdd rf_ram.memory\[263\]\[0\] clknet_leaf_195_clk vss _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09204__A1 vss _02805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_180_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10408_ vdd rf_ram.memory\[38\]\[0\] clknet_leaf_130_clk vss _00152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11388_ _01120_ vdd vss clknet_leaf_224_clk net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09755__A2 vss net21 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07766__A1 vss _03524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10339_ vdd rf_ram.memory\[285\]\[1\] clknet_leaf_180_clk vss _00083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06569__A2 vss _02752_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09507__A2 vss _03083_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07518__A1 vss _03319_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05880_ vss vdd rf_ram.memory\[79\]\[0\] _02019_ rf_ram.memory\[77\]\[0\] _01912_
+ _01755_ rf_ram.memory\[76\]\[0\] _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__08191__A1 vss _03787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07550_ vdd _03406_ _03404_ _00337_ _03393_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06501_ vdd vss _02692_ cpu.ctrl.pc cpu.ctrl.pc_plus_4_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07481_ vdd vss _03364_ rf_ram.memory\[328\]\[1\] _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09220_ vdd vss _04458_ rf_ram.memory\[349\]\[0\] _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09691__A1 vss _04740_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06432_ rf_ram.memory\[98\]\[1\] _02627_ vss vdd rf_ram.memory\[97\]\[1\] _01772_
+ rf_ram.memory\[99\]\[1\] _01857_ _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_115_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_506 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_2_0_clk_I vss clknet_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09151_ vdd vss _04415_ _02908_ _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08246__A2 vss _02946_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06363_ _01494_ vdd vss _02558_ _02555_ _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_185_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05420__B vss _01615_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_539 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09082_ vdd vss _04372_ net239 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10053__A2 vss _02894_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05314_ _01510_ _01509_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08102_ vdd _03750_ _03748_ _00545_ _03724_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_707 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06235__C vss _01670_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08033_ vdd vss _03708_ rf_ram.memory\[56\]\[1\] _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06294_ _01928_ vdd vss _02489_ _02487_ _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_114_477 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05245_ _01444_ vdd vss _01445_ cpu.bne_or_bge _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_943 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput60 vss net60 i_ibus_rdt[5] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05480__A2 vss _01543_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09746__A2 vss net18 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05176_ vdd vss _01377_ _01353_ rf_ram_if.rdata0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07757__A1 vss _02991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11648__I vss net129 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09984_ vdd vss _04957_ rf_ram.memory\[275\]\[1\] _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_122_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08935_ vdd vss _04281_ rf_ram.memory\[399\]\[0\] _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08866_ vdd _04238_ _04235_ _00821_ _04237_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input21_I vss i_dbus_rdt[27] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07817_ vdd vss _03573_ rf_ram.memory\[413\]\[0\] _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_228 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08797_ _04195_ vss vdd _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_07748_ vdd vss _03530_ rf_ram.memory\[377\]\[0\] _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07679_ vdd _03486_ _03485_ _00386_ _03455_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09682__A1 vss _04740_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10690_ vdd rf_ram.memory\[414\]\[0\] clknet_leaf_91_clk vss _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_547 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09418_ vss _01027_ _04584_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09349_ vdd vss _04545_ _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_383 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06426__B vss _01783_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_992 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07996__A1 vss _03651_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07101__I vss _03017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11311_ _01044_ vdd vss clknet_leaf_266_clk net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_120_403 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_792 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05471__A2 vss _01666_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11242_ vdd rf_ram.memory\[66\]\[0\] clknet_leaf_59_clk vss _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11173_ vdd rf_ram.memory\[97\]\[1\] clknet_leaf_70_clk vss _00909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10124_ vdd _05042_ _05040_ _01276_ _05017_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06161__B vss _01693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10055_ vdd _05000_ _04999_ _01249_ _04982_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08173__A1 vss _02881_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07920__A1 vss _02983_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_935 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10957_ vdd rf_ram.regzero clknet_leaf_281_clk vss _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_1097 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10888_ vdd rf_ram.memory\[217\]\[0\] clknet_leaf_301_clk vss _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_865 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_731 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09976__A2 vss _04951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11509_ vdd rf_ram.memory\[326\]\[0\] clknet_leaf_143_clk vss _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_58 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1025 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_1_clk_I vss clknet_5_1__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06411__A1 vss _01909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05466__I vss _01661_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08400__A2 vss _02761_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06981_ vdd _03048_ _03047_ _00126_ _03014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05932_ _02127_ vdd vss _02128_ _01350_ _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_08720_ vdd vss _04147_ rf_ram.memory\[89\]\[0\] _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06962__A2 vss _03009_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08164__A1 vss _03787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08651_ vdd _04104_ _04102_ _00740_ _04097_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05863_ rf_ram.memory\[231\]\[0\] _01959_ _01940_ rf_ram.memory\[230\]\[0\] _02059_
+ vss vdd rf_ram.memory\[229\]\[0\] _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07602_ vdd _03438_ _03436_ _00357_ _03425_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05794_ rf_ram.memory\[167\]\[0\] _01520_ _01989_ rf_ram.memory\[166\]\[0\] _01990_
+ vss vdd rf_ram.memory\[165\]\[0\] _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08582_ vdd _04060_ _04059_ _00715_ _04058_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07533_ vdd _03396_ _03395_ _00330_ _03389_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_1176 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_1238 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_330_clk_I vss clknet_5_1__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_823 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_300 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07464_ vdd vss _03352_ _02921_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_355 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_333 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06415_ _01790_ vdd vss _02610_ _02607_ _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09203_ vdd _04447_ _04445_ _00949_ _04434_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09416__A1 vss _04466_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09134_ vdd vss _04405_ rf_ram.memory\[91\]\[1\] _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07395_ _03309_ vss vdd _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_29_394 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_331 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06346_ _01805_ vdd vss _02541_ rf_ram.memory\[198\]\[1\] _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09065_ vdd vss _04361_ net237 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_71_194 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06277_ _01953_ rf_ram.memory\[147\]\[1\] vdd vss _02472_ rf_ram.memory\[146\]\[1\]
+ _01958_ _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06650__A1 vss _02743_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_868 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05228_ vdd vss _01428_ _01375_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_1200 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08016_ vdd vss _03698_ rf_ram.memory\[572\]\[0\] _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_778 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05159_ _01362_ _01361_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_21_1108 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09967_ vdd vss _04946_ rf_ram.memory\[295\]\[1\] _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08918_ vdd _04270_ _04267_ _00841_ _04269_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08687__I vss _04057_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09898_ vdd _04903_ _04902_ _01189_ _04884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08155__A1 vss _03757_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_414 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07902__A1 vss _03619_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06166__B1 vss _01688_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08849_ vdd _04227_ _04225_ _00815_ _04205_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09655__A1 vss net1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10811_ vdd rf_ram.memory\[551\]\[1\] clknet_leaf_324_clk vss _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10742_ vdd rf_ram.memory\[43\]\[0\] clknet_leaf_131_clk vss _00486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_916 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05677__C1 vss _01811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_949 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_675 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10673_ vdd rf_ram.memory\[376\]\[1\] clknet_leaf_109_clk vss _00417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_18__f_clk_I vss clknet_3_4_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05141__A1 vss _01343_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05692__A2 vss _01787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_399 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07969__A1 vss _03651_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06641__A1 vss _02748_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08630__A2 vss _03765_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11225_ vdd rf_ram.memory\[329\]\[1\] clknet_leaf_152_clk vss _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08394__A1 vss _03922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11156_ vdd rf_ram.memory\[102\]\[0\] clknet_leaf_63_clk vss _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10107_ vdd _05032_ _05031_ _01269_ _05014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11087_ vdd rf_ram.memory\[12\]\[0\] clknet_leaf_295_clk vss _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10038_ vdd vss _04990_ net248 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08146__A1 vss _02888_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09646__A1 vss _01409_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_300 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05668__C1 vss _01778_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07121__A2 vss _02911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_798 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_275 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06200_ rf_ram.memory\[457\]\[1\] _01725_ _01724_ rf_ram.memory\[456\]\[1\] _02395_
+ vss vdd rf_ram.memory\[459\]\[1\] _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09949__A2 vss _02815_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06880__A1 vss _02970_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05683__A2 vss _01845_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07180_ vdd vss _03176_ rf_ram.memory\[1\]\[0\] _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_171_678 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06131_ _01746_ vdd vss _02326_ _02323_ _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06062_ _01504_ vdd vss _02257_ rf_ram.memory\[374\]\[1\] _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06632__A1 vss _02743_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_389 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08385__A1 vss _02959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09821_ vdd _04856_ _04854_ _01158_ _04840_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_158_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09752_ vdd vss _04813_ _04804_ net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08703_ vdd _04136_ _04134_ _00760_ _04129_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06964_ vdd _03037_ _03036_ _00120_ _03014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06148__B1 vss _01810_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05915_ vdd vss _02111_ rf_ram.memory\[121\]\[0\] _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09885__A1 vss _04887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09683_ _04736_ vdd vss _04765_ net1 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08688__A2 vss _04078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06895_ vdd vss _02991_ _02716_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_179_756 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05846_ _01650_ vdd vss _02042_ rf_ram.memory\[192\]\[0\] _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_94_1275 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06699__A1 vss _02820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08634_ vdd _04093_ _04091_ _00734_ _04062_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09840__B vss _02714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08565_ vdd _04049_ _04048_ _00709_ _04023_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05777_ vdd vss _01973_ rf_ram.memory\[134\]\[0\] _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09637__A1 vss _04524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07516_ vdd vss _03385_ rf_ram.memory\[362\]\[1\] _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08496_ vdd vss _04003_ rf_ram.memory\[359\]\[1\] _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_344 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_461 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07447_ vdd vss _03342_ rf_ram.memory\[331\]\[1\] _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_170_clk vdd vss clknet_leaf_170_clk clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06320__B1 vss _01911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_437 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_284_clk_I vss clknet_5_18__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05674__A2 vss _01724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07378_ vdd vss _03299_ rf_ram.memory\[250\]\[1\] _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_150_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_481 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06329_ vdd vss _02524_ rf_ram.memory\[209\]\[1\] _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09117_ vdd vss _04393_ _02908_ _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05426__A2 vss _01614_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09048_ vdd vss _04351_ rf_ram.memory\[103\]\[1\] _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_299_clk_I vss clknet_5_7__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_356 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06423__C vss _01660_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_531 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_1091 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output175_I vss net175 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_518 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07179__A2 vss _02997_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_222_clk_I vss clknet_5_22__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08376__A1 vss _03919_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10183__A1 vss _02916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11010_ vdd rf_ram.memory\[157\]\[0\] clknet_leaf_3_clk vss _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_1006 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1275 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08128__A1 vss _03754_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09876__A1 vss _03309_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_406 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05898__C1 vss _01645_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_119 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09628__A1 vss _04643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08300__A1 vss _03852_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_264 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06665__I vss _02828_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_686 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10725_ vdd rf_ram.memory\[461\]\[1\] clknet_leaf_119_clk vss _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_746 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10656_ vdd rf_ram.memory\[380\]\[0\] clknet_leaf_106_clk vss _00400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_976 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10587_ vdd rf_ram.memory\[321\]\[1\] clknet_leaf_164_clk vss _00331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_140_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08603__A2 vss _04067_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1000 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_391 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06090__A2 vss _01709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11208_ vdd rf_ram.memory\[83\]\[0\] clknet_leaf_47_clk vss _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08367__A1 vss _03887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10174__A1 vss _05046_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11139_ vdd rf_ram.memory\[111\]\[1\] clknet_leaf_72_clk vss _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05744__I vss _01640_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08119__A1 vss _03757_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09867__A1 vss _02838_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05700_ rf_ram.memory\[412\]\[0\] _01896_ vss vdd rf_ram.memory\[415\]\[0\] _01608_
+ rf_ram.memory\[413\]\[0\] _01702_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_06680_ vdd _02841_ _02840_ _00032_ _02820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_155_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05631_ _01696_ rf_ram.memory\[483\]\[0\] vdd vss _01827_ rf_ram.memory\[482\]\[0\]
+ _01777_ _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_86_540 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08350_ vdd _03905_ _03904_ _00638_ _03884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10229__A2 vss _02844_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09619__A1 vss _04643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05562_ vss vdd rf_ram.memory\[265\]\[0\] _01715_ rf_ram.memory\[267\]\[0\] _01654_
+ _01652_ rf_ram.memory\[266\]\[0\] _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_07301_ vdd vss _03251_ rf_ram.memory\[258\]\[0\] _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_152_clk vdd vss clknet_leaf_152_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05493_ vdd vss _01689_ rf_ram.memory\[345\]\[0\] _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_129_675 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08281_ vdd vss _03862_ rf_ram.memory\[194\]\[1\] _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06302__B1 vss _01953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1145 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07232_ vdd vss _03208_ rf_ram.memory\[423\]\[0\] _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06853__A1 vss _02930_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05656__A2 vss _01787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1208 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_971 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_133 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07163_ vdd _03165_ _03163_ _00191_ _03161_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05408__A2 vss _01537_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06114_ _02308_ vdd vss _02309_ _01527_ _02307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_41_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_391 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07094_ vdd _03121_ _03120_ _00166_ _03087_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06045_ vdd vss _02240_ rf_ram.memory\[353\]\[1\] _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_164_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06081__A2 vss _01623_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_726 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08358__A1 vss net235 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09804_ vdd _04846_ _04845_ _01151_ _04837_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06369__B1 vss _01610_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_573 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07996_ vdd _03683_ _03682_ _00506_ _03651_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09735_ vdd vss _04801_ _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06947_ vdd vss _03027_ rf_ram.memory\[232\]\[0\] _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_119_1035 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09666_ _04736_ vdd vss _04751_ net1 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06878_ vdd vss _02980_ _02935_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07333__A2 vss _02917_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08530__A1 vss _04026_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08617_ vdd _04083_ _04082_ _00727_ _04058_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05829_ _01978_ vdd vss _02025_ _02022_ _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09597_ vdd vss _04707_ _03992_ net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08548_ vdd vss _04039_ net235 _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05895__A2 vss _01711_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_143_clk vdd vss clknet_leaf_143_clk clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_119_130 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08479_ _03992_ vss vdd _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_10510_ vdd rf_ram.memory\[271\]\[0\] clknet_leaf_194_clk vss _00254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11490_ vdd rf_ram.memory\[275\]\[1\] clknet_leaf_181_clk vss _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10441_ vdd rf_ram.memory\[485\]\[1\] clknet_leaf_224_clk vss _00185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06057__C1 vss _01646_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_998 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08597__A1 vss _04062_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_380 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10372_ vdd rf_ram.memory\[231\]\[0\] clknet_leaf_276_clk vss _00116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06072__A2 vss _01683_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_884 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10156__A1 vss _05049_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_41_clk_I vss clknet_5_13__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07021__A1 vss _03050_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_176_clk_I vss clknet_5_30__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09849__A1 vss _02713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_56_clk_I vss clknet_5_9__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_838 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08521__A1 vss _03953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_150_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_359 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05886__A2 vss _01537_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09077__A2 vss _02984_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_269 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_134_clk vdd vss clknet_leaf_134_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_55_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10708_ vdd rf_ram.memory\[430\]\[0\] clknet_leaf_101_clk vss _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05638__A2 vss _01644_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_554 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_114_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10639_ vdd rf_ram.memory\[403\]\[1\] clknet_leaf_96_clk vss _00383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_648 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06063__A2 vss _01536_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_129_clk_I vss clknet_5_13__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05810__A2 vss _01677_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10147__A1 vss _03672_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07850_ vdd _03593_ _03592_ _00450_ _03587_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05474__I vss rf_ram.i_raddr\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07012__A1 vss _02738_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07781_ vdd vss _03550_ rf_ram.memory\[437\]\[1\] _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06801_ _02927_ _02819_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_78_1067 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08760__A1 vss _01353_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 vss net3 i_dbus_rdt[10] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09520_ _02709_ vdd vss _04648_ _01419_ _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_06732_ vdd vss _02877_ rf_ram.memory\[518\]\[1\] _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_1219 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_326 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08512__A1 vss _01353_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06663_ vdd _02827_ _02823_ _00029_ _02826_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09451_ vss _01043_ _04601_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_545 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05614_ _01810_ _01714_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_87_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08402_ vdd _03937_ _03936_ _00658_ _03919_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09382_ vdd vss _04563_ _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06594_ vdd _02772_ _02770_ _00015_ _02748_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_188_1022 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_707 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_125_clk vdd vss clknet_leaf_125_clk clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05545_ rf_ram.memory\[275\]\[0\] _01740_ vdd vss _01741_ rf_ram.memory\[274\]\[0\]
+ _01623_ _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__07079__A1 vss _03087_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_370 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_532 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_74_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08333_ vdd _03894_ _03893_ _00632_ _03884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_426 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_228 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_781 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06826__A1 vss _02930_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_111 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05629__A2 vss _01692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06287__C1 vss _01610_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08815__A2 vss _04195_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08264_ vdd vss _03851_ rf_ram.memory\[205\]\[1\] _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05476_ _01659_ _01660_ _01671_ vdd vss _01672_ _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_116_122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1185 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07215_ vdd _03197_ _03195_ _00211_ _03193_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_105_829 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08195_ vdd vss _03809_ rf_ram.memory\[538\]\[0\] _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_851 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07146_ vdd vss _03154_ _02761_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_676 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_30_613 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_158 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07251__A1 vss _02752_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07077_ vdd vss _03111_ _02788_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input51_I vss i_ibus_rdt[26] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06028_ _01505_ vdd vss _02223_ rf_ram.memory\[566\]\[1\] _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05801__A2 vss _01664_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1033 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06211__C1 vss _01773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08751__A1 vss _04129_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07979_ vdd vss _03673_ _03672_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09718_ vdd vss _04789_ _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07306__A2 vss _03253_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10990_ vdd rf_ram.memory\[163\]\[0\] clknet_leaf_339_clk vss _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_523 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09649_ _04736_ vss vdd _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_167_534 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06429__B vss _02004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05868__A2 vss _01683_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05333__B vss _01528_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11611_ vss net164 net91 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_154_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_116_clk vdd vss clknet_leaf_116_clk clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_33_1173 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11542_ vdd rf_ram.memory\[373\]\[1\] clknet_leaf_111_clk vss _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07490__A1 vss _03356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11473_ vdd rf_ram.memory\[33\]\[0\] clknet_leaf_202_clk vss _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06164__B vss _01620_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06293__A2 vss _01606_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10424_ vdd rf_ram.memory\[48\]\[0\] clknet_leaf_208_clk vss _00168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05559__I vss _01613_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_613 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06045__A2 vss _01617_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10355_ vdd rf_ram.memory\[280\]\[1\] clknet_leaf_178_clk vss _00099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10286_ vdd rf_ram.memory\[455\]\[0\] clknet_leaf_112_clk vss _00030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10129__A1 vss _05017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1280 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05294__I vss _01409_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09298__A2 vss _04507_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05859__A2 vss _01664_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_830 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_107_clk vdd vss clknet_leaf_107_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06808__A1 vss _02801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_921 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07949__I vss _03359_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_885 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05330_ _01526_ vss vdd _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__06269__C1 vss _01953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1273 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_77 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_209 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06284__A2 vss _01799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05261_ vss _01460_ cpu.decode.op22 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_24_473 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_974 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07000_ vdd vss _03061_ rf_ram.memory\[225\]\[1\] _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05192_ vdd vss _01392_ _01391_ net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07233__A1 vss _03190_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1056 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_79 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06036__A2 vss _01544_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_999 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08951_ vdd _04290_ _04289_ _00854_ _04266_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08981__A1 vss _04301_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05795__A1 vss _01552_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08882_ vdd vss _04248_ net240 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07902_ vdd _03625_ _03624_ _00470_ _03619_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07536__A2 vss _03390_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07833_ vdd _03582_ _03581_ _00444_ _03554_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_5_25__f_clk vdd vss clknet_5_25__leaf_clk clknet_3_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07764_ vdd _03539_ _03538_ _00418_ _03521_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_1005 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07695_ vdd vss _03497_ _02917_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09503_ vdd _04636_ _04635_ _01060_ _04634_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_1173 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06715_ vdd vss _02864_ rf_ram.memory\[520\]\[1\] _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06646_ vdd vss _02814_ _02736_ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09434_ vss _01035_ _04592_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_228 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09365_ vdd vss _04554_ _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06577_ vdd vss _02759_ _02719_ _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_47_554 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05528_ _01724_ _01643_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_09296_ vdd vss _04513_ rf_ram.memory\[64\]\[1\] _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08316_ vdd vss _03883_ rf_ram.memory\[220\]\[1\] _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_513 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_640 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06763__I vss _02898_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_272 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_1101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_866 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05459_ _01655_ vss vdd _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_34_226 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08247_ vdd vss _03841_ rf_ram.memory\[528\]\[0\] _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06275__A2 vss _01846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08178_ vss _03798_ _02845_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_07129_ vdd vss _03144_ rf_ram.memory\[4\]\[1\] _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10140_ vdd vss _05053_ rf_ram.memory\[453\]\[1\] _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08972__A1 vss _03071_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06432__C1 vss _01772_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05786__A1 vss _01909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput170 o_ext_rs2[0] net170 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput192 o_ext_rs2[2] net192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_98_1218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10071_ vdd vss _05010_ rf_ram.memory\[508\]\[1\] _05008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput181 o_ext_rs2[1] net181 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08724__A1 vss _02971_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05538__A1 vss _01347_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_618 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10973_ vdd rf_ram.memory\[509\]\[1\] clknet_leaf_221_clk vss _00710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_337_clk vdd vss clknet_leaf_337_clk clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_183_868 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07463__A1 vss _03326_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11525_ vdd rf_ram.memory\[308\]\[0\] clknet_leaf_145_clk vss _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_259 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07215__A1 vss _03193_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09204__A2 vss _03035_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11456_ vdd rf_ram.memory\[18\]\[1\] clknet_leaf_283_clk vss _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06018__A2 vss _01511_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10407_ vdd rf_ram.memory\[390\]\[1\] clknet_leaf_121_clk vss _00151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11387_ _01119_ vdd vss clknet_leaf_224_clk net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10338_ vdd rf_ram.memory\[285\]\[0\] clknet_leaf_173_clk vss _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08963__A1 vss _04269_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07518__A2 vss _02894_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10269_ vdd rf_ram.memory\[241\]\[1\] clknet_leaf_282_clk vss _00013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_178_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06848__I vss _02959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_328_clk vdd vss clknet_leaf_328_clk clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07480_ vdd _03363_ _03362_ _00310_ _03356_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_487 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06500_ _02691_ net131 _01376_ vss _01400_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09140__A1 vss _04401_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1100 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_876 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09691__A2 vss net31 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05701__A1 vss _01603_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06431_ _01923_ vdd vss _02626_ rf_ram.memory\[96\]\[1\] _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09150_ vdd _04414_ _04412_ _00929_ _04401_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_727 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06362_ _01953_ rf_ram.memory\[227\]\[1\] vdd vss _02557_ rf_ram.memory\[226\]\[1\]
+ _01958_ _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07454__A1 vss _02775_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09081_ vdd _04371_ _04369_ _00903_ _04367_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06293_ rf_ram.memory\[138\]\[1\] _02488_ vss vdd rf_ram.memory\[137\]\[1\] _01610_
+ rf_ram.memory\[139\]\[1\] _01608_ _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_05313_ vdd vss _01509_ _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_08101_ vdd vss _03750_ rf_ram.memory\[556\]\[1\] _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08032_ vdd _03707_ _03706_ _00518_ _03686_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05244_ vdd _01342_ _01439_ _01444_ cpu.alu.i_rs1 vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_787 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_905 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput61 vss net61 i_ibus_rdt[6] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput50 vss net50 i_ibus_rdt[25] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05175_ vdd vss net130 _01375_ _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07757__A2 vss _03496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08954__A1 vss _02991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09983_ vdd _04956_ _04955_ _01221_ _04950_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08934_ vdd vss _04280_ _02953_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08706__A1 vss _04126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08865_ vdd vss _04238_ rf_ram.memory\[409\]\[1\] _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_157_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11664__I vss net115 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07816_ vdd vss _03572_ _02959_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08796_ vdd _04194_ _04192_ _00795_ _04170_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07747_ vdd vss _03529_ _02983_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input14_I vss i_dbus_rdt[20] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09131__A1 vss net244 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_319_clk vdd vss clknet_leaf_319_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07678_ vdd vss _03486_ rf_ram.memory\[402\]\[0\] _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07693__A1 vss _03491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06629_ vss _02801_ _02800_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_94_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09417_ _02707_ vdd vss _04584_ net87 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_852 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09348_ _04540_ net229 vdd vss _04545_ net228 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_65_1206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11310_ _01043_ vdd vss clknet_leaf_266_clk net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_7_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09279_ vss _00971_ _04501_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09198__A1 vss _04434_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11241_ vdd rf_ram.memory\[64\]\[1\] clknet_leaf_23_clk vss _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_max_cap251_I vss net252 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11172_ vdd rf_ram.memory\[97\]\[0\] clknet_leaf_70_clk vss _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06442__B vss _01563_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_640 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06405__C1 vss _01656_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output82_I vss net82 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05759__A1 vss _01951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10123_ vdd vss _05042_ rf_ram.memory\[438\]\[1\] _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06420__A2 vss _01770_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_0__f_clk_I vss clknet_3_0_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10054_ vdd vss _05000_ rf_ram.memory\[34\]\[0\] _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06184__A1 vss _01769_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08173__A2 vss _02917_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07920__A2 vss _03547_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05572__I vss _01660_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05392__C1 vss _01554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10956_ vdd rf_ram.memory\[188\]\[1\] clknet_leaf_6_clk vss _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06487__A2 vss _01661_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10887_ vdd rf_ram.memory\[21\]\[1\] clknet_leaf_207_clk vss _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07436__A1 vss _03323_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06239__A2 vss _01706_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11508_ vdd rf_ram.memory\[327\]\[1\] clknet_leaf_169_clk vss _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_551 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_538 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_549 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09189__A1 vss net242 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1030 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11439_ vdd cpu.mem_bytecnt\[0\] clknet_leaf_241_clk vss _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08936__A1 vss _04266_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_925 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06980_ vdd vss _03048_ rf_ram.memory\[426\]\[0\] _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input6_I vss i_dbus_rdt[13] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05931_ _02125_ _02126_ vdd vss _02127_ _02123_ _02124_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08650_ vdd vss _04104_ rf_ram.memory\[161\]\[1\] _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05862_ vdd vss _02058_ rf_ram.memory\[228\]\[0\] _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07601_ vdd vss _03438_ rf_ram.memory\[354\]\[1\] _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05482__I vss _01617_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05383__C1 vss _01517_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08581_ vdd vss _04060_ rf_ram.memory\[168\]\[0\] _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05793_ _01989_ vss vdd _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07532_ vdd vss _03396_ rf_ram.memory\[321\]\[0\] _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_113_1008 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_295 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_187_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07463_ vdd _03351_ _03349_ _00305_ _03326_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06414_ _01856_ _01857_ rf_ram.memory\[115\]\[1\] _02608_ vdd vss _02609_ rf_ram.memory\[114\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_09202_ vdd vss _04447_ rf_ram.memory\[70\]\[1\] _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07394_ vdd _03308_ _03306_ _00279_ _03292_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_710 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09133_ vdd _04404_ _04403_ _00922_ _04397_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06345_ _01860_ vdd vss _02540_ _02538_ _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08742__B vss _01506_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09064_ vdd _04360_ _04358_ _00897_ _04334_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05989__A1 vss net252 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_4_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06276_ vdd vss _02471_ rf_ram.memory\[145\]\[1\] _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_142_573 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_938 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05227_ vdd vss _01426_ _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08015_ vdd vss _03697_ _02839_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_1148 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05158_ _01354_ _01355_ _01360_ vdd vss _01361_ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_09966_ vdd _04945_ _04944_ _01215_ _04918_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06402__A2 vss _01785_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08968__I vss _04061_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08917_ vdd vss _04270_ rf_ram.memory\[439\]\[1\] _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09897_ vdd vss _04903_ rf_ram.memory\[263\]\[0\] _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_96_clk vdd vss clknet_leaf_96_clk clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08848_ vdd vss _04227_ rf_ram.memory\[133\]\[1\] _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_1021 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_58_1065 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output120_I vss net120 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09104__A1 vss _04364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08779_ vdd _04184_ _04183_ _00788_ _04167_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09655__A2 vss net2 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10810_ vdd rf_ram.memory\[551\]\[0\] clknet_leaf_324_clk vss _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07666__A1 vss _02866_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10741_ vdd rf_ram.memory\[457\]\[1\] clknet_leaf_51_clk vss _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06469__A2 vss _01605_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05677__B1 vss _01810_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_991 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07418__A1 vss _02866_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10672_ vdd rf_ram.memory\[376\]\[0\] clknet_leaf_114_clk vss _00416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_1026 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_20_clk vdd vss clknet_leaf_20_clk clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_180_679 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_253 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_91_994 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_1036 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11224_ vdd rf_ram.memory\[329\]\[0\] clknet_leaf_152_clk vss _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08918__A1 vss _04269_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06172__B vss _01756_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05567__I vss _01653_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_960 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11155_ vdd rf_ram.memory\[103\]\[1\] clknet_leaf_66_clk vss _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10106_ vdd vss _05032_ rf_ram.memory\[312\]\[0\] _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11086_ vdd rf_ram.memory\[130\]\[1\] clknet_leaf_24_clk vss _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05516__B vss _01602_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10037_ vdd _04989_ _04987_ _01242_ _04985_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08146__A2 vss _03765_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05365__C1 vss _01539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_424 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05380__A2 vss _01502_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10939_ rf_ram_if.rtrig0 vdd vss clknet_leaf_278_clk rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05668__B1 vss _01848_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06066__C vss _01670_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_1147 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05683__A3 vss _01878_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_11_clk vdd vss clknet_leaf_11_clk clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_182_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06130_ rf_ram.memory\[299\]\[1\] _02324_ vdd vss _02325_ rf_ram.memory\[298\]\[1\]
+ _01777_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_121_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_516 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08082__A1 vss _03724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06061_ _01658_ vdd vss _02256_ _02254_ _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_121_88 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_100_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_869 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08909__A1 vss _04234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_571 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_999 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09820_ vdd vss _04856_ rf_ram.memory\[259\]\[1\] _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08385__A2 vss _03903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06963_ vdd vss _03037_ rf_ram.memory\[22\]\[0\] _03036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09751_ vdd vss _04812_ _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05426__B vss _01615_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05914_ _01916_ vdd vss _02110_ rf_ram.memory\[120\]\[0\] _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_78_clk vdd vss clknet_leaf_78_clk clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08702_ vdd vss _04136_ rf_ram.memory\[39\]\[1\] _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06148__A1 vss rf_ram.memory\[312\]\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06894_ vdd _02990_ _02988_ _00097_ _02975_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09682_ vdd vss _04764_ _04740_ _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07896__A1 vss _03619_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05845_ rf_ram.memory\[196\]\[0\] _02041_ vss vdd rf_ram.memory\[199\]\[0\] _01713_
+ rf_ram.memory\[197\]\[0\] _01721_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_55_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08633_ vdd vss _04093_ rf_ram.memory\[549\]\[1\] _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05776_ _01972_ _01615_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08564_ vdd vss _04049_ rf_ram.memory\[509\]\[0\] _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07515_ vdd _03384_ _03383_ _00324_ _03356_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07648__A1 vss _03455_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09637__A2 vss net61 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1060 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08495_ vdd _04002_ _04001_ _00686_ _03953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_941 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_1141 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_1003 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_405 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07446_ vdd _03341_ _03340_ _00298_ _03323_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_844 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07377_ vdd _03298_ _03297_ _00272_ _03289_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09116_ vdd _04392_ _04390_ _00917_ _04367_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06328_ _01551_ vdd vss _02523_ rf_ram.memory\[208\]\[1\] _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08073__A1 vss _02761_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07820__A1 vss _03557_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09047_ vdd _04350_ _04349_ _00890_ _04331_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06259_ rf_ram.memory\[420\]\[1\] _02454_ vss vdd rf_ram.memory\[423\]\[1\] _01646_
+ rf_ram.memory\[421\]\[1\] _01810_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_142_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_746 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_102_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09949_ vdd vss _04935_ net248 _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__10183__A2 vss _03902_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09325__A1 vss _04463_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_69_clk vdd vss clknet_leaf_69_clk clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09876__A2 vss _02954_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07887__A1 vss _03590_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1063 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05898__B1 vss _01646_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_552 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05362__A2 vss _01532_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_0_clk_I vss clknet_5_1__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10724_ vdd rf_ram.memory\[461\]\[0\] clknet_leaf_118_clk vss _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_827 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_490 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06311__A1 vss _02494_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10655_ vdd rf_ram.memory\[3\]\[1\] clknet_leaf_40_clk vss _00399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07777__I vss _03039_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08064__A1 vss _03721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10586_ vdd rf_ram.memory\[321\]\[0\] clknet_leaf_164_clk vss _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_140_307 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07811__A1 vss net236 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_508 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05297__I vss rf_ram.i_raddr\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_576 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1154 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11207_ vdd rf_ram.memory\[179\]\[1\] clknet_leaf_16_clk vss _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06378__A1 vss _01600_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09564__A1 vss _03992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11138_ vdd rf_ram.memory\[111\]\[0\] clknet_leaf_71_clk vss _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_78_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_6__f_clk vdd vss clknet_5_6__leaf_clk clknet_3_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09867__A2 vss _02921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11069_ vdd rf_ram.memory\[135\]\[0\] clknet_leaf_15_clk vss _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_0_clk vdd vss clknet_leaf_0_clk clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07878__A1 vss _02916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05630_ vdd vss _01826_ rf_ram.memory\[481\]\[0\] _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_148_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06550__A1 vss cpu.immdec.imm11_7\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05353__A2 vss _01523_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05760__I vss _01526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_1226 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05561_ _01756_ vdd vss _01757_ rf_ram.memory\[264\]\[0\] _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_129_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07300_ vdd vss _03250_ net239 _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_574 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_1124 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_974 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05492_ _01688_ vss vdd _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08280_ vdd _03861_ _03860_ _00612_ _03852_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_449 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07231_ vdd vss _03207_ _02829_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07162_ vdd vss _03165_ rf_ram.memory\[496\]\[1\] _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06113_ vss vdd rf_ram.memory\[271\]\[1\] _01646_ rf_ram.memory\[269\]\[1\] _01645_
+ _01644_ rf_ram.memory\[268\]\[1\] _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_81_290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07093_ vdd vss _03121_ rf_ram.memory\[502\]\[0\] _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_997 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06044_ _01615_ vdd vss _02239_ rf_ram.memory\[352\]\[1\] _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08358__A2 vss _03903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09803_ vdd vss _04846_ rf_ram.memory\[75\]\[0\] _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07995_ vdd vss _03683_ rf_ram.memory\[466\]\[0\] _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09307__A1 vss _04466_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05592__A2 vss _01787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09734_ _04791_ _04800_ vdd vss _04801_ net110 _04790_ net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06946_ vdd vss _03026_ _02728_ _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06877_ vdd _02979_ _02977_ _00091_ _02975_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_817 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09665_ _04749_ _04740_ vdd vss _04750_ net123 _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_173_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_1095 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05828_ _02019_ rf_ram.memory\[211\]\[0\] vdd vss _02024_ rf_ram.memory\[210\]\[0\]
+ _01804_ _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08616_ vdd vss _04083_ rf_ram.memory\[163\]\[0\] _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06541__A1 vss _02716_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09596_ _04705_ _04706_ vdd vss _01083_ _04703_ _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08547_ _04038_ vss vdd _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_05759_ _01954_ vdd vss _01955_ _01951_ _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_119_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_511 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08478_ _03991_ vss vdd _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_175_782 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07429_ vdd vss _03331_ _02923_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_169_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_123 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10440_ vdd rf_ram.memory\[485\]\[0\] clknet_leaf_224_clk vss _00184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06057__B1 vss _01645_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_131_830 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_165 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_688 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10371_ vdd rf_ram.memory\[232\]\[1\] clknet_leaf_276_clk vss _00115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_395 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05568__C1 vss _01668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05583__A2 vss _01697_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06780__A1 vss _02909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_338 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05740__C1 vss _01811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_861 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08285__A1 vss _03852_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10707_ vdd rf_ram.memory\[410\]\[1\] clknet_leaf_88_clk vss _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_793 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10092__A1 vss _05014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_763 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_955 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_134 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08037__A1 vss _03686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10638_ vdd rf_ram.memory\[403\]\[0\] clknet_leaf_97_clk vss _00382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_329 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10569_ vdd rf_ram.memory\[365\]\[1\] clknet_leaf_172_clk vss _00313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09785__A1 vss _02787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_688 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_452 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_1139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_850 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10147__A2 vss _02889_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05755__I vss _01693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06360__B vss _01956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07012__A2 vss _02917_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_283_clk_I vss clknet_5_18__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07780_ vdd _03549_ _03548_ _00424_ _03521_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06800_ vdd _02926_ _02924_ _00067_ _02876_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06771__A1 vss _02881_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 vss net4 i_dbus_rdt[11] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_06731_ _02876_ _02825_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09450_ _04593_ vdd vss _04601_ net75 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05704__B vss _01629_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06662_ vdd vss _02827_ rf_ram.memory\[347\]\[1\] _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05490__I vss _01499_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08401_ vdd vss _03937_ rf_ram.memory\[209\]\[0\] _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_298_clk_I vss clknet_5_7__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05326__A2 vss _01511_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05613_ _01650_ vdd vss _01809_ rf_ram.memory\[314\]\[0\] _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09381_ _04552_ net214 vdd vss _04563_ net212 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06593_ vdd vss _02772_ rf_ram.memory\[233\]\[1\] _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05544_ vdd vss _01740_ rf_ram.memory\[273\]\[0\] _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08332_ vdd vss _03894_ rf_ram.memory\[217\]\[0\] _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_1056 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_221_clk_I vss clknet_5_22__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06287__B1 vss _01636_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08263_ vdd _03850_ _03849_ _00606_ _03820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05475_ _01665_ _01667_ _01669_ _01670_ vdd vss _01671_ _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_07214_ vdd vss _03197_ rf_ram.memory\[261\]\[1\] _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08194_ vdd vss _03808_ _02812_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07145_ vdd _03153_ _03151_ _00185_ _03126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_236_clk_I vss clknet_5_22__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07251__A2 vss _02869_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07076_ vdd _03110_ _03108_ _00159_ _03092_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_100_502 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11667__I vss net118 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06027_ _02221_ vdd vss _02222_ _01495_ _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_input44_I vss i_ibus_rdt[19] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1001 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06211__B1 vss _01772_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07978_ vss _03672_ _02831_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_96_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09581__B vss _04678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06929_ vdd vss _03015_ _02752_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05565__A2 vss _01509_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09717_ _04768_ _04788_ vdd vss _04789_ net104 _04767_ net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__06762__A1 vss _02750_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09700__A1 vss _04740_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06496__I vss _01376_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09648_ vdd vss _04735_ net1 _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06514__A1 vss _01388_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_308 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09579_ _01469_ _04646_ _04690_ vdd vss _04692_ _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_148_760 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08267__A1 vss _03230_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11610_ vss net163 net90 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11541_ vdd rf_ram.memory\[373\]\[0\] clknet_leaf_110_clk vss _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09600__I vss net48 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11472_ vdd rf_ram.memory\[340\]\[1\] clknet_leaf_169_clk vss _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_547 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08019__A1 vss _03690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10423_ vdd rf_ram.memory\[502\]\[1\] clknet_leaf_185_clk vss _00167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10354_ vdd rf_ram.memory\[280\]\[0\] clknet_leaf_177_clk vss _00098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_496 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05253__A1 vss _01385_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10285_ vdd rf_ram.memory\[347\]\[1\] clknet_leaf_142_clk vss _00029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06180__B vss _01660_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08742__A2 vss _04158_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05556__A2 vss _01631_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_636 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_513 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05524__B vss _01707_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06505__A1 vss _01409_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08258__A1 vss _03820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10065__A1 vss _04982_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_782 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06269__B1 vss _01968_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06808__A2 vss _02894_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_421 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_465 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05260_ vdd vss _01459_ _01436_ _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05191_ _01391_ vss vdd _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_3_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_150_991 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_1213 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06441__B1 vss _01607_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_291_clk vdd vss clknet_leaf_291_clk clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08430__A1 vss _03953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05244__A1 vss cpu.alu.i_rs1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08950_ vdd vss _04290_ rf_ram.memory\[121\]\[0\] _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06992__A1 vss _03055_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07901_ vdd vss _03625_ rf_ram.memory\[444\]\[0\] _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08881_ vdd _04247_ _04245_ _00827_ _04237_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07832_ vdd vss _03582_ rf_ram.memory\[432\]\[0\] _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05547__A2 vss _01692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06744__A1 vss _02873_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07763_ vdd vss _03539_ rf_ram.memory\[394\]\[0\] _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09502_ vdd vss _04636_ rf_ram.memory\[289\]\[0\] _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_811 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08497__A1 vss _03956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05434__B vss _01629_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07694_ _03496_ vss vdd _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_116_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_124 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06714_ vdd _02863_ _02862_ _00044_ _02820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_1065 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09433_ _02707_ vdd vss _04592_ net67 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06645_ _02813_ vss vdd _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_160_clk_I vss clknet_5_27__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_365 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09364_ _04552_ net205 vdd vss _04554_ net204 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08315_ vdd _03882_ _03881_ _00626_ _03852_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06576_ vdd vss _02758_ _02756_ _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05527_ _01602_ vdd vss _01723_ rf_ram.memory\[330\]\[0\] _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_443 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09295_ vdd _04512_ _04511_ _00976_ _04463_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_40_clk_I vss clknet_5_7__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_763 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05458_ vdd vss _01654_ _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_7_674 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08246_ vdd vss _03840_ _03798_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_175_clk_I vss clknet_5_31__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_435 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08177_ vdd _03797_ _03795_ _00573_ _03790_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_132_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_55_clk_I vss clknet_5_9__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07128_ vdd _03143_ _03142_ _00178_ _03123_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05389_ rf_ram.memory\[562\]\[0\] _01585_ vss vdd rf_ram.memory\[561\]\[0\] _01555_
+ rf_ram.memory\[563\]\[0\] _01554_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_31_945 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1265 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06983__A1 vss _03018_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08972__A2 vss _04303_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06432__B1 vss _01857_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07059_ vdd _03099_ _03097_ _00153_ _03092_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_282_clk vdd vss clknet_leaf_282_clk clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xoutput160 o_ext_rs1[2] net160 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput182 o_ext_rs2[20] net182 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10070_ vdd _05009_ _05008_ _01255_ _04982_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput193 o_ext_rs2[30] net193 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput171 o_ext_rs2[10] net171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09921__A1 vss _04887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08724__A2 vss _03945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_113_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08488__A1 vss net248 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10972_ vdd rf_ram.memory\[509\]\[0\] clknet_leaf_221_clk vss _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_124 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07115__I vss _03134_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_128_clk_I vss clknet_5_13__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10047__A1 vss _04985_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06175__B vss _01504_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_694 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09988__A1 vss _04950_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_823 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_124_903 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06266__A3 vss _02460_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11524_ vdd rf_ram.memory\[508\]\[1\] clknet_leaf_198_clk vss _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_969 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11455_ vdd rf_ram.memory\[18\]\[0\] clknet_leaf_283_clk vss _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_777 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_31__f_clk vdd vss clknet_5_31__leaf_clk clknet_3_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10406_ vdd rf_ram.memory\[390\]\[0\] clknet_leaf_121_clk vss _00150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_468 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_271 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_298 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_671 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08412__A1 vss _03919_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11386_ _01118_ vdd vss clknet_leaf_224_clk net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05226__A1 vss _01388_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06974__A1 vss _02781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10337_ vdd rf_ram.memory\[303\]\[1\] clknet_leaf_135_clk vss _00081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_181 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05777__A2 vss _01531_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_273_clk vdd vss clknet_leaf_273_clk clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_178_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10268_ vdd rf_ram.memory\[241\]\[0\] clknet_leaf_282_clk vss _00012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09912__A1 vss _04911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1130 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10199_ vdd vss _05089_ _02908_ _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06726__A1 vss _02826_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_321 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06430_ rf_ram.memory\[100\]\[1\] _02625_ vss vdd rf_ram.memory\[103\]\[1\] _01696_
+ rf_ram.memory\[101\]\[1\] _01848_ _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_75_127 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10038__A1 vss net248 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06864__I vss _02819_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06361_ vdd vss _02556_ rf_ram.memory\[225\]\[1\] _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07454__A2 vss _02815_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06292_ _01923_ vdd vss _02487_ rf_ram.memory\[136\]\[1\] _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09080_ vdd vss _04371_ rf_ram.memory\[57\]\[1\] _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05312_ vdd vss _01508_ _01496_ _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_08100_ vdd _03749_ _03748_ _00544_ _03721_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08651__A1 vss _04097_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_295 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08031_ vdd vss _03707_ rf_ram.memory\[56\]\[0\] _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput40 vss net40 i_ibus_rdt[15] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05243_ vdd vss _01443_ cpu.alu.i_rs1 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput51 vss net51 i_ibus_rdt[26] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput62 vss net62 i_ibus_rdt[7] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05174_ vss _01376_ cpu.state.i_ctrl_misalign vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__08954__A2 vss _04038_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06414__B1 vss _01857_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09982_ vdd vss _04956_ rf_ram.memory\[275\]\[0\] _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_264_clk vdd vss clknet_leaf_264_clk clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08933_ vdd _04279_ _04277_ _00847_ _04269_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05768__A2 vss _01664_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09903__A1 vss _04884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_696 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06178__C1 vss _01668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08864_ _04237_ vss vdd _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_58_1214 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06717__A1 vss _02779_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07815_ vdd _03571_ _03569_ _00437_ _03557_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07390__A1 vss _02752_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06193__A2 vss _01543_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05925__C1 vss _01679_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08795_ vdd vss _04194_ rf_ram.memory\[139\]\[1\] _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07746_ vdd _03528_ _03526_ _00411_ _03524_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09131__A2 vss _04005_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07677_ vdd vss _03485_ _02923_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09416_ vdd _04583_ _04581_ _01026_ _04466_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_181_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177_674 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10029__A1 vss _04982_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06628_ vdd vss _02800_ _02797_ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_165_858 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06559_ vdd _02744_ _02743_ _00008_ _02739_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09347_ vdd vss _04544_ _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08642__A1 vss _02828_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09278_ _04497_ vdd vss _04501_ cpu.genblk3.csr.mcause3_0\[1\] _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_1144 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08229_ vdd vss _03830_ rf_ram.memory\[532\]\[1\] _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_574 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11240_ vdd rf_ram.memory\[64\]\[0\] clknet_leaf_23_clk vss _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09442__I0 vss net71 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06405__B1 vss _01654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10201__A1 vss _05078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05339__B vss _01506_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_255_clk vdd vss clknet_leaf_255_clk clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11171_ vdd rf_ram.memory\[569\]\[1\] clknet_leaf_304_clk vss _00907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10122_ vdd _05041_ _05040_ _01275_ _05014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output75_I vss net75 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06956__A1 vss _02766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10053_ vdd vss _04999_ _02868_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1061 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05392__B1 vss _01555_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_775 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07133__A1 vss _03123_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10955_ vdd rf_ram.memory\[188\]\[0\] clknet_leaf_6_clk vss _00693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10886_ vdd rf_ram.memory\[21\]\[0\] clknet_leaf_208_clk vss _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06341__C1 vss _01925_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08881__A1 vss _04237_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06684__I vss _02843_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_992 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_661 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_374 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_508 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11507_ vdd rf_ram.memory\[327\]\[0\] clknet_5_30__leaf_clk vss _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_344 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_295 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09189__A2 vss _04418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09433__I0 vss net67 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11438_ _01170_ vdd vss clknet_leaf_241_clk cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11369_ _01101_ vdd vss clknet_leaf_218_clk cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06352__C vss _01362_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_246_clk vdd vss clknet_leaf_246_clk clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09436__S vss _04593_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05930_ rf_ram.memory\[98\]\[0\] _02126_ vss vdd rf_ram.memory\[97\]\[0\] _01772_
+ rf_ram.memory\[99\]\[0\] _01857_ _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_119_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_88 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05763__I vss _01695_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05861_ _01494_ vdd vss _02057_ _02054_ _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07600_ vdd _03437_ _03436_ _00356_ _03422_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07372__A1 vss _03289_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06175__A2 vss _01662_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08580_ vdd vss _04059_ net250 _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07531_ vdd vss _03395_ _03319_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05922__A2 vss _01641_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05383__B1 vss _01521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05792_ vdd vss _01988_ rf_ram.memory\[164\]\[0\] _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10259__A1 vss _02916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_652 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_797 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_85 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07462_ vdd vss _03351_ rf_ram.memory\[367\]\[1\] _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05712__B vss _01907_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08872__A1 vss _02787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_858 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05686__A1 vss _01769_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06413_ vdd vss _02608_ rf_ram.memory\[113\]\[1\] _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07393_ vdd vss _03308_ rf_ram.memory\[265\]\[1\] _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09201_ vdd _04446_ _04445_ _00948_ _04431_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_1218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_661 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_823 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_379 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09132_ vdd vss _04404_ rf_ram.memory\[91\]\[0\] _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06344_ rf_ram.memory\[202\]\[1\] _02539_ vss vdd rf_ram.memory\[201\]\[1\] _01645_
+ rf_ram.memory\[203\]\[1\] _01636_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_72_675 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08624__A1 vss _04062_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_541 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09063_ vdd vss _04360_ rf_ram.memory\[100\]\[1\] _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06275_ _01956_ vdd vss _02470_ rf_ram.memory\[144\]\[1\] _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_124_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05226_ vdd vss _01426_ _01388_ _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08014_ vdd _03696_ _03694_ _00511_ _03690_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06262__C vss _01717_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_764 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09854__B vss cpu.mem_bytecnt\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05157_ vdd vss _01360_ _01357_ _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06938__A1 vss _03014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09965_ vdd vss _04945_ rf_ram.memory\[295\]\[0\] _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09896_ vdd vss _04902_ _02828_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08916_ _04269_ _04061_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08847_ vdd _04226_ _04225_ _00814_ _04202_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09352__A2 vss _03991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06166__A2 vss _01623_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08778_ vdd vss _04184_ rf_ram.memory\[142\]\[0\] _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_135_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07729_ vdd _03517_ _03515_ _00405_ _03491_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_184_419 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08863__A1 vss _04234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07666__A2 vss _03089_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10740_ vdd rf_ram.memory\[457\]\[0\] clknet_leaf_51_clk vss _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_959 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10671_ vdd rf_ram.memory\[395\]\[1\] clknet_leaf_116_clk vss _00415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_299 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07418__A2 vss _03101_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08615__A1 vss _02888_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_105_221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11223_ vdd rf_ram.memory\[339\]\[1\] clknet_leaf_176_clk vss _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_228_clk vdd vss clknet_leaf_228_clk clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06929__A1 vss _02752_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09040__A1 vss net250 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_27__f_clk_I vss clknet_3_6_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11154_ vdd rf_ram.memory\[103\]\[0\] clknet_leaf_66_clk vss _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10105_ vdd vss _05031_ _02800_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_11085_ vdd rf_ram.memory\[130\]\[0\] clknet_leaf_27_clk vss _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10036_ vdd vss _04989_ rf_ram.memory\[326\]\[1\] _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06157__A2 vss _01683_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05365__B1 vss _01540_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07106__A1 vss _03123_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08854__A1 vss _04205_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10938_ vdd rf_ram.i_raddr\[0\] clknet_leaf_259_clk vss _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_931 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_1080 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_116_519 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10869_ vdd rf_ram.memory\[194\]\[1\] clknet_leaf_36_clk vss _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_823 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_834 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_327 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_483 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06363__B vss _01494_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06060_ rf_ram.memory\[379\]\[1\] _01763_ _01500_ rf_ram.memory\[378\]\[1\] _02255_
+ vss vdd rf_ram.memory\[377\]\[1\] _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__05840__A1 vss _01972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_219_clk vdd vss clknet_leaf_219_clk clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_583 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07593__A1 vss _02935_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06396__A2 vss _01770_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09582__A2 vss _04678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06962_ vdd vss _03036_ _03035_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09750_ _04791_ _04811_ vdd vss _04812_ net115 _04790_ net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_20_1121 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05913_ _01790_ vdd vss _02109_ _02106_ _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08701_ vdd _04135_ _04134_ _00759_ _04126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09681_ vdd vss cpu.bufreg2.o_sh_done_r _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06148__A2 vss _01666_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06893_ vdd vss _02990_ rf_ram.memory\[300\]\[1\] _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07345__A1 vss _03257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08632_ vdd _04092_ _04091_ _00733_ _04058_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05844_ _01805_ vdd vss _02040_ rf_ram.memory\[198\]\[0\] _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08563_ vdd vss _04048_ _02915_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05775_ _01966_ _01970_ vdd vss _01971_ _01955_ _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07514_ vdd vss _03384_ rf_ram.memory\[362\]\[0\] _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08494_ vdd vss _04002_ rf_ram.memory\[359\]\[0\] _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08845__A1 vss _02794_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06257__C vss _01658_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07445_ vdd vss _03341_ rf_ram.memory\[331\]\[0\] _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_975 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_828 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_368 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06320__A2 vss _01856_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_566 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_174_485 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_305 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_73_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07376_ vdd vss _03298_ rf_ram.memory\[250\]\[0\] _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09115_ vdd vss _04392_ rf_ram.memory\[93\]\[1\] _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06327_ _02521_ vdd vss _02522_ _01951_ _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08073__A2 vss _03729_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06258_ _01805_ vdd vss _02453_ rf_ram.memory\[422\]\[1\] _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09046_ vdd vss _04350_ rf_ram.memory\[103\]\[0\] _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05209_ cpu.state.cnt_r\[3\] cpu.state.cnt_r\[2\] vdd vss _01409_ cpu.state.cnt_r\[1\]
+ cpu.state.cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_4
X_06189_ _01783_ vdd vss _02384_ rf_ram.memory\[472\]\[1\] _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_1043 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_780 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_391 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09948_ vdd _04934_ _04932_ _01208_ _04921_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09879_ vdd vss _04892_ rf_ram.memory\[239\]\[1\] _04890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09089__A1 vss _04364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_520 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05352__B vss _01505_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10723_ vdd rf_ram.memory\[445\]\[1\] clknet_leaf_78_clk vss _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_316 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10654_ vdd rf_ram.memory\[3\]\[0\] clknet_leaf_40_clk vss _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10585_ vdd rf_ram.memory\[361\]\[1\] clknet_leaf_160_clk vss _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09261__A1 vss cpu.mem_bytecnt\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_500 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_280 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_336 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07811__A2 vss _03234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_544 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09013__A1 vss rf_ram.memory\[10\]\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11206_ vdd rf_ram.memory\[179\]\[0\] clknet_leaf_17_clk vss _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09564__A2 vss net51 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07575__A1 vss _03393_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05527__B vss _01602_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11137_ vdd rf_ram.memory\[112\]\[1\] clknet_leaf_75_clk vss _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07327__A1 vss _03260_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11068_ vdd rf_ram.memory\[136\]\[1\] clknet_leaf_13_clk vss _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07878__A2 vss _03234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10019_ vdd vss _04978_ rf_ram.memory\[505\]\[1\] _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_153_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05560_ _01756_ _01601_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06550__A2 vss _02730_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_211 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_780 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1148 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08827__A1 vss _04202_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05491_ _01687_ _01686_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_74_759 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06302__A2 vss _01958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07230_ vdd _03206_ _03204_ _00217_ _03193_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_183_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_171_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_444 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07161_ vdd _03164_ _03163_ _00190_ _03157_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06112_ vdd vss _02307_ rf_ram.memory\[270\]\[1\] _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05488__I vss _01550_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07092_ vdd vss _03120_ _02915_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_6 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_731 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06043_ _02237_ vdd vss _02238_ _01603_ _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09004__A1 vss _04298_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_555 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_391 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09555__A2 vss _02709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07566__A1 vss _02795_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09802_ vdd vss _04845_ net246 _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06369__A2 vss _01634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07994_ vdd vss _03682_ _03672_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07208__I vss _03017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07318__A1 vss _02958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09733_ vdd vss _04800_ _04781_ net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06945_ vdd _03025_ _03023_ _00113_ _03018_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06876_ vdd vss _02979_ rf_ram.memory\[282\]\[1\] _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09664_ vdd vss _04749_ _04737_ _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_555 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1074 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05827_ vdd vss _02023_ rf_ram.memory\[209\]\[0\] _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_55_1036 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08615_ vdd vss _04082_ _02888_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09595_ vdd vss _04706_ cpu.immdec.imm24_20\[1\] _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08546_ vdd vss _04037_ _02764_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05758_ rf_ram.memory\[157\]\[0\] _01516_ _01614_ rf_ram.memory\[156\]\[0\] _01954_
+ vss vdd rf_ram.memory\[159\]\[0\] _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_05689_ _01778_ rf_ram.memory\[395\]\[0\] vdd vss _01885_ rf_ram.memory\[394\]\[0\]
+ _01777_ _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_147_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09491__A1 vss cpu.alu.i_rs1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08477_ _03989_ net65 vdd vss _03990_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_0_49_299 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07428_ vdd _03330_ _03328_ _00291_ _03326_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_625 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05900__B vss _01707_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07359_ vdd vss _03287_ rf_ram.memory\[268\]\[0\] _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_781 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_617 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_155 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10370_ vdd rf_ram.memory\[232\]\[0\] clknet_leaf_276_clk vss _00114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09029_ _04339_ vss vdd _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_20_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05568__B1 vss _01763_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_133 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06780__A2 vss _02911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_328 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_542 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_1289 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06532__A2 vss _01525_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05740__B1 vss _01725_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_920 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08809__A1 vss net247 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_586 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_225 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10706_ vdd rf_ram.memory\[410\]\[0\] clknet_leaf_88_clk vss _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07788__I vss _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06296__A1 vss _01674_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_455 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10637_ vdd rf_ram.memory\[385\]\[1\] clknet_leaf_91_clk vss _00381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10568_ vdd rf_ram.memory\[365\]\[0\] clknet_leaf_172_clk vss _00312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07796__A1 vss _02908_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09785__A2 vss _04507_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10499_ vdd rf_ram.memory\[25\]\[1\] clknet_leaf_200_clk vss _00243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07548__A1 vss _03389_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09444__S vss _04593_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 vss net5 i_dbus_rdt[12] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_127_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06730_ vdd _02875_ _02874_ _00048_ _02873_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06771__A2 vss _02904_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06661_ _02826_ vss vdd _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07720__A1 vss _02971_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05612_ _01808_ vss vdd _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08400_ vdd vss _03936_ _03892_ _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05731__B1 vss _01925_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09380_ vdd vss _04562_ _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06592_ vdd _02771_ _02770_ _00014_ _02743_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_188_1013 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05543_ _01615_ vdd vss _01739_ rf_ram.memory\[272\]\[0\] _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08331_ vdd vss _03893_ _03892_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_145_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_636 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05474_ _01670_ rf_ram.i_raddr\[3\] vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08262_ vdd vss _03850_ rf_ram.memory\[205\]\[0\] _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07213_ vdd _03196_ _03195_ _00210_ _03190_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08193_ vdd _03807_ _03805_ _00579_ _03790_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06039__A1 vss _01351_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07787__A1 vss _03524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_691 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07144_ vdd vss _03153_ rf_ram.memory\[485\]\[1\] _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07075_ vdd vss _03110_ rf_ram.memory\[493\]\[1\] _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05798__B1 vss _01520_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06026_ _02219_ _02220_ vdd vss _02221_ _02217_ _02218_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__08200__A2 vss _03811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07977_ vdd _03671_ _03669_ _00499_ _03654_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input37_I vss i_ibus_rdt[12] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06928_ _03014_ vss vdd _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09716_ vdd vss _04788_ _04781_ net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06777__I vss _02908_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09700__A2 vss net3 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06859_ vdd vss _02967_ _02822_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09647_ vdd vss _04734_ _01401_ _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_132_1034 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09578_ _04690_ vdd vss _04691_ cpu.immdec.imm31 _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_139_249 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_901 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08267__A2 vss _02795_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08529_ vdd vss _04027_ rf_ram.memory\[49\]\[1\] _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11540_ vdd rf_ram.memory\[392\]\[1\] clknet_leaf_53_clk vss _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1205 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11471_ vdd rf_ram.memory\[340\]\[0\] clknet_leaf_169_clk vss _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09216__A1 vss _04431_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1238 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_680 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10422_ vdd rf_ram.memory\[502\]\[0\] clknet_leaf_185_clk vss _00166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07778__A1 vss _03547_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10353_ vdd rf_ram.memory\[300\]\[1\] clknet_leaf_137_clk vss _00097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_1103 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09519__A2 vss cpu.decode.opcode\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10284_ vdd rf_ram.memory\[347\]\[0\] clknet_leaf_142_clk vss _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05591__I vss _01514_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07702__A1 vss _03488_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1075 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07311__I vss _03013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_578 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_548 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11669_ vss net193 net121 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_792 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_937 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05190_ vdd vss cpu.branch_op _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07769__A1 vss _03521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_935 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_272 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06992__A2 vss _02894_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07900_ vdd vss _03624_ _02839_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08880_ vdd vss _04247_ rf_ram.memory\[128\]\[1\] _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_20_692 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07831_ vdd vss _03581_ _02945_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08194__A1 vss _02812_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06597__I vss net247 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07762_ vdd vss _03538_ _02775_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09501_ vdd vss _04635_ _03445_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07693_ vdd _03495_ _03493_ _00391_ _03491_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_91_1022 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09694__A1 vss _04740_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06713_ vdd vss _02863_ rf_ram.memory\[520\]\[0\] _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09432_ vss _01034_ _04591_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06644_ vdd vss _02812_ _02773_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_177_889 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06575_ vdd vss _02757_ _01562_ _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09363_ vdd vss _04553_ _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_523 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_517 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05526_ rf_ram.memory\[333\]\[0\] _01721_ _01709_ rf_ram.memory\[332\]\[0\] _01722_
+ vss vdd rf_ram.memory\[335\]\[0\] _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08314_ vdd vss _03882_ rf_ram.memory\[220\]\[0\] _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09294_ vdd vss _04512_ rf_ram.memory\[64\]\[0\] _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_455 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05457_ _01653_ vss vdd _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08245_ vdd _03839_ _03837_ _00599_ _03823_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09857__B vss _02690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06680__A1 vss _02820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05388_ _01552_ vdd vss _01584_ rf_ram.memory\[560\]\[0\] _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08176_ vdd vss _03797_ rf_ram.memory\[542\]\[1\] _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_149 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07127_ vdd vss _03143_ rf_ram.memory\[4\]\[0\] _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_480 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07058_ vdd vss _03099_ rf_ram.memory\[38\]\[1\] _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput161 o_ext_rs1[30] net161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput150 o_ext_rs1[20] net150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput194 o_ext_rs2[31] net194 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput183 o_ext_rs2[21] net183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput172 o_ext_rs2[11] net172 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06009_ _02202_ _02203_ vdd vss _02204_ _02200_ _02201_ _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09592__B vss _01491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_399 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07932__A1 vss _03619_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05943__B1 vss _01624_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05625__B vss _01684_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08488__A2 vss _03496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10971_ vdd rf_ram.memory\[499\]\[1\] clknet_leaf_185_clk vss _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06499__A1 vss _01375_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05171__A1 vss _01368_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06456__B vss _01562_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_331 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_731 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11408__CLK vss clknet_5_28__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11523_ vdd rf_ram.memory\[508\]\[0\] clknet_leaf_211_clk vss _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1035 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_282_clk_I vss clknet_5_19__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_594 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_222 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06671__A1 vss _02820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1079 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11454_ vdd rf_ram.memory\[219\]\[1\] clknet_leaf_298_clk vss _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10405_ vdd rf_ram.memory\[391\]\[1\] clknet_leaf_118_clk vss _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_378 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_570 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05586__I vss _01682_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11385_ _01117_ vdd vss clknet_leaf_219_clk net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10336_ vdd rf_ram.memory\[303\]\[0\] clknet_leaf_135_clk vss _00080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_297_clk_I vss clknet_5_7__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_467 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06974__A2 vss _03040_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10267_ vdd rf_ram.memory\[201\]\[1\] clknet_leaf_37_clk vss _00011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09912__A2 vss _02992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_220_clk_I vss clknet_5_22__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06187__B1 vss _01778_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10198_ vdd _05088_ _05086_ _01304_ _05081_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_79_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_834 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_235_clk_I vss clknet_5_22__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05162__A1 vss cpu.genblk3.csr.o_new_irq vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10038__A2 vss _02801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09979__A2 vss _04951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07041__I vss _03013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08100__A1 vss _03721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06360_ _01956_ vdd vss _02555_ rf_ram.memory\[224\]\[1\] _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06291_ _02485_ vdd vss _02486_ _01909_ _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_05311_ _01506_ vdd vss _01507_ rf_ram.memory\[526\]\[0\] _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput30 vss net30 i_dbus_rdt[6] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_126_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_414 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_86_1146 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08030_ vdd vss _03706_ _03668_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05242_ _01442_ vss vdd cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_114_469 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput41 vss net41 i_ibus_rdt[16] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput52 vss net52 i_ibus_rdt[27] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput63 vss net63 i_ibus_rdt[8] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05496__I vss _01682_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05173_ vss _01375_ net138 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09981_ vdd vss _04955_ _02865_ _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05217__A2 vss cpu.mem_bytecnt\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08932_ vdd vss _04279_ rf_ram.memory\[123\]\[1\] _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_95 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08167__A1 vss _03790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08863_ vdd _04236_ _04235_ _00820_ _04234_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07914__A1 vss _03622_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06178__B1 vss _01763_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07814_ vdd vss _03571_ rf_ram.memory\[434\]\[1\] _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05925__B1 vss _01793_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08794_ vdd _04193_ _04192_ _00794_ _04167_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07745_ vdd vss _03528_ rf_ram.memory\[396\]\[1\] _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07390__A2 vss _03253_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07676_ vdd _03484_ _03482_ _00385_ _03458_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09415_ vdd vss _04583_ rf_ram.memory\[299\]\[1\] _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06627_ _02730_ vdd vss _02799_ _02798_ cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_0_137_539 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06558_ vdd vss _02744_ rf_ram.memory\[200\]\[0\] _02739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_662 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09346_ _04540_ net228 vdd vss _04544_ net227 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_940 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_364 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_369 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05509_ _01700_ _01704_ vdd vss _01705_ _01681_ _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__06102__B1 vss _01625_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_753 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06489_ _02683_ vdd vss _02684_ _01348_ _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09277_ _04499_ vdd vss _04500_ _01365_ _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08642__A2 vss _02881_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08228_ vdd _03829_ _03828_ _00592_ _03820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_71_890 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09442__I1 vss net72 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08159_ vdd vss _03786_ rf_ram.memory\[545\]\[1\] _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11170_ vdd rf_ram.memory\[569\]\[0\] clknet_leaf_305_clk vss _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1133 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10121_ vdd vss _05041_ rf_ram.memory\[438\]\[0\] _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_1253 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1096 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_max_cap237_I vss _02903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06956__A2 vss _02806_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10052_ vdd _04998_ _04996_ _01248_ _04985_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08158__A1 vss _03754_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07905__A1 vss _02787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05916__B1 vss _01911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1050 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10954_ vdd rf_ram.memory\[172\]\[1\] clknet_leaf_3_clk vss _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_191_clk vdd vss clknet_leaf_191_clk clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06341__B1 vss _01912_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10885_ vdd rf_ram.memory\[242\]\[1\] clknet_leaf_215_clk vss _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05695__A2 vss _01846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06892__A1 vss _02970_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_865 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_537 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11506_ vdd rf_ram.memory\[246\]\[1\] clknet_leaf_212_clk vss _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06644__A1 vss _02773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_767 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_69 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05852__C1 vss _01959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11437_ vdd cpu.ctrl.i_jump clknet_leaf_239_clk vss _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_940 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_1039 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08397__A1 vss _03919_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_776 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11368_ vdd cpu.decode.opcode\[0\] clknet_5_20__leaf_clk vss _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10319_ vdd rf_ram.memory\[511\]\[1\] clknet_leaf_211_clk vss _00063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_798 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_1196 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11299_ _01032_ vdd vss clknet_leaf_251_clk net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_05860_ _01953_ rf_ram.memory\[227\]\[0\] vdd vss _02056_ rf_ram.memory\[226\]\[0\]
+ _01958_ _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA_clkbuf_leaf_174_clk_I vss clknet_5_31__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05791_ _01986_ _01362_ vdd vss _01987_ _01351_ _01971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09452__S vss _04593_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07530_ vdd _03394_ _03391_ _00329_ _03393_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10259__A2 vss _03692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_54_clk_I vss clknet_5_9__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08321__A1 vss _03884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07461_ vdd _03350_ _03349_ _00304_ _03323_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05712__C vss net254 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_182_clk vdd vss clknet_leaf_182_clk clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08872__A2 vss _03945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06412_ _01916_ vdd vss _02607_ rf_ram.memory\[112\]\[1\] _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07392_ vdd _03307_ _03306_ _00278_ _03289_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_189_clk_I vss clknet_5_29__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09200_ vdd vss _04446_ rf_ram.memory\[70\]\[0\] _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_29_342 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06883__A1 vss _02750_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_550 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_69_clk_I vss clknet_5_8__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09131_ vdd vss _04403_ net244 _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06343_ _01916_ vdd vss _02538_ rf_ram.memory\[200\]\[1\] _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_8_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09821__A1 vss _04840_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09062_ vdd _04359_ _04358_ _00896_ _04331_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06635__A1 vss _02773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_112_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_976 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06274_ _01564_ vdd vss _02469_ _02466_ _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_115_789 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_998 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05225_ vdd vss _01425_ _01398_ _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08013_ vdd vss _03696_ rf_ram.memory\[573\]\[1\] _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05156_ vdd vss _01359_ _01337_ _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07060__A1 vss _02764_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_127_clk_I vss clknet_5_13__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09964_ vdd vss _04944_ _03445_ _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05610__A2 vss _01804_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08915_ vdd _04268_ _04267_ _00840_ _04266_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_494 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09895_ vdd _04901_ _04899_ _01188_ _04887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09888__A1 vss _04884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08330__I vss _02737_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08846_ vdd vss _04226_ rf_ram.memory\[133\]\[0\] _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_406 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08560__A1 vss _04023_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06020__C1 vss _01517_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05374__A1 vss _01351_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05989_ _02184_ vdd vss _02185_ net252 _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_08777_ vdd vss _04183_ _02971_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07728_ vdd vss _03517_ rf_ram.memory\[37\]\[1\] _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08312__A1 vss _03855_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07659_ vdd vss _03474_ rf_ram.memory\[404\]\[1\] _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_173_clk vdd vss clknet_leaf_173_clk clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10670_ vdd rf_ram.memory\[395\]\[0\] clknet_leaf_116_clk vss _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05677__A2 vss _01666_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09329_ vdd vss _04534_ rf_ram.memory\[309\]\[0\] _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_369 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_470 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06087__C1 vss _01715_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09812__A1 vss _02828_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08615__A2 vss _04067_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_520 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_304 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_895 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11222_ vdd rf_ram.memory\[339\]\[0\] clknet_leaf_176_clk vss _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08379__A1 vss _03922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06929__A2 vss _02801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09040__A2 vss _04339_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11153_ vdd rf_ram.memory\[104\]\[1\] clknet_leaf_68_clk vss _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11084_ vdd rf_ram.memory\[409\]\[1\] clknet_leaf_88_clk vss _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10104_ vdd _05030_ _05028_ _01268_ _05017_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05601__A2 vss _01719_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10035_ vdd _04988_ _04987_ _01241_ _04982_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06011__C1 vss _01554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08303__A1 vss _03230_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_164_clk vdd vss clknet_leaf_164_clk clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05532__C vss _01658_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10110__A1 vss net250 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10937_ vdd rf_ram_if.wdata0_r\[1\] clknet_leaf_261_clk vss cpu.o_wdata0 vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05668__A2 vss _01863_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_267 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06865__A1 vss _02773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_604 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10868_ vdd rf_ram.memory\[194\]\[0\] clknet_leaf_36_clk vss _00612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_301 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_637 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10799_ vdd rf_ram.memory\[557\]\[1\] clknet_leaf_333_clk vss _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_334 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_879 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06617__A1 vss _02743_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07290__A1 vss _02836_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_575 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07042__A1 vss _02830_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10177__A1 vss _03892_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07593__A2 vss _02822_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06250__C1 vss _01857_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06961_ vss _03035_ _02996_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__09319__C2 vss cpu.immdec.imm11_7\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05912_ _01856_ _01857_ rf_ram.memory\[115\]\[0\] _02107_ vdd vss _02108_ rf_ram.memory\[114\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_08700_ vdd vss _04135_ rf_ram.memory\[39\]\[0\] _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09680_ vdd vss _04762_ _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06892_ vdd _02989_ _02988_ _00096_ _02970_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06002__C1 vss _01539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08631_ vdd vss _04092_ rf_ram.memory\[549\]\[0\] _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05843_ _01860_ vdd vss _02039_ _02037_ _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_178_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08562_ vdd _04047_ _04045_ _00708_ _04026_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05774_ _01969_ vdd vss _01970_ _01951_ _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_155_clk vdd vss clknet_leaf_155_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07513_ vdd vss _03383_ _02775_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08493_ vdd vss _04001_ _02829_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_426 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07444_ vdd vss _03340_ _02781_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06856__A1 vss _02927_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05659__A2 vss _01782_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_705 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08845__A2 vss _04195_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1095 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07375_ vdd vss _03297_ _03055_ _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_868 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09114_ vdd _04391_ _04390_ _00916_ _04364_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72_473 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06326_ vss vdd rf_ram.memory\[213\]\[1\] _01968_ rf_ram.memory\[215\]\[1\] _02019_
+ _01804_ rf_ram.memory\[214\]\[1\] _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__06608__A1 vss _02743_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06257_ _02449_ _02450_ _02451_ _01658_ vdd vss _02452_ _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__06084__A2 vss _01706_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09045_ vdd vss _04349_ _02828_ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05831__A2 vss _01515_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05208_ vdd vss _01408_ _01399_ _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06188_ _01790_ vdd vss _02383_ _02380_ _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07033__A1 vss _03053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09156__I vss _04004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05139_ _01342_ cpu.csr_d_sel vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05617__C vss _01658_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09947_ vdd vss _04934_ rf_ram.memory\[338\]\[1\] _04932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08781__A1 vss _04170_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08533__A1 vss _04023_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09878_ vdd _04891_ _04890_ _01181_ _04884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08829_ vdd _04215_ _04213_ _00807_ _04205_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05898__A2 vss _01801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_146_clk vdd vss clknet_leaf_146_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_166_921 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10722_ vdd rf_ram.memory\[445\]\[0\] clknet_leaf_78_clk vss _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06847__A1 vss _02750_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_442 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_656 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_738 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10653_ vdd rf_ram.memory\[381\]\[1\] clknet_leaf_107_clk vss _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10584_ vdd rf_ram.memory\[361\]\[0\] clknet_leaf_160_clk vss _00328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1182 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09261__A2 vss _01385_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_134 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_1161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06480__C1 vss _01653_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10159__A1 vss _05046_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05822__A2 vss _01523_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1280 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_1058 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05594__I vss _01493_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11205_ vdd rf_ram.memory\[84\]\[1\] clknet_leaf_49_clk vss _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07024__A1 vss _02738_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06232__C1 vss _01763_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11136_ vdd rf_ram.memory\[112\]\[0\] clknet_leaf_75_clk vss _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08772__A1 vss _02953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11067_ vdd rf_ram.memory\[136\]\[0\] clknet_leaf_12_clk vss _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_512 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10018_ vdd _04977_ _04976_ _01235_ _04950_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05543__B vss _01615_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_532 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06838__A1 vss _02930_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_137_clk vdd vss clknet_leaf_137_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_50_1104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05490_ _01686_ vss vdd _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_46_429 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_979 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07160_ vdd vss _03164_ rf_ram.memory\[496\]\[0\] _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_87_1060 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_771 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06093__C vss _01658_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06111_ _02302_ _02305_ vdd vss _02306_ _02294_ _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_07091_ vdd _03119_ _03117_ _00165_ _03092_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07263__A1 vss _02738_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_955 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06042_ rf_ram.memory\[359\]\[1\] _01608_ _01606_ rf_ram.memory\[358\]\[1\] _02237_
+ vss vdd rf_ram.memory\[357\]\[1\] _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_125_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_189 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07566__A2 vss _03390_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09801_ vdd _04844_ _04842_ _01150_ _04840_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_1239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_1010 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07993_ vdd _03681_ _03679_ _00505_ _03654_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09732_ vdd vss _04799_ _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07318__A2 vss _02946_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06944_ vdd vss _03025_ rf_ram.memory\[206\]\[1\] _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06875_ vdd _02978_ _02977_ _00090_ _02970_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09663_ vdd vss _04748_ net120 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08614_ vdd _04081_ _04079_ _00726_ _04062_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05826_ _01551_ vdd vss _02022_ rf_ram.memory\[208\]\[0\] _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_1184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09594_ vdd vss _04705_ _04526_ net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_132_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08545_ vdd _04036_ _04034_ _00702_ _04026_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_49_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06829__A1 vss _02935_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_128_clk vdd vss clknet_leaf_128_clk clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05757_ _01953_ vss vdd _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05688_ vdd vss _01884_ rf_ram.memory\[393\]\[0\] _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08476_ _03989_ _02695_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07427_ vdd vss _03330_ rf_ram.memory\[333\]\[1\] _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_1025 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07358_ vdd vss _03286_ _02788_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_760 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06057__A2 vss _01666_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_467 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_169 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06309_ rf_ram.memory\[173\]\[1\] _01516_ _01683_ rf_ram.memory\[172\]\[1\] _02504_
+ vss vdd rf_ram.memory\[175\]\[1\] _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_32_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_681 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07289_ vdd _03243_ _03241_ _00239_ _03225_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_501 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_300_clk vdd vss clknet_leaf_300_clk clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_130_331 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09028_ vdd _04338_ _04336_ _00883_ _04334_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output173_I vss net173 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05804__A2 vss _01501_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05628__B vss _01746_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07006__A1 vss _03053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08506__A1 vss cpu.immdec.imm11_7\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06459__B vss _01525_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1115 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_119_clk vdd vss clknet_leaf_119_clk clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08809__A2 vss _04195_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_896 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10705_ vdd rf_ram.memory\[431\]\[1\] clknet_leaf_99_clk vss _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07493__A1 vss _02788_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_475 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_1171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10636_ vdd rf_ram.memory\[385\]\[0\] clknet_leaf_92_clk vss _00380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05589__I vss _01686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07245__A1 vss _03193_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_787 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06048__A2 vss _01614_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_793 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1165 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10567_ vdd rf_ram.memory\[328\]\[1\] clknet_leaf_151_clk vss _00311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07796__A2 vss _03559_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10498_ vdd rf_ram.memory\[25\]\[0\] clknet_leaf_199_clk vss _00242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_5_14__f_clk vdd vss clknet_5_14__leaf_clk clknet_3_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06205__C1 vss _01810_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1120 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08745__A1 vss _01495_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_11__f_clk_I vss clknet_3_2_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11119_ vdd rf_ram.memory\[121\]\[1\] clknet_leaf_84_clk vss _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput6 vss net6 i_dbus_rdt[13] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_1059 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06660_ _02825_ vss vdd _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_188_342 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05611_ rf_ram.memory\[316\]\[0\] _01807_ vss vdd rf_ram.memory\[319\]\[0\] _01726_
+ rf_ram.memory\[317\]\[0\] _01725_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__06088__C vss _01717_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_176_537 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_217 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_863 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06591_ vdd vss _02771_ rf_ram.memory\[233\]\[0\] _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_143_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05542_ _01737_ vdd vss _01738_ _01675_ _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08330_ vss _03892_ _02737_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_05473_ rf_ram.memory\[370\]\[0\] _01669_ vss vdd rf_ram.memory\[369\]\[0\] _01668_
+ rf_ram.memory\[371\]\[0\] _01519_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__06287__A2 vss _01662_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08261_ vdd vss _03849_ _03230_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_941 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07212_ vdd vss _03196_ rf_ram.memory\[261\]\[0\] _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05499__I vss _01518_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1098 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07236__A1 vss _02806_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_765 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_782 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08192_ vdd vss _03807_ rf_ram.memory\[53\]\[1\] _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_473 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07143_ vdd _03152_ _03151_ _00184_ _03123_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08984__A1 vss _04298_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07074_ vdd _03109_ _03108_ _00158_ _03087_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_627 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06025_ rf_ram.memory\[546\]\[1\] _02220_ vss vdd rf_ram.memory\[545\]\[1\] _01517_
+ rf_ram.memory\[547\]\[1\] _01521_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_58_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08736__A1 vss _02713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06211__A2 vss _01711_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07976_ vdd vss _03671_ rf_ram.memory\[46\]\[1\] _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06927_ _03013_ _02742_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09715_ vdd vss _04787_ _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09161__A1 vss _04401_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09646_ _04732_ vdd vss _04733_ _01409_ _04731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06858_ vdd _02966_ _02964_ _00085_ _02930_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06789_ vdd vss _02919_ rf_ram.memory\[510\]\[0\] _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05809_ _02004_ vdd vss _02005_ rf_ram.memory\[190\]\[0\] _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09577_ cpu.decode.opcode\[1\] vdd vss _04690_ _01399_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_92_310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08528_ _04026_ vss vdd _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_93_866 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08459_ _03975_ vdd vss _03976_ net120 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_33_1154 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_248 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11470_ vdd rf_ram.memory\[341\]\[1\] clknet_leaf_170_clk vss _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_922 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05202__I vss cpu.state.stage_two_req vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10421_ vdd rf_ram.memory\[490\]\[1\] clknet_leaf_183_clk vss _00165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_832 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_448 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07778__A2 vss _03072_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10352_ vdd rf_ram.memory\[300\]\[0\] clknet_leaf_137_clk vss _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_320 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output98_I vss net98 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06461__C vss rf_ram.i_raddr\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10283_ vdd rf_ram.memory\[346\]\[1\] clknet_leaf_141_clk vss _00027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_695 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1272 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06968__I vss _03039_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06202__A2 vss _01804_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06189__B vss _01783_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05961__A1 vss _01599_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_537 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07466__A1 vss _03323_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_181 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_866 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06269__A2 vss _01614_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_581 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_905 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11668_ vss net191 net119 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10619_ vdd rf_ram.memory\[313\]\[1\] clknet_leaf_154_clk vss _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07218__A1 vss _03190_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_292 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11599_ vdd rf_ram.memory\[574\]\[0\] clknet_leaf_306_clk vss _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_796 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_465 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06441__A2 vss _01605_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08718__A1 vss _04129_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07830_ vdd _03580_ _03578_ _00443_ _03557_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08194__A2 vss _02846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07761_ vdd _03537_ _03535_ _00417_ _03524_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05782__I vss _01493_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1035 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09500_ _04634_ _04396_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09143__A1 vss _04397_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06712_ vdd vss _02862_ _02728_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07692_ vdd vss _03495_ rf_ram.memory\[401\]\[1\] _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_504 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_95_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_56_1132 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_172 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09431_ _02707_ vdd vss _04591_ net96 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06643_ vdd vss _02811_ _02719_ _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09362_ _04552_ net204 vdd vss _04553_ net203 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06574_ vdd vss _02756_ _02720_ _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_118_913 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05525_ vdd vss _01721_ _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_74_321 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08313_ vdd vss _03881_ _03230_ _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09293_ vdd vss _04511_ net237 _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_62_505 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_144_231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_618 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05456_ _01652_ _01499_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_62_549 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08244_ vdd vss _03839_ rf_ram.memory\[52\]\[1\] _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_933 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09857__C vss _01391_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_966 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05387_ rf_ram.memory\[564\]\[0\] _01583_ vss vdd rf_ram.memory\[567\]\[0\] _01554_
+ rf_ram.memory\[565\]\[0\] _01555_ _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_31_903 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08175_ vdd _03796_ _03795_ _00572_ _03787_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07126_ vdd vss _03142_ _02883_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06432__A2 vss _01785_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07057_ vdd _03098_ _03097_ _00152_ _03087_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xoutput151 o_ext_rs1[21] net151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput140 o_ext_rs1[11] net140 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08709__A1 vss net235 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput184 o_ext_rs2[22] net184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput173 o_ext_rs2[12] net173 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_11_682 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput162 o_ext_rs1[31] net162 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput195 o_ext_rs2[3] net195 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06008_ rf_ram.memory\[530\]\[1\] _02203_ vss vdd rf_ram.memory\[529\]\[1\] _01555_
+ rf_ram.memory\[531\]\[1\] _01554_ _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__06196__A1 vss _02379_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1102 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07959_ vdd _03660_ _03659_ _00492_ _03651_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output136_I vss net136 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10970_ vdd rf_ram.memory\[499\]\[0\] clknet_leaf_185_clk vss _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06499__A2 vss _02690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09629_ vdd vss _04723_ _04524_ net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_502 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07448__A1 vss _03326_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_693 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05171__A2 vss _01371_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_50_clk vdd vss clknet_leaf_50_clk clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11522_ vdd rf_ram.memory\[307\]\[1\] clknet_leaf_151_clk vss _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_163_551 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11453_ vdd rf_ram.memory\[219\]\[0\] clknet_leaf_298_clk vss _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08948__A1 vss _04269_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10404_ vdd rf_ram.memory\[391\]\[0\] clknet_leaf_118_clk vss _00148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09339__I vss _04539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_413 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_796 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11384_ _01116_ vdd vss clknet_leaf_218_clk net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10335_ vdd rf_ram.memory\[286\]\[1\] clknet_leaf_175_clk vss _00079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_470 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05631__B1 vss _01696_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10266_ vdd rf_ram.memory\[201\]\[0\] clknet_leaf_37_clk vss _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05816__B vss _01923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09074__I vss _04061_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10197_ vdd vss _05088_ rf_ram.memory\[210\]\[1\] _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05551__B vss _01746_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1041 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_682 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_185_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_158_378 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07439__A1 vss _02921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_326 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139_570 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_41_clk vdd vss clknet_leaf_41_clk clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_17_719 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1035 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_1103 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06290_ rf_ram.memory\[140\]\[1\] _02485_ vss vdd rf_ram.memory\[143\]\[1\] _01857_
+ rf_ram.memory\[141\]\[1\] _01931_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_56_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05310_ vss _01506_ _01505_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xinput20 vss net20 i_dbus_rdt[26] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput31 vss net31 i_dbus_rdt[7] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05241_ vdd vss _01441_ _01343_ _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_763 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1109 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08939__A1 vss net245 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput42 vss net42 i_ibus_rdt[17] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05172_ _01374_ vdd vss _00007_ _01351_ _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xinput53 vss net53 i_ibus_rdt[28] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_796 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput64 vss net64 i_ibus_rdt[9] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_969 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06414__A2 vss _01856_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09980_ vdd _04954_ _04951_ _01220_ _04953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05217__A3 vss _01385_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08931_ vdd _04278_ _04277_ _00846_ _04266_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_852 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08862_ vdd vss _04236_ rf_ram.memory\[409\]\[0\] _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_58_85 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07813_ vdd _03570_ _03569_ _00436_ _03554_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09116__A1 vss _04367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08793_ vdd vss _04193_ rf_ram.memory\[139\]\[0\] _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07744_ vdd _03527_ _03526_ _00410_ _03521_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07675_ vdd vss _03484_ rf_ram.memory\[384\]\[1\] _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05689__B1 vss _01778_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09414_ vdd _04582_ _04581_ _01025_ _04463_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_95_928 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06626_ vdd vss cpu.immdec.imm11_7\[3\] _02798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_48_811 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05153__A2 vss _01343_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_32_clk vdd vss clknet_leaf_32_clk clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09345_ vdd vss _04543_ _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06557_ _02743_ vss vdd _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_48_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05508_ _01703_ vdd vss _01704_ _01603_ _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06488_ _02681_ _02682_ vdd vss _02683_ _02679_ _02680_ rf_ram.i_raddr\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09276_ vdd vss _04499_ _01364_ cpu.genblk3.csr.mcause3_0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07850__A1 vss _03587_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_275 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05439_ _01635_ vss vdd _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_16_730 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08227_ vdd vss _03829_ rf_ram.memory\[532\]\[0\] _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06292__B vss _01923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_880 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08158_ vdd _03785_ _03784_ _00566_ _03754_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07602__A1 vss _03425_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06405__A2 vss _01652_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07109_ vdd vss _03131_ _02728_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08089_ vdd vss _03743_ rf_ram.memory\[558\]\[0\] _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10120_ vdd vss _05040_ _03008_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_99_clk vdd vss clknet_leaf_99_clk clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10051_ vdd vss _04998_ rf_ram.memory\[306\]\[1\] _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07905__A2 vss _02832_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09107__A1 vss _02916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05392__A2 vss _01538_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10953_ vdd rf_ram.memory\[172\]\[0\] clknet_leaf_4_clk vss _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_654 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_168_643 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06467__B vss _01601_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_287 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_490 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10884_ vdd rf_ram.memory\[242\]\[0\] clknet_leaf_215_clk vss _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_23_clk vdd vss clknet_leaf_23_clk clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_66_641 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_652 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_264 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11505_ vdd rf_ram.memory\[246\]\[0\] clknet_leaf_213_clk vss _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_195 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05597__I vss _01617_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05852__B1 vss _01968_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11436_ _01168_ cpu.state.cnt_r\[3\] vdd vss clknet_leaf_242_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_0_46_1131 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11367_ vdd cpu.csr_d_sel clknet_leaf_235_clk vss _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09594__A1 vss _04526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10318_ vdd rf_ram.memory\[511\]\[0\] clknet_leaf_211_clk vss _00062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11298_ _01031_ vdd vss clknet_leaf_251_clk net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09346__A1 vss net227 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05546__B vss _01620_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10249_ vdd vss _05119_ _02838_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05790_ _01982_ _01985_ vdd vss _01986_ _01975_ _01979_ _01349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__05383__A2 vss _01544_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_473 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_602 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07460_ vdd vss _03350_ rf_ram.memory\[367\]\[0\] _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_1119 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1091 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07391_ vdd vss _03307_ rf_ram.memory\[265\]\[0\] _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06411_ _02605_ vdd vss _02606_ _01909_ _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_151_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_540 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09130_ vdd _04402_ _04398_ _00921_ _04401_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_14_clk vdd vss clknet_leaf_14_clk clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06342_ _02536_ vdd vss _02537_ _01972_ _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08085__A1 vss _03721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_370 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09061_ vdd vss _04359_ rf_ram.memory\[100\]\[0\] _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_127_595 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06273_ _01959_ rf_ram.memory\[155\]\[1\] vdd vss _02468_ rf_ram.memory\[154\]\[1\]
+ _01958_ _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08012_ vdd _03695_ _03694_ _00510_ _03686_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_170_885 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05224_ vdd _01423_ _01383_ _01424_ _01412_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_941 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05155_ vdd vss _01358_ cpu.decode.op26 cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09963_ vdd _04943_ _04941_ _01214_ _04921_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07060__A2 vss _02799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08914_ vdd vss _04268_ rf_ram.memory\[439\]\[0\] _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09337__A1 vss _04466_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_484 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_462 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_682 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09894_ vdd vss _04901_ rf_ram.memory\[18\]\[1\] _04899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07899__A1 vss _03622_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08845_ vdd vss _04225_ _02794_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08776_ vdd _04182_ _04180_ _00787_ _04170_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_281_clk_I vss clknet_5_19__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06020__B1 vss _01521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input12_I vss i_dbus_rdt[19] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07727_ vdd _03516_ _03515_ _00404_ _03488_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05988_ _02183_ net254 vdd vss _02184_ _01349_ _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06571__A1 vss _02743_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_120 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07658_ vdd _03473_ _03472_ _00378_ _03455_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_94_224 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_296_clk_I vss clknet_5_7__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06323__A1 vss _01768_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07589_ vdd vss _03431_ rf_ram.memory\[355\]\[0\] _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05531__C1 vss _01726_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06609_ vdd vss _02784_ rf_ram.memory\[235\]\[1\] _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09328_ vdd vss _04533_ _03445_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07897__I vss _03359_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06087__B1 vss _01654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09812__A2 vss _03035_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_869 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1078 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07823__A1 vss _03554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_986 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09259_ vdd vss cpu.genblk3.csr.mie_mtie _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_181_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11221_ vdd rf_ram.memory\[349\]\[1\] clknet_leaf_176_clk vss _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_738 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11152_ vdd rf_ram.memory\[104\]\[0\] clknet_leaf_68_clk vss _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_1040 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output80_I vss net80 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09328__A1 vss _03445_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10103_ vdd vss _05030_ rf_ram.memory\[311\]\[1\] _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05598__C1 vss _01793_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11083_ vdd rf_ram.memory\[409\]\[0\] clknet_leaf_89_clk vss _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10034_ vdd vss _04988_ rf_ram.memory\[326\]\[0\] _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_249_clk_I vss clknet_5_21__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06011__B1 vss _01555_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_716 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05365__A2 vss _01544_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06197__B vss _01707_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_202 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05813__C vss _01860_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08303__A2 vss _02960_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10110__A2 vss _03088_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_747 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10936_ vdd rf_ram_if.wdata0_r\[0\] clknet_leaf_261_clk vss net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10867_ vdd rf_ram.memory\[195\]\[1\] clknet_leaf_46_clk vss _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_1139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06078__B1 vss _01696_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_441 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10798_ vdd rf_ram.memory\[557\]\[0\] clknet_leaf_333_clk vss _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07290__A2 vss _03135_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_749 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11419_ vdd rf_ram.memory\[75\]\[0\] clknet_leaf_24_clk vss _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10177__A2 vss _02775_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07042__A2 vss _02939_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09319__A1 vss _04526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06250__B1 vss _01931_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07047__I vss _03017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_3_clk vdd vss clknet_leaf_3_clk clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06960_ vdd _03034_ _03032_ _00119_ _03018_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09319__B2 vss cpu.immdec.imm11_7\[4\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05911_ vdd vss _02107_ rf_ram.memory\[113\]\[0\] _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06891_ vdd vss _02989_ rf_ram.memory\[300\]\[0\] _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input4_I vss i_dbus_rdt[11] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09463__S vss _04604_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05842_ rf_ram.memory\[202\]\[0\] _02038_ vss vdd rf_ram.memory\[201\]\[0\] _01645_
+ rf_ram.memory\[203\]\[0\] _01636_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__06002__B1 vss _01540_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08630_ vdd vss _04091_ _02794_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06553__A1 vss _02728_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08561_ vdd vss _04047_ rf_ram.memory\[499\]\[1\] _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_7_1006 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05773_ rf_ram.memory\[151\]\[0\] _01953_ _01958_ rf_ram.memory\[150\]\[0\] _01969_
+ vss vdd rf_ram.memory\[149\]\[0\] _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07512_ vdd _03382_ _03380_ _00323_ _03360_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08492_ vdd _04000_ _03998_ _00685_ _03956_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_596 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_410 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07443_ vdd _03339_ _03337_ _00297_ _03326_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_257 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_123 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08058__A1 vss _03721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_476 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07374_ vdd _03296_ _03294_ _00271_ _03292_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_128_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09113_ vdd vss _04391_ rf_ram.memory\[93\]\[0\] _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07805__A1 vss _03557_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06325_ vdd vss _02520_ rf_ram.memory\[212\]\[1\] _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06256_ rf_ram.memory\[424\]\[1\] _02451_ vss vdd rf_ram.memory\[427\]\[1\] _01811_
+ rf_ram.memory\[425\]\[1\] _01810_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09044_ vdd _04348_ _04346_ _00889_ _04334_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_60_647 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_587 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05292__A1 vss cpu.alu.i_rs1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05207_ _01405_ _01406_ vdd vss _01407_ _01390_ _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_06187_ _01778_ rf_ram.memory\[467\]\[1\] vdd vss _02382_ rf_ram.memory\[466\]\[1\]
+ _01777_ _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_25_1001 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_102_1213 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_1102 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05138_ _01340_ vdd vss _01341_ cpu.state.genblk1.misalign_trap_sync_r cpu.genblk3.csr.o_new_irq
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__08230__A1 vss _03823_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09946_ vdd _04933_ _04932_ _01207_ _04918_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06792__A1 vss _02876_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09730__A1 vss _04781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09877_ vdd vss _04891_ rf_ram.memory\[239\]\[0\] _04890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05914__B vss _01916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08828_ vdd vss _04215_ rf_ram.memory\[135\]\[1\] _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06544__A1 vss _01347_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output216_I vss net216 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08759_ vdd vss _04172_ _01363_ _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_178_771 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08297__A1 vss _03855_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_224 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_410 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10721_ vdd rf_ram.memory\[462\]\[1\] clknet_leaf_120_clk vss _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_819 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08049__A1 vss _03690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10652_ vdd rf_ram.memory\[381\]\[0\] clknet_leaf_107_clk vss _00396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_465 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_482 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10583_ vdd rf_ram.memory\[322\]\[1\] clknet_leaf_163_clk vss _00327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_893 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09797__A1 vss net245 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09261__A3 vss cpu.decode.co_ebreak vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_173_clk_I vss clknet_5_31__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1173 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06480__B1 vss _01655_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_53_clk_I vss clknet_5_12__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11204_ vdd rf_ram.memory\[84\]\[0\] clknet_leaf_49_clk vss _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07024__A2 vss _02813_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08221__A1 vss _03798_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06232__B1 vss _01668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11135_ vdd rf_ram.memory\[113\]\[1\] clknet_5_10__leaf_clk vss _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_188_clk_I vss clknet_5_29__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08772__A2 vss _04152_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11066_ vdd rf_ram.memory\[137\]\[1\] clknet_leaf_11_clk vss _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_68_clk_I vss clknet_5_8__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10017_ vdd vss _04977_ rf_ram.memory\[505\]\[0\] _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09721__A1 vss _04781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_111_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_546 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08288__A1 vss _03230_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10095__A1 vss _02814_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_126_clk_I vss clknet_5_13__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10919_ vdd rf_ram.memory\[177\]\[1\] clknet_leaf_16_clk vss _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_936 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27_622 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_660 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06110_ _02304_ vdd vss _02305_ _01603_ _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07090_ vdd vss _03119_ rf_ram.memory\[490\]\[1\] _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07263__A2 vss _02883_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06041_ vdd vss _02236_ rf_ram.memory\[356\]\[1\] _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_989 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_568 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_112_535 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07992_ vdd vss _03681_ rf_ram.memory\[477\]\[1\] _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09800_ vdd vss _04844_ rf_ram.memory\[58\]\[1\] _04842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09731_ _04791_ _04798_ vdd vss _04799_ net108 _04790_ net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06943_ vdd _03024_ _03023_ _00112_ _03014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06874_ vdd vss _02978_ rf_ram.memory\[282\]\[0\] _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_809 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_1021 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09662_ vdd vss net120 _04747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_94_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08613_ vdd vss _04081_ rf_ram.memory\[129\]\[1\] _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05825_ _02020_ vdd vss _02021_ _01951_ _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09593_ vdd vss _04704_ _04477_ cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08544_ vdd vss _04036_ rf_ram.memory\[171\]\[1\] _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05756_ vdd vss _01952_ rf_ram.memory\[158\]\[0\] _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_82_95 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09720__I vss _04760_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06829__A2 vss _02946_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05687_ _01693_ vdd vss _01883_ rf_ram.memory\[392\]\[0\] _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_599 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08475_ vdd vss _00680_ _01436_ _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_402 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07426_ vdd _03329_ _03328_ _00290_ _03323_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_238 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_295 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09779__A1 vss _04637_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07357_ vdd _03285_ _03283_ _00265_ _03260_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_614 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06308_ vdd vss _02503_ rf_ram.memory\[174\]\[1\] _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08451__A1 vss _02714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_636 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_693 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_811 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07288_ vdd vss _03243_ rf_ram.memory\[471\]\[1\] _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09027_ vdd vss _04338_ rf_ram.memory\[107\]\[1\] _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06239_ rf_ram.memory\[438\]\[1\] _02434_ vss vdd rf_ram.memory\[437\]\[1\] _01931_
+ rf_ram.memory\[439\]\[1\] _01911_ _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_130_321 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09400__B1 vss _04564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08203__A1 vss _03790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09951__A1 vss _04918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10010__A1 vss _04953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05568__A2 vss _01500_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09929_ vdd vss _04923_ _04911_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09703__A1 vss _04740_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08506__A2 vss cpu.immdec.imm11_7\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06517__A1 vss _02703_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05740__A2 vss _01724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10077__A1 vss _04985_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10704_ vdd rf_ram.memory\[431\]\[0\] clknet_leaf_99_clk vss _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07493__A2 vss _03101_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08690__A1 vss _04126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_181_755 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_273 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10635_ vdd rf_ram.memory\[404\]\[1\] clknet_leaf_114_clk vss _00379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_435 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_413 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_649 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_126 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_441 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_964 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_975 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_159 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10566_ vdd rf_ram.memory\[328\]\[0\] clknet_leaf_157_clk vss _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_967 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10497_ vdd rf_ram.memory\[468\]\[1\] clknet_leaf_53_clk vss _00241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06205__B1 vss _01811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11118_ vdd rf_ram.memory\[121\]\[0\] clknet_leaf_84_clk vss _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput7 vss net7 i_dbus_rdt[14] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11049_ vdd rf_ram.memory\[143\]\[0\] clknet_leaf_10_clk vss _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05610_ _01805_ vdd vss _01806_ rf_ram.memory\[318\]\[0\] _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_118_1050 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07181__A1 vss _03157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_376 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05731__A2 vss _01719_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10068__A1 vss _02838_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06590_ vdd vss _02770_ _02752_ _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_1004 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05541_ vss vdd rf_ram.memory\[277\]\[0\] _01678_ rf_ram.memory\[279\]\[0\] _01679_
+ _01687_ rf_ram.memory\[278\]\[0\] _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__06141__C1 vss _01713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05472_ _01668_ _01655_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_15_1066 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08681__A1 vss _04097_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08260_ vdd _03848_ _03846_ _00605_ _03823_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_166_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07211_ vdd vss _03195_ _02795_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08191_ vdd _03806_ _03805_ _00578_ _03787_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_7_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_446 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07142_ vdd vss _03152_ rf_ram.memory\[485\]\[0\] _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07236__A2 vss _03040_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_287 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08433__A1 vss _03956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09481__I0 vss net89 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07073_ vdd vss _03109_ rf_ram.memory\[493\]\[0\] _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_294_clk vdd vss clknet_leaf_294_clk clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05798__A2 vss _01958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06024_ _01528_ vdd vss _02219_ rf_ram.memory\[544\]\[1\] _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09933__A1 vss _04921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07975_ vdd _03670_ _03669_ _00498_ _03651_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06926_ vdd _03012_ _03010_ _00107_ _02975_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09714_ _04768_ _04786_ vdd vss _04787_ net103 _04767_ net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06857_ vdd vss _02966_ rf_ram.memory\[284\]\[1\] _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05970__A2 vss _01514_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09645_ _01376_ _04732_ cpu.mem_bytecnt\[1\] _01375_ _01385_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_05808_ _02004_ _01504_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_171_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06788_ vdd vss _02918_ _02915_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09576_ vss _01080_ _04689_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05739_ _01805_ vdd vss _01935_ rf_ram.memory\[430\]\[0\] _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08527_ vdd _04025_ _04024_ _00695_ _04023_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_925 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08458_ vdd vss _03975_ _03973_ _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08672__A1 vss _02838_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_20__f_clk vdd vss clknet_5_20__leaf_clk clknet_3_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07409_ vdd vss _03318_ rf_ram.memory\[372\]\[1\] _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_344 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_964 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_619 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10420_ vdd rf_ram.memory\[490\]\[0\] clknet_leaf_183_clk vss _00164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08389_ vdd _03929_ _03927_ _00653_ _03922_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08424__A1 vss _03919_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05238__A1 vss net134 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10351_ vdd rf_ram.memory\[281\]\[1\] clknet_leaf_180_clk vss _00095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10231__A1 vss _05078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_285_clk vdd vss clknet_leaf_285_clk clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10282_ vdd rf_ram.memory\[346\]\[0\] clknet_leaf_141_clk vss _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06738__A1 vss _02876_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05946__C1 vss _01609_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_3__f_clk_I vss clknet_3_0_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_606 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_1060 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09561__S vss _04678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07163__A1 vss _03161_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_650 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06984__I vss _03013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06371__C1 vss _01702_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_897 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05477__A1 vss _01600_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_344 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_446 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11667_ net190 vss vdd net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10618_ vdd rf_ram.memory\[313\]\[0\] clknet_leaf_105_clk vss _00362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_405 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_682 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05229__A1 vss cpu.alu.i_rs1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11598_ vdd rf_ram.rdata\[1\] clknet_leaf_281_clk vss _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09463__I0 vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10549_ vdd rf_ram.memory\[370\]\[1\] clknet_leaf_149_clk vss _00293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_276_clk vdd vss clknet_leaf_276_clk clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_110_825 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_696 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_195 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07760_ vdd vss _03537_ rf_ram.memory\[376\]\[1\] _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05401__A1 vss _01369_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05952__A2 vss _01613_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06711_ vdd _02861_ _02859_ _00043_ _02826_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09471__S vss _04604_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07691_ vdd _03494_ _03493_ _00390_ _03488_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_200_clk vdd vss clknet_leaf_200_clk clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09430_ vss _01033_ _04590_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_177_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06901__A1 vss _02975_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05165__B1 vss _01367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06642_ vdd vss _02810_ _02756_ _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_177_869 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06573_ vdd _02755_ _02753_ _00011_ _02748_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09361_ _04552_ vss vdd _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_05524_ _01707_ vdd vss _01720_ rf_ram.memory\[334\]\[0\] _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09292_ vdd _04510_ _04508_ _00975_ _04466_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08312_ vdd _03880_ _03878_ _00625_ _03855_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08654__A1 vss _04094_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_547 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08243_ vdd _03838_ _03837_ _00598_ _03820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05455_ _01650_ vdd vss _01651_ rf_ram.memory\[376\]\[0\] _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_145_777 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_826 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1240 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09454__I0 vss net77 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05386_ _01505_ vdd vss _01582_ rf_ram.memory\[566\]\[0\] _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08174_ vdd vss _03796_ rf_ram.memory\[542\]\[0\] _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10213__A1 vss _05081_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07125_ vdd _03141_ _03139_ _00177_ _03126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_267_clk vdd vss clknet_leaf_267_clk clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_31_937 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07056_ vdd vss _03098_ rf_ram.memory\[38\]\[0\] _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_61 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09906__A1 vss _03445_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput152 o_ext_rs1[22] net152 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput141 o_ext_rs1[12] net141 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput130 o_dbus_sel[0] net130 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08709__A2 vss _04078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06007_ _01552_ vdd vss _02202_ rf_ram.memory\[528\]\[1\] _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput185 o_ext_rs2[23] net185 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput174 o_ext_rs2[13] net174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_input42_I vss i_ibus_rdt[17] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput163 o_ext_rs1[3] net163 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05928__C1 vss _01696_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05906__C vss _01362_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput196 o_ext_rs2[4] net196 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_177_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07958_ vdd vss _03660_ rf_ram.memory\[480\]\[0\] _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05943__A2 vss _01605_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07889_ vdd vss _03617_ rf_ram.memory\[445\]\[0\] _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06909_ vdd vss _03001_ _02822_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07145__A1 vss _03126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output129_I vss net129 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05922__B vss _02004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09628_ vdd _04663_ _01447_ _01099_ _04643_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_683 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09559_ vdd vss _04677_ _01491_ _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05171__A3 vss _01372_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_761 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11521_ vdd rf_ram.memory\[307\]\[0\] clknet_leaf_150_clk vss _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_777 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06120__A2 vss _01644_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11452_ vdd rf_ram.memory\[229\]\[1\] clknet_leaf_281_clk vss _01184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11383_ _01115_ vdd vss clknet_5_23__leaf_clk net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10403_ vdd rf_ram.memory\[215\]\[1\] clknet_leaf_301_clk vss _00147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10204__A1 vss _03892_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_258_clk vdd vss clknet_leaf_258_clk clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10334_ vdd rf_ram.memory\[286\]\[0\] clknet_leaf_174_clk vss _00078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1237 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_308 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_103_162 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10265_ vdd rf_ram.memory\[200\]\[1\] clknet_leaf_33_clk vss _00009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05919__C1 vss _01786_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10196_ vdd _05087_ _05086_ _01303_ _05078_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07384__A1 vss _03292_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06187__A2 vss _01777_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05934__A2 vss _01530_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07136__A1 vss _02915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08884__A1 vss _04234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06344__C1 vss _01645_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_119 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_519 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_69 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07439__A2 vss _02883_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_675 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08636__A1 vss _02893_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_574 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_777 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput10 vss net10 i_dbus_rdt[17] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 vss net21 i_dbus_rdt[27] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_859 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05240_ _01439_ vdd vss _01440_ _01430_ _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__08939__A2 vss _04038_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput32 vss net32 i_dbus_rdt[8] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05171_ _01372_ _01373_ vdd vss _01374_ _01368_ _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xinput54 vss net54 i_ibus_rdt[29] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_249_clk vdd vss clknet_leaf_249_clk clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_24_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput43 vss net43 i_ibus_rdt[18] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput65 net65 vss vdd i_rst vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08930_ vdd vss _04278_ rf_ram.memory\[123\]\[0\] _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05793__I vss _01640_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08861_ vdd vss _04235_ _02983_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07812_ vdd vss _03570_ rf_ram.memory\[434\]\[0\] _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06178__A2 vss _01500_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07375__A1 vss _03055_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05925__A2 vss _01863_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_30 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08792_ vdd vss _04192_ net246 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07743_ vdd vss _03527_ rf_ram.memory\[396\]\[0\] _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07127__A1 vss rf_ram.memory\[4\]\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07674_ vdd _03483_ _03482_ _00384_ _03455_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08609__I vss _04077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09413_ vdd vss _04582_ rf_ram.memory\[299\]\[0\] _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06625_ vdd vss _02797_ _02796_ _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09344_ _04540_ net227 vdd vss _04543_ net224 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08627__A1 vss _04058_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06556_ _02742_ vss vdd _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_168_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05507_ vss vdd rf_ram.memory\[341\]\[0\] _01702_ rf_ram.memory\[343\]\[0\] _01688_
+ _01623_ rf_ram.memory\[342\]\[0\] _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__06102__A2 vss _01623_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06487_ rf_ram.memory\[3\]\[1\] _01635_ _01661_ rf_ram.memory\[2\]\[1\] _02682_ vss
+ vdd rf_ram.memory\[1\]\[1\] _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_09275_ vss _00970_ _04498_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_160_511 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05438_ _01634_ _01633_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09427__I0 vss net94 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08226_ vdd vss _03828_ _03798_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08157_ vdd vss _03785_ rf_ram.memory\[545\]\[0\] _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09052__A1 vss _04331_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07108_ vdd _03130_ _03128_ _00171_ _03126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05369_ _01561_ _01564_ vdd vss _01565_ _01558_ _01559_ _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08088_ vdd vss _03742_ _02971_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_1065 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05917__B vss _01928_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07039_ vdd vss _03086_ rf_ram.memory\[215\]\[1\] _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_1210 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10050_ vdd _04997_ _04996_ _01247_ _04982_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06169__A2 vss _01631_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07366__A1 vss _03289_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1287 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05916__A2 vss _01706_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09107__A2 vss _04005_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07118__A1 vss _03123_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08866__A1 vss _04237_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06326__C1 vss _01968_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10952_ vdd rf_ram_if.wen0_r clknet_leaf_259_clk vss _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_1183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_299 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06341__A2 vss _01649_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10883_ vdd rf_ram.memory\[220\]\[1\] clknet_leaf_31_clk vss _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_839 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_517 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_360 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11504_ vdd rf_ram.memory\[505\]\[1\] clknet_leaf_198_clk vss _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_336 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_80_166 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_712 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11435_ _01167_ vdd vss clknet_leaf_242_clk cpu.state.cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_85_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11366_ _01098_ vdd vss clknet_leaf_235_clk cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09594__A2 vss net46 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11297_ _01030_ vdd vss clknet_leaf_252_clk net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_0_138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10317_ vdd rf_ram.memory\[512\]\[1\] clknet_leaf_268_clk vss _00061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10248_ vdd _05118_ _05116_ _01324_ _02825_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09346__A2 vss _03991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07357__A1 vss _03260_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05907__A2 vss _01510_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10179_ vdd _05076_ _05075_ _01297_ _05046_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07109__A1 vss _02728_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08857__A1 vss _04202_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06377__C vss _01860_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06410_ rf_ram.memory\[118\]\[1\] _02605_ vss vdd rf_ram.memory\[117\]\[1\] _01931_
+ rf_ram.memory\[119\]\[1\] _01911_ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__06332__A2 vss _01537_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07390_ vdd vss _03306_ _02752_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06341_ rf_ram.memory\[204\]\[1\] _02536_ vss vdd rf_ram.memory\[207\]\[1\] _01925_
+ rf_ram.memory\[205\]\[1\] _01912_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__06096__A1 vss _01368_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_574 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09060_ vdd vss _04358_ net241 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_634 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06272_ vdd vss _02467_ rf_ram.memory\[153\]\[1\] _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_53_870 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05223_ vdd _01383_ _01422_ _01423_ _01421_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08011_ vdd vss _03695_ rf_ram.memory\[573\]\[0\] _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09034__A1 vss _04334_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_391 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_756 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_531 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05154_ vdd vss _01357_ _01347_ _01356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09962_ vdd vss _04943_ rf_ram.memory\[335\]\[1\] _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06399__A2 vss _01683_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08913_ vdd vss _04267_ _03039_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07348__A1 vss _02813_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09893_ vdd _04900_ _04899_ _01187_ _04884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08844_ vdd _04224_ _04222_ _00813_ _04205_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05987_ _02182_ vdd vss _02183_ _01348_ _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08775_ vdd vss _04182_ rf_ram.memory\[143\]\[1\] _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07726_ vdd vss _03516_ rf_ram.memory\[37\]\[0\] _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_931 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07520__A1 vss _03356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07657_ vdd vss _03473_ rf_ram.memory\[404\]\[0\] _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07588_ vdd vss _03430_ _02889_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05531__B1 vss _01725_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_176 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06608_ vdd _02783_ _02782_ _00018_ _02743_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09327_ vdd _04532_ _04530_ _00988_ _04466_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_303 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06539_ vdd vss _02725_ _02723_ _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_168_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09258_ _04482_ _04483_ _04485_ vdd vss _00966_ _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_44_870 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_706 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09189_ vdd vss _04439_ net242 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08209_ vdd vss _03817_ _03798_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11220_ vdd rf_ram.memory\[349\]\[0\] clknet_leaf_192_clk vss _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07587__A1 vss _03425_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11151_ vdd rf_ram.memory\[105\]\[1\] clknet_leaf_68_clk vss _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_max_cap242_I vss _02865_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09328__A2 vss _03072_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10102_ vdd _05029_ _05028_ _01267_ _05014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05598__B1 vss _01778_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output73_I vss net73 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11082_ vdd rf_ram.memory\[131\]\[1\] clknet_leaf_28_clk vss _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10033_ vdd vss _04987_ _02805_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05382__B vss _01528_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_942 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08839__A1 vss _04205_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_575 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06314__A2 vss _01989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10935_ vdd rf_ram_if.wdata1_r\[2\] clknet_leaf_261_clk vss cpu.o_wdata1 vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_151_1061 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10866_ vdd rf_ram.memory\[195\]\[0\] clknet_leaf_46_clk vss _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_781 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_124_500 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_133 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10797_ vdd rf_ram.memory\[558\]\[1\] clknet_leaf_319_clk vss _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_511 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05825__A1 vss _01951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_509 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_358 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09016__A1 vss _04301_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11418_ vdd rf_ram.memory\[58\]\[1\] clknet_leaf_287_clk vss _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11349_ vdd cpu.immdec.imm30_25\[5\] clknet_leaf_254_clk vss _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09319__A2 vss net35 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05910_ _01916_ vdd vss _02106_ rf_ram.memory\[112\]\[0\] _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06890_ vdd vss _02988_ _02788_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05841_ _01916_ vdd vss _02037_ rf_ram.memory\[200\]\[0\] _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06388__B vss _01551_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06553__A2 vss _02738_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08560_ vdd _04046_ _04045_ _00707_ _04023_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05772_ _01968_ vss vdd _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_187_761 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07511_ vdd vss _03382_ rf_ram.memory\[323\]\[1\] _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07502__A1 vss _03360_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08491_ vdd vss _04000_ rf_ram.memory\[369\]\[1\] _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06305__A2 vss _01664_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07442_ vdd vss _03339_ rf_ram.memory\[36\]\[1\] _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_76_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_1__f_clk vdd vss clknet_5_1__leaf_clk clknet_3_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07373_ vdd vss _03296_ rf_ram.memory\[267\]\[1\] _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09112_ vdd vss _04390_ _02959_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_965 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06324_ _02518_ vdd vss _02519_ net251 _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_06255_ _01650_ vdd vss _02450_ rf_ram.memory\[426\]\[1\] _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09007__A1 vss _02971_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09043_ vdd vss _04348_ rf_ram.memory\[104\]\[1\] _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_497 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06186_ vdd vss _02381_ rf_ram.memory\[465\]\[1\] _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05206_ vdd vss _01406_ cpu.decode.co_mem_word _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_309_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05137_ _01339_ vdd vss _01340_ cpu.decode.op21 _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__05467__B vss _01504_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_1035 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09945_ vdd vss _04933_ rf_ram.memory\[338\]\[0\] _04932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09876_ vdd vss _04890_ _03309_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09730__A2 vss net12 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08827_ vdd _04214_ _04213_ _00806_ _04202_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07741__A1 vss _03524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06544__A2 vss _01366_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08758_ vdd _04171_ _04168_ _00780_ _04170_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07709_ vdd _03505_ _03503_ _00397_ _03491_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08689_ vdd vss _04128_ rf_ram.memory\[154\]\[0\] _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_36_1131 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10720_ vdd rf_ram.memory\[462\]\[0\] clknet_leaf_50_clk vss _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_177_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10651_ vdd rf_ram.memory\[400\]\[1\] clknet_leaf_115_clk vss _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_850 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09246__A1 vss _02714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10582_ vdd rf_ram.memory\[322\]\[0\] clknet_leaf_163_clk vss _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09797__A2 vss _02921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_784 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_272 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09261__A4 vss _01460_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06480__B2 vss rf_ram.memory\[13\]\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1027 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11203_ vdd rf_ram.memory\[85\]\[1\] clknet_leaf_50_clk vss _00939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08221__A2 vss _03072_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05377__B vss _01528_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11134_ vdd rf_ram.memory\[113\]\[0\] clknet_leaf_74_clk vss _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_794 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11065_ vdd rf_ram.memory\[137\]\[0\] clknet_leaf_11_clk vss _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10016_ vdd vss _04976_ _02910_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09721__A2 vss net9 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07732__A1 vss _03488_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06001__B vss _01528_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08288__A2 vss _02904_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_361 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09485__A1 vss _01411_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_400 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10095__A2 vss _02909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10918_ vdd rf_ram.memory\[177\]\[0\] clknet_leaf_16_clk vss _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06299__A1 vss _01552_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_69 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10849_ vdd rf_ram.memory\[532\]\[1\] clknet_leaf_310_clk vss _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_280_clk_I vss clknet_5_19__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_125_897 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06040_ vdd vss _02235_ _02211_ _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06223__A1 vss _01675_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07991_ vdd _03680_ _03679_ _00504_ _03651_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_295_clk_I vss clknet_5_7__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1219 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07971__A1 vss _03654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09730_ vdd vss _04798_ _04781_ net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06942_ vdd vss _03024_ rf_ram.memory\[206\]\[0\] _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_589 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06873_ vdd vss _02977_ _02813_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09661_ _04745_ _04746_ vdd vss _01108_ _03974_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_1142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08612_ vdd _04080_ _04079_ _00725_ _04058_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05824_ rf_ram.memory\[215\]\[0\] _02019_ _01940_ rf_ram.memory\[214\]\[0\] _02020_
+ vss vdd rf_ram.memory\[213\]\[0\] _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__05306__I vss _01501_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09592_ vdd _01491_ _04698_ _04703_ _01469_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_171_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_512 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05755_ _01951_ _01693_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08543_ vdd _04035_ _04034_ _00701_ _04023_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_106_81 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_85 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_233_clk_I vss clknet_5_23__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05686_ _01881_ vdd vss _01882_ _01769_ _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08474_ rf_ram.rdata\[1\] vdd vss _03988_ _01378_ rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_174_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07425_ vdd vss _03329_ rf_ram.memory\[333\]\[0\] _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_989 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09228__A1 vss _04434_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_617 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_559 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_781 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_959 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07356_ vdd vss _03285_ rf_ram.memory\[252\]\[1\] _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07287_ vdd _03242_ _03241_ _00238_ _03222_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_1102 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_248_clk_I vss clknet_5_21__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_689 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_497 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06307_ _01564_ vdd vss _02502_ _02499_ _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06238_ vdd vss _02433_ rf_ram.memory\[436\]\[1\] _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09026_ vdd _04337_ _04336_ _00882_ _04331_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_115_374 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05265__A2 vss cpu.decode.co_ebreak vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06169_ vdd vss _02364_ rf_ram.memory\[510\]\[1\] _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08203__A2 vss _03811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09928_ vdd _04922_ _04919_ _01200_ _04921_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07962__A1 vss _02836_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1066 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_125 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07714__A1 vss _03491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09703__A2 vss net4 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09859_ vdd _04870_ _04879_ _04880_ _04878_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09911__I vss _02814_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10703_ vdd rf_ram.memory\[411\]\[1\] clknet_leaf_90_clk vss _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09219__A1 vss _03319_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_617 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10634_ vdd rf_ram.memory\[404\]\[0\] clknet_leaf_102_clk vss _00378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10565_ vdd rf_ram.memory\[366\]\[1\] clknet_leaf_171_clk vss _00309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_992 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_84_1235 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06453__A1 vss _01526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_480 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10496_ vdd rf_ram.memory\[468\]\[0\] clknet_leaf_53_clk vss _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_856 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_467 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_121_344 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10001__A2 vss _02992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11117_ vdd rf_ram.memory\[449\]\[1\] clknet_leaf_113_clk vss _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07705__A1 vss _02960_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 vss net8 i_dbus_rdt[15] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11048_ vdd rf_ram.memory\[144\]\[1\] clknet_leaf_337_clk vss _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_832 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05192__A1 vss _01391_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05570__B vss _01349_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05540_ vdd vss _01736_ rf_ram.memory\[276\]\[0\] _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10068__A2 vss _03158_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1102 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_1023 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08130__A1 vss _03757_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_20__f_clk_I vss clknet_3_5_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05471_ _01526_ vdd vss _01667_ rf_ram.memory\[368\]\[0\] _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06141__B1 vss _01715_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07210_ vdd _03194_ _03191_ _00209_ _03193_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08190_ vdd vss _03806_ rf_ram.memory\[53\]\[0\] _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06692__A1 vss _02788_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09469__S vss _04604_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_244 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07141_ vdd vss _03151_ _02795_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_497 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09630__A1 vss _04643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07072_ vdd vss _03108_ _02844_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_489 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06023_ rf_ram.memory\[549\]\[1\] _01539_ _01538_ rf_ram.memory\[548\]\[1\] _02218_
+ vss vdd rf_ram.memory\[551\]\[1\] _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_2_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09394__B1 vss _04564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08736__A3 vss _03984_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07944__A1 vss _03622_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05745__B vss _01805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07974_ vdd vss _03670_ rf_ram.memory\[46\]\[0\] _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_1139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06925_ vdd vss _03012_ rf_ram.memory\[278\]\[1\] _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09713_ vdd vss _04786_ _04781_ net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__09697__A1 vss _04740_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06856_ vdd _02965_ _02964_ _00084_ _02927_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09644_ vdd vss _04731_ cpu.mem_bytecnt\[1\] _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_172_clk_I vss clknet_5_30__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1031 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05807_ _01999_ _02002_ vdd vss _02003_ _01991_ _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09575_ _04678_ vdd vss _04689_ cpu.immdec.imm30_25\[4\] _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06787_ _02917_ vss vdd _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05738_ _01929_ _01933_ vdd vss _01934_ _01914_ _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA_clkbuf_leaf_52_clk_I vss clknet_5_9__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_364 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08347__I vss _03902_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08526_ vdd vss _04025_ rf_ram.memory\[49\]\[0\] _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_175_550 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05669_ _01864_ vdd vss _01865_ _01769_ _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_93_835 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06295__C vss _01349_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08457_ vdd vss net109 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08672__A2 vss _04078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07408_ vdd _03317_ _03316_ _00284_ _03289_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_187_clk_I vss clknet_5_28__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_976 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06683__A1 vss _02750_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05891__C1 vss _01912_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08388_ vdd vss _03929_ rf_ram.memory\[189\]\[1\] _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07339_ vdd vss _03275_ rf_ram.memory\[270\]\[0\] _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_116_672 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_67_clk_I vss clknet_5_8__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09621__A1 vss _02828_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_110_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10350_ vdd rf_ram.memory\[281\]\[0\] clknet_leaf_180_clk vss _00094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06435__A1 vss _01569_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_776 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05238__A2 vss _01436_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10281_ vdd rf_ram.memory\[294\]\[1\] clknet_leaf_143_clk vss _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09009_ vdd _04326_ _04325_ _00876_ _04298_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_344 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_692 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_163 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08188__A1 vss _03790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07935__A1 vss _02752_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_125_clk_I vss clknet_5_13__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05655__B vss _01693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05946__B1 vss _01607_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1149 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09688__A1 vss _04740_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05374__C vss _01569_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08360__A1 vss _03884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06486__B vss _01525_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_128 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06371__B1 vss _01625_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_731 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_504 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11383__CLK vss clknet_5_23__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_762 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11666_ net189 vss vdd net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_4_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10617_ vdd rf_ram.memory\[353\]\[1\] clknet_leaf_156_clk vss _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09612__A1 vss _04637_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11597_ vdd rf_ram.rdata\[0\] clknet_leaf_282_clk vss _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09463__I1 vss net82 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_283 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_220 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10548_ vdd rf_ram.memory\[370\]\[0\] clknet_leaf_149_clk vss _00292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_940 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_160 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05634__C1 vss _01678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10479_ vdd rf_ram.memory\[421\]\[1\] clknet_leaf_104_clk vss _00223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_651 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08179__A1 vss _03798_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09679__A1 vss net1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06710_ vdd vss _02861_ rf_ram.memory\[521\]\[1\] _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07690_ vdd vss _03494_ rf_ram.memory\[401\]\[0\] _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06641_ vdd _02809_ _02807_ _00025_ _02748_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05165__A1 vss _01353_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06362__B1 vss _01953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06572_ vdd vss _02755_ rf_ram.memory\[201\]\[1\] _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08103__A1 vss _02780_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09360_ vdd vss _04551_ _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_164_509 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09291_ vdd vss _04510_ rf_ram.memory\[65\]\[1\] _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05523_ _01719_ _01686_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08311_ vdd vss _03880_ rf_ram.memory\[243\]\[1\] _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_274 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05454_ _01650_ _01601_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08242_ vdd vss _03838_ rf_ram.memory\[52\]\[0\] _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09851__A1 vss _02713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_726 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09603__A1 vss _04643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05385_ _01580_ vdd vss _01581_ _01495_ _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_6_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09454__I1 vss net78 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08173_ vdd vss _03795_ _02881_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07124_ vdd vss _03141_ rf_ram.memory\[487\]\[1\] _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07055_ vdd vss _03097_ _02806_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_140_472 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05640__A2 vss _01755_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput131 o_dbus_sel[1] net131 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput142 o_ext_rs1[13] net142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput120 o_dbus_dat[2] net120 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06006_ rf_ram.memory\[532\]\[1\] _02201_ vss vdd rf_ram.memory\[535\]\[1\] _01520_
+ rf_ram.memory\[533\]\[1\] _01516_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__09906__A2 vss _02883_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput186 o_ext_rs2[24] net186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07917__A1 vss _03619_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput175 o_ext_rs2[14] net175 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput153 o_ext_rs1[23] net153 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput164 o_ext_rs1[4] net164 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05928__B1 vss _01848_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput197 o_ext_rs2[5] net197 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_07957_ vdd vss _03659_ _02903_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_103_1183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input35_I vss i_ibus_rdt[10] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06908_ vdd _03000_ _02998_ _00101_ _02975_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07888_ vdd vss _03616_ _02959_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_168_837 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09627_ vdd _04660_ _01400_ _01098_ _04643_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06839_ vdd vss _02953_ _02779_ _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_167_336 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09558_ _02711_ vdd vss _04676_ _01469_ _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_183_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05171__A4 vss _01373_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08509_ _01469_ _04012_ _01399_ vdd vss _04013_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_182_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_108_414 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11520_ vdd rf_ram.memory\[507\]\[1\] clknet_leaf_199_clk vss _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09489_ _04624_ _04616_ vdd vss _01058_ _02690_ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09842__A1 vss _02714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_559 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09410__B vss _04539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_710 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11451_ vdd rf_ram.memory\[229\]\[0\] clknet_leaf_281_clk vss _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06408__A1 vss _01768_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11382_ _01114_ vdd vss clknet_leaf_229_clk net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_61_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10204__A2 vss _02866_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10402_ vdd rf_ram.memory\[215\]\[0\] clknet_leaf_301_clk vss _00146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05369__C vss _01564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05616__C1 vss _01811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10333_ vdd rf_ram.memory\[304\]\[1\] clknet_leaf_146_clk vss _00077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_951 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07081__A1 vss _03092_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_984 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05631__A2 vss _01777_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10264_ vdd rf_ram.memory\[200\]\[0\] clknet_leaf_33_clk vss _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05919__B1 vss _01931_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10195_ vdd vss _05087_ rf_ram.memory\[210\]\[0\] _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07156__I vss _03017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09572__S vss _04678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07136__A2 vss _02923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08333__A1 vss _03884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08884__A2 vss _04248_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_194_clk vdd vss clknet_leaf_194_clk clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06344__B1 vss _01636_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06895__A1 vss _02716_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05404__I vss _01599_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08636__A2 vss _04067_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_378 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_895 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput11 vss net11 i_dbus_rdt[18] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11649_ vss net171 net99 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput22 vss net22 i_dbus_rdt[28] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09436__I1 vss net69 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_69 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput33 vss net33 i_dbus_rdt[9] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05170_ cpu.immdec.imm19_12_20\[8\] _01367_ cpu.immdec.imm24_20\[4\] vdd vss _01373_
+ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
Xinput55 vss net55 i_ibus_rdt[2] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput44 vss net44 i_ibus_rdt[19] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_122_450 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07072__A1 vss _02844_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput66 vss net66 i_timer_irq vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_656 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05622__A2 vss _01543_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06280__C1 vss _01968_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08860_ _04234_ _04057_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_0_876 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07811_ vdd vss _03569_ net236 _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07375__A2 vss _02813_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08572__A1 vss _04026_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08791_ vdd _04191_ _04189_ _00793_ _04170_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_165_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07742_ vdd vss _03526_ _02788_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08324__A1 vss _03887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07673_ vdd vss _03483_ rf_ram.memory\[384\]\[0\] _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10131__A1 vss _02805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_185_clk vdd vss clknet_leaf_185_clk clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05138__A1 vss cpu.state.genblk1.misalign_trap_sync_r vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05689__A2 vss _01777_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09412_ vdd vss _04581_ net246 _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06624_ vdd vss _02796_ cpu.immdec.imm11_7\[2\] _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05314__I vss _01509_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09343_ vdd vss _04542_ _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_176_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_164_339 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09824__A1 vss _04837_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06555_ vdd _02740_ rf_ram_if.wdata1_r\[0\] _02741_ _01353_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_356 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_868 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_81 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06486_ _01525_ vdd vss _02681_ rf_ram.memory\[0\]\[1\] _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05506_ _01702_ _01609_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_12
X_09274_ _04497_ vdd vss _04498_ cpu.genblk3.csr.mcause3_0\[0\] _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05437_ _01633_ vss vdd _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08225_ vdd _03827_ _03825_ _00591_ _03823_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08156_ vdd vss _03784_ net238 _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05368_ vss _01564_ _01563_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_07107_ vdd vss _03130_ rf_ram.memory\[501\]\[1\] _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_1060 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10198__A1 vss _05081_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1033 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_792 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08087_ vdd _03741_ _03739_ _00539_ _03724_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09456__I vss _01411_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_234 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05299_ _01495_ _01494_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05613__A2 vss _01808_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06810__A1 vss _02927_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07038_ vdd _03085_ _03084_ _00146_ _03050_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_470 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_1255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08563__A1 vss _02915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06023__C1 vss _01540_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08989_ vdd _04314_ _04313_ _00868_ _04298_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05933__B vss net251 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08315__A1 vss _03852_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_176_clk vdd vss clknet_leaf_176_clk clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10122__A1 vss _05014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10951_ vdd rf_ram.memory\[79\]\[1\] clknet_leaf_18_clk vss _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06326__B1 vss _02019_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06877__A1 vss _02975_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10130__I vss _02742_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_79_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10882_ vdd rf_ram.memory\[220\]\[0\] clknet_leaf_32_clk vss _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_301 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_637 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_131 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_462 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_884 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11503_ vdd rf_ram.memory\[505\]\[0\] clknet_leaf_199_clk vss _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06483__C vss _01562_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05852__A2 vss _01614_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11434_ vdd cpu.state.cnt_r\[1\] clknet_leaf_242_clk vss _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07054__A1 vss _03092_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_100_clk vdd vss clknet_leaf_100_clk clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11365_ _01097_ vdd vss clknet_leaf_235_clk cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05604__A2 vss _01799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11296_ _01029_ vdd vss clknet_leaf_253_clk net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10316_ vdd rf_ram.memory\[512\]\[0\] clknet_leaf_271_clk vss _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10247_ vdd vss _05118_ rf_ram.memory\[264\]\[1\] _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10178_ vdd vss _05076_ rf_ram.memory\[202\]\[0\] _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07109__A2 vss _02911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05843__B vss _01860_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_167_clk vdd vss clknet_leaf_167_clk clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_187_976 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09806__A1 vss _04840_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_996 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06340_ vdd vss _02535_ rf_ram.memory\[206\]\[1\] _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06271_ _01956_ vdd vss _02466_ rf_ram.memory\[152\]\[1\] _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_25_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05222_ cpu.mem_bytecnt\[1\] vdd vss _01422_ _01385_ cpu.state.o_cnt\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08010_ vdd vss _03694_ _02959_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_865 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_167_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_898 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05153_ _01336_ vdd vss _01356_ cpu.decode.op21 _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_09961_ vdd _04942_ _04941_ _01213_ _04918_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08912_ _04266_ _04057_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07348__A2 vss _02997_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05309__I vss _01504_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09892_ vdd vss _04900_ rf_ram.memory\[18\]\[0\] _04899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08545__A1 vss _04026_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08843_ vdd vss _04224_ rf_ram.memory\[134\]\[1\] _04222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05986_ _02181_ _01493_ vdd vss _02182_ _02178_ _02179_ _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08774_ vdd _04181_ _04180_ _00786_ _04167_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06020__A2 vss _01532_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07524__I vss _03100_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10104__A1 vss _05017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07725_ vdd vss _03515_ _02795_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_158_clk vdd vss clknet_leaf_158_clk clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06859__A1 vss _02822_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_965 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07656_ vdd vss _03472_ _03088_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_80 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07587_ vdd _03429_ _03427_ _00351_ _03425_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06607_ vdd vss _02783_ rf_ram.memory\[235\]\[0\] _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09326_ vdd vss _04532_ rf_ram.memory\[109\]\[1\] _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06538_ vdd vss _02724_ rf_ram.i_raddr\[3\] _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__06087__A2 vss _01652_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_309 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07284__A1 vss _03225_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09257_ vdd vss _04485_ _04484_ _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06469_ _01624_ rf_ram.memory\[19\]\[1\] vdd vss _02664_ rf_ram.memory\[18\]\[1\]
+ _01605_ _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xclkbuf_leaf_330_clk vdd vss clknet_leaf_330_clk clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08208_ vdd _03816_ _03814_ _00585_ _03790_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output189_I vss net189 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_556 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09188_ vdd _04438_ _04436_ _00943_ _04434_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05834__A2 vss _01501_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_893 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_269 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08139_ vdd vss _03774_ rf_ram.memory\[54\]\[1\] _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07036__A1 vss _02738_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11150_ vdd rf_ram.memory\[105\]\[0\] clknet_leaf_67_clk vss _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08784__A1 vss _04167_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10101_ vdd vss _05029_ rf_ram.memory\[311\]\[0\] _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05647__C vss _01670_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_max_cap235_I vss _03082_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08536__A1 vss _02865_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11081_ vdd rf_ram.memory\[131\]\[0\] clknet_leaf_27_clk vss _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10032_ vdd _04986_ _04983_ _01240_ _04985_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06011__A2 vss _01538_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_149_clk vdd vss clknet_leaf_149_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10934_ vdd rf_ram_if.wdata1_r\[1\] clknet_leaf_261_clk vss net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_306 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10865_ vdd rf_ram.memory\[197\]\[1\] clknet_leaf_42_clk vss _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1200 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07275__A1 vss _02899_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06078__A2 vss _01687_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1079 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_112 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10796_ vdd rf_ram.memory\[558\]\[0\] clknet_leaf_320_clk vss _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_321_clk vdd vss clknet_leaf_321_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11417_ vdd rf_ram.memory\[58\]\[0\] clknet_leaf_287_clk vss _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_532 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11348_ vdd cpu.immdec.imm30_25\[4\] clknet_leaf_254_clk vss _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06250__A2 vss _01799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08527__A1 vss _04023_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11279_ _01014_ vdd vss clknet_leaf_244_clk net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_158_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05840_ _02035_ vdd vss _02036_ _01972_ _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__06002__A2 vss _01544_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_1259 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07510_ vdd _03381_ _03380_ _00322_ _03356_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05771_ vdd vss _01967_ rf_ram.memory\[148\]\[0\] _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08490_ vdd _03999_ _03998_ _00684_ _03953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07441_ vdd _03338_ _03337_ _00296_ _03323_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_1076 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07372_ vdd _03295_ _03294_ _00270_ _03289_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_119_328 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06069__A2 vss _01543_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09111_ vdd _04389_ _04387_ _00915_ _04367_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06323_ _02517_ _01569_ vdd vss _02518_ _01768_ _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__09255__A2 vss _01356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_312_clk vdd vss clknet_leaf_312_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06254_ rf_ram.memory\[428\]\[1\] _02449_ vss vdd rf_ram.memory\[431\]\[1\] _01726_
+ rf_ram.memory\[429\]\[1\] _01725_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_170_640 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09007__A2 vss _04303_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09042_ vdd _04347_ _04346_ _00888_ _04331_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05816__A2 vss _01922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_893 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06185_ _01693_ vdd vss _02380_ rf_ram.memory\[464\]\[1\] _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05205_ vdd vss _01405_ cpu.decode.co_mem_word cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06226__C1 vss _01608_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_397 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05136_ vdd vss _01339_ cpu.decode.opcode\[2\] cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_29_1183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08766__A1 vss _04170_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09944_ vdd vss _04932_ _04911_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06241__A2 vss _01782_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08518__A1 vss _03956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1259 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09875_ vdd vss _01180_ _02713_ _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09191__A1 vss _04431_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08826_ vdd vss _04214_ rf_ram.memory\[135\]\[0\] _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_1051 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_169_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05752__A1 vss net252 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05969_ _01550_ vdd vss _02165_ rf_ram.memory\[24\]\[0\] _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08757_ vdd vss _04171_ rf_ram.memory\[146\]\[1\] _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07708_ vdd vss _03505_ rf_ram.memory\[381\]\[1\] _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_71_1034 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08688_ vdd vss _04127_ _02812_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_913 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07639_ vdd vss _03462_ rf_ram.memory\[406\]\[1\] _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output104_I vss net104 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_434 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10650_ vdd rf_ram.memory\[400\]\[0\] clknet_leaf_115_clk vss _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07257__A1 vss _02894_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09309_ _04013_ vdd vss _04521_ _04477_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_10581_ vdd rf_ram.memory\[362\]\[1\] clknet_leaf_162_clk vss _00325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_303_clk vdd vss clknet_leaf_303_clk clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_133_342 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06465__C1 vss _01617_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_476 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_1174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05658__B vss _01790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_578 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07009__A1 vss _03050_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06480__A2 vss _01643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_392 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_126 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11202_ vdd rf_ram.memory\[85\]\[0\] clknet_leaf_49_clk vss _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06232__A2 vss _01509_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11133_ vdd rf_ram.memory\[114\]\[1\] clknet_leaf_74_clk vss _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11064_ vdd rf_ram.memory\[138\]\[1\] clknet_leaf_11_clk vss _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10015_ vdd _04975_ _04973_ _01234_ _04953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05991__A1 vss _02017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05393__B vss _01528_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09485__A2 vss _03989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10917_ vdd rf_ram.memory\[178\]\[1\] clknet_leaf_16_clk vss _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_760 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_1074 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_618 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05412__I vss _01607_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_955 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10848_ vdd rf_ram.memory\[532\]\[0\] clknet_leaf_311_clk vss _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07248__A1 vss _03190_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_415 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_117 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_679 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10779_ vdd rf_ram.memory\[567\]\[1\] clknet_leaf_328_clk vss _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08996__A1 vss _04301_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_498 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06471__A2 vss _01682_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_857 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07420__A1 vss _03323_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07990_ vdd vss _03680_ rf_ram.memory\[477\]\[0\] _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06941_ vdd vss _03023_ _02738_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06399__B vss _01684_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09660_ _04736_ vdd vss _04746_ net1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06872_ vdd _02976_ _02973_ _00089_ _02975_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_119_1019 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_1045 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08611_ vdd vss _04080_ rf_ram.memory\[129\]\[0\] _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1056 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05823_ _02019_ _01695_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09591_ vss _01082_ _04702_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_173_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05754_ _01949_ vdd vss _01950_ _01373_ _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_08542_ vdd vss _04035_ rf_ram.memory\[171\]\[0\] _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_570 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07487__A1 vss _03360_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08473_ vss _00679_ _03987_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07424_ vdd vss _03328_ _03319_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05685_ rf_ram.memory\[397\]\[0\] _01772_ _01711_ rf_ram.memory\[396\]\[0\] _01881_
+ vss vdd rf_ram.memory\[399\]\[0\] _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_175_798 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07355_ vdd _03284_ _03283_ _00264_ _03257_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_169_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08987__A1 vss net236 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07286_ vdd vss _03242_ rf_ram.memory\[471\]\[0\] _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06306_ _01520_ rf_ram.memory\[171\]\[1\] vdd vss _02501_ rf_ram.memory\[170\]\[1\]
+ _01989_ _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06237_ _02419_ _02431_ net254 vdd vss _02432_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_09025_ vdd vss _04337_ rf_ram.memory\[107\]\[0\] _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_868 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input65_I vss i_rst vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06168_ _02355_ _02359_ _02362_ vdd vss _02363_ _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_13_384 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06214__A2 vss _01697_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06099_ _02293_ vdd vss _02294_ _01675_ _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_106_1170 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09927_ vdd vss _04922_ rf_ram.memory\[342\]\[1\] _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07962__A2 vss _03009_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09164__A1 vss _04397_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08911__A1 vss _04237_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09858_ _02710_ vdd vss _04879_ _01399_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09789_ vdd _04836_ _04834_ _01146_ _04637_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08809_ vdd vss _04203_ net247 _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05941__B vss _01550_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_811 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08808__I vss _04057_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07478__A1 vss _02728_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10702_ vdd rf_ram.memory\[411\]\[0\] clknet_leaf_89_clk vss _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_80_clk vdd vss clknet_leaf_80_clk clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06150__A1 vss _01600_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09219__A2 vss _02960_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_538 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10633_ vdd rf_ram.memory\[386\]\[1\] clknet_leaf_80_clk vss _00377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10564_ vdd rf_ram.memory\[366\]\[0\] clknet_leaf_171_clk vss _00308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_1135 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07650__A1 vss _03458_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10495_ vdd rf_ram.memory\[471\]\[1\] clknet_leaf_54_clk vss _00239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_800 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05388__B vss _01552_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09575__S vss _04678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_660 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1091 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06205__A2 vss _01801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_866 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11116_ vdd rf_ram.memory\[449\]\[0\] clknet_leaf_113_clk vss _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05964__A1 vss _01903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09155__A1 vss _04401_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07705__A2 vss _03496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05407__I vss _01602_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08902__A1 vss _02916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06012__B vss _01552_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11047_ vdd rf_ram.memory\[144\]\[0\] clknet_leaf_337_clk vss _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput9 vss net9 i_dbus_rdt[16] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_308_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05192__A2 vss net134 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_434 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_71_clk vdd vss clknet_leaf_71_clk clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_157_754 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_467 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05470_ _01666_ _01643_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_15_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06692__A2 vss _02846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07140_ vdd _03150_ _03148_ _00183_ _03126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_125_651 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09630__A2 vss _01382_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07641__A1 vss _02889_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06444__A2 vss _01513_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07071_ vdd _03107_ _03105_ _00157_ _03092_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06022_ _01506_ vdd vss _02217_ rf_ram.memory\[550\]\[1\] _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_61_1066 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07973_ vdd vss _03669_ _03668_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09146__A1 vss net250 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09712_ vdd vss _04785_ _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06924_ vdd _03011_ _03010_ _00106_ _02970_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09697__A2 vss net33 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06855_ vdd vss _02965_ rf_ram.memory\[284\]\[0\] _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09643_ vdd _04730_ _04728_ _01106_ _04637_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_96_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05806_ _02001_ vdd vss _02002_ _01552_ _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09574_ _03967_ vdd vss _04688_ cpu.immdec.imm30_25\[5\] net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__05761__B vss _01956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08525_ vdd vss _04024_ net248 _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06380__A1 vss _01368_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06786_ vdd vss _02916_ _02773_ _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_148_721 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05737_ _01932_ vdd vss _01933_ _01909_ _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_62_clk vdd vss clknet_leaf_62_clk clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_93_803 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05668_ vss vdd rf_ram.memory\[479\]\[0\] _01778_ rf_ram.memory\[477\]\[0\] _01848_
+ _01863_ rf_ram.memory\[476\]\[0\] _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_93_858 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_92_302 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08456_ vdd vss net98 _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_175_595 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07407_ vdd vss _03317_ rf_ram.memory\[372\]\[0\] _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07880__A1 vss _03587_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08387_ vdd _03928_ _03927_ _00652_ _03919_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05599_ _01794_ vdd vss _01795_ _01675_ _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07338_ vdd vss _03274_ _02958_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05891__B1 vss _01925_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09621__A2 vss _04507_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07632__A1 vss _03455_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1112 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06435__A2 vss _02618_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07269_ vdd vss _03231_ _03230_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05238__A3 vss _01437_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10280_ vdd rf_ram.memory\[294\]\[0\] clknet_leaf_145_clk vss _00024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09008_ vdd vss _04326_ rf_ram.memory\[110\]\[0\] _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output171_I vss net171 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_991 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_687 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07935__A2 vss _02832_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09688__A2 vss net30 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07699__A1 vss _03491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05671__B vss _01707_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_53_clk vdd vss clknet_leaf_53_clk clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05390__C vss _01495_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_294_clk_I vss clknet_5_7__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1246 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11665_ net188 vss vdd net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_22_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10616_ vdd rf_ram.memory\[353\]\[0\] clknet_leaf_156_clk vss _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_554 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_571 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_251 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_960 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11596_ vdd rf_ram.memory\[9\]\[1\] clknet_leaf_38_clk vss _01328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07623__A1 vss _03425_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10547_ vdd rf_ram.memory\[333\]\[1\] clknet_leaf_167_clk vss _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06426__A2 vss _01989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06007__B vss _01552_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10478_ vdd rf_ram.memory\[421\]\[0\] clknet_leaf_104_clk vss _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05634__B1 vss _01688_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05846__B vss _01650_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08179__A2 vss _02960_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_232_clk_I vss clknet_5_23__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_247_clk_I vss clknet_5_21__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06640_ vdd vss _02809_ rf_ram.memory\[294\]\[1\] _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_95_1184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_44_clk vdd vss clknet_leaf_44_clk clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06571_ vdd _02754_ _02753_ _00010_ _02743_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05522_ _01712_ _01716_ vdd vss _01718_ _01708_ _01710_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06114__A1 vss _01527_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09290_ vdd _04509_ _04508_ _00974_ _04463_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09300__A1 vss _04463_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08310_ vdd _03879_ _03878_ _00624_ _03852_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08103__A2 vss _03729_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07862__A1 vss _03590_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05453_ _01649_ vss vdd _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08241_ vdd vss _03837_ _03668_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_925 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_576 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_705 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05384_ _01578_ _01579_ vdd vss _01580_ _01576_ _01577_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_28_796 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08172_ vdd _03794_ _03792_ _00571_ _03790_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07614__A1 vss _03445_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06417__A2 vss _01918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07123_ vdd _03140_ _03139_ _00176_ _03123_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_1106 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07054_ vdd _03096_ _03094_ _00151_ _03092_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_665 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput110 o_dbus_dat[20] net110 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput121 o_dbus_dat[30] net121 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput143 o_ext_rs1[14] net143 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06005_ _01505_ vdd vss _02200_ rf_ram.memory\[534\]\[1\] _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput132 o_dbus_sel[2] net132 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput176 o_ext_rs2[15] net176 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_56_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput154 o_ext_rs1[24] net154 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput165 o_ext_rs1[5] net165 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05475__C vss _01670_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput187 o_ext_rs2[25] net187 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput198 o_ext_rs2[6] net198 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05389__C1 vss _01555_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09119__A1 vss _04364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06050__B1 vss _01608_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07956_ vdd _03658_ _03656_ _00491_ _03654_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06907_ vdd vss _03000_ rf_ram.memory\[2\]\[1\] _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input28_I vss i_dbus_rdt[4] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07887_ vdd _03615_ _03613_ _00465_ _03590_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_928 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06838_ vdd _02952_ _02950_ _00079_ _02930_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_69_118 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09626_ vdd _04658_ _01452_ _01097_ _04643_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09557_ _03967_ vdd vss _04675_ cpu.immdec.imm30_25\[1\] net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06769_ vdd vss _02903_ _02716_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xclkbuf_leaf_35_clk vdd vss clknet_leaf_35_clk clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09488_ _04622_ vdd vss _04624_ net87 _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08508_ vdd vss _04012_ _01469_ net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_109_927 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08439_ vdd vss _03961_ _02953_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07853__A1 vss _02971_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05510__I vss _01686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_530 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11450_ vdd rf_ram.memory\[239\]\[1\] clknet_leaf_284_clk vss _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07605__A1 vss _03422_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11381_ _01113_ vdd vss clknet_leaf_229_clk net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10401_ vdd rf_ram.memory\[216\]\[1\] clknet_leaf_300_clk vss _00145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05616__B1 vss _01810_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10332_ vdd rf_ram.memory\[304\]\[0\] clknet_leaf_146_clk vss _00076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10263_ vdd _05127_ _05125_ _01330_ _02825_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08030__A1 vss _03668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10194_ vdd vss _05086_ _03892_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09652__I vss net1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06592__A1 vss _02743_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_337 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_26_clk vdd vss clknet_leaf_26_clk clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08097__A1 vss _03724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_324 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07844__A1 vss _03587_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput12 vss net12 i_dbus_rdt[19] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11648_ vss net201 net129 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_163_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput23 vss net23 i_dbus_rdt[29] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11579_ vdd rf_ram.memory\[207\]\[0\] clknet_leaf_34_clk vss _01311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput45 vss net45 i_ibus_rdt[20] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09597__A1 vss _03992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput34 net34 vss vdd i_ibus_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__07072__A2 vss _02911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput56 vss net56 i_ibus_rdt[30] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_171_clk_I vss clknet_5_30__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06280__B1 vss _01959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_51_clk_I vss clknet_5_12__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07810_ vdd _03568_ _03566_ _00435_ _03557_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08790_ vdd vss _04191_ rf_ram.memory\[149\]\[1\] _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07741_ vdd _03525_ _03522_ _00409_ _03524_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_186_clk_I vss clknet_5_28__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06583__A1 vss _02731_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05386__A2 vss _01532_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_66_clk_I vss clknet_5_8__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09521__A1 vss _03967_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07672_ vdd vss _03482_ _02904_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10131__A2 vss _02832_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_438 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08178__I vss _02845_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05138__A2 vss cpu.genblk3.csr.o_new_irq vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09411_ vdd vss _01024_ _04576_ _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06623_ _02795_ _02794_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_181_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_17_clk vdd vss clknet_leaf_17_clk clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09342_ _04540_ net224 vdd vss _04542_ net213 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08088__A1 vss _02971_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06554_ vdd vss _02740_ _01369_ rf_ram_if.wdata0_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05505_ vdd vss _01701_ rf_ram.memory\[340\]\[0\] _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07835__A1 vss _03557_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_124_clk_I vss clknet_5_13__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06485_ rf_ram.memory\[5\]\[1\] _01714_ _01643_ rf_ram.memory\[4\]\[1\] _02680_ vss
+ vdd rf_ram.memory\[7\]\[1\] _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_75_688 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_817 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_508 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09273_ _04481_ vdd vss _01387_ _04497_ _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_05436_ vdd vss _01632_ rf_ram.memory\[366\]\[0\] _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_267 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05330__I vss _01525_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_722 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_454 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08224_ vdd vss _03827_ rf_ram.memory\[533\]\[1\] _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05367_ _01563_ vss vdd _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09588__A1 vss _02709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08155_ vdd _03783_ _03781_ _00565_ _03757_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07106_ vdd _03129_ _03128_ _00170_ _03123_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_714 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_139_clk_I vss clknet_5_27__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08086_ vdd vss _03741_ rf_ram.memory\[55\]\[1\] _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08260__A1 vss _03823_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05298_ _01494_ _01493_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_19_clk_I vss clknet_5_2__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07037_ vdd vss _03085_ rf_ram.memory\[215\]\[0\] _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08012__A1 vss _03686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08563__A2 vss _02960_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06023__B1 vss _01539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1000 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08988_ vdd vss _04314_ rf_ram.memory\[114\]\[0\] _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05377__A2 vss _01524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07939_ vdd _03647_ _03645_ _00485_ _03622_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_39_1130 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output134_I vss net134 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10950_ vdd rf_ram.memory\[79\]\[0\] clknet_leaf_18_clk vss _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09609_ vdd vss _04715_ rf_ram.memory\[73\]\[0\] _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10881_ vdd rf_ram.memory\[243\]\[1\] clknet_leaf_282_clk vss _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_1196 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_931 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_724 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_633 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07826__A1 vss _02839_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11502_ vdd rf_ram.memory\[348\]\[1\] clknet_leaf_191_clk vss _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1014 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_1183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_151_524 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1015 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_204 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11433_ vdd cpu.state.cnt_r\[0\] clknet_leaf_238_clk vss _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09579__A1 vss _01391_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10189__A2 vss _02972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_585 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11364_ vdd rf_ram.memory\[71\]\[1\] clknet_leaf_63_clk vss _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_1183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_1014 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_909 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08251__A1 vss _02845_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_966 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11295_ _01028_ vdd vss clknet_leaf_250_clk net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10315_ vdd rf_ram.memory\[513\]\[1\] clknet_leaf_267_clk vss _00059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05396__B vss _01351_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10246_ vdd _05117_ _05116_ _01323_ _02819_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08003__A1 vss _03686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10177_ vdd vss _05075_ _03892_ _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05773__C1 vss _01968_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09503__A1 vss _04634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05540__A2 vss _01735_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_975 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08490__A1 vss _03953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05828__B1 vss _02019_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06270_ _02464_ vdd vss _02465_ _01951_ _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_170_833 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05221_ vdd vss _01421_ _01416_ _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_170_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_894 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05152_ _01344_ vdd vss _01355_ cpu.immdec.imm24_20\[1\] _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09960_ vdd vss _04942_ rf_ram.memory\[335\]\[0\] _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09990__A1 vss _04953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_6_clk vdd vss clknet_leaf_6_clk clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08911_ vdd _04265_ _04263_ _00839_ _04237_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_95 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09891_ vdd vss _04899_ _02922_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08842_ vdd _04223_ _04222_ _00812_ _04202_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_1005 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05985_ rf_ram.memory\[3\]\[0\] _01635_ _01661_ rf_ram.memory\[2\]\[0\] _02181_ vss
+ vdd rf_ram.memory\[1\]\[0\] _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08773_ vdd vss _04181_ rf_ram.memory\[143\]\[0\] _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07724_ vdd _03514_ _03512_ _00403_ _03491_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_1098 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07655_ vdd _03471_ _03469_ _00377_ _03458_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06859__A2 vss _02941_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05325__I vss _01520_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06606_ vdd vss _02782_ _02766_ _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07586_ vdd vss _03429_ rf_ram.memory\[316\]\[1\] _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05531__A2 vss _01724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07808__A1 vss _03554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09325_ vdd _04531_ _04530_ _00987_ _04463_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06537_ vdd vss _02723_ _02720_ _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_0_118_543 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06468_ vdd vss _02663_ rf_ram.memory\[17\]\[1\] _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09256_ vdd vss _01356_ _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_146_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_80 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_749 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05419_ _01615_ vss vdd _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08207_ vdd vss _03816_ rf_ram.memory\[536\]\[1\] _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06399_ _01684_ vdd vss _02594_ rf_ram.memory\[88\]\[1\] _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09187_ vdd vss _04438_ rf_ram.memory\[179\]\[1\] _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08138_ vdd _03773_ _03772_ _00558_ _03754_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07036__A2 vss _03083_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08233__A1 vss _03820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10040__A1 vss _04982_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09981__A1 vss _02865_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08069_ vdd vss _03731_ rf_ram.memory\[562\]\[0\] _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10100_ vdd vss _05028_ _02800_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05598__A2 vss _01777_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11080_ vdd rf_ram.memory\[132\]\[1\] clknet_leaf_15_clk vss _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10031_ vdd vss _04986_ rf_ram.memory\[327\]\[1\] _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09733__A1 vss _04781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1091 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08536__A2 vss _03945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05944__B vss _01493_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_26__f_clk vdd vss clknet_5_26__leaf_clk clknet_3_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05507__C1 vss _01702_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_408 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10933_ vdd rf_ram_if.wdata1_r\[0\] clknet_leaf_261_clk vss rf_ram_if.wdata1_r\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10864_ vdd rf_ram.memory\[197\]\[0\] clknet_leaf_42_clk vss _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_1096 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_975 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10795_ vdd rf_ram.memory\[55\]\[1\] clknet_leaf_298_clk vss _00539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07275__A2 vss _03234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_660 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_433 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08472__A1 vss _01369_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_811 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_855 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11416_ vdd rf_ram.memory\[80\]\[1\] clknet_leaf_48_clk vss _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_717 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_555 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11347_ vdd cpu.immdec.imm30_25\[3\] clknet_leaf_264_clk vss _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06015__B vss _01351_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06786__A1 vss _02773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09724__A1 vss _04781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11278_ vdd net214 clknet_leaf_243_clk vss _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10229_ vdd vss _05107_ _02765_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06538__A1 vss rf_ram.i_raddr\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1137 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05854__B vss _01956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05746__C1 vss _01646_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_14__f_clk_I vss clknet_3_3_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xhold1 vdd rf_ram_if.wdata1_r\[2\] vss net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_179_719 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05770_ _01494_ vdd vss _01966_ _01963_ _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_706 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1060 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05761__A2 vss _01735_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_920 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_1071 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07440_ vdd vss _03338_ rf_ram.memory\[36\]\[0\] _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_69_290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08456__I vss net98 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_446 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07371_ vdd vss _03295_ rf_ram.memory\[267\]\[0\] _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_468 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09110_ vdd vss _04389_ rf_ram.memory\[94\]\[1\] _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06322_ _02516_ vdd vss _02517_ _01600_ _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_57_496 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09041_ vdd vss _04347_ rf_ram.memory\[104\]\[0\] _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06253_ _01805_ vdd vss _02448_ rf_ram.memory\[430\]\[1\] _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09287__I vss _04004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11610__I vss net90 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06184_ _02378_ vdd vss _02379_ _01769_ _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_115_579 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05204_ _01341_ vdd vss _01404_ cpu.state.init_done _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__08215__A1 vss _03798_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_696 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06226__B1 vss _01702_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09963__A1 vss _04921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05135_ vdd vss _01338_ _01334_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_09943_ vdd _04931_ _04929_ _01206_ _04921_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_1138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05985__C1 vss _01714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06529__A1 vss _02714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09874_ vdd _04471_ _01418_ _04889_ cpu.state.init_done vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08825_ vdd vss _04213_ _02828_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_1183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_80 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input10_I vss i_dbus_rdt[17] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10089__A1 vss _05017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05968_ _01493_ vdd vss _02164_ _02161_ _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08756_ vss _04170_ _04061_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_07707_ vdd _03504_ _03503_ _00396_ _03488_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05899_ _01746_ vdd vss _02095_ _02093_ _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08687_ _04126_ _04057_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_178_763 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_402 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07638_ vdd _03461_ _03460_ _00370_ _03455_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06701__A1 vss _02826_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07569_ vdd vss _03418_ rf_ram.memory\[357\]\[1\] _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_181_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_411 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09308_ vdd vss cpu.immdec.imm11_7\[1\] _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10580_ vdd rf_ram.memory\[362\]\[0\] clknet_leaf_162_clk vss _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07257__A2 vss _03040_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_800 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09239_ vdd vss _04470_ rf_ram.memory\[319\]\[1\] _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_170 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06465__B1 vss _01624_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10261__A1 vss _02819_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06614__I vss _02787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08206__A1 vss _03787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1240 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09954__A1 vss _04911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10013__A1 vss _04950_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11201_ vdd rf_ram.memory\[86\]\[1\] clknet_leaf_45_clk vss _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11132_ vdd rf_ram.memory\[114\]\[0\] clknet_leaf_74_clk vss _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06768__A1 vss _02876_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11063_ vdd rf_ram.memory\[138\]\[0\] clknet_leaf_11_clk vss _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09557__I1 vss net50 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10014_ vdd vss _04975_ rf_ram.memory\[348\]\[1\] _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07193__A1 vss _03161_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_153_1114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06940__A1 vss _03018_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10916_ vdd rf_ram.memory\[178\]\[0\] clknet_leaf_16_clk vss _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08693__A1 vss _04129_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_958 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_750 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10847_ vdd rf_ram.memory\[533\]\[1\] clknet_leaf_310_clk vss _00591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10778_ vdd rf_ram.memory\[567\]\[0\] clknet_leaf_329_clk vss _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_164_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05849__B vss _01350_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_466 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06759__A1 vss _02873_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06940_ vdd _03022_ _03020_ _00111_ _03018_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_181_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06871_ vdd vss _02976_ rf_ram.memory\[302\]\[1\] _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05982__A2 vss _01640_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I vss i_dbus_rdt[0] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07184__A1 vss _02738_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_230_clk vdd vss clknet_leaf_230_clk clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08610_ vdd vss _04079_ net238 _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05822_ vdd vss _02018_ rf_ram.memory\[212\]\[0\] _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05734__A2 vss _01531_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06931__A1 vss _03014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09590_ _04701_ vdd vss _04702_ _04697_ cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05753_ _01948_ vdd vss _01949_ _01372_ _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_89_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08541_ vdd vss _04034_ net246 _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05684_ vdd vss _01880_ rf_ram.memory\[398\]\[0\] _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_89_396 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08472_ rf_ram.rdata\[1\] vdd vss _03987_ _01369_ _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__08684__A1 vss _04094_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07423_ vdd _03327_ _03324_ _00289_ _03326_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_273 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_94 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05603__I vss _01613_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07354_ vdd vss _03284_ rf_ram.memory\[252\]\[0\] _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08436__A1 vss _03953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08987__A2 vss _04303_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07285_ vdd vss _03241_ _02836_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_797 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_297_clk vdd vss clknet_leaf_297_clk clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06305_ vdd vss _02500_ rf_ram.memory\[169\]\[1\] _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10243__A1 vss _02825_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06236_ _02425_ _01660_ _02430_ vdd vss _02431_ _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_09024_ vdd vss _04336_ net246 _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_86_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09936__A1 vss _04918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05670__A1 vss _01850_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08739__A2 vss _04158_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06167_ _02361_ vdd vss _02362_ _01603_ _02360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_130_379 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06098_ vss vdd rf_ram.memory\[277\]\[1\] _01678_ rf_ram.memory\[279\]\[1\] _01679_
+ _01687_ rf_ram.memory\[278\]\[1\] _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA_input58_I vss i_ibus_rdt[3] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05958__C1 vss _01655_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09926_ _04921_ _04400_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05973__A2 vss _01530_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1109 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_221_clk vdd vss clknet_leaf_221_clk clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_77_1222 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09857_ _02690_ _01391_ vdd vss _04878_ _01382_ _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__06922__A1 vss _02958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09788_ vdd vss _04836_ rf_ram.memory\[76\]\[1\] _04834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08808_ _04202_ _04057_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08739_ vdd vss _04159_ _01497_ _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07478__A2 vss _02815_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10701_ vdd rf_ram.memory\[432\]\[1\] clknet_leaf_81_clk vss _00445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_435 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05513__I vss _01508_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_254 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_265 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_939 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_405 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10632_ vdd rf_ram.memory\[386\]\[0\] clknet_leaf_93_clk vss _00376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_118 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09475__I0 vss net88 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_170 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10563_ vdd rf_ram.memory\[32\]\[1\] clknet_leaf_203_clk vss _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_288_clk vdd vss clknet_leaf_288_clk clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10234__A1 vss _02737_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_972 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_162 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10494_ vdd rf_ram.memory\[471\]\[0\] clknet_leaf_54_clk vss _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_672 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_182 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11115_ vdd rf_ram.memory\[122\]\[1\] clknet_leaf_86_clk vss _00851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11046_ vdd rf_ram.memory\[145\]\[1\] clknet_leaf_336_clk vss _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07166__A1 vss _03157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_212_clk vdd vss clknet_leaf_212_clk clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08902__A2 vss _04038_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06913__A1 vss _02975_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06374__C1 vss _01625_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06126__C1 vss _01773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08666__A1 vss _04097_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06141__A2 vss _01709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08418__A1 vss _03919_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_279_clk vdd vss clknet_leaf_279_clk clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09091__A1 vss _04367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07070_ vdd vss _03107_ rf_ram.memory\[494\]\[1\] _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07641__A2 vss _03089_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1182 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06021_ _02214_ _02215_ vdd vss _02216_ _02212_ _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_140_655 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07972_ vss _03668_ _02868_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__09146__A2 vss _03035_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09711_ _04768_ _04784_ vdd vss _04785_ net102 _04767_ net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__05955__A2 vss _01661_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1089 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06923_ vdd vss _03011_ rf_ram.memory\[278\]\[0\] _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06854_ vdd vss _02964_ _02839_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_203_clk vdd vss clknet_leaf_203_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09642_ vdd vss _04730_ rf_ram.memory\[78\]\[1\] _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06904__A1 vss _02894_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06365__C1 vss _01968_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_1022 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06785_ vss _02915_ _02910_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_78_823 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05805_ rf_ram.memory\[173\]\[0\] _01516_ _01692_ rf_ram.memory\[172\]\[0\] _02001_
+ vss vdd rf_ram.memory\[175\]\[0\] _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_09573_ vss _01079_ _04687_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05736_ vss vdd rf_ram.memory\[447\]\[0\] _01857_ rf_ram.memory\[445\]\[0\] _01931_
+ _01799_ rf_ram.memory\[444\]\[0\] _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__06380__A2 vss _02547_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08524_ _04023_ vss vdd _03685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__05183__A3 vss _01382_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08657__A1 vss _02953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_901 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_1114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06132__A2 vss _01782_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05667_ _01863_ _01633_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08455_ _01401_ vdd vss _03972_ _01408_ _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07406_ vdd vss _03316_ _03100_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05598_ vss vdd rf_ram.memory\[293\]\[0\] _01793_ rf_ram.memory\[295\]\[0\] _01778_
+ _01777_ rf_ram.memory\[294\]\[0\] _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_136_939 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08409__A1 vss _03922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08386_ vdd vss _03928_ rf_ram.memory\[189\]\[0\] _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_433 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09457__I0 vss net78 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05489__B vss _01684_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09082__A1 vss net239 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10216__A1 vss _05078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07337_ vdd _03273_ _03271_ _00257_ _03260_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_723 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07268_ vss _03230_ _02737_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_14_650 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06219_ _01786_ rf_ram.memory\[387\]\[1\] vdd vss _02414_ rf_ram.memory\[386\]\[1\]
+ _01785_ _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07199_ vdd vss _03187_ _02761_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09007_ vdd vss _04325_ _02971_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06199__A2 vss _01706_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07396__A1 vss _03309_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05946__A2 vss _01661_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09909_ vdd vss _04910_ rf_ram.memory\[292\]\[1\] _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07148__A1 vss _03123_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08896__A1 vss _04237_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05952__B vss _01601_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05254__S0 vss _01376_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06371__A2 vss _01606_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07320__A1 vss _03257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11664_ net187 vss vdd net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09448__I0 vss net74 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1034 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10615_ vdd rf_ram.memory\[314\]\[1\] clknet_leaf_105_clk vss _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_1080 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1035 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09073__A1 vss _04364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11595_ vdd rf_ram.memory\[9\]\[0\] clknet_leaf_38_clk vss _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10546_ vdd rf_ram.memory\[333\]\[0\] clknet_leaf_142_clk vss _00290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08820__A1 vss net250 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10477_ vdd rf_ram.memory\[422\]\[1\] clknet_leaf_101_clk vss _00221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_195 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07387__A1 vss _03289_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05937__A2 vss _01682_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05418__I vss _01613_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08887__A1 vss _03672_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06347__C1 vss _01713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1130 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08729__I vss _04077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11029_ vdd rf_ram.memory\[150\]\[1\] clknet_leaf_2_clk vss _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07633__I vss _03359_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177_828 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06362__A2 vss _01958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06570_ vdd vss _02754_ rf_ram.memory\[201\]\[0\] _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_333 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_176_349 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05521_ _01717_ _01493_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_47_539 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05452_ _01647_ vdd vss _01648_ _01527_ _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08240_ vdd _03836_ _03834_ _00597_ _03823_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_117_427 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_818 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08171_ vdd vss _03794_ rf_ram.memory\[543\]\[1\] _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09064__A1 vss _04334_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07122_ vdd vss _03140_ rf_ram.memory\[487\]\[0\] _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_414 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05383_ rf_ram.memory\[547\]\[0\] _01521_ _01544_ rf_ram.memory\[546\]\[0\] _01579_
+ vss vdd rf_ram.memory\[545\]\[0\] _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__07614__A2 vss _02984_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08811__A1 vss _04202_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07053_ vdd vss _03096_ rf_ram.memory\[390\]\[1\] _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_88_53 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput100 o_dbus_dat[11] net100 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_70_586 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_986 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_828 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput111 o_dbus_dat[21] net111 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput122 o_dbus_dat[31] net122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06004_ _02198_ vdd vss _02199_ _01495_ _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput133 o_dbus_sel[3] net133 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput177 o_ext_rs2[16] net177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput155 o_ext_rs1[25] net155 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput166 o_ext_rs1[6] net166 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput144 o_ext_rs1[15] net144 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput188 o_ext_rs2[26] net188 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput199 o_ext_rs2[7] net199 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05928__A2 vss _01863_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_7__f_clk vdd vss clknet_5_7__leaf_clk clknet_3_1_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05389__B1 vss _01554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05328__I vss _01523_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07955_ vdd vss _03658_ rf_ram.memory\[481\]\[1\] _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11002__CLK vss clknet_5_0__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06906_ vdd _02999_ _02998_ _00100_ _02970_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08639__I vss _04061_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07886_ vdd vss _03615_ rf_ram.memory\[462\]\[1\] _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09625_ vdd _04722_ _04720_ _01096_ _04637_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06837_ vdd vss _02952_ rf_ram.memory\[286\]\[1\] _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07550__A1 vss _03393_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06353__A2 vss _01501_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06768_ vdd _02902_ _02900_ _00059_ _02876_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09556_ _04523_ vdd vss _01075_ _04673_ _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05719_ _01915_ _01536_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06105__A2 vss _01626_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07302__A1 vss _03222_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06699_ vdd _02854_ _02853_ _00038_ _02820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09487_ vdd _04623_ _04622_ _01057_ _02690_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08507_ cpu.immdec.imm11_7\[4\] vdd vss _04011_ cpu.immdec.imm11_7\[0\] cpu.immdec.imm11_7\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_175_360 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_859 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08438_ vdd _03960_ _03958_ _00671_ _03956_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07853__A2 vss _03234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_701 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05864__A1 vss _01951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_268 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09055__A1 vss _02794_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08369_ vdd vss _03917_ rf_ram.memory\[185\]\[0\] _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10400_ vdd rf_ram.memory\[216\]\[0\] clknet_leaf_300_clk vss _00144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08802__A1 vss _04170_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11380_ _01112_ vdd vss clknet_leaf_232_clk cpu.bufreg2.o_sh_done_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_33_255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xwire249 net249 vss vdd _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__05616__A1 vss rf_ram.memory\[312\]\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10331_ vdd rf_ram.memory\[287\]\[1\] clknet_leaf_174_clk vss _00075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output89_I vss net89 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_307_clk_I vss clknet_5_4__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10262_ vdd vss _05127_ rf_ram.memory\[574\]\[1\] _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_108_1096 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07369__A1 vss _03292_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05919__A2 vss _01799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08030__A2 vss _02992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10193_ vdd _05085_ _05083_ _01302_ _05081_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08869__A1 vss _04234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07541__A1 vss _03319_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06344__A2 vss _01662_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_541 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_1022 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_339 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11647_ vss net200 net128 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_892 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput13 vss net13 i_dbus_rdt[1] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11578_ vdd rf_ram.memory\[442\]\[1\] clknet_leaf_56_clk vss _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_983 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput24 vss net24 i_dbus_rdt[2] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09597__A2 vss net47 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput46 vss net46 i_ibus_rdt[21] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput35 vss net35 i_ibus_rdt[10] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10529_ vdd rf_ram.memory\[250\]\[1\] clknet_leaf_217_clk vss _00273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_417 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05857__B vss _01564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput57 vss net57 i_ibus_rdt[31] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_299 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05148__I vss _01350_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07740_ vdd vss _03525_ rf_ram.memory\[378\]\[1\] _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07780__A1 vss _03521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_22 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06583__A2 vss _02764_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07363__I vss _03013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07671_ vss _03481_ _03088_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09410_ vdd _04539_ _04579_ _04580_ _04578_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06622_ vdd vss _02794_ _02750_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_06553_ vdd vss _02739_ _02728_ _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09341_ vdd vss _04541_ _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08088__A2 vss _03729_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_861 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05504_ _01620_ vdd vss _01700_ _01694_ _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06099__A1 vss _01675_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06484_ _01503_ vdd vss _02679_ rf_ram.memory\[6\]\[1\] _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_7_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09272_ vdd vss _04496_ _01365_ _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09037__A1 vss _04331_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05435_ _01631_ vss vdd _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_62_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08223_ vdd _03826_ _03825_ _00590_ _03820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_173_897 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05366_ vdd _01562_ rf_ram.i_raddr\[3\] vss vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_08154_ vdd vss _03783_ rf_ram.memory\[546\]\[1\] _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_85 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07105_ vdd vss _03129_ rf_ram.memory\[501\]\[0\] _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_70_350 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08085_ vdd _03740_ _03739_ _00538_ _03721_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05767__B vss _01956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07036_ vdd vss _03084_ _02738_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05297_ _01493_ vss vdd rf_ram.i_raddr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_140_271 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_485 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_1149 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_91 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_293_clk_I vss clknet_5_7__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input40_I vss i_ibus_rdt[15] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07771__A1 vss _03524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08987_ vdd vss _04313_ net236 _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07938_ vdd vss _03647_ rf_ram.memory\[457\]\[1\] _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07869_ vdd vss _03605_ rf_ram.memory\[408\]\[0\] _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_1078 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06326__A2 vss _01804_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09608_ vdd vss _04714_ net249 _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10880_ vdd rf_ram.memory\[243\]\[0\] clknet_leaf_282_clk vss _00624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1207 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_601 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09539_ _04662_ _04663_ vdd vss _01069_ _04648_ _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_clkbuf_leaf_231_clk_I vss clknet_5_23__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09276__A1 vss _01364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07826__A2 vss _03559_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05521__I vss _01493_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_829 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_509 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11501_ vdd rf_ram.memory\[348\]\[0\] clknet_leaf_177_clk vss _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09028__A1 vss _04334_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11432_ vdd rf_ram.memory\[61\]\[1\] clknet_leaf_293_clk vss _01164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1048 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_246_clk_I vss clknet_5_21__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_704 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11363_ vdd rf_ram.memory\[71\]\[0\] clknet_leaf_64_clk vss _01095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08251__A2 vss _02954_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_496 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10314_ vdd rf_ram.memory\[513\]\[0\] clknet_leaf_268_clk vss _00058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11294_ _01027_ vdd vss clknet_leaf_250_clk net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10245_ vdd vss _05117_ rf_ram.memory\[264\]\[0\] _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10176_ vdd _05074_ _05072_ _01296_ _05049_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07762__A1 vss _02775_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06565__A2 vss _02748_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05773__B1 vss _01953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1133 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06317__A2 vss _01631_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_159_636 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_159_658 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_69 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_308 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_792 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06527__I vss _02713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_683 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_823 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_514 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_553 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05220_ _01419_ vdd vss _01420_ cpu.immdec.imm31 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_163_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05151_ vss _01354_ cpu.immdec.imm19_12_20\[5\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_150_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05461__C1 vss _01656_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08910_ vdd vss _04265_ rf_ram.memory\[125\]\[1\] _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09890_ vdd _04898_ _04896_ _01186_ _04887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08841_ vdd vss _04223_ rf_ram.memory\[134\]\[0\] _04222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1044 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05984_ _01525_ vdd vss _02180_ rf_ram.memory\[0\]\[0\] _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08772_ vdd vss _04180_ _02953_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07505__A1 vss _03356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07723_ vdd vss _03514_ rf_ram.memory\[398\]\[1\] _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06308__A2 vss _01501_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07654_ vdd vss _03471_ rf_ram.memory\[386\]\[1\] _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06605_ _02781_ _02780_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_07585_ vdd _03428_ _03427_ _00350_ _03422_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05341__I vss _01536_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09324_ vdd vss _04531_ rf_ram.memory\[109\]\[0\] _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_731 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06536_ _01341_ vdd vss _02722_ _01352_ _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_111_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05819__A1 vss _01600_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06467_ _01601_ vdd vss _02662_ rf_ram.memory\[16\]\[1\] _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09255_ _04482_ _01341_ vdd vss _04483_ cpu.genblk3.csr.mstatus_mpie _01356_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_172_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_385 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_92 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05418_ _01614_ _01613_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06492__A1 vss _02603_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_531 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08206_ vdd _03815_ _03814_ _00584_ _03787_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06398_ _02592_ vdd vss _02593_ _01769_ _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09186_ vdd _04437_ _04436_ _00942_ _04431_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_16_553 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07268__I vss _02737_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08137_ vdd vss _03773_ rf_ram.memory\[54\]\[0\] _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05349_ rf_ram.memory\[514\]\[0\] _01545_ vss vdd rf_ram.memory\[513\]\[0\] _01539_
+ rf_ram.memory\[515\]\[0\] _01540_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__09981__A2 vss _02958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_794 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08068_ vdd vss _03730_ net236 _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07019_ vdd vss _03073_ _03055_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10030_ _04985_ _04400_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_175_1009 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07744__A1 vss _03521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09733__A2 vss net14 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05960__B vss _01599_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10932_ vdd rf_ram_if.rreq_r clknet_leaf_254_clk vss _00676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05507__B1 vss _01688_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_170_clk_I vss clknet_5_31__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10863_ vdd rf_ram.memory\[205\]\[1\] clknet_leaf_31_clk vss _00607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_820 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_50_clk_I vss clknet_5_12__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1195 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10794_ vdd rf_ram.memory\[55\]\[0\] clknet_leaf_297_clk vss _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_1161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_261 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_185_clk_I vss clknet_5_28__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_350 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11415_ vdd rf_ram.memory\[80\]\[0\] clknet_leaf_48_clk vss _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_65_clk_I vss clknet_5_8__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_681 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_929 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11346_ vdd cpu.immdec.imm30_25\[2\] clknet_leaf_260_clk vss _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07983__A1 vss _03654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11277_ vdd net212 clknet_leaf_245_clk vss _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08511__B vss _01366_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09724__A2 vss net10 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10228_ vdd _05106_ _05104_ _01316_ _05081_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05746__B1 vss _01810_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_123_clk_I vss clknet_5_13__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10159_ vdd _05064_ _05063_ _01289_ _05046_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xhold2 vdd rf_ram_if.wdata0_r\[1\] vss net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__05210__A2 vss _01409_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09488__A1 vss net87 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_138_clk_I vss clknet_5_25__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_217 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08160__A1 vss _03757_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_959 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07370_ vdd vss _03294_ _02781_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_18_clk_I vss clknet_5_2__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05161__I vss cpu.state.genblk1.misalign_trap_sync_r vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06321_ _02514_ _02515_ vdd vss _02516_ _02512_ _02513_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_06252_ _02439_ _02443_ _02446_ vdd vss _02447_ _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_0_127_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09040_ vdd vss _04346_ net250 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09660__A1 vss net1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_694 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_193 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_3_5_0_clk_I vss clknet_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05203_ cpu.state.init_done _01402_ vdd vss _01403_ _01342_ cpu.bufreg2.o_sh_done_r
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_06183_ vss vdd rf_ram.memory\[469\]\[1\] _01848_ rf_ram.memory\[471\]\[1\] _01786_
+ _01785_ rf_ram.memory\[470\]\[1\] _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__09412__A1 vss net246 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08215__A2 vss _03009_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_84 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05134_ vdd vss _01337_ _01335_ _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_187_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09942_ vdd vss _04931_ rf_ram.memory\[33\]\[1\] _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_111_764 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1076 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05985__B1 vss _01635_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09873_ _03989_ vdd vss _01179_ _02713_ _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08824_ vdd _04212_ _04210_ _00805_ _04205_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05336__I vss _01531_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08755_ vdd _04169_ _04168_ _00779_ _04167_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07706_ vdd vss _03504_ rf_ram.memory\[381\]\[0\] _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05780__B vss _01923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05967_ _01624_ rf_ram.memory\[19\]\[0\] vdd vss _02163_ rf_ram.memory\[18\]\[0\]
+ _01605_ _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09479__A1 vss cpu.bufreg.i_sh_signed vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05898_ rf_ram.memory\[91\]\[0\] _01646_ _01801_ rf_ram.memory\[90\]\[0\] _02094_
+ vss vdd rf_ram.memory\[89\]\[0\] _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__08151__A1 vss _02893_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08686_ vdd _04125_ _04123_ _00754_ _04097_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07637_ vdd vss _03461_ rf_ram.memory\[406\]\[0\] _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07568_ vdd _03417_ _03416_ _00344_ _03389_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_70 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_146_650 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09307_ vdd _04519_ _04517_ _00981_ _04466_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06519_ vdd vss _02707_ _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07499_ vdd vss _03375_ rf_ram.memory\[324\]\[0\] _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09651__A1 vss net98 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09238_ vdd _04469_ _04468_ _00962_ _04463_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output194_I vss net194 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09169_ vdd _04426_ _04425_ _00936_ _04397_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_181_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_1008 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09954__A2 vss _02946_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11200_ vdd rf_ram.memory\[86\]\[0\] clknet_leaf_45_clk vss _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11131_ vdd rf_ram.memory\[115\]\[1\] clknet_leaf_74_clk vss _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_max_cap240_I vss _02888_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05955__B vss _01503_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output71_I vss net71 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07717__A1 vss _03488_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11062_ vdd rf_ram.memory\[13\]\[1\] clknet_leaf_31_clk vss _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10013_ vdd _04974_ _04973_ _01233_ _04950_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08390__A1 vss _03892_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_6__f_clk_I vss clknet_3_1_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05690__B vss _01746_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_764 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10915_ vdd rf_ram.memory\[209\]\[1\] clknet_leaf_29_clk vss _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09890__A1 vss _04887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10846_ vdd rf_ram.memory\[533\]\[0\] clknet_leaf_299_clk vss _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_823 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05259__A2 vss _01382_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10777_ vdd rf_ram.memory\[568\]\[1\] clknet_leaf_307_clk vss _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_642 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_694 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06805__I vss _02825_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_355 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_1076 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_697 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06208__A1 vss _01674_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_377 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07956__A1 vss _03654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11329_ vdd rf_ram.memory\[289\]\[1\] clknet_leaf_123_clk vss _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05967__B1 vss _01624_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05431__A2 vss _01626_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06870_ _02975_ _02825_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_174_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07184__A2 vss _02806_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05821_ _02016_ vdd vss _02017_ net251 _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_05752_ _01947_ vdd vss _01948_ net252 _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_08540_ vdd _04033_ _04031_ _00700_ _04026_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08133__A1 vss _03754_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05683_ _01878_ vdd vss _01879_ _01368_ _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_89_386 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08471_ vdd vss _00678_ _02714_ _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07422_ vdd vss _03327_ rf_ram.memory\[371\]\[1\] _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05498__A2 vss _01692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09881__A1 vss _03309_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_272 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07353_ vdd vss _03283_ _03055_ _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09633__A1 vss _04524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11621__I vss net71 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1019 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07284_ vdd _03240_ _03238_ _00237_ _03225_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06304_ _01956_ vdd vss _02499_ rf_ram.memory\[168\]\[1\] _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_170_450 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06235_ _02427_ _02428_ _02429_ _01670_ vdd vss _02430_ _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_09023_ vdd _04335_ _04332_ _00881_ _04334_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_388 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06166_ rf_ram.memory\[486\]\[1\] _02361_ vss vdd rf_ram.memory\[485\]\[1\] _01702_
+ rf_ram.memory\[487\]\[1\] _01688_ _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_40_150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1041 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06097_ vdd vss _02292_ rf_ram.memory\[276\]\[1\] _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05958__B1 vss _01653_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05422__A2 vss _01617_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09925_ vdd _04920_ _04919_ _01199_ _04918_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_102_1025 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09856_ vdd vss _04877_ cpu.state.genblk1.misalign_trap_sync_r _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08372__A1 vss _03887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08807_ vdd _04201_ _04199_ _00799_ _04170_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06922__A2 vss _03009_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09787_ vdd _04835_ _04834_ _01145_ _04634_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05186__A1 vss cpu.mem_bytecnt\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06999_ vdd _03060_ _03059_ _00132_ _03050_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08124__A1 vss _03757_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08738_ vdd vss _04158_ _01369_ _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08669_ vdd _04115_ _04114_ _00747_ _04094_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09321__C2 vss cpu.immdec.imm11_7\[4\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10700_ vdd rf_ram.memory\[432\]\[0\] clknet_leaf_81_clk vss _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05489__A2 vss _01683_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09872__A1 vss _04887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06150__A3 vss _02344_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10631_ vdd rf_ram.memory\[405\]\[1\] clknet_leaf_115_clk vss _00375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_650 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09475__I1 vss net89 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06438__A1 vss _01903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10562_ vdd rf_ram.memory\[32\]\[0\] clknet_leaf_205_clk vss _00306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10234__A2 vss _02946_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_404 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_193 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05646__C1 vss _01668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10493_ vdd rf_ram.memory\[472\]\[1\] clknet_leaf_126_clk vss _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09388__B1 vss _04564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_336 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11114_ vdd rf_ram.memory\[122\]\[0\] clknet_leaf_86_clk vss _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06610__A1 vss _02748_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11045_ vdd rf_ram.memory\[145\]\[0\] clknet_leaf_336_clk vss _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08363__A1 vss _02991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06374__B1 vss _01678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06126__B1 vss _01848_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08115__A1 vss _02751_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_86_334 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09863__A1 vss _04837_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09615__A1 vss _04634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10829_ vdd rf_ram.memory\[542\]\[1\] clknet_leaf_274_clk vss _00573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_992 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_776 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06020_ rf_ram.memory\[555\]\[1\] _01521_ _01532_ rf_ram.memory\[554\]\[1\] _02215_
+ vss vdd rf_ram.memory\[553\]\[1\] _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_23_640 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07929__A1 vss _03622_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1111 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05595__B vss _01790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07971_ vdd _03667_ _03665_ _00497_ _03654_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06922_ vdd vss _03010_ _02958_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09710_ vdd vss _04784_ _04781_ net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06853_ vdd _02963_ _02961_ _00083_ _02930_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10161__A1 vss _05049_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09641_ vdd _04729_ _04728_ _01105_ _04634_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05168__A1 vss _01369_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06365__B1 vss _01959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06904__A2 vss _02997_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06784_ vdd _02914_ _02912_ _00063_ _02876_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05804_ vdd vss _02000_ rf_ram.memory\[174\]\[0\] _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09572_ _04678_ vdd vss _04687_ cpu.immdec.imm30_25\[3\] _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05735_ _01931_ _01626_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05614__I vss _01714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08523_ vdd _04022_ _04020_ _00694_ _03956_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_1251 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_701 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_868 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_356 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08657__A2 vss _03945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09854__A1 vss _01385_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_542 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05666_ vdd vss _01862_ rf_ram.memory\[478\]\[0\] _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_1305 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_827 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08454_ vdd net126 _03970_ _03971_ _01401_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_406 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05597_ _01793_ _01617_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_07405_ vdd _03315_ _03313_ _00283_ _03292_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08385_ vdd vss _03927_ _02959_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09457__I1 vss net79 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05891__A2 vss _01719_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07336_ vdd vss _03273_ rf_ram.memory\[254\]\[1\] _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09082__A2 vss _04339_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_623 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09006_ vdd _04324_ _04322_ _00875_ _04301_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_116_697 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07267_ vdd _03229_ _03227_ _00231_ _03225_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_640 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06218_ vdd vss _02413_ rf_ram.memory\[385\]\[1\] _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_147_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07198_ vdd _03186_ _03184_ _00205_ _03161_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_336 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05643__A2 vss _01662_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1211 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06149_ _02341_ _02342_ _02343_ _01658_ vdd vss _02344_ _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_130_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06053__C1 vss _01636_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07396__A2 vss _02992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08593__A1 vss _02805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09908_ vdd _04909_ _04908_ _01193_ _04884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08345__A1 vss _03887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09839_ vdd _02709_ _03984_ _04868_ rf_ram_if.rgnt vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_154_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05254__S1 vss _01375_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_829 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06659__A1 vss _02820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09845__A1 vss _01413_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_838 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_1237 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_512 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11663_ net186 vss vdd net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05867__C1 vss _01636_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09448__I1 vss net75 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10614_ vdd rf_ram.memory\[314\]\[0\] clknet_leaf_105_clk vss _00358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05882__A2 vss _01922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07084__A1 vss _03087_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11594_ vdd rf_ram.memory\[28\]\[1\] clknet_leaf_204_clk vss _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10545_ vdd rf_ram.memory\[371\]\[1\] clknet_leaf_153_clk vss _00289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_792 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_152 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_130_clk vdd vss clknet_leaf_130_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08820__A2 vss _04195_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10476_ vdd rf_ram.memory\[422\]\[0\] clknet_leaf_101_clk vss _00220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06831__A1 vss _02927_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05634__A2 vss _01623_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_676 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06304__B vss _01956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1110 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08336__A1 vss _03309_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_197_clk vdd vss clknet_leaf_197_clk clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06347__B1 vss _01721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11028_ vdd rf_ram.memory\[150\]\[0\] clknet_leaf_327_clk vss _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08887__A2 vss _02909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09836__A1 vss _04840_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05520_ rf_ram.memory\[322\]\[0\] _01716_ vss vdd rf_ram.memory\[321\]\[0\] _01715_
+ rf_ram.memory\[323\]\[0\] _01713_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_05451_ rf_ram.memory\[380\]\[0\] _01647_ vss vdd rf_ram.memory\[383\]\[0\] _01646_
+ rf_ram.memory\[381\]\[0\] _01645_ _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_137_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05873__A2 vss _01989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_540 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08170_ vdd _03793_ _03792_ _00570_ _03787_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_103_63 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07121_ vdd vss _03139_ _02829_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_83_882 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05382_ _01528_ vdd vss _01578_ rf_ram.memory\[544\]\[0\] _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_121_clk vdd vss clknet_leaf_121_clk clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06822__A1 vss _02909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07052_ vdd _03095_ _03094_ _00150_ _03087_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05625__A2 vss _01683_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput101 o_dbus_dat[12] net101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_42_278 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput112 o_dbus_dat[22] net112 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput123 o_dbus_dat[3] net123 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06003_ _02196_ _02197_ vdd vss _02198_ _02194_ _02195_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xoutput134 o_dbus_we net134 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05609__I vss _01503_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08575__A1 vss _04023_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput145 o_ext_rs1[16] net145 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput167 o_ext_rs1[7] net167 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput156 o_ext_rs1[26] net156 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput189 o_ext_rs2[27] net189 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput178 o_ext_rs2[17] net178 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06050__A2 vss _01606_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07954_ vdd _03657_ _03656_ _00490_ _03651_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08327__A1 vss _03884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07885_ vdd _03614_ _03613_ _00464_ _03587_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_188_clk vdd vss clknet_leaf_188_clk clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06905_ vdd vss _02999_ rf_ram.memory\[2\]\[0\] _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06836_ vdd _02951_ _02950_ _00078_ _02927_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06889__A1 vss _02975_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09624_ vdd vss _04722_ rf_ram.memory\[71\]\[1\] _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05344__I vss _01520_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_328 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09827__A1 vss _03668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06767_ vdd vss _02902_ rf_ram.memory\[513\]\[1\] _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09555_ _04526_ vdd vss _04674_ cpu.immdec.imm7 _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05718_ _01913_ vdd vss _01914_ _01909_ _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06698_ vdd vss _02854_ rf_ram.memory\[523\]\[0\] _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09486_ vdd vss _04623_ _01375_ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08506_ vdd vss _04010_ cpu.immdec.imm11_7\[2\] cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_136_715 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05649_ _01832_ _01844_ net253 vdd vss _01845_ _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_66_849 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08437_ vdd vss _03960_ rf_ram.memory\[174\]\[1\] _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09055__A2 vss _04339_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08368_ vdd vss _03916_ _02983_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xwire239 net239 _02893_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_112_clk vdd vss clknet_leaf_112_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07066__A1 vss _03092_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07319_ vdd vss _03263_ rf_ram.memory\[272\]\[0\] _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08299_ vdd vss _03873_ rf_ram.memory\[244\]\[0\] _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_554 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05616__A2 vss _01666_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10330_ vdd rf_ram.memory\[287\]\[0\] clknet_leaf_174_clk vss _00074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10261_ vdd _05126_ _05125_ _01329_ _02819_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05519__I vss _01714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10192_ vdd vss _05085_ rf_ram.memory\[238\]\[1\] _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06041__A2 vss _01537_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_179_clk vdd vss clknet_leaf_179_clk clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05682__C vss _01362_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10125__A1 vss net244 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07541__A2 vss _02904_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_657 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_1034 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_940 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11646_ net199 vss vdd net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_71_329 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05855__A2 vss _01515_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_103_clk vdd vss clknet_leaf_103_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput14 vss net14 i_dbus_rdt[20] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput25 vss net25 i_dbus_rdt[30] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11577_ vdd rf_ram.memory\[442\]\[0\] clknet_leaf_56_clk vss _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07057__A1 vss _03087_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_223 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput36 vss net36 i_ibus_rdt[11] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__06813__I vss _02800_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06804__A1 vss _02927_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput58 vss net58 i_ibus_rdt[3] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10528_ vdd rf_ram.memory\[250\]\[0\] clknet_leaf_217_clk vss _00272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput47 net47 vss vdd i_ibus_rdt[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_122_442 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06280__A2 vss _01940_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_497 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08557__A1 vss _04026_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10459_ vdd rf_ram.memory\[473\]\[1\] clknet_leaf_43_clk vss _00203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05429__I vss _01624_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_868 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05873__B vss _01783_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05791__A1 vss _01351_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07670_ vdd _03480_ _03478_ _00383_ _03458_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09809__A1 vss _04837_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06621_ vdd vss _02793_ _02785_ _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_59_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06552_ vss _02738_ _02737_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09340_ _04540_ net213 vdd vss _04541_ cpu.ctrl.pc _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05503_ rf_ram.memory\[339\]\[0\] _01698_ vdd vss _01699_ rf_ram.memory\[338\]\[0\]
+ _01687_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_74_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09271_ vdd vss _04495_ _01364_ cpu.genblk3.csr.mcause3_0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_512 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06483_ _02676_ _02677_ vdd vss _02678_ _02674_ _02675_ _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08222_ vdd vss _03826_ rf_ram.memory\[533\]\[0\] _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05434_ _01629_ vdd vss _01630_ _01622_ _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05846__A2 vss _01649_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08153_ vdd _03782_ _03781_ _00564_ _03754_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05365_ rf_ram.memory\[539\]\[0\] _01540_ _01544_ rf_ram.memory\[538\]\[0\] _01561_
+ vss vdd rf_ram.memory\[537\]\[0\] _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__06256__C1 vss _01811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1220 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07104_ vdd vss _03128_ _02915_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08796__A1 vss _04170_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1074 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08084_ vdd vss _03740_ rf_ram.memory\[55\]\[0\] _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_1025 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_751 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05296_ vss _00003_ _01492_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07035_ _03083_ vss vdd net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_140_261 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08548__A1 vss net235 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_475 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06271__A2 vss _01735_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06008__C1 vss _01555_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_484 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1236 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08986_ vdd _04312_ _04310_ _00867_ _04301_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07220__A1 vss _03193_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05783__B vss _01978_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06023__A2 vss _01538_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07937_ vdd _03646_ _03645_ _00484_ _03619_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input33_I vss i_dbus_rdt[9] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10107__A1 vss _05014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1170 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07868_ vdd vss _03604_ _02991_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07799_ vdd vss _03562_ rf_ram.memory\[415\]\[1\] _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05534__A1 vss _01674_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06819_ vdd vss _02939_ _02796_ _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09607_ vdd _04681_ _01331_ _01087_ _04643_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_167_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09538_ vdd vss _04663_ _04526_ net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_607 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07287__A1 vss _03222_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_955 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11500_ vdd rf_ram.memory\[277\]\[1\] clknet_leaf_179_clk vss _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_819 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_333_clk vdd vss clknet_leaf_333_clk clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09469_ _04604_ vdd vss _04611_ net84 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_184_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_370 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11431_ vdd rf_ram.memory\[61\]\[0\] clknet_leaf_291_clk vss _01163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_149_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11362_ _01094_ vdd vss clknet_leaf_257_clk cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08787__A1 vss _03071_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10313_ vdd rf_ram.memory\[514\]\[1\] clknet_leaf_267_clk vss _00057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11293_ vdd rf_ram.memory\[299\]\[1\] clknet_leaf_133_clk vss _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10244_ vdd vss _05116_ _02727_ _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07211__A1 vss _02795_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10175_ vdd vss _05074_ rf_ram.memory\[20\]\[1\] _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_1210 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08711__A1 vss _04126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_618 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_361 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_465 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_324_clk vdd vss clknet_leaf_324_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_72_616 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05828__A2 vss _01804_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_893 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05868__B vss _01684_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11629_ vss net152 net79 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_1214 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06543__I vss cpu.immdec.imm11_7\[4\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_727 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05150_ _01353_ vss vdd _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__06253__A2 vss _01804_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05159__I vss _01361_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05461__B1 vss _01654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08840_ vdd vss _04222_ _02805_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06005__A2 vss _01532_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06410__C1 vss _01931_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05983_ rf_ram.memory\[5\]\[0\] _01714_ _01643_ rf_ram.memory\[4\]\[0\] _02179_ vss
+ vdd rf_ram.memory\[7\]\[0\] _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA_clkbuf_3_1_0_clk_I vss clknet_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08771_ vdd _04179_ _04177_ _00785_ _04170_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07722_ vdd _03513_ _03512_ _00402_ _03488_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07653_ vdd _03470_ _03469_ _00376_ _03455_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11624__I vss net74 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_306_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06604_ vdd vss _02780_ _02779_ _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_07584_ vdd vss _03428_ rf_ram.memory\[316\]\[0\] _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_125_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09323_ vdd vss _04530_ net243 _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06718__I vss _02865_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07269__A1 vss _03230_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_454 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_315_clk vdd vss clknet_leaf_315_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06535_ vdd vss cpu.immdec.imm11_7\[0\] _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_1241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06466_ _02660_ vdd vss _02661_ _01903_ _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_34_1095 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09254_ _04481_ vdd vss _04482_ _01356_ _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_146_887 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_364 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06492__A2 vss _02630_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09185_ vdd vss _04437_ rf_ram.memory\[179\]\[0\] _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05417_ _01613_ vss vdd _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_28_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08205_ vdd vss _03815_ rf_ram.memory\[536\]\[0\] _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06229__C1 vss _01721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06397_ rf_ram.memory\[92\]\[1\] _02592_ vss vdd rf_ram.memory\[95\]\[1\] _01773_
+ rf_ram.memory\[93\]\[1\] _01772_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_08136_ vdd vss _03772_ _03668_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08769__A1 vss _04167_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_378 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05348_ _01544_ _01543_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07441__A1 vss _03323_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08067_ _03729_ vss vdd _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_05279_ vdd _01477_ _01475_ cpu.o_wdata0 _01366_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_109_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07018_ _03072_ vss vdd _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_3_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09194__A1 vss net236 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08941__A1 vss _04266_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06402__B vss _01707_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08969_ vdd vss _04302_ rf_ram.memory\[118\]\[1\] _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_902 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10931_ vdd rf_ram.memory\[176\]\[1\] clknet_leaf_12_clk vss _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10862_ vdd rf_ram.memory\[205\]\[0\] clknet_leaf_30_clk vss _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_501 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10793_ vdd rf_ram.memory\[560\]\[1\] clknet_leaf_325_clk vss _00537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_123 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_306_clk vdd vss clknet_leaf_306_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_81_413 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_898 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_887 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11414_ vdd rf_ram.memory\[76\]\[1\] clknet_leaf_21_clk vss _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_660 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11345_ vdd cpu.immdec.imm30_25\[1\] clknet_leaf_260_clk vss _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11276_ vdd net211 clknet_leaf_246_clk vss _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10227_ vdd vss _05106_ rf_ram.memory\[212\]\[1\] _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_1231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05707__I vss _01525_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06312__B vss _02004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10158_ vdd vss _05064_ rf_ram.memory\[44\]\[0\] _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_94_1207 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10089_ vdd _05021_ _05019_ _01262_ _05017_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05870__C vss _01620_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09488__A2 vss _03989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06171__A1 vss _01527_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_903 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08999__A1 vss _04298_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1149 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06320_ rf_ram.memory\[178\]\[1\] _02515_ vss vdd rf_ram.memory\[177\]\[1\] _01931_
+ rf_ram.memory\[179\]\[1\] _01911_ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA_clkbuf_leaf_292_clk_I vss clknet_5_24__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_23__f_clk_I vss clknet_3_5_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06251_ _02445_ vdd vss _02446_ _01909_ _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_5_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10935__D vss cpu.o_wdata1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05202_ vdd vss cpu.state.stage_two_req _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06182_ vdd vss _02377_ rf_ram.memory\[468\]\[1\] _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09412__A2 vss _02801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_384 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07423__A1 vss _03326_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06226__A2 vss _01634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06206__C vss _01717_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1033 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05133_ vdd vss _01336_ cpu.decode.opcode\[2\] cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_09941_ vdd _04930_ _04929_ _01205_ _04918_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09176__A1 vss _04401_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11619__I vss net69 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08923__A1 vss _04269_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09872_ vdd _04888_ _04885_ _01178_ _04887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_230_clk_I vss clknet_5_23__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05737__A1 vss _01909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08823_ vdd vss _04212_ rf_ram.memory\[136\]\[1\] _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05966_ vdd vss _02162_ rf_ram.memory\[17\]\[0\] _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08754_ vdd vss _04169_ rf_ram.memory\[146\]\[0\] _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07705_ vdd vss _03503_ _02960_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_245_clk_I vss clknet_5_21__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09479__A2 vss net89 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_721 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_92_clk vdd vss clknet_leaf_92_clk clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05897_ _01684_ vdd vss _02093_ rf_ram.memory\[88\]\[0\] _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08685_ vdd vss _04125_ rf_ram.memory\[155\]\[1\] _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08151__A2 vss _03765_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07636_ vdd vss _03460_ _03008_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07567_ vdd vss _03417_ rf_ram.memory\[357\]\[0\] _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09306_ vdd vss _04519_ rf_ram.memory\[63\]\[1\] _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06518_ _02707_ _01411_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09237_ vdd vss _04469_ rf_ram.memory\[319\]\[0\] _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07498_ vdd vss _03374_ _03319_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06449_ _02643_ vdd vss _02644_ _01903_ _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06465__A2 vss _01605_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_800 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output187_I vss net187 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09168_ vdd vss _04426_ rf_ram.memory\[86\]\[0\] _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_896 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07414__A1 vss _03289_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06217__A2 vss _01782_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09099_ vdd _04382_ _04381_ _00910_ _04364_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08119_ vdd _03761_ _03759_ _00551_ _03757_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_32_866 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11130_ vdd rf_ram.memory\[115\]\[0\] clknet_leaf_73_clk vss _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09167__A1 vss _03008_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06132__B vss _01783_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11061_ vdd rf_ram.memory\[13\]\[0\] clknet_leaf_31_clk vss _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10012_ vdd vss _04974_ rf_ram.memory\[348\]\[0\] _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08390__A2 vss _02829_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_321 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_83_clk vdd vss clknet_leaf_83_clk clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_93_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_505 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06153__A1 vss _01597_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10914_ vdd rf_ram.memory\[209\]\[0\] clknet_leaf_28_clk vss _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10845_ vdd rf_ram.memory\[534\]\[1\] clknet_leaf_308_clk vss _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_936 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10776_ vdd rf_ram.memory\[568\]\[0\] clknet_leaf_324_clk vss _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_164_470 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07653__A1 vss _03455_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_939 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06307__B vss _01564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_298 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07405__A1 vss _03292_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06026__C vss _01495_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11328_ vdd rf_ram.memory\[289\]\[0\] clknet_leaf_123_clk vss _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05437__I vss _01508_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11259_ _00994_ vdd vss clknet_leaf_250_clk net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_101_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05820_ _02015_ _01569_ vdd vss _02016_ _01768_ _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_167_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_94_1037 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_74_clk vdd vss clknet_leaf_74_clk clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05751_ _01946_ _01569_ vdd vss _01947_ _01674_ _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_187_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09330__A1 vss _04463_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05682_ _01877_ _01362_ vdd vss _01878_ _01674_ _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08470_ vdd vss rf_ram_if.rreq_r _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_49_229 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07892__A1 vss _03590_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07421_ _03326_ _03017_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_58_741 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09881__A2 vss _02795_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_92_519 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07352_ vdd _03282_ _03280_ _00263_ _03260_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_605 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1032 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_418 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06303_ _01494_ vdd vss _02498_ _02495_ _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09633__A2 vss net59 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_941 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06217__B vss _01783_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07283_ vdd vss _03240_ rf_ram.memory\[472\]\[1\] _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06447__A2 vss _01536_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06234_ rf_ram.memory\[402\]\[1\] _02429_ vss vdd rf_ram.memory\[401\]\[1\] _01656_
+ rf_ram.memory\[403\]\[1\] _01763_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_143_665 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09022_ vdd vss _04335_ rf_ram.memory\[108\]\[1\] _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_32_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_143_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06165_ vdd vss _02360_ rf_ram.memory\[484\]\[1\] _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06096_ _02290_ vdd vss _02291_ _01368_ _02263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__06731__I vss _02825_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09924_ vdd vss _04920_ rf_ram.memory\[342\]\[0\] _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05347__I vss _01530_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09855_ _04876_ vdd vss _01172_ _02713_ _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_08806_ vdd vss _04201_ rf_ram.memory\[13\]\[1\] _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_184_clk_I vss clknet_5_29__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06383__A1 vss _01972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09786_ vdd vss _04835_ rf_ram.memory\[76\]\[0\] _04834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05186__A2 vss _01385_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06998_ vdd vss _03060_ rf_ram.memory\[225\]\[0\] _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_65_clk vdd vss clknet_leaf_65_clk clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_64_clk_I vss clknet_5_8__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05949_ vdd vss _02145_ rf_ram.memory\[62\]\[0\] _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_505 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08737_ vdd vss _00773_ _01369_ _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08668_ vdd vss _04115_ rf_ram.memory\[157\]\[0\] _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09321__B2 vss cpu.immdec.imm30_25\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09321__A1 vss _04526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07619_ vdd vss _03449_ _02904_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_404 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07883__A1 vss _02836_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_199_clk_I vss clknet_5_25__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_869 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10630_ vdd rf_ram.memory\[405\]\[0\] clknet_leaf_102_clk vss _00374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_245 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08599_ vdd vss _04072_ rf_ram.memory\[165\]\[0\] _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_79_clk_I vss clknet_5_11__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_796 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10561_ vdd rf_ram.memory\[367\]\[1\] clknet_leaf_163_clk vss _00305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07635__A1 vss _03458_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_122_clk_I vss clknet_5_15__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_963 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10492_ vdd rf_ram.memory\[472\]\[0\] clknet_leaf_126_clk vss _00236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05646__B1 vss _01763_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_799 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_298 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_367 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09388__A1 vss net216 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_137_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1083 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11113_ vdd rf_ram.memory\[399\]\[1\] clknet_leaf_93_clk vss _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_1104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_17_clk_I vss clknet_5_2__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11044_ vdd rf_ram_if.wen1_r clknet_leaf_259_clk vss _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08363__A2 vss _03903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_56_clk vdd vss clknet_leaf_56_clk clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_162 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_302 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_1043 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08115__A2 vss _03729_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_1196 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_746 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_508 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_1038 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_903 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05720__I vss _01550_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10828_ vdd rf_ram.memory\[542\]\[0\] clknet_leaf_274_clk vss _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07626__A1 vss _03422_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10759_ vdd rf_ram.memory\[467\]\[1\] clknet_leaf_125_clk vss _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06429__A2 vss _01641_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_643 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_36_991 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_696 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1145 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07970_ vdd vss _03667_ rf_ram.memory\[47\]\[1\] _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_1009 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06921_ _03009_ vss vdd _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09551__A1 vss _01391_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06852_ vdd vss _02963_ rf_ram.memory\[285\]\[1\] _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09640_ vdd vss _04729_ rf_ram.memory\[78\]\[0\] _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06783_ vdd vss _02914_ rf_ram.memory\[511\]\[1\] _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09571_ _03967_ vdd vss _04686_ cpu.immdec.imm30_25\[4\] net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05803_ _01564_ vdd vss _01999_ _01996_ _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05734_ vdd vss _01930_ rf_ram.memory\[446\]\[0\] _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_47_clk vdd vss clknet_leaf_47_clk clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09303__A1 vss _03668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08522_ vdd vss _04022_ rf_ram.memory\[188\]\[1\] _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_713 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08453_ vdd vss _03970_ _01418_ _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_148_768 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07865__A1 vss _03587_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05665_ _01860_ vdd vss _01861_ _01855_ _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07404_ vdd vss _03315_ rf_ram.memory\[247\]\[1\] _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11632__I vss net82 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05596_ vdd vss _01792_ rf_ram.memory\[292\]\[0\] _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_133_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08384_ vdd _03926_ _03924_ _00651_ _03922_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07335_ vdd _03272_ _03271_ _00256_ _03257_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07266_ vdd vss _03229_ rf_ram.memory\[196\]\[1\] _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08290__A1 vss _03852_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_287 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06217_ _01783_ vdd vss _02412_ rf_ram.memory\[384\]\[1\] _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09005_ vdd vss _04324_ rf_ram.memory\[111\]\[1\] _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07197_ vdd vss _03186_ rf_ram.memory\[474\]\[1\] _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input63_I vss i_ibus_rdt[8] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06148_ rf_ram.memory\[312\]\[1\] _02343_ vss vdd rf_ram.memory\[315\]\[1\] _01811_
+ rf_ram.memory\[313\]\[1\] _01810_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__08042__A1 vss _03686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06053__B1 vss _01610_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06079_ _01620_ vdd vss _02274_ _02271_ _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_111_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08593__A2 vss _04067_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09907_ vdd vss _04909_ rf_ram.memory\[292\]\[0\] _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09542__A1 vss _04478_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10152__A2 vss _02894_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09838_ vdd vss _04867_ cpu.state.cnt_r\[3\] _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09769_ vdd vss _04824_ _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_38_clk vdd vss clknet_leaf_38_clk clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_150_1119 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09845__A2 vss _03989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_407 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11662_ vss net185 net113 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05867__B1 vss _01610_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06636__I vss _02805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10613_ vdd rf_ram.memory\[354\]\[1\] clknet_leaf_156_clk vss _00357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07608__A1 vss _02898_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11593_ vdd rf_ram.memory\[28\]\[0\] clknet_leaf_210_clk vss _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10544_ vdd rf_ram.memory\[371\]\[0\] clknet_leaf_153_clk vss _00288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_654 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_991 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_771 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10475_ vdd rf_ram.memory\[423\]\[1\] clknet_leaf_103_clk vss _00219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_102_370 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08336__A2 vss _02946_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1019 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09533__A1 vss _04478_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11027_ vdd rf_ram.memory\[151\]\[1\] clknet_leaf_2_clk vss _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_1176 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05715__I vss _01695_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_622 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_29_clk vdd vss clknet_leaf_29_clk clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_644 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07847__A1 vss _03590_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1030 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05450_ _01646_ _01635_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05450__I vss _01635_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05381_ rf_ram.memory\[549\]\[0\] _01539_ _01538_ rf_ram.memory\[548\]\[0\] _01577_
+ vss vdd rf_ram.memory\[551\]\[0\] _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_28_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_568 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07120_ vdd _03138_ _03136_ _00175_ _03126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_55_596 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_265 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08272__A1 vss _03855_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06822__A2 vss _02941_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07051_ vdd vss _03095_ rf_ram.memory\[390\]\[0\] _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput113 o_dbus_dat[23] net113 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput102 o_dbus_dat[13] net102 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06002_ rf_ram.memory\[514\]\[1\] _02197_ vss vdd rf_ram.memory\[513\]\[1\] _01539_
+ rf_ram.memory\[515\]\[1\] _01540_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
Xoutput124 o_dbus_dat[4] net124 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08024__A1 vss _03690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09772__A1 vss _04634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput135 o_ext_funct3[0] net135 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput168 o_ext_rs1[8] net168 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput146 o_ext_rs1[17] net146 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_2_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput157 o_ext_rs1[27] net157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput179 o_ext_rs2[18] net179 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05389__A2 vss _01544_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07953_ vdd vss _03657_ rf_ram.memory\[481\]\[0\] _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11627__I vss net77 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05794__C1 vss _01516_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06230__B vss _01629_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07884_ vdd vss _03614_ rf_ram.memory\[462\]\[0\] _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06904_ vdd vss _02998_ _02894_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06338__A1 vss _01972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06835_ vdd vss _02951_ rf_ram.memory\[286\]\[0\] _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09623_ vdd _04721_ _04720_ _01095_ _04634_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_167_307 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05561__A2 vss _01755_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09827__A2 vss _02917_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06766_ vdd _02901_ _02900_ _00058_ _02873_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09554_ _01419_ vdd vss _04673_ cpu.immdec.imm31 _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__07838__A1 vss _03554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05717_ rf_ram.memory\[439\]\[0\] _01911_ _01706_ rf_ram.memory\[438\]\[0\] _01913_
+ vss vdd rf_ram.memory\[437\]\[0\] _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_66_817 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06697_ vdd vss _02853_ _02781_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09485_ _04621_ vdd vss _04622_ _01411_ _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_38_508 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08505_ vdd vss _04009_ _01369_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_110_1103 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_919 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_407 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05648_ _01838_ _01660_ _01843_ vdd vss _01844_ _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_08436_ vdd _03959_ _03958_ _00670_ _03953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06510__A1 vss _01382_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_535 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08367_ vdd _03915_ _03913_ _00645_ _03887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_50_1271 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05579_ _01774_ vdd vss _01775_ _01769_ _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07318_ vdd vss _03262_ _02958_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_117_941 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_360 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_473 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08298_ vdd vss _03872_ _03309_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08263__A1 vss _03820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07249_ vdd vss _03218_ rf_ram.memory\[420\]\[1\] _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10070__A1 vss _04982_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10260_ vdd vss _05126_ rf_ram.memory\[574\]\[0\] _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08015__A1 vss _02839_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06124__C vss _01361_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10191_ vdd _05084_ _05083_ _01301_ _05078_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05785__C1 vss _01857_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06140__B vss _01707_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10125__A2 vss _02832_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05552__A2 vss _01543_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1172 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_441 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_1160 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_338 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_373 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06501__A1 vss cpu.ctrl.pc vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_168 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11645_ vss net198 net126 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput15 vss net15 i_dbus_rdt[21] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_190 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput26 vss net26 i_dbus_rdt[31] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11576_ vdd rf_ram.memory\[211\]\[1\] clknet_leaf_29_clk vss _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput37 vss net37 i_ibus_rdt[12] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10527_ vdd rf_ram.memory\[267\]\[1\] clknet_leaf_140_clk vss _00271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput48 vss net48 i_ibus_rdt[23] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput59 vss net59 i_ibus_rdt[4] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_165_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_122_465 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10458_ vdd rf_ram.memory\[473\]\[0\] clknet_leaf_44_clk vss _00202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_942 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1045 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_1165 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_69 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10389_ vdd rf_ram.memory\[225\]\[1\] clknet_leaf_273_clk vss _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09506__A1 vss _04637_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05445__I vss _01640_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05791__A2 vss _01971_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06620_ vdd vss _02792_ _02723_ _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_177_605 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05543__A2 vss _01683_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_290 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08756__I vss _04061_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06740__A1 vss _02716_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06551_ vdd vss _02737_ _02731_ _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08493__A1 vss _02829_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05502_ vdd vss _01698_ rf_ram.memory\[337\]\[0\] _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06482_ rf_ram.memory\[9\]\[1\] _01714_ _01643_ rf_ram.memory\[8\]\[1\] _02677_ vss
+ vdd rf_ram.memory\[11\]\[1\] _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_87_496 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09270_ _04494_ _01485_ vdd vss _00969_ _04492_ _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05433_ _01629_ _01563_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08221_ vdd vss _03825_ _03798_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05700__C1 vss _01608_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_500 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08245__A1 vss _03823_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08152_ vdd vss _03782_ rf_ram.memory\[546\]\[0\] _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05364_ _01552_ vdd vss _01560_ rf_ram.memory\[536\]\[0\] _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06256__B1 vss _01810_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10052__A1 vss _04985_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09993__A1 vss _04950_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07103_ vdd _03127_ _03124_ _00169_ _03126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05295_ _01491_ vdd vss _01492_ _01486_ _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08083_ vdd vss _03739_ _03668_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_9_clk vdd vss clknet_leaf_9_clk clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_5_15__f_clk vdd vss clknet_5_15__leaf_clk clknet_3_3_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07034_ vdd vss _03082_ _02779_ _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08548__A2 vss _04038_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_696 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06008__B1 vss _01554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08985_ vdd vss _04312_ rf_ram.memory\[115\]\[1\] _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09255__C vss _01341_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07936_ vdd vss _03646_ rf_ram.memory\[457\]\[0\] _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05231__A1 vss cpu.bufreg.i_sh_signed vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05355__I vss _01550_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input26_I vss i_dbus_rdt[31] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1069 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07867_ vdd _03603_ _03601_ _00457_ _03590_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07798_ vdd _03561_ _03560_ _00430_ _03554_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06818_ vdd _02938_ _02936_ _00073_ _02930_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09606_ vdd vss _01086_ _04712_ _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_35_1008 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09537_ vdd vss _04662_ cpu.csr_imm _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06749_ _02889_ vss vdd _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_182_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_513 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06495__B1 vss _02462_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09468_ vss _01051_ _04610_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08419_ vdd vss _03948_ rf_ram.memory\[29\]\[1\] _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09399_ vdd vss _04572_ _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_188_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11430_ vdd rf_ram.memory\[62\]\[1\] clknet_leaf_289_clk vss _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08236__A1 vss _03798_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06247__B1 vss _01925_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10043__A1 vss _02812_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11361_ _01093_ vdd vss clknet_leaf_258_clk cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_46_1115 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08787__A2 vss _04152_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06135__B vss _01790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06798__A1 vss _02873_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output94_I vss net94 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10312_ vdd rf_ram.memory\[514\]\[0\] clknet_leaf_262_clk vss _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11292_ vdd rf_ram.memory\[299\]\[0\] clknet_leaf_133_clk vss _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09736__A1 vss _04781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10243_ vdd _05115_ _05113_ _01322_ _02825_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07211__A2 vss _02941_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10174_ vdd _05073_ _05072_ _01295_ _05046_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05758__C1 vss _01953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_794 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05222__A1 vss _01385_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05773__A2 vss _01958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1109 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06183__C1 vss _01848_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06722__A1 vss _02866_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05930__C1 vss _01772_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_496 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1075 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85_967 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08475__A1 vss _01436_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11628_ vss net151 net78 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_154_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09975__A1 vss _02922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_782 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_886 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11559_ vdd rf_ram.memory\[448\]\[0\] clknet_leaf_112_clk vss _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_588 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_69_79 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05997__C1 vss _01517_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09727__A1 vss _04781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06410__B1 vss _01911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_260_clk vdd vss clknet_leaf_260_clk clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05982_ _01503_ vdd vss _02178_ rf_ram.memory\[6\]\[0\] _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05764__A2 vss _01515_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08770_ vdd vss _04179_ rf_ram.memory\[144\]\[1\] _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07721_ vdd vss _03513_ rf_ram.memory\[398\]\[0\] _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_402 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05516__A2 vss _01711_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07652_ vdd vss _03470_ rf_ram.memory\[386\]\[0\] _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07583_ vdd vss _03427_ _02935_ _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_149_104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_1091 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_901 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06603_ vdd vss _02779_ _01496_ _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_177_479 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_159 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06534_ _01366_ _02720_ _01332_ vss _01347_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09322_ vdd vss _04529_ _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_164_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07269__A2 vss _02899_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_948 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06465_ rf_ram.memory\[23\]\[1\] _01624_ _01605_ rf_ram.memory\[22\]\[1\] _02660_
+ vss vdd rf_ram.memory\[21\]\[1\] _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_09253_ vdd vss _04481_ _01366_ _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05416_ _01611_ vdd vss _01612_ _01603_ _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_146_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06396_ vdd vss _02591_ rf_ram.memory\[94\]\[1\] _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09184_ vdd vss _04436_ net242 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_959 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08204_ vdd vss _03814_ _03798_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06229__B1 vss _01726_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09966__A1 vss _04918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10025__A1 vss _04953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05347_ _01543_ vss vdd _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_7_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08135_ vdd _03771_ _03769_ _00557_ _03757_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_70_160 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_925 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08066_ vdd _03728_ _03726_ _00531_ _03724_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05278_ _01476_ _01366_ vdd vss _01477_ _01381_ _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__05452__A1 vss _01527_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1024 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07017_ vdd vss _03071_ _02750_ _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__09194__A2 vss _04418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_45_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_251_clk vdd vss clknet_leaf_251_clk clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08968_ _04301_ _04061_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08899_ vdd _04258_ _04257_ _00834_ _04234_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07919_ vdd _03635_ _03633_ _00477_ _03622_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output132_I vss net132 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10930_ vdd rf_ram.memory\[176\]\[0\] clknet_leaf_6_clk vss _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05507__A2 vss _01623_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1131 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06704__A1 vss _02820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_969 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_79_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10861_ vdd rf_ram.memory\[526\]\[1\] clknet_leaf_315_clk vss _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_939 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10792_ vdd rf_ram.memory\[560\]\[0\] clknet_leaf_323_clk vss _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_321 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05969__B vss _01550_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_343 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_296 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_959 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08209__A1 vss _03798_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_847 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11413_ vdd rf_ram.memory\[76\]\[0\] clknet_leaf_21_clk vss _01145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_741 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_503 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11344_ vdd cpu.immdec.imm30_25\[0\] clknet_leaf_260_clk vss _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11275_ vdd net210 clknet_leaf_246_clk vss _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07475__I vss _03359_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1179 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10226_ vdd _05105_ _05104_ _01315_ _05078_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05994__A2 vss _01502_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07196__A1 vss _03157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_242_clk vdd vss clknet_leaf_242_clk clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05746__A2 vss _01666_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10157_ vdd vss _05063_ _02787_ _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06943__A1 vss _03014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10088_ vdd vss _05021_ rf_ram.memory\[30\]\[1\] _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08696__A1 vss _04126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1220 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05903__C1 vss _01715_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08448__A1 vss _03956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07120__A1 vss _03126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_786 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06250_ rf_ram.memory\[444\]\[1\] _02445_ vss vdd rf_ram.memory\[447\]\[1\] _01857_
+ rf_ram.memory\[445\]\[1\] _01931_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_26_831 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_471 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09948__A1 vss _04921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05682__A1 vss _01674_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05201_ vdd vss _01401_ _01399_ _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_25_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06181_ _02363_ _02375_ net253 vdd vss _02376_ _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_41_823 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05132_ cpu.csr_d_sel vdd vss _01335_ cpu.decode.co_mem_word cpu.bne_or_bge vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__08620__A1 vss _02760_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09940_ vdd vss _04930_ rf_ram.memory\[33\]\[0\] _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_889 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05985__A2 vss _01661_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_964 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_975 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_580 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09871_ vdd vss _04888_ rf_ram.memory\[60\]\[1\] _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_233_clk vdd vss clknet_leaf_233_clk clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08822_ vdd _04211_ _04210_ _00804_ _04202_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05965_ _01601_ vdd vss _02161_ rf_ram.memory\[16\]\[0\] _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08753_ vdd vss _04168_ net236 _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07704_ vdd _03502_ _03500_ _00395_ _03491_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_1130 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09479__A3 vss _03989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05896_ _02091_ vdd vss _02092_ _01769_ _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_17_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08684_ vdd _04124_ _04123_ _00753_ _04094_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07635_ vdd _03459_ _03456_ _00369_ _03458_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06162__A2 vss _01697_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07566_ vdd vss _03416_ _02795_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08439__A1 vss _02953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10246__A1 vss _02819_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09305_ vdd _04518_ _04517_ _00980_ _04463_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05789__B vss _01928_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06517_ vdd vss _02706_ _02703_ _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_180_419 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07497_ vdd _03373_ _03371_ _00317_ _03360_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09236_ vdd vss _04468_ _03445_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_119_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07111__A1 vss _03123_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06448_ rf_ram.memory\[39\]\[1\] _01607_ _01661_ rf_ram.memory\[38\]\[1\] _02643_
+ vss vdd rf_ram.memory\[37\]\[1\] _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_09167_ vdd vss _04425_ _03008_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06379_ _02573_ _01569_ vdd vss _02574_ _01768_ _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09098_ vdd vss _04382_ rf_ram.memory\[96\]\[0\] _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08118_ vdd vss _03761_ rf_ram.memory\[553\]\[1\] _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_344 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_390 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08049_ vdd _03717_ _03715_ _00525_ _03690_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09167__A2 vss _04418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05808__I vss _01504_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11060_ vdd rf_ram.memory\[140\]\[1\] clknet_leaf_10_clk vss _00797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10011_ vdd vss _04973_ _04911_ _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07178__A1 vss _03161_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05728__A2 vss _01922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_224_clk vdd vss clknet_leaf_224_clk clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_99_834 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07350__A1 vss _03257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10913_ vdd rf_ram.memory\[17\]\[1\] clknet_leaf_288_clk vss _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_742 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10844_ vdd rf_ram.memory\[534\]\[0\] clknet_leaf_312_clk vss _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_641 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05900__A2 vss _01785_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_200 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07102__A1 vss rf_ram.memory\[48\]\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10775_ vdd rf_ram.memory\[56\]\[1\] clknet_leaf_294_clk vss _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08850__A1 vss net241 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1089 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08602__A1 vss _04062_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_182 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05416__A1 vss _01603_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11327_ vdd cpu.alu.cmp_r clknet_leaf_233_clk vss _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05967__A2 vss _01605_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_305_clk_I vss clknet_5_4__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07169__A1 vss _02915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11258_ _00993_ vdd vss clknet_leaf_248_clk cpu.ctrl.pc vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06916__A1 vss _02970_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10209_ vdd vss _05095_ net245 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_215_clk vdd vss clknet_leaf_215_clk clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11189_ vdd rf_ram.memory\[169\]\[1\] clknet_leaf_8_clk vss _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05750_ _01945_ vdd vss _01946_ _01350_ _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__06392__A2 vss _01510_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05195__A3 vss cpu.decode.opcode\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05453__I vss _01613_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08669__A1 vss _04094_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05681_ _01876_ vdd vss _01877_ _01350_ _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_77_528 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07420_ vdd _03325_ _03324_ _00288_ _03323_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_159_265 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09469__I0 vss net84 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07351_ vdd vss _03282_ rf_ram.memory\[26\]\[1\] _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10228__A1 vss _05081_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_279 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09094__A1 vss _04364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06302_ _01953_ rf_ram.memory\[163\]\[1\] vdd vss _02497_ rf_ram.memory\[162\]\[1\]
+ _01958_ _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_155_471 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07282_ vdd _03239_ _03238_ _00236_ _03222_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_182_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06233_ _01903_ vdd vss _02428_ rf_ram.memory\[400\]\[1\] _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09021_ vss _04334_ _04061_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_66_1118 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_683 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06164_ _01620_ vdd vss _02359_ _02356_ _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_180_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06233__B vss _01903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06095_ _02289_ _01361_ vdd vss _02290_ _01350_ _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__05958__A2 vss _01499_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_185 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09923_ vdd vss _04919_ _04911_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08004__I vss _02747_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_206_clk vdd vss clknet_leaf_206_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09854_ cpu.mem_bytecnt\[1\] vdd vss _04876_ _01385_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08805_ vdd _04200_ _04199_ _00798_ _04167_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05791__C vss _01362_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09785_ vdd vss _04834_ _02787_ _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_1247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06997_ vdd vss _03059_ _03055_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05948_ _02140_ _02143_ vdd vss _02144_ _02132_ _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08736_ _03984_ vdd vss _04157_ _02713_ _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__07332__A1 vss _03260_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05879_ vdd vss _02075_ rf_ram.memory\[78\]\[0\] _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08667_ vdd vss _04114_ _02959_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09321__A2 vss net36 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07618_ vdd _03448_ _03446_ _00363_ _03425_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07883__A2 vss _02972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08598_ vdd vss _04071_ _02794_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07549_ vdd vss _03406_ rf_ram.memory\[35\]\[1\] _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10560_ vdd rf_ram.memory\[367\]\[0\] clknet_leaf_162_clk vss _00304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_931 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08832__A1 vss _04202_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_469 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10491_ vdd rf_ram.memory\[417\]\[1\] clknet_leaf_98_clk vss _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09219_ vdd vss _04457_ _03319_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_815 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06071__A1 vss _01675_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_541 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05949__A2 vss _01530_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11112_ vdd rf_ram.memory\[399\]\[0\] clknet_leaf_93_clk vss _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08899__A1 vss _04234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05982__B vss _01503_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11043_ vdd rf_ram.memory\[146\]\[1\] clknet_leaf_336_clk vss _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_291_clk_I vss clknet_5_18__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07571__A1 vss _02935_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06374__A2 vss _01677_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06126__A2 vss _01863_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07323__A1 vss _03055_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08584__I vss _04061_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1175 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_230 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09076__A1 vss _04367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10827_ vdd rf_ram.memory\[543\]\[1\] clknet_leaf_312_clk vss _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07626__A2 vss _03452_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_780 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10758_ vdd rf_ram.memory\[467\]\[0\] clknet_leaf_125_clk vss _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05222__B vss cpu.mem_bytecnt\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06037__C vss _01564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10689_ vdd rf_ram.memory\[435\]\[1\] clknet_leaf_82_clk vss _00433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_164_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_164_1065 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_1174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_244_clk_I vss clknet_5_21__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05448__I vss _01643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06920_ vdd vss _03008_ _02773_ _03007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA_clkbuf_leaf_259_clk_I vss clknet_5_17__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06851_ vdd _02962_ _02961_ _00082_ _02927_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06365__A2 vss _01940_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06782_ vdd _02913_ _02912_ _00062_ _02873_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09570_ vdd _04685_ _04678_ _01078_ _04680_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05802_ _01520_ rf_ram.memory\[171\]\[0\] vdd vss _01998_ rf_ram.memory\[170\]\[0\]
+ _01989_ _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_05733_ _01928_ vdd vss _01929_ _01924_ _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09303__A2 vss _02909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_815 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08521_ vdd _04021_ _04020_ _00693_ _03953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07314__A1 vss _03257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08452_ vdd vss _03969_ _01369_ _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_33_1106 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_870 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05876__A1 vss _01600_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07403_ vdd _03314_ _03313_ _00282_ _03289_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05664_ _01860_ vss vdd _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_175_566 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06228__B vss _01615_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_909 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05595_ _01790_ vdd vss _01791_ _01784_ _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09067__A1 vss _04331_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_328 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08383_ vdd vss _03926_ rf_ram.memory\[180\]\[1\] _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_948 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07617__A2 vss _03446_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_994 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07334_ vdd vss _03272_ rf_ram.memory\[254\]\[0\] _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08814__A1 vss _04205_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07265_ vdd _03228_ _03227_ _00230_ _03222_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06216_ _01746_ vdd vss _02411_ _02408_ _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09004_ vdd _04323_ _04322_ _00874_ _04298_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_84_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07196_ vdd _03185_ _03184_ _00204_ _03157_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06147_ _01650_ vdd vss _02342_ rf_ram.memory\[314\]\[1\] _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__05358__I vss _01520_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_483 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06078_ rf_ram.memory\[339\]\[1\] _02272_ vdd vss _02273_ rf_ram.memory\[338\]\[1\]
+ _01687_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_input56_I vss i_ibus_rdt[30] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09906_ vdd vss _04908_ _03445_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07553__A1 vss _03389_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09542__A2 vss net41 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09837_ cpu.state.o_cnt\[2\] vdd vss _04866_ cpu.mem_bytecnt\[1\] _01385_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06356__A2 vss _01735_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09768_ _04760_ _04823_ vdd vss _04824_ net122 _04766_ _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_08719_ vdd vss _04146_ _02983_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06108__A2 vss _01543_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09699_ vdd vss _04776_ _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_68_325 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11661_ vss net184 net112 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10612_ vdd rf_ram.memory\[354\]\[0\] clknet_leaf_160_clk vss _00356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07608__A2 vss _03390_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11592_ vdd rf_ram.memory\[264\]\[1\] clknet_leaf_139_clk vss _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08805__A1 vss _04167_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10543_ vdd rf_ram.memory\[334\]\[1\] clknet_leaf_143_clk vss _00287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05619__A1 vss _01768_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_441 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05977__B vss _01503_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_417 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_474 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10474_ vdd rf_ram.memory\[423\]\[0\] clknet_leaf_103_clk vss _00218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09230__A1 vss net249 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08579__I vss _04057_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06347__A2 vss _01709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11026_ vdd rf_ram.memory\[151\]\[0\] clknet_leaf_328_clk vss _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09297__A1 vss _04466_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1080 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09049__A1 vss _04334_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06048__B vss _01615_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05380_ _01506_ vdd vss _01576_ rf_ram.memory\[550\]\[0\] _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07050_ vdd vss _03094_ _02806_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_141_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_183_clk_I vss clknet_5_29__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_299 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06001_ _01528_ vdd vss _02196_ rf_ram.memory\[512\]\[1\] _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_42_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09221__A1 vss _04431_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput114 o_dbus_dat[24] net114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_leaf_63_clk_I vss clknet_5_8__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput103 o_dbus_dat[14] net103 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput125 o_dbus_dat[5] net125 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput136 o_ext_funct3[1] net136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput158 o_ext_rs1[28] net158 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput147 o_ext_rs1[18] net147 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07783__A1 vss net237 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_198_clk_I vss clknet_5_28__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput169 o_ext_rs1[9] net169 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_leaf_78_clk_I vss clknet_5_11__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07952_ vdd vss _03656_ _02898_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05794__B1 vss _01520_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07535__A1 vss _03393_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07883_ vdd vss _03613_ _02836_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06903_ vss _02997_ _02996_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06834_ vdd vss _02950_ _02917_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_121_clk_I vss clknet_5_13__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09622_ vdd vss _04721_ rf_ram.memory\[71\]\[0\] _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09553_ _04672_ vdd vss _01074_ _04654_ _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09288__A1 vss net238 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08504_ vdd _04008_ _04006_ _00689_ _03956_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_656 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06765_ vdd vss _02901_ rf_ram.memory\[513\]\[0\] _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_511 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_136_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05716_ _01912_ vss vdd _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06696_ vdd _02852_ _02850_ _00037_ _02826_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09484_ _01387_ _03989_ vdd vss _04621_ _04620_ _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_175_341 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05647_ _01840_ _01841_ _01842_ _01670_ vdd vss _01843_ _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_93_648 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_339 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08435_ vdd vss _03959_ rf_ram.memory\[174\]\[0\] _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_16_clk_I vss clknet_5_2__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08366_ vdd vss _03915_ rf_ram.memory\[184\]\[1\] _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06510__A2 vss cpu.decode.opcode\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05578_ vss vdd rf_ram.memory\[303\]\[0\] _01773_ rf_ram.memory\[301\]\[0\] _01772_
+ _01711_ rf_ram.memory\[300\]\[0\] _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_07317_ vdd _03261_ _03258_ _00249_ _03260_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_1245 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_975 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08297_ vdd _03871_ _03869_ _00619_ _03855_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_6_661 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07248_ vdd _03217_ _03216_ _00224_ _03190_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_146 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07179_ vdd vss _03175_ _02899_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08015__A2 vss _03693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10190_ vdd vss _05084_ rf_ram.memory\[238\]\[0\] _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output162_I vss net162 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07774__A1 vss _03521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05785__B1 vss _01931_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06329__A2 vss _01515_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1140 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_69_623 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06647__I vss _02814_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_500 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_68_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11644_ vss net197 cpu.bufreg2.o_sh_done_r vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_107_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput16 vss net16 i_dbus_rdt[22] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11575_ vdd rf_ram.memory\[211\]\[0\] clknet_leaf_29_clk vss _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput27 vss net27 i_dbus_rdt[3] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10526_ vdd rf_ram.memory\[267\]\[0\] clknet_leaf_140_clk vss _00270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06265__A1 vss net252 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput38 vss net38 i_ibus_rdt[13] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput49 vss net49 i_ibus_rdt[24] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__05473__C1 vss _01668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10457_ vdd rf_ram.memory\[198\]\[1\] clknet_leaf_45_clk vss _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09203__A1 vss _04434_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10388_ vdd rf_ram.memory\[225\]\[0\] clknet_leaf_274_clk vss _00132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05726__I vss _01536_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06331__B vss _01978_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07517__A1 vss _03360_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11009_ vdd rf_ram.memory\[158\]\[1\] clknet_leaf_1_clk vss _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_17__f_clk_I vss clknet_3_4_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_987 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06550_ _02735_ vdd vss _02736_ cpu.immdec.imm11_7\[2\] _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XANTENNA__06557__I vss _02742_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05501_ vss _01697_ _01514_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06481_ _01525_ vdd vss _02676_ rf_ram.memory\[10\]\[1\] _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08493__A2 vss _03496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05432_ _01625_ rf_ram.memory\[363\]\[0\] vdd vss _01628_ rf_ram.memory\[362\]\[0\]
+ _01623_ _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_90_607 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08220_ vdd _03824_ _03821_ _00589_ _03823_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_184_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05700__B1 vss _01702_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08151_ vdd vss _03781_ _02893_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05363_ vss vdd rf_ram.memory\[543\]\[0\] _01554_ rf_ram.memory\[541\]\[0\] _01555_
+ _01538_ rf_ram.memory\[540\]\[0\] _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_113_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_77 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07102_ vdd vss _03127_ rf_ram.memory\[48\]\[1\] _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08082_ vdd _03738_ _03736_ _00537_ _03724_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05294_ _01491_ vss vdd _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_141_742 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07033_ vdd _03081_ _03079_ _00145_ _03053_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07756__A1 vss _03524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06559__A2 vss _02743_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11638__I vss net89 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06241__B vss _01916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08984_ vdd _04311_ _04310_ _00866_ _04298_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07935_ vdd vss _03645_ _02752_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05231__A2 vss net134 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07508__A1 vss _03319_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07866_ vdd vss _03603_ rf_ram.memory\[42\]\[1\] _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1194 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09605_ _04701_ cpu.immdec.imm24_20\[4\] vdd vss _04713_ _04524_ net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_3_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08181__A1 vss _03787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07797_ vdd vss _03561_ rf_ram.memory\[415\]\[0\] _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06817_ vdd vss _02938_ rf_ram.memory\[288\]\[1\] _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input19_I vss i_dbus_rdt[25] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_976 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09536_ _04660_ _04661_ vdd vss _01068_ _04653_ _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06748_ vdd vss _02888_ _02779_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_149_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09467_ _04604_ vdd vss _04610_ net83 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_164_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06679_ vdd vss _02841_ rf_ram.memory\[476\]\[0\] _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_109_717 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08418_ vdd _03947_ _03946_ _00664_ _03919_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06495__A1 vss _01371_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_478 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09398_ _04564_ net222 vdd vss _04572_ net221 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_117_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08349_ vdd vss _03905_ rf_ram.memory\[181\]\[0\] _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08236__A2 vss _02923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06416__B vss _01916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10043__A2 vss _03158_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1097 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11360_ vdd cpu.decode.op22 clknet_leaf_257_clk vss _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10311_ vdd rf_ram.memory\[515\]\[1\] clknet_leaf_271_clk vss _00055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output87_I vss net87 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11291_ vdd cpu.ctrl.pc_plus_offset_cy_r clknet_leaf_239_clk vss _00006_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07747__A1 vss _02983_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10242_ vdd vss _05115_ rf_ram.memory\[213\]\[1\] _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_661 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10173_ vdd vss _05073_ rf_ram.memory\[20\]\[0\] _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05758__B1 vss _01516_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05990__B vss _01372_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08172__A1 vss _03790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06183__B1 vss _01786_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05930__B1 vss _01857_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06722__A2 vss _02869_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_784 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_946 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_21__f_clk vdd vss clknet_5_21__leaf_clk clknet_3_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06486__A1 vss rf_ram.memory\[0\]\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08592__I vss _03902_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_832 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11627_ vss net150 net77 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09975__A2 vss _03253_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11558_ vdd rf_ram.memory\[44\]\[1\] clknet_leaf_127_clk vss _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_764 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07986__A1 vss _03651_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10509_ vdd rf_ram.memory\[255\]\[1\] clknet_leaf_217_clk vss _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_578 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11489_ vdd rf_ram.memory\[275\]\[0\] clknet_leaf_189_clk vss _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05997__B1 vss _01521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07738__A1 vss _03521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05461__A2 vss _01652_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09727__A2 vss net11 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1060 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06840__I vss _02953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06061__B vss _01658_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05456__I vss _01499_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05213__A2 vss cpu.mem_bytecnt\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07720_ vdd vss _03512_ _02971_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05981_ _02175_ _02176_ vdd vss _02177_ _02173_ _02174_ _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07671__I vss _03088_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1169 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07651_ vdd vss _03469_ net239 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07582_ vdd _03426_ _03423_ _00349_ _03425_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07910__A1 vss _02822_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06602_ vdd _02778_ _02776_ _00017_ _02748_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_935 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09321_ cpu.immdec.imm30_25\[0\] _04521_ net36 _04526_ _04529_ vss vdd cpu.immdec.imm11_7\[4\]
+ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_06533_ _02718_ vdd vss _02719_ _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_4
XANTENNA__06477__A1 vss _01903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09663__A1 vss net120 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08466__A2 vss _01364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_182 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06464_ vdd vss _02659_ rf_ram.memory\[20\]\[1\] _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_916 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09252_ vdd vss cpu.genblk3.csr.mstatus_mie _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_47_158 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05415_ rf_ram.memory\[359\]\[0\] _01608_ _01606_ rf_ram.memory\[358\]\[0\] _01611_
+ vss vdd rf_ram.memory\[357\]\[0\] _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__05685__C1 vss _01773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09183_ vdd _04435_ _04432_ _00941_ _04434_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06395_ _02586_ _02589_ vdd vss _02590_ _02578_ _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_84_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08203_ vdd _03813_ _03811_ _00583_ _03790_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_160_336 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06236__B vss _01660_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_377 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08134_ vdd vss _03771_ rf_ram.memory\[550\]\[1\] _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05346_ _01528_ vdd vss _01542_ rf_ram.memory\[512\]\[0\] _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_126_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07977__A1 vss _03654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_583 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08065_ vdd vss _03728_ rf_ram.memory\[563\]\[1\] _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05277_ vdd vss _01476_ _01381_ _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07729__A1 vss _03491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07016_ vdd _03070_ _03068_ _00139_ _03053_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05366__I vss rf_ram.i_raddr\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08967_ vdd _04300_ _04299_ _00860_ _04298_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08898_ vdd vss _04258_ rf_ram.memory\[429\]\[0\] _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07918_ vdd vss _03635_ rf_ram.memory\[45\]\[1\] _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07849_ vdd vss _03593_ rf_ram.memory\[410\]\[0\] _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_169_926 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10860_ vdd rf_ram.memory\[526\]\[0\] clknet_leaf_315_clk vss _00604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05912__B1 vss _01857_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09519_ cpu.decode.opcode\[1\] _04647_ _01399_ vss _01450_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_66_445 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_1115 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10791_ vdd rf_ram.memory\[561\]\[1\] clknet_leaf_332_clk vss _00535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_164_620 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_94_765 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_309 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08209__A2 vss _03083_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05691__A2 vss _01782_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10016__A2 vss _02984_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11412_ vdd rf_ram.memory\[187\]\[1\] clknet_leaf_18_clk vss _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11343_ vdd cpu.immdec.imm7 clknet_leaf_236_clk vss _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11274_ vdd net209 clknet_leaf_246_clk vss _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06660__I vss _02747_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1147 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10182__I vss _02742_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10225_ vdd vss _05105_ rf_ram.memory\[212\]\[0\] _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10156_ vdd _05062_ _05060_ _01288_ _05049_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10087_ vdd _05020_ _05019_ _01261_ _05014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08145__A1 vss _03757_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_734 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09893__A1 vss _04884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05903__B1 vss _01654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_70_1231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10989_ vdd rf_ram.memory\[129\]\[1\] clknet_leaf_28_clk vss _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09645__A1 vss cpu.mem_bytecnt\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06459__A1 vss rf_ram.memory\[48\]\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_949 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05200_ vdd _01400_ cpu.decode.co_mem_word vss vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_170_656 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1025 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07959__A1 vss _03651_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06180_ _02369_ _01660_ _02374_ vdd vss _02375_ _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_4_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_111_76 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08620__A2 vss _02881_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05131_ cpu.decode.op26 cpu.decode.co_ebreak vdd vss _01334_ _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__06092__C1 vss _01713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1057 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09870_ _04887_ _04400_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_110_233 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_299 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08384__A1 vss _03922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08821_ vdd vss _04211_ rf_ram.memory\[136\]\[0\] _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10191__A1 vss _05078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_174_1001 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05964_ _02159_ vdd vss _02160_ _01903_ _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08752_ vss _04167_ _04057_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__08136__A1 vss _03668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07703_ vdd vss _03502_ rf_ram.memory\[400\]\[1\] _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08683_ vdd vss _04124_ rf_ram.memory\[155\]\[0\] _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07634_ vdd vss _03459_ rf_ram.memory\[388\]\[1\] _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05895_ rf_ram.memory\[92\]\[0\] _02091_ vss vdd rf_ram.memory\[95\]\[0\] _01773_
+ rf_ram.memory\[93\]\[0\] _01772_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_07565_ vdd _03415_ _03413_ _00343_ _03393_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11651__I vss net101 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08439__A2 vss _03949_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09636__A1 vss _04524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07496_ vdd vss _03373_ rf_ram.memory\[364\]\[1\] _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09304_ vdd vss _04518_ rf_ram.memory\[63\]\[0\] _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06516_ vdd vss _02705_ cpu.bufreg.c_r _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09235_ vdd _04467_ _04464_ _00961_ _04466_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_366 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06447_ vdd vss _02642_ rf_ram.memory\[36\]\[1\] _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_286 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_483 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05673__A2 vss _01719_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09166_ vdd _04424_ _04422_ _00935_ _04401_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09939__A2 vss _02899_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06378_ _02572_ vdd vss _02573_ _01600_ _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_160_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_142_881 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_870 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09097_ vdd vss _04381_ net237 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05329_ _01525_ rf_ram.i_raddr\[2\] vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08117_ vdd _03760_ _03759_ _00550_ _03754_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07576__I vss _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08048_ vdd vss _03717_ rf_ram.memory\[566\]\[1\] _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06622__A1 vss _02750_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1288 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_778 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10010_ vdd _04972_ _04970_ _01232_ _04953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09999_ vdd vss _04966_ rf_ram.memory\[276\]\[1\] _04964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06386__B1 vss _01925_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_99_868 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10912_ vdd rf_ram.memory\[17\]\[0\] clknet_leaf_288_clk vss _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06689__A1 vss _02820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09875__A1 vss _02713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_401 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09627__A1 vss _04643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10843_ vdd rf_ram.memory\[535\]\[1\] clknet_leaf_299_clk vss _00587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10774_ vdd rf_ram.memory\[56\]\[0\] clknet_leaf_294_clk vss _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_160_clk vdd vss clknet_leaf_160_clk clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_137_686 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08850__A2 vss _04195_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06861__A1 vss _02927_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_369 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11326_ vdd cpu.bufreg.c_r clknet_leaf_255_clk vss _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06613__A1 vss _02716_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06323__C vss _01569_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11257_ vdd rf_ram.memory\[99\]\[1\] clknet_leaf_77_clk vss _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07169__A2 vss _02954_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1090 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11188_ vdd rf_ram.memory\[169\]\[0\] clknet_leaf_9_clk vss _00924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10208_ vdd _05094_ _05092_ _01308_ _05081_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_175_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10139_ vdd _05052_ _05051_ _01281_ _05046_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_1305 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_1286 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_553 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05680_ _01874_ _01875_ vdd vss _01876_ _01872_ _01873_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_187_586 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09618__A1 vss _04643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07350_ vdd _03281_ _03280_ _00262_ _03257_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_1061 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06301_ vdd vss _02496_ rf_ram.memory\[161\]\[1\] _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_151_clk vdd vss clknet_leaf_151_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_122_53 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09020_ vdd _04333_ _04332_ _00880_ _04331_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07281_ vdd vss _03239_ rf_ram.memory\[472\]\[0\] _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_442 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06232_ rf_ram.memory\[404\]\[1\] _02427_ vss vdd rf_ram.memory\[407\]\[1\] _01763_
+ rf_ram.memory\[405\]\[1\] _01668_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__05655__A2 vss _01782_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_556 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06163_ _01687_ _01696_ rf_ram.memory\[483\]\[1\] _02357_ vdd vss _02358_ rf_ram.memory\[482\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__06065__C1 vss _01664_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_339 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06604__A1 vss _02779_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06094_ _02288_ vdd vss _02289_ _01349_ _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_141_1033 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_531 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05812__C1 vss _01773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06080__A2 vss _01537_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09922_ _04918_ _04396_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08357__A1 vss _03887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10164__A1 vss _05046_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1099 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09853_ vdd vss _01171_ _02713_ _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_147_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09784_ vdd _04833_ _04831_ _01144_ _04637_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08804_ vdd vss _04200_ rf_ram.memory\[13\]\[0\] _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08109__A1 vss net247 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06996_ vdd _03058_ _03056_ _00131_ _03053_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08735_ vdd vss _03968_ _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05947_ _02142_ vdd vss _02143_ _01903_ _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09857__A1 vss _01382_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05878_ vdd _02074_ _01597_ _01368_ _02046_ vss _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_08666_ vdd _04113_ _04111_ _00746_ _04097_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07617_ vdd vss _03448_ rf_ram.memory\[313\]\[1\] _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_80 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08597_ vdd _04070_ _04068_ _00720_ _04062_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05894__A2 vss _01770_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07548_ vdd _03405_ _03404_ _00336_ _03389_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10219__A2 vss _03082_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_962 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07096__A1 vss _03092_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06408__C vss _01362_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07479_ vdd vss _03363_ rf_ram.memory\[328\]\[0\] _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_142_clk vdd vss clknet_leaf_142_clk clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10490_ vdd rf_ram.memory\[417\]\[0\] clknet_leaf_95_clk vss _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06843__A1 vss _02927_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output192_I vss net192 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_859 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09218_ vdd _04456_ _04454_ _00955_ _04434_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05646__A2 vss _01500_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1219 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_155 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09149_ vdd vss _04414_ rf_ram.memory\[8\]\[1\] _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06424__B vss _02004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11111_ vdd rf_ram.memory\[123\]\[1\] clknet_leaf_86_clk vss _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08348__A1 vss _03071_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11042_ vdd rf_ram.memory\[146\]\[0\] clknet_leaf_336_clk vss _00779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08899__A2 vss _04257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07571__A2 vss _02960_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_676 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_553 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07323__A2 vss _02909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10826_ vdd rf_ram.memory\[543\]\[0\] clknet_leaf_312_clk vss _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_729 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10757_ vdd rf_ram.memory\[478\]\[1\] clknet_leaf_123_clk vss _00501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_133_clk vdd vss clknet_leaf_133_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07087__A1 vss _02775_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_420 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10688_ vdd rf_ram.memory\[435\]\[0\] clknet_leaf_81_clk vss _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06834__A1 vss _02917_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05637__A2 vss _01631_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1033 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_1142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_1006 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05729__I vss _01695_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1103 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08587__A1 vss _02828_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1039 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06062__A2 vss _01662_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09645__B vss _01375_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11309_ _01042_ vdd vss clknet_leaf_266_clk net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__10146__A1 vss _05049_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06850_ vdd vss _02962_ rf_ram.memory\[285\]\[0\] _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07011__A1 vss _03053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05464__I vss _01599_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05801_ vdd vss _01997_ rf_ram.memory\[169\]\[0\] _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06781_ vdd vss _02913_ rf_ram.memory\[511\]\[0\] _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08520_ vdd vss _04021_ rf_ram.memory\[188\]\[0\] _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05732_ _01928_ _01563_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05663_ _01857_ rf_ram.memory\[475\]\[0\] vdd vss _01859_ rf_ram.memory\[474\]\[0\]
+ _01856_ _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08451_ vdd vss _00676_ _02714_ _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08511__A1 vss _03989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07402_ vdd vss _03314_ rf_ram.memory\[247\]\[0\] _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05594_ _01790_ _01493_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08382_ vdd _03925_ _03924_ _00650_ _03919_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_124_clk vdd vss clknet_leaf_124_clk clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07333_ vdd vss _03271_ _03055_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_543 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_483 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07264_ vdd vss _03228_ rf_ram.memory\[196\]\[0\] _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_960 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1242 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06215_ _01778_ rf_ram.memory\[395\]\[1\] vdd vss _02410_ rf_ram.memory\[394\]\[1\]
+ _01777_ _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_131_615 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09003_ vdd vss _04323_ rf_ram.memory\[111\]\[0\] _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06244__B vss _01790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07195_ vdd vss _03185_ rf_ram.memory\[474\]\[0\] _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06146_ rf_ram.memory\[316\]\[1\] _02341_ vss vdd rf_ram.memory\[319\]\[1\] _01726_
+ rf_ram.memory\[317\]\[1\] _01725_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__07250__A1 vss _03193_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06053__A2 vss _01644_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06077_ vdd vss _02272_ rf_ram.memory\[337\]\[1\] _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09555__B vss _04526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09905_ vdd _04907_ _04905_ _01192_ _04887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10137__A1 vss _02794_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input49_I vss i_ibus_rdt[24] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05800__A2 vss _01510_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07002__A1 vss _03055_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09836_ vdd _04865_ _04863_ _01164_ _04840_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06979_ vdd vss _03047_ _02775_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09767_ vdd vss _04823_ _04804_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09698_ _04768_ _04775_ vdd vss _04776_ net129 _04767_ net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_08718_ vdd _04145_ _04143_ _00766_ _04129_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08502__A1 vss _03953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_2__f_clk vdd vss clknet_5_2__leaf_clk clknet_3_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08649_ vdd _04103_ _04102_ _00739_ _04094_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06419__B vss _01928_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1090 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_304_clk_I vss clknet_5_4__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11660_ net183 vss vdd net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05867__A2 vss _01634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10611_ vdd rf_ram.memory\[315\]\[1\] clknet_leaf_105_clk vss _00355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_589 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_115_clk vdd vss clknet_leaf_115_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11591_ vdd rf_ram.memory\[264\]\[0\] clknet_leaf_139_clk vss _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07069__A1 vss _03087_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10542_ vdd rf_ram.memory\[334\]\[0\] clknet_leaf_143_clk vss _00286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_146_280 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06816__A1 vss _02927_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06933__I vss _03017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_924 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06292__A2 vss _01922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_319_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1147 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10473_ vdd rf_ram.memory\[424\]\[1\] clknet_leaf_104_clk vss _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06029__C1 vss _01554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09230__A2 vss _02815_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_613 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07241__A1 vss _02795_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06044__A2 vss _01614_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_681 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11025_ vdd rf_ram.memory\[152\]\[1\] clknet_leaf_328_clk vss _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_832 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_258 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_329 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_724 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05858__A2 vss _01846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_106_clk vdd vss clknet_leaf_106_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_126_921 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10809_ vdd rf_ram.memory\[552\]\[1\] clknet_leaf_320_clk vss _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06807__A1 vss _02930_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_874 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07480__A1 vss _03356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06064__B vss _01526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06283__A2 vss _01531_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05459__I vss _01513_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06000_ rf_ram.memory\[517\]\[1\] _01539_ _01538_ rf_ram.memory\[516\]\[1\] _02195_
+ vss vdd rf_ram.memory\[519\]\[1\] _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_24_974 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput104 o_dbus_dat[15] net104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput115 o_dbus_dat[25] net115 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_10_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_782 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput137 o_ext_funct3[2] net137 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput126 o_dbus_dat[6] net126 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput159 o_ext_rs1[29] net159 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput148 o_ext_rs1[19] net148 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06035__A2 vss _01524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07783__A2 vss _03234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07951_ vdd _03655_ _03652_ _00489_ _03654_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10119__A1 vss _05017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1167 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06902_ vdd vss _02996_ _02867_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07882_ vdd _03612_ _03610_ _00463_ _03590_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06833_ vdd _02949_ _02947_ _00077_ _02930_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09621_ vdd vss _04720_ _02828_ _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08732__A1 vss _04126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09552_ net44 _04650_ cpu.immdec.imm19_12_20\[8\] vdd vss _04672_ _04478_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06764_ vdd vss _02900_ _02881_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07299__A1 vss _03225_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09288__A2 vss _04507_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08503_ vdd vss _04008_ rf_ram.memory\[79\]\[1\] _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05715_ _01911_ _01695_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_77_123 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06695_ vdd vss _02852_ rf_ram.memory\[524\]\[1\] _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09483_ vdd vss cpu.state.cnt_r\[1\] _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05646_ rf_ram.memory\[498\]\[0\] _01842_ vss vdd rf_ram.memory\[497\]\[0\] _01668_
+ rf_ram.memory\[499\]\[0\] _01763_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_08434_ vdd vss _03958_ _02971_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05143__B vss _01341_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05577_ _01773_ _01695_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08365_ vdd _03914_ _03913_ _00644_ _03884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06259__C1 vss _01646_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07316_ vdd vss _03261_ rf_ram.memory\[256\]\[1\] _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08454__B vss net126 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_727 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08296_ vdd vss _03871_ rf_ram.memory\[203\]\[1\] _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_290_clk_I vss clknet_5_24__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_546 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07247_ vdd vss _03217_ rf_ram.memory\[420\]\[0\] _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_581 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07471__A1 vss _02972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1061 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07178_ vdd _03174_ _03172_ _00197_ _03161_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_44_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07223__A1 vss _03190_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06129_ vdd vss _02324_ rf_ram.memory\[297\]\[1\] _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_121_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output155_I vss net155 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09819_ vdd _04855_ _04854_ _01157_ _04837_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08723__A1 vss _04129_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06928__I vss _03013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_692 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_243_clk_I vss clknet_5_21__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_336_clk vdd vss clknet_leaf_336_clk clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11643_ vss net196 net124 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_182_868 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_671 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_811 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_362 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_258_clk_I vss clknet_5_17__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput17 vss net17 i_dbus_rdt[23] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11574_ vdd rf_ram.memory\[191\]\[1\] clknet_leaf_27_clk vss _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput28 vss net28 i_dbus_rdt[4] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10525_ vdd rf_ram.memory\[251\]\[1\] clknet_leaf_215_clk vss _00269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput39 vss net39 i_ibus_rdt[14] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__05473__B1 vss _01519_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10456_ vdd rf_ram.memory\[198\]\[0\] clknet_leaf_44_clk vss _00200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_1144 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06017__A2 vss _01502_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_421 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10387_ vdd rf_ram.memory\[226\]\[1\] clknet_leaf_272_clk vss _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11008_ vdd rf_ram.memory\[158\]\[0\] clknet_leaf_1_clk vss _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08714__A1 vss _03008_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06059__B vss _01650_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_327_clk vdd vss clknet_leaf_327_clk clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06480_ rf_ram.memory\[12\]\[1\] _02675_ vss vdd rf_ram.memory\[15\]\[1\] _01653_
+ rf_ram.memory\[13\]\[1\] _01655_ _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_05500_ _01696_ _01695_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_05431_ vdd vss _01627_ rf_ram.memory\[361\]\[0\] _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_135_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_65 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_510 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_228 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08150_ vdd _03780_ _03778_ _00563_ _03757_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07101_ vss _03126_ _03017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_55_373 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_587 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05362_ _01505_ vdd vss _01558_ rf_ram.memory\[542\]\[0\] _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06256__A2 vss _01666_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07453__A1 vss _03326_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_795 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05293_ vdd _01490_ _01489_ _01430_ _01487_ vss _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_08081_ vdd vss _03738_ rf_ram.memory\[560\]\[1\] _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07032_ vdd vss _03081_ rf_ram.memory\[216\]\[1\] _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_30_218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05189__I vss cpu.ctrl.pc vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_776 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07205__A1 vss _02806_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_955 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_933 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06008__A2 vss _01501_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08953__A1 vss _04269_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_454 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08983_ vdd vss _04311_ rf_ram.memory\[115\]\[0\] _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07934_ vdd _03644_ _03642_ _00483_ _03622_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07508__A2 vss _02889_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07865_ vdd _03602_ _03601_ _00456_ _03587_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11654__I vss net104 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09604_ _04700_ vdd vss _04712_ _04478_ cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07796_ vdd vss _03560_ _02908_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06816_ vdd _02937_ _02936_ _00072_ _02927_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05652__I vss _01617_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09535_ vdd vss _04661_ cpu.immdec.imm19_12_20\[2\] _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_318_clk vdd vss clknet_leaf_318_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06747_ vdd vss _02887_ _02719_ _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06678_ vdd vss _02840_ _02836_ _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09130__A1 vss _04401_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09466_ vss _01050_ _04609_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05629_ _01693_ vdd vss _01825_ rf_ram.memory\[480\]\[0\] _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_93_446 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08417_ vdd vss _03947_ rf_ram.memory\[29\]\[0\] _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06495__A2 vss _02235_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_857 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_74_660 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09397_ vdd vss _04571_ _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05601__B vss _01707_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08348_ vdd vss _03904_ _03071_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_693 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_395 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07444__A1 vss _02781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1178 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06247__A2 vss _01719_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ vdd vss _03861_ rf_ram.memory\[194\]\[0\] _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_220 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10310_ vdd rf_ram.memory\[515\]\[0\] clknet_leaf_272_clk vss _00054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11290_ vdd cpu.ctrl.pc_plus_4_cy_r clknet_leaf_242_clk vss _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10241_ vdd _05114_ _05113_ _01321_ _02819_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07747__A2 vss _03496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08944__A1 vss _03672_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1020 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10172_ vdd vss _05072_ _02996_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06151__C vss net253 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_1161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_9__f_clk_I vss clknet_3_2_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_182_clk_I vss clknet_5_29__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_62_clk_I vss clknet_5_8__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_903 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_309_clk vdd vss clknet_leaf_309_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_9_1066 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09121__A1 vss _04367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_197_clk_I vss clknet_5_28__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07683__A1 vss _02908_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1193 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06486__A2 vss _01613_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_77_clk_I vss clknet_5_8__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11626_ vss net148 net76 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_167_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_378 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06238__A2 vss _01510_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_120_clk_I vss clknet_5_13__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11557_ vdd rf_ram.memory\[44\]\[0\] clknet_leaf_129_clk vss _01289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_546 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10508_ vdd rf_ram.memory\[255\]\[0\] clknet_leaf_219_clk vss _00252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_719 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11488_ vdd rf_ram.memory\[274\]\[1\] clknet_leaf_181_clk vss _01220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09188__A1 vss _04434_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10439_ vdd rf_ram.memory\[498\]\[1\] clknet_leaf_222_clk vss _00183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_135_clk_I vss clknet_5_24__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06410__A2 vss _01856_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05980_ rf_ram.memory\[9\]\[0\] _01714_ _01643_ rf_ram.memory\[8\]\[0\] _02176_ vss
+ vdd rf_ram.memory\[11\]\[0\] _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__05213__A3 vss _01385_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_15_clk_I vss clknet_5_2__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07650_ vdd _03468_ _03466_ _00375_ _03458_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05472__I vss _01655_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06568__I vss _02751_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07581_ vdd vss _03426_ rf_ram.memory\[356\]\[1\] _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07910__A2 vss _03547_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_730 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06601_ vdd vss _02778_ rf_ram.memory\[234\]\[1\] _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_149_128 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_86 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09112__A1 vss _02959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06532_ vdd vss _02718_ _01497_ _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_09320_ vdd vss _04528_ _00985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09251_ vdd vss _00965_ _04476_ _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08466__A3 vss _02709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07674__A1 vss _03455_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06463_ _02657_ _01568_ vdd vss _02658_ _01599_ _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_7_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08202_ vdd vss _03813_ rf_ram.memory\[537\]\[1\] _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05685__B1 vss _01772_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09182_ vdd vss _04435_ rf_ram.memory\[84\]\[1\] _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06394_ _02588_ vdd vss _02589_ _01972_ _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_05414_ _01610_ _01609_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06229__A2 vss _01801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07426__A1 vss _03323_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08133_ vdd _03770_ _03769_ _00556_ _03754_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05345_ rf_ram.memory\[517\]\[0\] _01539_ _01538_ rf_ram.memory\[516\]\[0\] _01541_
+ vss vdd rf_ram.memory\[519\]\[0\] _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_44_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_941 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08064_ vdd _03727_ _03726_ _00530_ _03721_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05988__A1 vss _01349_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11649__I vss net99 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07015_ vdd vss _03070_ rf_ram.memory\[222\]\[1\] _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05276_ _01449_ _01451_ vdd vss _01475_ _01383_ _01427_ _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_101_415 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08926__A1 vss _04266_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05204__A3 vss _01341_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08966_ vdd vss _04300_ rf_ram.memory\[118\]\[0\] _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input31_I vss i_dbus_rdt[7] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_95_clk vdd vss clknet_leaf_95_clk clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08897_ vdd vss _04257_ net243 _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07917_ vdd _03634_ _03633_ _00476_ _03619_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07848_ vdd vss _03592_ _02813_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_151_1002 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output118_I vss net118 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07779_ vdd vss _03549_ rf_ram.memory\[437\]\[0\] _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_763 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09518_ vdd vss cpu.immdec.imm19_12_20\[0\] _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_91_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xserv_rf_top_255 o_dbus_adr[0] vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_66_424 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10790_ vdd rf_ram.memory\[561\]\[0\] clknet_leaf_332_clk vss _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07665__A1 vss _03458_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06468__A2 vss _01514_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09449_ vss _01042_ _04600_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_163_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_136_367 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09406__A2 vss _03991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11411_ vdd rf_ram.memory\[187\]\[0\] clknet_leaf_18_clk vss _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11342_ vdd cpu.immdec.imm19_12_20\[8\] clknet_leaf_216_clk vss _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_105_765 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05979__A1 vss rf_ram.memory\[10\]\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08090__A1 vss _03721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_858 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11273_ vdd net208 clknet_leaf_246_clk vss _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09029__I vss _04037_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10224_ vdd vss _05104_ _03892_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10155_ vdd vss _05062_ rf_ram.memory\[450\]\[1\] _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_86_clk vdd vss clknet_leaf_86_clk clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10086_ vdd vss _05020_ rf_ram.memory\[30\]\[0\] _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06156__A1 vss _01675_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1092 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09342__B2 vss net224 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09342__A1 vss net213 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_582 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_755 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10988_ vdd rf_ram.memory\[129\]\[0\] clknet_leaf_27_clk vss _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09645__A2 vss _01376_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07656__A1 vss _03088_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06459__A2 vss _01643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_507 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_613 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07408__A1 vss _03289_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11609_ net160 vss vdd net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_108_581 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_10_clk vdd vss clknet_leaf_10_clk clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_26_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05130_ vdd vss cpu.decode.op21 _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_123_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06092__B1 vss _01721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06072__B vss _01615_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_584 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_410 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_180_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08820_ vdd vss _04210_ net250 _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09581__A1 vss _03992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07682__I vss _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_77_clk vdd vss clknet_leaf_77_clk clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05963_ rf_ram.memory\[23\]\[0\] _01624_ _01605_ rf_ram.memory\[22\]\[0\] _02159_
+ vss vdd rf_ram.memory\[21\]\[0\] _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08751_ vdd _04166_ _04164_ _00778_ _04129_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07702_ vdd _03501_ _03500_ _00394_ _03488_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09333__A1 vss net240 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05894_ vdd vss _02090_ rf_ram.memory\[94\]\[0\] _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08136__A2 vss _03009_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08682_ vdd vss _04123_ _02821_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07633_ _03458_ vss vdd _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_136_96 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_508 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07564_ vdd vss _03415_ rf_ram.memory\[318\]\[1\] _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07495_ vdd _03372_ _03371_ _00316_ _03356_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09303_ vdd vss _04517_ _03668_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06515_ vdd vss _02704_ cpu.alu.i_rs1 _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09234_ vdd vss _04467_ rf_ram.memory\[329\]\[1\] _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_118_334 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06446_ _01493_ vdd vss _02641_ _02638_ _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_63_438 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_833 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09165_ vdd vss _04424_ rf_ram.memory\[87\]\[1\] _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_185_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06377_ _02570_ _02571_ vdd vss _02572_ _02568_ _02569_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08116_ vdd vss _03760_ rf_ram.memory\[553\]\[0\] _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09096_ vdd _04380_ _04378_ _00909_ _04367_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_9_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08072__A1 vss _03724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05328_ vss _01524_ _01523_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_05259_ _01456_ _01173_ vdd vss _01458_ _01380_ _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08047_ vdd _03716_ _03715_ _00524_ _03686_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09998_ vdd _04965_ _04964_ _01227_ _04950_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08949_ vdd vss _04289_ _02983_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06138__A1 vss _01675_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_68_clk vdd vss clknet_leaf_68_clk clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_169_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10911_ vdd rf_ram.memory\[199\]\[1\] clknet_leaf_39_clk vss _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10842_ vdd rf_ram.memory\[535\]\[0\] clknet_leaf_298_clk vss _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07638__A1 vss _03455_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10773_ vdd rf_ram.memory\[570\]\[1\] clknet_leaf_305_clk vss _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06157__B vss _01684_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06310__A1 vss _01552_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05996__B vss _01528_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_551 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07810__A1 vss _03557_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06074__B1 vss _01688_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11325_ vdd cpu.state.i_ctrl_misalign clknet_leaf_249_clk vss _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11256_ vdd rf_ram.memory\[99\]\[0\] clknet_leaf_77_clk vss _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11187_ vdd rf_ram.memory\[91\]\[1\] clknet_leaf_57_clk vss _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10207_ vdd vss _05094_ rf_ram.memory\[211\]\[1\] _05092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10138_ vdd vss _05052_ rf_ram.memory\[453\]\[0\] _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_59_clk vdd vss clknet_leaf_59_clk clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10069_ vdd vss _05009_ rf_ram.memory\[508\]\[0\] _05008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_187_510 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_82_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_543 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07877__A1 vss _03590_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05337__C1 vss _01517_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05888__B1 vss _02019_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05352__A2 vss _01532_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09618__A2 vss _01460_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06067__B vss _01599_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_952 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07280_ vdd vss _03238_ _02836_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06300_ _01956_ vdd vss _02495_ rf_ram.memory\[160\]\[1\] _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06231_ _01504_ vdd vss _02426_ rf_ram.memory\[406\]\[1\] _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_142_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06162_ vdd vss _02357_ rf_ram.memory\[481\]\[1\] _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08054__A1 vss _03690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_487 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06065__B1 vss _01519_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06093_ _02286_ _02287_ vdd vss _02288_ _02284_ _02285_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07801__A1 vss _02866_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09921_ vdd _04917_ _04915_ _01198_ _04887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_145_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05812__B1 vss _01848_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_240 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09852_ vdd vss _04875_ _01385_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09783_ vdd vss _04833_ rf_ram.memory\[187\]\[1\] _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08803_ vdd vss _04199_ net243 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08109__A2 vss _03729_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06995_ vdd vss _03058_ rf_ram.memory\[226\]\[1\] _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08734_ vdd _04155_ _04153_ _00772_ _04129_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05946_ rf_ram.memory\[39\]\[0\] _01607_ _01661_ rf_ram.memory\[38\]\[0\] _02142_
+ vss vdd rf_ram.memory\[37\]\[0\] _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_22_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07868__A1 vss _02991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05877_ _02072_ _01569_ vdd vss _02073_ _01768_ _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08665_ vdd vss _04113_ rf_ram.memory\[158\]\[1\] _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07616_ vdd _03447_ _03446_ _00362_ _03422_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_163_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05660__I vss _01686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08596_ vdd vss _04070_ rf_ram.memory\[166\]\[1\] _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06756__I vss _02893_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07547_ vdd vss _03405_ rf_ram.memory\[35\]\[0\] _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_181_719 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_119_643 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_585 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07478_ vdd vss _03362_ _02728_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08971__I vss _04037_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08293__A1 vss _03230_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1119 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_646 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09217_ vdd vss _04456_ rf_ram.memory\[67\]\[1\] _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06429_ _02004_ vdd vss _02624_ rf_ram.memory\[102\]\[1\] _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_output185_I vss net185 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09148_ vdd _04413_ _04412_ _00928_ _04397_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_791 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08045__A1 vss _03008_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09793__A1 vss _04837_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09079_ vdd _04370_ _04369_ _00902_ _04364_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11110_ vdd rf_ram.memory\[123\]\[0\] clknet_leaf_86_clk vss _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_688 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08348__A2 vss _03903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11041_ vdd rf_ram.memory\[147\]\[1\] clknet_leaf_337_clk vss _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_644 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09848__A2 vss _01413_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1058 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10825_ vdd rf_ram.memory\[544\]\[1\] clknet_leaf_314_clk vss _00569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_259 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10756_ vdd rf_ram.memory\[478\]\[0\] clknet_leaf_123_clk vss _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07087__A2 vss _02911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_213 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10687_ vdd rf_ram.memory\[415\]\[1\] clknet_leaf_90_clk vss _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_933 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_432 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06834__A2 vss _02941_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_616 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09784__A1 vss _04637_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08587__A2 vss _03949_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_964 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_688 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06598__A1 vss _02766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09645__C vss _01385_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11308_ _01041_ vdd vss clknet_leaf_265_clk net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11239_ vdd rf_ram.memory\[65\]\[1\] clknet_leaf_60_clk vss _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05800_ _01527_ vdd vss _01996_ rf_ram.memory\[168\]\[0\] _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06780_ vdd vss _02912_ _02909_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09839__A2 vss _03984_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05731_ _01925_ rf_ram.memory\[443\]\[0\] vdd vss _01927_ rf_ram.memory\[442\]\[0\]
+ _01719_ _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_188_852 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05662_ vdd vss _01858_ rf_ram.memory\[473\]\[0\] _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_72_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08450_ _03967_ vdd vss _03968_ cpu.state.genblk1.misalign_trap_sync_r cpu.state.stage_two_req
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08381_ vdd vss _03925_ rf_ram.memory\[180\]\[0\] _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07401_ vdd vss _03313_ _03309_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06522__B2 vss _01375_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_708 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05593_ _01786_ rf_ram.memory\[291\]\[0\] vdd vss _01789_ rf_ram.memory\[290\]\[0\]
+ _01785_ _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_129_963 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_440 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07332_ vdd _03270_ _03268_ _00255_ _03260_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08275__A1 vss _03852_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07263_ vdd vss _03227_ _02738_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_972 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06214_ vdd vss _02409_ rf_ram.memory\[393\]\[1\] _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09002_ vdd vss _04322_ _02953_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07194_ vdd vss _03184_ _02813_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08027__A1 vss _03686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06145_ _01805_ vdd vss _02340_ rf_ram.memory\[318\]\[1\] _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_108_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09775__A1 vss net243 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06589__A1 vss _02748_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06076_ _01684_ vdd vss _02271_ rf_ram.memory\[336\]\[1\] _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_44_1259 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09904_ vdd vss _04907_ rf_ram.memory\[345\]\[1\] _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11657__I vss net107 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06260__B vss _01756_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10137__A2 vss _02836_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09127__I vss _02747_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09835_ vdd vss _04865_ rf_ram.memory\[61\]\[1\] _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07002__A2 vss _02904_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06978_ vdd _03046_ _03044_ _00125_ _03018_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05564__A2 vss _01662_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09766_ vdd vss _04822_ _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06761__A1 vss _02876_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05929_ _01923_ vdd vss _02125_ rf_ram.memory\[96\]\[0\] _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_1202 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09697_ vdd vss _04775_ _04740_ net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08717_ vdd vss _04145_ rf_ram.memory\[150\]\[1\] _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05604__B vss _01602_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08648_ vdd vss _04103_ rf_ram.memory\[161\]\[0\] _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_658 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_146 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06513__A1 vss _01391_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_395 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_360 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08579_ _04058_ _04057_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_10610_ vdd rf_ram.memory\[315\]\[0\] clknet_leaf_105_clk vss _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11590_ vdd rf_ram.memory\[213\]\[1\] clknet_leaf_303_clk vss _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10073__A1 vss _03445_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10541_ vdd rf_ram.memory\[372\]\[1\] clknet_leaf_146_clk vss _00285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_693 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06277__B1 vss _01953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06435__B vss net251 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_1006 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10472_ vdd rf_ram.memory\[424\]\[0\] clknet_leaf_104_clk vss _00216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06029__B1 vss _01555_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_986 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07241__A2 vss _03040_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1040 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05788__C1 vss _01702_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11024_ vdd rf_ram.memory\[152\]\[0\] clknet_leaf_327_clk vss _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_99_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06752__A1 vss _02873_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08741__A2 vss _04158_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_614 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_103_34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10808_ vdd rf_ram.memory\[552\]\[0\] clknet_leaf_321_clk vss _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_909 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10739_ vdd rf_ram.memory\[440\]\[1\] clknet_leaf_55_clk vss _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_341 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_1185 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_454 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06345__B vss _01860_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput105 o_dbus_dat[16] net105 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput116 o_dbus_dat[26] net116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput127 o_dbus_dat[7] net127 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_23_496 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput149 o_ext_rs1[1] net149 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput138 o_ext_rs1[0] net138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09509__A1 vss _04634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07950_ vdd vss _03655_ rf_ram.memory\[456\]\[1\] _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_290_clk vdd vss clknet_leaf_290_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05243__A1 vss cpu.alu.i_rs1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06901_ vdd _02995_ _02993_ _00099_ _02975_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05794__A2 vss _01989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07881_ vdd vss _03612_ rf_ram.memory\[446\]\[1\] _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_53 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06832_ vdd vss _02949_ rf_ram.memory\[304\]\[1\] _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09620_ vdd _04651_ _01393_ _01094_ _04643_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09551_ _04670_ vdd vss _04671_ _01391_ cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06763_ _02899_ vss vdd _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05714_ vdd vss _01910_ rf_ram.memory\[436\]\[0\] _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08502_ vdd _04007_ _04006_ _00688_ _03953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_682 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06694_ vdd _02851_ _02850_ _00036_ _02820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09482_ vss _01056_ _04619_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_188_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05703__C1 vss _01721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05645_ _01526_ vdd vss _01841_ rf_ram.memory\[496\]\[0\] _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08433_ vdd _03957_ _03954_ _00669_ _03956_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_894 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_714 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_505 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05576_ _01772_ _01617_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08364_ vdd vss _03914_ rf_ram.memory\[184\]\[0\] _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08248__A1 vss _03820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06259__B1 vss _01810_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10055__A1 vss _04982_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07315_ _03260_ _03017_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_73_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06255__B vss _01650_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_292 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08295_ vdd _03870_ _03869_ _00618_ _03852_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_61_514 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07246_ vdd vss _03216_ _02882_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07471__A2 vss _03101_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_413 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07177_ vdd vss _03174_ rf_ram.memory\[482\]\[1\] _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_15_975 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06128_ _01693_ vdd vss _02323_ rf_ram.memory\[296\]\[1\] _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08420__A1 vss _03922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input61_I vss i_ibus_rdt[6] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06059_ _01650_ vdd vss _02254_ rf_ram.memory\[376\]\[1\] _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_80 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_281_clk vdd vss clknet_leaf_281_clk clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_100_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05785__A2 vss _01799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09818_ vdd vss _04855_ rf_ram.memory\[259\]\[0\] _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05537__A2 vss _01367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06734__A1 vss _02795_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09749_ vdd vss _04811_ _04804_ net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__08487__A1 vss _03956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06149__C vss _01658_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05988__C vss net254 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05170__B1 vss _01367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11642_ vss net195 net123 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_37_544 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput18 vss net18 i_dbus_rdt[24] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11573_ vdd rf_ram.memory\[191\]\[0\] clknet_leaf_27_clk vss _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_182 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10524_ vdd rf_ram.memory\[251\]\[0\] clknet_leaf_215_clk vss _00268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput29 vss net29 i_dbus_rdt[5] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_122_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10455_ vdd rf_ram.memory\[1\]\[1\] clknet_leaf_39_clk vss _00199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_799 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_794 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_272_clk vdd vss clknet_leaf_272_clk clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10386_ vdd rf_ram.memory\[226\]\[0\] clknet_leaf_277_clk vss _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06973__A1 vss _03018_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11007_ vdd rf_ram.memory\[15\]\[1\] clknet_leaf_295_clk vss _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08714__A2 vss _04078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_90_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07150__A1 vss _03126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_685 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05430_ _01626_ vss vdd _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__05700__A2 vss _01634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10037__A1 vss _04985_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_538 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_864 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05361_ _01553_ _01556_ vdd vss _01557_ _01548_ _01549_ _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA_clkbuf_5_26__f_clk_I vss clknet_3_6_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06075__B vss _01629_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07100_ vdd _03125_ _03124_ _00168_ _03123_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05292_ vdd vss _01489_ cpu.alu.i_rs1 cpu.alu.add_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08080_ vdd _03737_ _03736_ _00536_ _03721_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_183_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07031_ vdd _03080_ _03079_ _00144_ _03050_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07205__A2 vss _02941_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08402__A1 vss _03919_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_260 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_23_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09450__I0 vss net75 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_263_clk vdd vss clknet_leaf_263_clk clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_41_1218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05216__A1 vss _01413_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08982_ vdd vss _04310_ net242 _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06964__A1 vss _03014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_303_clk_I vss clknet_5_6__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05767__A2 vss _01846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07933_ vdd vss _03644_ rf_ram.memory\[440\]\[1\] _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_177_1044 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07864_ vdd vss _03602_ rf_ram.memory\[42\]\[0\] _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06815_ vdd vss _02937_ rf_ram.memory\[288\]\[0\] _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09603_ _04710_ _04711_ vdd vss _01085_ _04643_ _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__06716__A1 vss _02826_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07795_ vss _03559_ _03088_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_97_219 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_318_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09534_ vdd vss _04660_ _04526_ net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06746_ vdd _02886_ _02884_ _00053_ _02876_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08469__A1 vss _02714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07141__A1 vss _02795_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09465_ _04604_ vdd vss _04609_ net82 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06677_ _02839_ _02838_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_171_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_164_825 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05628_ _01746_ vdd vss _01824_ _01821_ _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08416_ vdd vss _03946_ _02959_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09969__A1 vss _03672_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09396_ _04564_ net221 vdd vss _04571_ net220 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_05559_ _01755_ vss vdd _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08347_ _03903_ vss vdd _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_11_1044 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07444__A2 vss _02815_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08278_ vdd vss _03860_ _03230_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08641__A1 vss _04097_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07229_ vdd vss _03206_ rf_ram.memory\[424\]\[1\] _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_446 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_15_750 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_254 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10240_ vdd vss _05114_ rf_ram.memory\[213\]\[0\] _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_254_clk vdd vss clknet_leaf_254_clk clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08944__A2 vss _02899_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10171_ vdd _05071_ _05069_ _01294_ _05049_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05758__A2 vss _01614_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06955__A1 vss _03018_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06707__A1 vss _02752_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07380__A1 vss _02775_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06183__A2 vss _01785_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_400 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11135__CLK vss clknet_5_10__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05930__A2 vss _01785_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05999__B vss _01506_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_127 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_831 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07683__A2 vss _03390_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11625_ vss net147 net75 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11556_ vdd rf_ram.memory\[450\]\[1\] clknet_leaf_112_clk vss _01288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08632__A1 vss _04058_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_582 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10507_ vdd rf_ram.memory\[272\]\[1\] clknet_leaf_190_clk vss _00251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11487_ vdd rf_ram.memory\[274\]\[0\] clknet_leaf_183_clk vss _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05997__A2 vss _01532_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07199__A1 vss _02761_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_427 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_79 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10438_ vdd rf_ram.memory\[498\]\[0\] clknet_leaf_222_clk vss _00182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_614 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05749__A2 vss _01942_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10369_ vdd rf_ram.memory\[206\]\[1\] clknet_leaf_38_clk vss _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_245_clk vdd vss clknet_leaf_245_clk clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06946__A1 vss _02728_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1284 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08699__A1 vss _02828_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_939 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07580_ vss _03425_ _03359_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06600_ vdd _02777_ _02776_ _00016_ _02743_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09112__A2 vss _04005_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10258__A1 vss _02825_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06531_ vdd vss _02717_ _01498_ _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05702__B vss _01615_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07123__A1 vss _03123_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09250_ vdd vss _04479_ _04478_ cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_173_611 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06462_ _01599_ _02656_ vdd vss _02657_ _02648_ _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__08871__A1 vss _04237_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08201_ vdd _03812_ _03811_ _00582_ _03787_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_133_508 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09181_ _04434_ _04400_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05413_ _01609_ vss vdd _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06393_ rf_ram.memory\[71\]\[1\] _01925_ _01719_ rf_ram.memory\[70\]\[1\] _02588_
+ vss vdd rf_ram.memory\[69\]\[1\] _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08132_ vdd vss _03770_ rf_ram.memory\[550\]\[0\] _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05344_ _01540_ vss vdd _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08063_ vdd vss _03727_ rf_ram.memory\[563\]\[0\] _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05275_ _01473_ vdd vss _01474_ _01458_ _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_144_1043 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_141_541 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_917 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07014_ vdd _03069_ _03068_ _00138_ _03050_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_720 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1076 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_242_clk_I vss clknet_5_21__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_961 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_236_clk vdd vss clknet_leaf_236_clk clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08965_ vdd vss _04299_ _03008_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_52_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07916_ vdd vss _03634_ rf_ram.memory\[45\]\[0\] _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11665__I vss net116 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08896_ vdd _04256_ _04254_ _00833_ _04237_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input24_I vss i_dbus_rdt[2] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_257_clk_I vss clknet_5_20__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07847_ vdd _03591_ _03588_ _00449_ _03590_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07362__A1 vss _03260_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06165__A2 vss _01735_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07778_ vdd vss _03548_ _03547_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05912__A2 vss _01856_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10249__A1 vss _02838_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_701 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09517_ vdd _04645_ _04644_ _01065_ _04643_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06729_ vdd vss _02875_ rf_ram.memory\[518\]\[0\] _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xserv_rf_top_256 o_dbus_adr[1] vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_67_959 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07114__A1 vss _02716_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09448_ _04593_ vdd vss _04600_ net74 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_549 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09379_ _04552_ net212 vdd vss _04562_ net211 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_19_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_160 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_699 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_519 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11410_ vdd rf_ram.memory\[77\]\[1\] clknet_leaf_20_clk vss _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08614__A1 vss _04062_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_675 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11341_ vdd cpu.immdec.imm19_12_20\[7\] clknet_leaf_216_clk vss _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_366 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_377 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06443__B vss _01601_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05979__A2 vss _01686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_697 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11272_ vdd net207 clknet_leaf_246_clk vss _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10223_ vdd _05103_ _05101_ _01314_ _05081_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_227_clk vdd vss clknet_leaf_227_clk clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10154_ vdd _05061_ _05060_ _01287_ _05046_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05573__I vss _01650_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10085_ vdd vss _05019_ _02916_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07353__A1 vss _03055_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09342__A2 vss _03991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05903__A2 vss _01652_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_414 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10987_ vdd rf_ram.memory\[164\]\[1\] clknet_leaf_330_clk vss _00724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07656__A2 vss _03135_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06313__C1 vss _01679_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_858 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_823 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11608_ vss net149 cpu.state.i_ctrl_misalign vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08605__A1 vss _04058_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_815 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11539_ vdd rf_ram.memory\[392\]\[0\] clknet_leaf_117_clk vss _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_528 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09030__A1 vss net247 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_218_clk vdd vss clknet_leaf_218_clk clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_0_444 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_279 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07592__A1 vss _03425_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05962_ vdd vss _02158_ rf_ram.memory\[20\]\[0\] _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05483__I vss _01624_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06579__I vss _02760_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08750_ vdd vss _04166_ rf_ram.memory\[147\]\[1\] _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06147__A2 vss _01808_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07701_ vdd vss _03501_ rf_ram.memory\[400\]\[0\] _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_1167 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09333__A2 vss _04037_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05893_ _02085_ _02088_ vdd vss _02089_ _02077_ _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_08681_ vdd _04122_ _04120_ _00752_ _04097_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_714 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07632_ vdd _03457_ _03456_ _00368_ _03455_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_747 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07563_ vdd _03414_ _03413_ _00342_ _03389_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09097__A1 vss net237 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09302_ vdd _04516_ _04514_ _00979_ _04466_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_572 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07494_ vdd vss _03372_ rf_ram.memory\[364\]\[0\] _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_622 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08844__A1 vss _04205_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_609 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06514_ _02702_ _01399_ _01421_ vdd vss _02703_ _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_119_869 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09233_ _04466_ _04400_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06445_ _01607_ rf_ram.memory\[35\]\[1\] vdd vss _02640_ rf_ram.memory\[34\]\[1\]
+ _01605_ _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_1_1104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09839__B vss _02709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09164_ vdd _04423_ _04422_ _00934_ _04397_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_951 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_694 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06376_ rf_ram.memory\[249\]\[1\] _01793_ _01863_ rf_ram.memory\[248\]\[1\] _02571_
+ vss vdd rf_ram.memory\[251\]\[1\] _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08115_ vdd vss _03759_ _02751_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_181_clk_I vss clknet_5_29__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09095_ vdd vss _04380_ rf_ram.memory\[97\]\[1\] _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72_995 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05327_ _01523_ _01509_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05258_ vdd _01173_ _01455_ _01442_ _01457_ vss _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_08046_ vdd vss _03716_ rf_ram.memory\[566\]\[0\] _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_61_clk_I vss clknet_5_9__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_209_clk vdd vss clknet_leaf_209_clk clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_3_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05189_ vdd vss cpu.ctrl.pc _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07583__A1 vss _02935_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09997_ vdd vss _04965_ rf_ram.memory\[276\]\[0\] _04964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_196_clk_I vss clknet_5_25__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06386__A2 vss _01808_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08948_ vdd _04288_ _04286_ _00853_ _04269_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_76_clk_I vss clknet_5_10__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08879_ vdd _04246_ _04245_ _00826_ _04234_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output130_I vss net130 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10910_ vdd rf_ram.memory\[199\]\[0\] clknet_leaf_39_clk vss _00654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07335__A1 vss _03257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_369 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10841_ vdd rf_ram.memory\[536\]\[1\] clknet_leaf_311_clk vss _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_728 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08835__A1 vss _03672_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1083 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10772_ vdd rf_ram.memory\[570\]\[0\] clknet_leaf_305_clk vss _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_134_clk_I vss clknet_5_24__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05649__A1 vss _01600_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_87_1037 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_14_clk_I vss clknet_5_2__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_149_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_509 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11324_ vdd net138 clknet_leaf_249_clk vss _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09012__A1 vss _02774_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11255_ vdd cpu.alu.add_cy_r clknet_leaf_218_clk vss _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05821__A1 vss net251 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_29_clk_I vss clknet_5_1__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10206_ vdd _05093_ _05092_ _01307_ _05078_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11186_ vdd rf_ram.memory\[91\]\[0\] clknet_leaf_57_clk vss _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_1133 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10137_ vdd vss _05051_ _02794_ _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_1244 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_1008 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10068_ vdd vss _05008_ _02838_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06129__A2 vss _01697_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_45 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05337__B1 vss _01521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06348__B vss _01650_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09079__A1 vss _04364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_553 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06230_ _01629_ vdd vss _02425_ _02423_ _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__06301__A2 vss _01664_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06161_ _01693_ vdd vss _02356_ rf_ram.memory\[480\]\[1\] _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06092_ rf_ram.memory\[328\]\[1\] _02287_ vss vdd rf_ram.memory\[331\]\[1\] _01713_
+ rf_ram.memory\[329\]\[1\] _01721_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__07801__A2 vss _03234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05478__I vss _01349_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09920_ vdd vss _04917_ rf_ram.memory\[343\]\[1\] _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_145_1171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_382 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07565__A1 vss _03393_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06368__A2 vss _01989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_274 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09851_ _04874_ vdd vss _01170_ _02713_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__09554__A2 vss _01491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09782_ vdd _04832_ _04831_ _01143_ _04634_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08802_ vdd _04198_ _04196_ _00797_ _04170_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06994_ vdd _03057_ _03056_ _00130_ _03050_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05945_ vdd vss _02141_ rf_ram.memory\[36\]\[0\] _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08733_ vdd vss _04155_ rf_ram.memory\[148\]\[1\] _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07317__A1 vss _03260_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07868__A2 vss _03559_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_306 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05876_ _02071_ vdd vss _02072_ _01600_ _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_15_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08664_ vdd _04112_ _04111_ _00745_ _04094_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07615_ vdd vss _03447_ rf_ram.memory\[313\]\[0\] _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_117_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08595_ vdd _04069_ _04068_ _00719_ _04058_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06258__B vss _01805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07546_ vdd vss _03404_ _02921_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08817__A1 vss _04202_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_48_255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07477_ vdd _03361_ _03357_ _00309_ _03360_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_162_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_614 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_666 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09216_ vdd _04455_ _04454_ _00954_ _04431_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08293__A2 vss _02781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_620 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09569__B vss _04678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_161_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06428_ _02621_ _02622_ vdd vss _02623_ _02619_ _02620_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_09147_ vdd vss _04413_ rf_ram.memory\[8\]\[0\] _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08045__A2 vss _03693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_494 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06359_ _01564_ vdd vss _02554_ _02551_ _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09078_ vdd vss _04370_ rf_ram.memory\[57\]\[0\] _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_188_70 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output178_I vss net178 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08029_ vdd _03705_ _03703_ _00517_ _03690_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07556__A1 vss _02806_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11040_ vdd rf_ram.memory\[147\]\[0\] clknet_leaf_0_clk vss _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_308 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07308__A1 vss _03222_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1112 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_1167 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10824_ vdd rf_ram.memory\[544\]\[0\] clknet_leaf_314_clk vss _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06531__A2 vss _01503_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_931 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_750 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10755_ vdd rf_ram.memory\[46\]\[1\] clknet_leaf_203_clk vss _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10686_ vdd rf_ram.memory\[415\]\[0\] clknet_leaf_90_clk vss _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_485 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05800__B vss _01527_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_753 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_861 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1080 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_797 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05298__I vss _01493_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11307_ _01040_ vdd vss clknet_leaf_265_clk net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_10_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_22_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06598__A2 vss _02775_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1198 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11238_ vdd rf_ram.memory\[65\]\[0\] clknet_leaf_61_clk vss _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_5_27__f_clk vdd vss clknet_5_27__leaf_clk clknet_3_6_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11169_ vdd rf_ram.memory\[98\]\[1\] clknet_leaf_62_clk vss _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06350__C vss _01717_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07018__I vss _03071_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1115 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1148 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05730_ vdd vss _01926_ rf_ram.memory\[441\]\[0\] _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_187_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_158_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05661_ _01857_ _01695_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_188_886 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08380_ vdd vss _03924_ _03134_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07400_ vdd _03312_ _03310_ _00281_ _03292_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06522__A2 vss _01376_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05592_ vdd vss _01788_ rf_ram.memory\[289\]\[0\] _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_07331_ vdd vss _03270_ rf_ram.memory\[271\]\[1\] _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_1170 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_720 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07262_ vdd _03226_ _03223_ _00229_ _03225_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_170_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_455 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09224__A1 vss _03319_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06213_ _01693_ vdd vss _02408_ rf_ram.memory\[392\]\[1\] _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09001_ vdd _04321_ _04319_ _00873_ _04301_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07193_ vdd _03183_ _03181_ _00203_ _03161_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_182_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06144_ _02337_ _02338_ vdd vss _02339_ _02335_ _02336_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_124_680 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09775__A2 vss _04507_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06075_ _01629_ vdd vss _02270_ _02267_ _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_112_864 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09903_ vdd _04906_ _04905_ _01191_ _04884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07538__A1 vss _03389_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05549__B1 vss _01696_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09834_ vdd _04864_ _04863_ _01163_ _04837_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06977_ vdd vss _03046_ rf_ram.memory\[427\]\[1\] _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09765_ _04760_ _04821_ vdd vss _04822_ net121 _04766_ net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__08468__B vss _03984_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05928_ rf_ram.memory\[100\]\[0\] _02124_ vss vdd rf_ram.memory\[103\]\[0\] _01696_
+ rf_ram.memory\[101\]\[0\] _01848_ _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09696_ vdd vss _04774_ _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08716_ vdd _04144_ _04143_ _00765_ _04126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08647_ vdd vss _04102_ net238 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05859_ vdd vss _02055_ rf_ram.memory\[225\]\[0\] _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07710__A1 vss net240 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08578_ _04057_ _02742_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_187_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07529_ vdd vss _03394_ rf_ram.memory\[361\]\[1\] _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1064 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_528 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10540_ vdd rf_ram.memory\[372\]\[0\] clknet_leaf_147_clk vss _00284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10073__A2 vss _03134_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10471_ vdd rf_ram.memory\[425\]\[1\] clknet_leaf_100_clk vss _00215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_831 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05788__B1 vss _01608_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_659 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11023_ vdd rf_ram.memory\[39\]\[1\] clknet_leaf_41_clk vss _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_1068 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05581__I vss _01686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_604 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06677__I vss _02838_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_86_125 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_184_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_1072 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10807_ vdd rf_ram.memory\[553\]\[1\] clknet_leaf_322_clk vss _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_125_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10738_ vdd rf_ram.memory\[440\]\[0\] clknet_leaf_55_clk vss _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_556 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_989 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09206__A1 vss _04431_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_589 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10669_ vdd rf_ram.memory\[377\]\[1\] clknet_leaf_108_clk vss _00413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput106 o_dbus_dat[17] net106 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput128 o_dbus_dat[8] net128 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput117 o_dbus_dat[27] net117 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput139 o_ext_rs1[10] net139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06900_ vdd vss _02995_ rf_ram.memory\[280\]\[1\] _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07880_ vdd _03611_ _03610_ _00462_ _03587_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08193__A1 vss _03790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09390__B1 vss _04564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06831_ vdd _02948_ _02947_ _00076_ _02927_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05705__B vss _01504_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05491__I vss _01686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07940__A1 vss _02781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09550_ _04669_ vdd vss _04670_ _01391_ _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06762_ vdd vss _02898_ _02750_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05713_ _01909_ _01756_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08501_ vdd vss _04007_ rf_ram.memory\[79\]\[0\] _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09481_ _01411_ vdd vss _04619_ net89 _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08432_ vdd vss _03957_ rf_ram.memory\[59\]\[1\] _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06693_ vdd vss _02851_ rf_ram.memory\[524\]\[0\] _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_867 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05703__B1 vss _01726_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05644_ rf_ram.memory\[500\]\[0\] _01840_ vss vdd rf_ram.memory\[503\]\[0\] _01519_
+ rf_ram.memory\[501\]\[0\] _01668_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_05575_ vdd vss _01771_ rf_ram.memory\[302\]\[0\] _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_129_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08363_ vdd vss _03913_ _02991_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_128_260 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09996__A2 vss _03135_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07314_ vdd _03259_ _03258_ _00248_ _03257_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08294_ vdd vss _03870_ rf_ram.memory\[203\]\[0\] _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_1237 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07245_ vdd _03215_ _03213_ _00223_ _03193_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09847__B vss _01391_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07759__A1 vss _03521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07176_ vdd _03173_ _03172_ _00196_ _03157_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11668__I vss net119 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06127_ _02321_ vdd vss _02322_ _01769_ _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_30_935 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06271__B vss _01956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06058_ _02252_ vdd vss _02253_ _01527_ _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA_input54_I vss i_ibus_rdt[29] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05234__A2 vss _01418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_681 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08184__A1 vss _02838_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_10__f_clk vdd vss clknet_5_10__leaf_clk clknet_3_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09817_ vdd vss _04854_ net240 _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09748_ vdd vss _04810_ _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06734__A2 vss _02846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06498__A1 vss _02690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09679_ _04736_ net124 vdd vss _04762_ net1 net28 _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_178_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_333 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_670 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_309 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1099 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11641_ net192 vss vdd net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__05170__A1 vss _01353_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_512 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06446__B vss _01493_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_876 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11572_ vdd rf_ram.memory\[210\]\[1\] clknet_leaf_30_clk vss _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07998__A1 vss _03654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10523_ vdd rf_ram.memory\[268\]\[1\] clknet_leaf_194_clk vss _00267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput19 vss net19 i_dbus_rdt[25] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_load_slew244_I vss _02821_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05473__A2 vss _01500_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10454_ vdd rf_ram.memory\[1\]\[0\] clknet_leaf_41_clk vss _00198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_818 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10385_ vdd rf_ram.memory\[227\]\[1\] clknet_leaf_277_clk vss _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05576__I vss _01617_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06422__A1 vss _01909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1266 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08175__A1 vss _03787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11006_ vdd rf_ram.memory\[15\]\[0\] clknet_leaf_295_clk vss _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07922__A1 vss _03619_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06489__A1 vss _01348_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_158 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_114_89 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05360_ rf_ram.memory\[531\]\[0\] _01554_ _01501_ rf_ram.memory\[530\]\[0\] _01556_
+ vss vdd rf_ram.memory\[529\]\[0\] _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__06356__B vss _01551_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_753 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07989__A1 vss _03672_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_414 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_334 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05291_ _01438_ vdd vss _01488_ _01486_ _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__06870__I vss _02825_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07030_ vdd vss _03080_ rf_ram.memory\[216\]\[0\] _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06091__B vss _01602_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05486__I vss _01508_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09450__I1 vss net76 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08981_ vdd _04309_ _04307_ _00865_ _04301_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_478 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07932_ vdd _03643_ _03642_ _00482_ _03619_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08797__I vss _04077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07863_ vdd vss _03601_ _02774_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_78_1131 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_155_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06814_ vdd vss _02936_ _02935_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09602_ _04526_ vdd vss _04711_ cpu.immdec.imm24_20\[3\] _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07794_ vdd _03558_ _03555_ _00429_ _03557_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09533_ vdd vss _04659_ _04478_ cpu.immdec.imm19_12_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_968 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09666__A1 vss net1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06745_ vdd vss _02886_ rf_ram.memory\[516\]\[1\] _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09464_ vss _01049_ _04608_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_309 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06676_ vdd vss _02838_ _02716_ _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05627_ _01688_ rf_ram.memory\[491\]\[0\] vdd vss _01823_ rf_ram.memory\[490\]\[0\]
+ _01687_ _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07141__A2 vss _02911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08415_ vss _03945_ _02996_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09395_ vdd vss _04570_ _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_149_1114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08346_ vdd vss _03902_ _02731_ _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__09969__A2 vss _02946_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05558_ _01753_ vdd vss _01754_ _01527_ _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_50_1094 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_870 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05489_ _01684_ vdd vss _01685_ rf_ram.memory\[344\]\[0\] _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_117_764 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08277_ vdd _03859_ _03857_ _00611_ _03855_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_1089 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09577__B vss cpu.decode.opcode\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07228_ vdd _03205_ _03204_ _00216_ _03190_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05455__A2 vss _01649_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06652__A1 vss _02748_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_583 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07159_ vdd vss _03163_ _02915_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05207__A2 vss _01382_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ vdd vss _05071_ rf_ram.memory\[447\]\[1\] _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output160_I vss net160 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_675 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07904__A1 vss _03622_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1226 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06707__A2 vss _02846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07380__A2 vss _03253_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09657__A1 vss net98 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05679__C1 vss _01810_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_333 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_798 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_938 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09409__A1 vss _01436_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_190_clk vdd vss clknet_leaf_190_clk clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11624_ vss net146 net74 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_182_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_731 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11555_ vdd rf_ram.memory\[450\]\[0\] clknet_leaf_113_clk vss _01287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_892 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05446__A2 vss _01641_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11486_ vdd rf_ram.memory\[464\]\[1\] clknet_leaf_134_clk vss _01218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10506_ vdd rf_ram.memory\[272\]\[0\] clknet_leaf_189_clk vss _00250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10437_ vdd rf_ram.memory\[486\]\[1\] clknet_leaf_223_clk vss _00181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07199__A2 vss _02941_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10368_ vdd rf_ram.memory\[206\]\[0\] clknet_leaf_38_clk vss _00112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_648 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06946__A2 vss _02766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10299_ vdd rf_ram.memory\[521\]\[1\] clknet_leaf_316_clk vss _00043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06159__B1 vss _01688_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08148__A1 vss _03754_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09896__A1 vss _02828_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08699__A2 vss _02921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09442__S vss _04593_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09648__A1 vss net1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06530_ vdd vss _02716_ _01512_ _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_140_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06461_ _02654_ _02655_ vdd vss _02656_ _02652_ _02653_ rf_ram.i_raddr\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06086__B vss _01602_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_675 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_181_clk vdd vss clknet_leaf_181_clk clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_118_517 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05412_ _01608_ _01607_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_56_651 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08200_ vdd vss _03812_ rf_ram.memory\[537\]\[0\] _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05685__A2 vss _01711_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06882__A1 vss _02975_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09180_ vdd _04433_ _04432_ _00940_ _04431_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06392_ vdd vss _02587_ rf_ram.memory\[68\]\[1\] _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_172_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05343_ _01539_ vss vdd _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08131_ vdd vss _03769_ _02805_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__06634__A1 vss _02748_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08062_ vdd vss _03726_ net242 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05274_ _01472_ vdd vss _01473_ _01381_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_144_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_244 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05842__C1 vss _01645_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07013_ vdd vss _03069_ rf_ram.memory\[222\]\[0\] _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08387__A1 vss _03919_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1130 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10194__A1 vss _03892_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_798 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08964_ _04298_ _04057_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07915_ vdd vss _03633_ _02844_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08895_ vdd vss _04256_ rf_ram.memory\[127\]\[1\] _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07846_ vdd vss _03591_ rf_ram.memory\[431\]\[1\] _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09860__B vss _02714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07777_ vss _03547_ _03039_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__09639__A1 vss _02971_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input17_I vss i_dbus_rdt[23] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10249__A2 vss _03035_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09516_ vdd vss _04645_ _04524_ net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06728_ vdd vss _02874_ _02806_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xserv_rf_top_257 o_mdu_valid vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09447_ vss _01041_ _04599_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_172_clk vdd vss clknet_leaf_172_clk clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06659_ vdd _02824_ _02823_ _00028_ _02820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_164_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_185 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05676__A2 vss _01804_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06873__A1 vss _02813_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09378_ _04561_ vss vdd _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__09811__A1 vss _04840_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08329_ vdd _03891_ _03889_ _00631_ _03887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11340_ vdd cpu.immdec.imm19_12_20\[6\] clknet_leaf_215_clk vss _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1253 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_175 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11271_ vdd net206 clknet_leaf_247_clk vss _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10222_ vdd vss _05103_ rf_ram.memory\[23\]\[1\] _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10185__A1 vss _05078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ vdd vss _05061_ rf_ram.memory\[450\]\[0\] _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07050__A1 vss _02806_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_8__f_clk vdd vss clknet_5_8__leaf_clk clknet_3_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_101_962 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10084_ vdd _05018_ _05015_ _01260_ _05017_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09878__A1 vss _04884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1023 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08550__A1 vss _04023_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07353__A2 vss _02839_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1007 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05803__B vss _01564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168_951 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08302__A1 vss _03855_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10986_ vdd rf_ram.memory\[164\]\[0\] clknet_leaf_331_clk vss _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_163_clk vdd vss clknet_leaf_163_clk clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05522__C vss _01717_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_826 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_314 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06313__B1 vss _01793_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_645 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_302_clk_I vss clknet_5_6__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_678 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11607_ vss net137 cpu.csr_d_sel vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_154_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_128_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09802__A1 vss net246 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_153 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_345 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11538_ vdd rf_ram.memory\[312\]\[1\] clknet_leaf_110_clk vss _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05824__C1 vss _01968_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_317_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06092__A2 vss _01724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11469_ vdd rf_ram.memory\[341\]\[0\] clknet_leaf_170_clk vss _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_1049 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_748 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09030__A2 vss _04339_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10176__A1 vss _05049_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_478 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_188_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input9_I vss i_dbus_rdt[16] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07700_ vdd vss _03500_ _02945_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_1135 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05961_ _02156_ _01568_ vdd vss _02157_ _01599_ _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__09869__A1 vss _04884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1071 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05892_ _02087_ vdd vss _02088_ _01972_ _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08680_ vdd vss _04122_ rf_ram.memory\[559\]\[1\] _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07631_ vdd vss _03457_ rf_ram.memory\[388\]\[0\] _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08541__A1 vss net246 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07562_ vdd vss _03414_ rf_ram.memory\[318\]\[0\] _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_540 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09097__A2 vss _04339_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09301_ vdd vss _04516_ rf_ram.memory\[66\]\[1\] _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06513_ vdd vss _02702_ _01391_ _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_154_clk vdd vss clknet_leaf_154_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07493_ vdd vss _03371_ _02788_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10100__A1 vss _02800_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09232_ vdd _04465_ _04464_ _00960_ _04463_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_150_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06444_ vdd vss _02639_ rf_ram.memory\[33\]\[1\] _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_185_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09163_ vdd vss _04423_ rf_ram.memory\[87\]\[0\] _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_90_215 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06375_ _01783_ vdd vss _02570_ rf_ram.memory\[250\]\[1\] _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_5_10__f_clk_I vss clknet_3_2_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05326_ rf_ram.memory\[525\]\[0\] _01517_ _01511_ rf_ram.memory\[524\]\[0\] _01522_
+ vss vdd rf_ram.memory\[527\]\[0\] _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08114_ vdd _03758_ _03755_ _00549_ _03757_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_142_862 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_391 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09094_ vdd _04379_ _04378_ _00908_ _04364_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05815__C1 vss _01786_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_304 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07280__A1 vss _02836_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05257_ vdd vss cpu.mem_if.signbit _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08045_ vdd vss _03715_ _03008_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10167__A1 vss _02908_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05830__A2 vss _01537_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05188_ vdd vss _01388_ _01384_ _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_177_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07583__A2 vss _02839_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09996_ vdd vss _04964_ _02940_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05607__C vss _01717_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08947_ vdd vss _04288_ rf_ram.memory\[449\]\[1\] _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08878_ vdd vss _04246_ rf_ram.memory\[128\]\[0\] _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07829_ vdd vss _03580_ rf_ram.memory\[412\]\[1\] _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_93_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10840_ vdd rf_ram.memory\[536\]\[0\] clknet_leaf_312_clk vss _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05897__A2 vss _01683_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_145_clk vdd vss clknet_leaf_145_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08835__A2 vss _03072_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1049 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10771_ vdd rf_ram.memory\[571\]\[1\] clknet_leaf_305_clk vss _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_118_881 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06454__B vss _01601_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_147 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06074__A2 vss _01623_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07271__A1 vss _03222_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11323_ _01056_ vdd vss clknet_leaf_254_clk net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11254_ vdd rf_ram.memory\[309\]\[1\] clknet_leaf_150_clk vss _00990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_1094 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09012__A2 vss _03945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07023__A1 vss _03053_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10205_ vdd vss _05093_ rf_ram.memory\[211\]\[0\] _05092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09484__C vss _03989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11185_ vdd rf_ram.memory\[92\]\[1\] clknet_leaf_56_clk vss _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08771__A1 vss _04170_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10136_ vdd _05050_ _05047_ _01280_ _05049_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10067_ vdd _05007_ _05005_ _01254_ _04985_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_101_1278 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08523__A1 vss _03956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_68 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05888__A2 vss _01804_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_136_clk vdd vss clknet_leaf_136_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10969_ vdd rf_ram.memory\[489\]\[1\] clknet_leaf_188_clk vss _00706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_241_clk_I vss clknet_5_21__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06298__C1 vss _01516_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09659__C vss _04740_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_256_clk_I vss clknet_5_20__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06160_ _01746_ vdd vss _02355_ _02352_ _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_103_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_40_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07262__A1 vss _03225_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06065__A2 vss _01500_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06091_ _01602_ vdd vss _02286_ rf_ram.memory\[330\]\[1\] _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__05812__A2 vss _01711_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10149__A1 vss _05046_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_556 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07014__A1 vss _03050_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05708__B vss _01903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09850_ vdd vss _04874_ cpu.state.cnt_r\[3\] cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08762__A1 vss _02760_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06222__C1 vss _01793_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09781_ vdd vss _04832_ rf_ram.memory\[187\]\[0\] _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08801_ vdd vss _04198_ rf_ram.memory\[140\]\[1\] _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06993_ vdd vss _03057_ rf_ram.memory\[226\]\[0\] _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05944_ _01493_ vdd vss _02140_ _02137_ _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08732_ vdd _04154_ _04153_ _00771_ _04126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08514__A1 vss _02787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08663_ vdd vss _04112_ rf_ram.memory\[158\]\[0\] _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05875_ _02068_ _02069_ _02070_ _01860_ vdd vss _02071_ _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_07614_ vdd vss _03446_ _03445_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05879__A2 vss _01531_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_209_clk_I vss clknet_5_25__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08594_ vdd vss _04069_ rf_ram.memory\[166\]\[0\] _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07545_ vdd _03403_ _03401_ _00335_ _03393_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_127_clk vdd vss clknet_leaf_127_clk clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07476_ vdd vss _03361_ rf_ram.memory\[366\]\[1\] _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_165_228 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_280 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_576 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06427_ rf_ram.memory\[104\]\[1\] _02622_ vss vdd rf_ram.memory\[107\]\[1\] _01679_
+ rf_ram.memory\[105\]\[1\] _01793_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09215_ vdd vss _04455_ rf_ram.memory\[67\]\[0\] _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_91_524 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_475 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06274__B vss _01564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09146_ vdd vss _04412_ net250 _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_933 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06358_ _01959_ rf_ram.memory\[235\]\[1\] vdd vss _02553_ rf_ram.memory\[234\]\[1\]
+ _01940_ _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__06056__A2 vss _01641_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07253__A1 vss _03190_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05309_ vss _01505_ _01504_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09077_ vdd vss _04369_ _03668_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_06289_ vdd vss _02484_ rf_ram.memory\[142\]\[1\] _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08028_ vdd vss _03705_ rf_ram.memory\[570\]\[1\] _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_191 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07556__A2 vss _03390_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09979_ vdd vss _04954_ rf_ram.memory\[274\]\[1\] _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08753__A1 vss net236 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08505__A1 vss _01369_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_118_clk vdd vss clknet_leaf_118_clk clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_129_409 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_1059 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10823_ vdd rf_ram.memory\[545\]\[1\] clknet_leaf_321_clk vss _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_976 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10754_ vdd rf_ram.memory\[46\]\[0\] clknet_leaf_132_clk vss _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_598 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07492__A1 vss _03360_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_957 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10685_ vdd rf_ram.memory\[436\]\[1\] clknet_leaf_80_clk vss _00429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_166 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_1111 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08992__A1 vss net248 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06452__C1 vss _01635_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11306_ _01039_ vdd vss clknet_leaf_265_clk net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11237_ vdd cpu.genblk3.csr.mcause3_0\[3\] clknet_leaf_257_clk vss _00973_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05558__A1 vss _01527_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11168_ vdd rf_ram.memory\[98\]\[0\] clknet_leaf_77_clk vss _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08744__A1 vss _04157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10119_ vdd _05039_ _05037_ _01274_ _05017_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11099_ vdd rf_ram.memory\[429\]\[1\] clknet_leaf_99_clk vss _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09514__I vss _03992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06359__B vss _01564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_180_clk_I vss clknet_5_31__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_89 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05660_ _01856_ _01686_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_1235 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_109_clk vdd vss clknet_leaf_109_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05591_ vss _01787_ _01514_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__09450__S vss _04593_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07330_ vdd _03269_ _03268_ _00254_ _03257_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_60_clk_I vss clknet_5_9__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_524 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07483__A1 vss _02844_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07261_ vdd vss _03226_ rf_ram.memory\[418\]\[1\] _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05710__C vss _01670_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09000_ vdd vss _04321_ rf_ram.memory\[112\]\[1\] _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_195_clk_I vss clknet_5_25__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06286__A2 vss _01915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05494__B1 vss _01688_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06212_ _02406_ vdd vss _02407_ _01769_ _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09224__A2 vss _02866_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_75_clk_I vss clknet_5_10__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_7_0_clk clknet_3_7_0_clk vss vdd clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07192_ vdd vss _03183_ rf_ram.memory\[473\]\[1\] _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07235__A1 vss _03193_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06143_ rf_ram.memory\[306\]\[1\] _02338_ vss vdd rf_ram.memory\[305\]\[1\] _01721_
+ rf_ram.memory\[307\]\[1\] _01726_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_83_1255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06074_ _01688_ rf_ram.memory\[347\]\[1\] vdd vss _02269_ rf_ram.memory\[346\]\[1\]
+ _01623_ _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_1_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09902_ vdd vss _04906_ rf_ram.memory\[345\]\[0\] _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_133_clk_I vss clknet_5_24__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09833_ vdd vss _04864_ rf_ram.memory\[61\]\[0\] _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06210__A2 vss _01770_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06976_ vdd _03045_ _03044_ _00124_ _03014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_13_clk_I vss clknet_5_2__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09764_ vdd vss _04821_ _04804_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_154_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05927_ _02004_ vdd vss _02123_ rf_ram.memory\[102\]\[0\] _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09695_ _04768_ _04773_ vdd vss _04774_ net128 _04767_ net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_08715_ vdd vss _04144_ rf_ram.memory\[150\]\[0\] _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_148_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08646_ vdd _04101_ _04099_ _00738_ _04097_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05858_ _01956_ vdd vss _02054_ rf_ram.memory\[224\]\[0\] _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07710__A2 vss _02997_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_28_clk_I vss clknet_5_3__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_548 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08577_ vdd _04056_ _04054_ _00714_ _04026_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05789_ _01928_ vdd vss _01985_ _01983_ _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07528_ _03393_ _03359_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_147_762 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_395 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07459_ vdd vss _03349_ _02954_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_92_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_866 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06277__A2 vss _01958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1106 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10470_ vdd rf_ram.memory\[425\]\[0\] clknet_leaf_100_clk vss _00214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output190_I vss net190 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07226__A1 vss _02728_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_253 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09129_ vdd vss _04402_ rf_ram.memory\[92\]\[1\] _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_60_741 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06029__A2 vss _01538_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08974__A1 vss _04298_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_640 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_690 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1064 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11022_ vdd rf_ram.memory\[39\]\[0\] clknet_leaf_41_clk vss _00759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08726__A1 vss _04126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_339_clk vdd vss clknet_leaf_339_clk clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09151__A1 vss _02908_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05712__A1 vss _01768_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1046 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_885 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_716 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05811__B vss _01916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10806_ vdd rf_ram.memory\[553\]\[0\] clknet_leaf_322_clk vss _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_412 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10737_ vdd rf_ram.memory\[458\]\[1\] clknet_leaf_50_clk vss _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06268__A2 vss _01501_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_957 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10668_ vdd rf_ram.memory\[377\]\[0\] clknet_leaf_108_clk vss _00412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10599_ vdd rf_ram.memory\[318\]\[1\] clknet_leaf_106_clk vss _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08965__A1 vss _03008_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput107 o_dbus_dat[18] net107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput118 o_dbus_dat[28] net118 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06425__C1 vss _01625_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput129 o_dbus_dat[9] net129 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05779__A1 vss _01972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06440__A2 vss _01513_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_43_1250 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06830_ vdd vss _02948_ rf_ram.memory\[304\]\[0\] _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05772__I vss _01918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07940__A2 vss _02869_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05951__A1 vss _01526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06761_ vdd _02897_ _02895_ _00057_ _02876_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06089__B vss _01707_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05712_ _01907_ net254 vdd vss _01908_ _01768_ _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08500_ vdd vss _04006_ _02953_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06692_ vdd vss _02850_ _02788_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09480_ vdd vss _04618_ _04616_ _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05643_ _01504_ vdd vss _01839_ rf_ram.memory\[502\]\[0\] _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_77_115 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08431_ _03956_ vss vdd _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__05721__B vss _01916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08362_ vdd _03912_ _03910_ _00643_ _03887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05574_ _01770_ _01530_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_50_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06259__A2 vss _01666_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07456__A1 vss _03323_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07313_ vdd vss _03259_ rf_ram.memory\[256\]\[0\] _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08293_ vdd vss _03869_ _03230_ _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_73_332 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07244_ vdd vss _03215_ rf_ram.memory\[421\]\[1\] _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_171_540 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_990 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07175_ vdd vss _03173_ rf_ram.memory\[482\]\[0\] _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_75_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08956__A1 vss _04266_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06126_ rf_ram.memory\[301\]\[1\] _01848_ _01863_ rf_ram.memory\[300\]\[1\] _02321_
+ vss vdd rf_ram.memory\[303\]\[1\] _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_06057_ rf_ram.memory\[380\]\[1\] _02252_ vss vdd rf_ram.memory\[383\]\[1\] _01646_
+ rf_ram.memory\[381\]\[1\] _01645_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__06431__A2 vss _01915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_868 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input47_I vss i_ibus_rdt[22] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08708__A1 vss _04129_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08184__A2 vss _02846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06195__A1 vss _01769_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09816_ vdd _04853_ _04851_ _01156_ _04840_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09747_ _04791_ _04809_ vdd vss _04810_ net114 _04790_ net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06959_ vdd vss _03034_ rf_ram.memory\[230\]\[1\] _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09133__A1 vss _04397_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_684 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_137 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09678_ _04759_ _04760_ vdd vss _04761_ _04737_ _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__07695__A1 vss _02917_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1176 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_1138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08629_ vdd _04090_ _04088_ _00732_ _04062_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11640_ vss net181 net109 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_321 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11571_ vdd rf_ram.memory\[210\]\[0\] clknet_leaf_30_clk vss _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05350__C vss _01495_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10522_ vdd rf_ram.memory\[268\]\[0\] clknet_leaf_194_clk vss _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_584 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10453_ vdd rf_ram.memory\[482\]\[1\] clknet_leaf_187_clk vss _00197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06462__B vss _01599_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1201 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10384_ vdd rf_ram.memory\[227\]\[0\] clknet_leaf_277_clk vss _00128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06181__C vss net253 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11005_ vdd rf_ram.memory\[160\]\[1\] clknet_leaf_338_clk vss _00742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05933__A1 vss _01569_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05394__C1 vss _01539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09124__A1 vss _02838_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_273 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_936 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_133_1108 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1243 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07438__A1 vss _03326_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07989__A2 vss _02960_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_40_clk vdd vss clknet_leaf_40_clk clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_153_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06110__A1 vss _01603_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_787 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05290_ _01486_ vdd vss _01487_ _01434_ _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_180_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1204 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1009 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08938__A1 vss _04269_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_925 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07610__A1 vss _03422_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06413__A2 vss _01787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08980_ vdd vss _04309_ rf_ram.memory\[116\]\[1\] _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_121_481 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07931_ vdd vss _03643_ rf_ram.memory\[440\]\[0\] _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07862_ vdd _03600_ _03598_ _00455_ _03590_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06813_ vss _02935_ _02800_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09601_ vdd vss _04710_ cpu.immdec.imm24_20\[4\] _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07793_ vdd vss _03558_ rf_ram.memory\[436\]\[1\] _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09532_ _04658_ vdd vss _01067_ _04656_ _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09666__A2 vss net24 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06744_ vdd _02885_ _02884_ _00052_ _02873_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07677__A1 vss _02923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06675_ vdd vss _02837_ _02785_ _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09463_ _04604_ vdd vss _04608_ net81 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_175_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05626_ vdd vss _01822_ rf_ram.memory\[489\]\[0\] _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_94_939 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08414_ vdd _03944_ _03942_ _00663_ _03922_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_65_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09394_ _04564_ net220 vdd vss _04570_ net219 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07429__A1 vss _02923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05557_ vss vdd rf_ram.memory\[271\]\[0\] _01636_ rf_ram.memory\[269\]\[0\] _01645_
+ _01644_ rf_ram.memory\[268\]\[0\] _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_08345_ vdd _03901_ _03899_ _00637_ _03887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_184_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_31_clk vdd vss clknet_leaf_31_clk clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08276_ vdd vss _03859_ rf_ram.memory\[195\]\[1\] _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05488_ _01684_ _01550_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_6_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07227_ vdd vss _03205_ rf_ram.memory\[424\]\[0\] _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_415 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08929__A1 vss net244 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07158_ vdd _03162_ _03159_ _00189_ _03161_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05860__B1 vss _01953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06109_ vss vdd rf_ram.memory\[287\]\[1\] _01625_ rf_ram.memory\[285\]\[1\] _01678_
+ _01634_ rf_ram.memory\[284\]\[1\] _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_113_993 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06404__A2 vss _01863_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_1012 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07089_ vdd _03118_ _03117_ _00164_ _03087_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_98_clk vdd vss clknet_leaf_98_clk clknet_5_14__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_1142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_96_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09354__B2 vss net232 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09106__A1 vss _04367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05376__C1 vss _01521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05391__A2 vss _01502_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07668__A1 vss _03455_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_405 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_1058 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05679__B1 vss _01646_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06457__B vss _01503_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_304 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09409__A2 vss _01437_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11623_ vss net145 net73 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_844 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_22_clk vdd vss clknet_leaf_22_clk clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11554_ vdd rf_ram.memory\[451\]\[1\] clknet_leaf_113_clk vss _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08093__A1 vss _02843_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07840__A1 vss _03557_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11485_ vdd rf_ram.memory\[464\]\[0\] clknet_leaf_124_clk vss _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10505_ vdd rf_ram.memory\[256\]\[1\] clknet_leaf_197_clk vss _00249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06192__B vss _01860_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05587__I vss _01550_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10436_ vdd rf_ram.memory\[486\]\[0\] clknet_leaf_223_clk vss _00180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_891 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_576 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10367_ vdd rf_ram.memory\[228\]\[1\] clknet_leaf_275_clk vss _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10298_ vdd rf_ram.memory\[521\]\[0\] clknet_leaf_316_clk vss _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_89_clk vdd vss clknet_leaf_89_clk clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09896__A2 vss _03253_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05906__A1 vss _01768_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05382__A2 vss _01524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_941 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06460_ rf_ram.memory\[51\]\[1\] _01518_ _01499_ rf_ram.memory\[50\]\[1\] _02655_
+ vss vdd rf_ram.memory\[49\]\[1\] _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_172_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05411_ _01607_ _01518_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06391_ _01978_ vdd vss _02586_ _02583_ _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_13_clk vdd vss clknet_leaf_13_clk clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08130_ vdd _03768_ _03766_ _00555_ _03757_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_141_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_482 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05342_ _01538_ vss vdd _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_28_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07831__A1 vss _02945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_201 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05273_ vdd vss _01472_ _01470_ _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_08061_ vdd _03725_ _03722_ _00529_ _03724_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05497__I vss _01550_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05842__B1 vss _01636_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07012_ vdd vss _03068_ _02738_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_999 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06398__A1 vss _01769_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10194__A2 vss _02923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08963_ vdd _04297_ _04295_ _00859_ _04269_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_1099 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07914_ vdd _03632_ _03630_ _00475_ _03622_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08894_ vdd _04255_ _04254_ _00832_ _04234_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_75_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_50 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07845_ _03590_ _03359_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07776_ vdd _03546_ _03544_ _00423_ _03524_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09639__A2 vss _04507_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09515_ vdd vss cpu.immdec.imm31 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_6_1209 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06727_ _02873_ _02819_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_177_974 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_91_1184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_788 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09446_ _04593_ vdd vss _04599_ net73 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06658_ vdd vss _02824_ rf_ram.memory\[347\]\[0\] _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06322__A1 vss _01600_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_849 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06873__A2 vss _02941_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05609_ _01805_ _01503_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06589_ vdd _02769_ _02767_ _00013_ _02748_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09377_ vdd vss _04560_ _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_46_140 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08328_ vdd vss _03891_ rf_ram.memory\[21\]\[1\] _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08075__A1 vss _03721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08259_ vdd vss _03848_ rf_ram.memory\[526\]\[1\] _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_105_757 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_519 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_891 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11270_ vdd net205 clknet_leaf_247_clk vss _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10221_ vdd _05102_ _05101_ _01313_ _05078_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_max_cap247_I vss _02774_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10152_ vdd vss _05060_ _02831_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07050__A2 vss _03089_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output78_I vss net78 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10083_ vdd vss _05018_ rf_ram.memory\[350\]\[1\] _05015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09327__A1 vss _04466_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_508 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05349__C1 vss _01539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06561__A1 vss _01353_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05364__A2 vss _01511_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_574 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10985_ vdd rf_ram.memory\[165\]\[1\] clknet_leaf_339_clk vss _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_473 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_613 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_438 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11606_ vss net136 cpu.decode.co_mem_word vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08066__A1 vss _03724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_858 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11537_ _01269_ vdd vss clknet_leaf_110_clk rf_ram.memory\[312\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__07813__A1 vss _03554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_893 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1007 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09802__A2 vss _04004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_368 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05824__B1 vss _02019_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1137 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11468_ vdd rf_ram.memory\[342\]\[1\] clknet_leaf_174_clk vss _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10419_ vdd rf_ram.memory\[491\]\[1\] clknet_leaf_183_clk vss _00163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11399_ _01131_ vdd vss clknet_leaf_227_clk net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08421__I vss _03902_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1114 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05960_ _01599_ _02155_ vdd vss _02156_ _02147_ _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xclkbuf_leaf_2_clk vdd vss clknet_leaf_2_clk clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05891_ rf_ram.memory\[71\]\[0\] _01925_ _01719_ rf_ram.memory\[70\]\[0\] _02087_
+ vss vdd rf_ram.memory\[69\]\[0\] _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07630_ vdd vss _03456_ _02882_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08541__A2 vss _03949_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_727 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07561_ vdd vss _03413_ _02935_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_941 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09300_ vdd _04515_ _04514_ _00978_ _04463_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06512_ vdd vss _02701_ _01469_ cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_07492_ vdd _03370_ _03368_ _00315_ _03360_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10100__A2 vss _03083_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_432 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09231_ vdd vss _04465_ rf_ram.memory\[329\]\[0\] _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06443_ _01601_ vdd vss _02638_ rf_ram.memory\[32\]\[1\] _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_90_205 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_535 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09162_ vdd vss _04422_ net235 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06374_ rf_ram.memory\[252\]\[1\] _02569_ vss vdd rf_ram.memory\[255\]\[1\] _01625_
+ rf_ram.memory\[253\]\[1\] _01678_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_145_178 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08113_ vdd vss _03758_ rf_ram.memory\[554\]\[1\] _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_858 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05325_ _01521_ vss vdd _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09093_ vdd vss _04379_ rf_ram.memory\[97\]\[0\] _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05815__B1 vss _01772_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_154 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07280__A2 vss _02992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05256_ vdd vss _01456_ _01342_ _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08044_ vdd _03714_ _03712_ _00523_ _03690_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05187_ vss _01387_ _01386_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XANTENNA__10167__A2 vss _03547_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09995_ vdd _04963_ _04961_ _01226_ _04953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_980 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08946_ vdd _04287_ _04286_ _00852_ _04266_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_305 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08877_ vdd vss _04245_ net237 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_07828_ vdd _03579_ _03578_ _00442_ _03554_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05346__A2 vss _01524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07759_ vdd _03536_ _03535_ _00416_ _03521_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output116_I vss net116 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_149_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10770_ vdd rf_ram.memory\[571\]\[0\] clknet_leaf_304_clk vss _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09429_ _02707_ vdd vss _04590_ net95 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_180_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_151_104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09796__A1 vss _04840_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_249 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_390 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11322_ _01055_ vdd vss clknet_leaf_253_clk net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_22_349 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11253_ vdd rf_ram.memory\[309\]\[0\] clknet_leaf_150_clk vss _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06470__B vss _01493_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10204_ vdd vss _05092_ _03892_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08220__A1 vss _03823_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11184_ vdd rf_ram.memory\[92\]\[0\] clknet_leaf_56_clk vss _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10135_ vdd vss _05050_ rf_ram.memory\[454\]\[1\] _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_100_281 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06782__A1 vss _02873_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10066_ vdd vss _05007_ rf_ram.memory\[307\]\[1\] _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05814__B vss _01505_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__I1 vss net53 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_861 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05337__A2 vss _01532_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05742__C1 vss _01811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1066 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10968_ vdd rf_ram.memory\[489\]\[0\] clknet_leaf_188_clk vss _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08287__A1 vss _03855_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10094__A1 vss _05017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06298__B1 vss _01520_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_134 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10899_ vdd rf_ram.memory\[183\]\[1\] clknet_leaf_14_clk vss _00643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08039__A1 vss _03690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09787__A1 vss _04634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_5_2__f_clk_I vss clknet_3_0_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_479 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06090_ rf_ram.memory\[333\]\[1\] _01715_ _01709_ rf_ram.memory\[332\]\[1\] _02285_
+ vss vdd rf_ram.memory\[335\]\[1\] _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09448__S vss _04593_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06380__B vss _01597_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08211__A1 vss _03787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06222__B1 vss _01778_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08800_ vdd _04197_ _04196_ _00796_ _04167_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09780_ vdd vss _04831_ net244 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06773__A1 vss _02873_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06992_ vdd vss _03056_ _03055_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08762__A2 vss _04152_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05943_ _01624_ rf_ram.memory\[35\]\[0\] vdd vss _02139_ rf_ram.memory\[34\]\[0\]
+ _01605_ _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08731_ vdd vss _04154_ rf_ram.memory\[148\]\[0\] _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09711__B2 vss net103 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08514__A2 vss _03949_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08662_ vdd vss _04111_ _02916_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07613_ _03445_ _02800_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05874_ rf_ram.memory\[248\]\[0\] _02070_ vss vdd rf_ram.memory\[251\]\[0\] _01696_
+ rf_ram.memory\[249\]\[0\] _01793_ _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_156_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08593_ vdd vss _04068_ _02805_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07544_ vdd vss _03403_ rf_ram.memory\[320\]\[1\] _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08278__A1 vss _03230_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1203 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07475_ vss _03360_ _03359_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10085__A1 vss _02916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_292 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06426_ _01783_ vdd vss _02621_ rf_ram.memory\[106\]\[1\] _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09214_ vdd vss _04454_ net240 _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_174_785 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_8_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09145_ vdd _04411_ _04409_ _00927_ _04401_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_72_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_688 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06357_ vdd vss _02552_ rf_ram.memory\[233\]\[1\] _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09242__A3 vss net66 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_811 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09076_ vdd _04368_ _04365_ _00901_ _04367_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05308_ _01504_ vss vdd _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06288_ _01978_ vdd vss _02483_ _02481_ _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__08450__A1 vss cpu.state.genblk1.misalign_trap_sync_r vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_130_844 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_535 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05239_ vdd vss _01439_ _01434_ _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08027_ vdd _03704_ _03703_ _00516_ _03686_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09978_ _04953_ _04400_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_301_clk_I vss clknet_5_6__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06764__A1 vss _02881_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08753__A2 vss _04152_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08929_ vdd vss _04277_ net244 _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output233_I vss net233 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08505__A2 vss _01491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1032 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_316_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08269__A1 vss _03852_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10822_ vdd rf_ram.memory\[545\]\[0\] clknet_leaf_321_clk vss _00566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_224 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10753_ vdd rf_ram.memory\[47\]\[1\] clknet_leaf_129_clk vss _00497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_566 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_39_246 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10684_ vdd rf_ram.memory\[436\]\[0\] clknet_leaf_80_clk vss _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_1113 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_1004 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_603 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08441__A1 vss _03953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08992__A2 vss _04303_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_321 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06452__B1 vss _01609_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11305_ _01038_ vdd vss clknet_leaf_252_clk net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_26_1129 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05809__B vss _02004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10000__A1 vss _04953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11236_ vdd cpu.genblk3.csr.mcause3_0\[2\] clknet_leaf_257_clk vss _00972_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09941__A1 vss _04918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11167_ vdd rf_ram.memory\[57\]\[1\] clknet_leaf_296_clk vss _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06755__A1 vss _02773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10118_ vdd vss _05039_ rf_ram.memory\[373\]\[1\] _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11098_ vdd rf_ram.memory\[429\]\[0\] clknet_leaf_99_clk vss _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05963__C1 vss _01617_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10049_ vdd vss _04997_ rf_ram.memory\[306\]\[0\] _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07315__I vss _03017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05590_ _01786_ vss vdd _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10067__A1 vss _04985_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05730__A2 vss _01918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_955 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06375__B vss _01783_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07483__A2 vss _03101_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07260_ _03225_ _03017_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06211_ rf_ram.memory\[397\]\[1\] _01772_ _01711_ rf_ram.memory\[396\]\[1\] _02406_
+ vss vdd rf_ram.memory\[399\]\[1\] _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07191_ vdd _03182_ _03181_ _00202_ _03157_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06142_ _01602_ vdd vss _02337_ rf_ram.memory\[304\]\[1\] _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_130_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_1208 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_271 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06073_ vdd vss _02268_ rf_ram.memory\[345\]\[1\] _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_293_clk vdd vss clknet_leaf_293_clk clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09901_ vdd vss _04905_ _03319_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05797__A2 vss _01664_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06994__A1 vss _03050_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05549__A2 vss _01687_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09832_ vdd vss _04863_ _03668_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06746__A1 vss _02876_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09763_ vdd vss _04820_ _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06975_ vdd vss _03045_ rf_ram.memory\[427\]\[0\] _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08714_ vdd vss _04143_ _03008_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05926_ _02120_ _02121_ vdd vss _02122_ _02118_ _02119_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_83_50 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09694_ vdd vss _04773_ _04740_ net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05706__C1 vss _01763_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07171__A1 vss _03157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08645_ vdd vss _04101_ rf_ram.memory\[519\]\[1\] _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05857_ _01564_ vdd vss _02053_ _02050_ _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_179_899 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08576_ vdd vss _04056_ rf_ram.memory\[16\]\[1\] _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07527_ vdd _03392_ _03391_ _00328_ _03389_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05721__A2 vss _01915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10058__A1 vss _02821_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05788_ rf_ram.memory\[139\]\[0\] _01608_ _01606_ rf_ram.memory\[138\]\[0\] _01984_
+ vss vdd rf_ram.memory\[137\]\[0\] _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07458_ vdd _03348_ _03346_ _00303_ _03326_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08671__A1 vss _04097_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_953 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05485__A1 vss _01675_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06409_ vdd vss _02604_ rf_ram.memory\[116\]\[1\] _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_107_638 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07389_ vdd _03305_ _03303_ _00277_ _03292_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_901 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07226__A2 vss _03040_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output183_I vss net183 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09128_ _04401_ _04400_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_284_clk vdd vss clknet_leaf_284_clk clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_128_1190 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_114_181 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05629__B vss _01693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_321 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09059_ vdd _04357_ _04355_ _00895_ _04334_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05788__A2 vss _01606_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06985__A1 vss _02766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_240_clk_I vss clknet_5_21__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09923__A1 vss _04911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06198__C1 vss _01713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11021_ vdd rf_ram.memory\[153\]\[1\] clknet_leaf_330_clk vss _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_1138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_255_clk_I vss clknet_5_20__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05364__B vss _01552_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06179__C vss _01670_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09151__A2 vss _04077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10805_ vdd rf_ram.memory\[554\]\[1\] clknet_leaf_321_clk vss _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10736_ vdd rf_ram.memory\[458\]\[0\] clknet_leaf_50_clk vss _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_333 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08662__A1 vss _02916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10667_ vdd rf_ram.memory\[396\]\[1\] clknet_leaf_96_clk vss _00411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08414__A1 vss _03922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10598_ vdd rf_ram.memory\[318\]\[0\] clknet_leaf_106_clk vss _00342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06425__B1 vss _01702_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10221__A1 vss _05078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05228__A1 vss _01375_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_275_clk vdd vss clknet_leaf_275_clk clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06976__A1 vss _03014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08965__A2 vss _04038_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput108 o_dbus_dat[19] net108 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput119 o_dbus_dat[29] net119 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_50_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_208_clk_I vss clknet_5_19__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09914__A1 vss _04884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11219_ vdd rf_ram.memory\[67\]\[1\] clknet_leaf_60_clk vss _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput90 o_dbus_adr[3] net90 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06728__A1 vss _02806_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06760_ vdd vss _02897_ rf_ram.memory\[514\]\[1\] _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05711_ _01900_ _01660_ _01906_ vdd vss _01907_ _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_06691_ vdd _02849_ _02847_ _00035_ _02826_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09461__S vss _04604_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07153__A1 vss _02883_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05642_ _01629_ vdd vss _01838_ _01836_ _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08430_ vdd _03955_ _03954_ _00668_ _03953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06884__I vss _02983_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05703__A2 vss _01801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_148_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_609 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_368 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05573_ _01769_ _01650_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08361_ vdd vss _03912_ rf_ram.memory\[183\]\[1\] _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_514 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_796 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06113__C1 vss _01646_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07312_ vdd vss _03258_ _02904_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08292_ vdd _03868_ _03866_ _00617_ _03855_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07243_ vdd _03214_ _03213_ _00222_ _03190_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_143_232 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08405__A1 vss net236 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_596 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07174_ vdd vss _03172_ _02894_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_15_967 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_266_clk vdd vss clknet_leaf_266_clk clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_160_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06125_ vdd vss _02320_ rf_ram.memory\[302\]\[1\] _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06967__A1 vss _02797_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06056_ vdd vss _02251_ rf_ram.memory\[382\]\[1\] _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09905__A1 vss _04887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09815_ vdd vss _04853_ rf_ram.memory\[7\]\[1\] _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09435__I vss _01411_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07392__A1 vss _03289_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09746_ vdd vss _04809_ _04804_ net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06958_ vdd _03033_ _03032_ _00118_ _03014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05909_ _02104_ vdd vss _02105_ _01909_ _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__05942__A2 vss _01513_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09677_ vdd vss _04760_ _04739_ _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_06889_ vdd _02987_ _02985_ _00095_ _02975_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08628_ vdd vss _04090_ rf_ram.memory\[539\]\[1\] _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07695__A2 vss _03496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08892__A1 vss _02908_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1008 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08559_ vdd vss _04046_ rf_ram.memory\[499\]\[0\] _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11570_ vdd rf_ram.memory\[238\]\[1\] clknet_leaf_285_clk vss _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08644__A1 vss _04094_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10521_ vdd rf_ram.memory\[252\]\[1\] clknet_leaf_219_clk vss _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_788 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10452_ vdd rf_ram.memory\[482\]\[0\] clknet_leaf_187_clk vss _00196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10203__A1 vss _05081_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09444__I0 vss net72 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10383_ vdd rf_ram.memory\[426\]\[1\] clknet_leaf_101_clk vss _00127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_161_1029 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_950 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_403 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_926 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_257_clk vdd vss clknet_leaf_257_clk clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06958__A1 vss _03014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11004_ vdd rf_ram.memory\[160\]\[0\] clknet_leaf_338_clk vss _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_194_clk_I vss clknet_5_28__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06186__A2 vss _01697_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_6_0_clk clknet_3_6_0_clk vss vdd clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__05394__B1 vss _01540_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_74_clk_I vss clknet_5_10__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09124__A2 vss _04005_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05933__A2 vss _02117_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07135__A1 vss _03126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05697__A1 vss _01675_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_89_clk_I vss clknet_5_11__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_869 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_344 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10719_ vdd rf_ram.memory\[446\]\[1\] clknet_leaf_78_clk vss _00463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_132_clk_I vss clknet_5_24__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_12_clk_I vss clknet_5_2__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06372__C vss _01620_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_358 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_753 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_147_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_141_758 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09060__A1 vss net241 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_248_clk vdd vss clknet_leaf_248_clk clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05621__A1 vss _01597_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07930_ vdd vss _03642_ _02991_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_27_clk_I vss clknet_5_3__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_99 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_1036 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07374__A1 vss _03292_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1009 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07861_ vdd vss _03600_ rf_ram.memory\[40\]\[1\] _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06177__A2 vss _01644_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07792_ _03557_ vss vdd _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06812_ vdd _02934_ _02932_ _00071_ _02930_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09600_ vdd vss net48 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05924__A2 vss _01989_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09531_ vdd vss _04658_ _04526_ net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06743_ vdd vss _02885_ rf_ram.memory\[516\]\[0\] _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07126__A1 vss _02883_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_302 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06674_ _02836_ vss vdd _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__08874__A1 vss _04234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_447 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09462_ vss _01048_ _04607_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05625_ _01684_ vdd vss _01821_ rf_ram.memory\[488\]\[0\] _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08413_ vdd vss _03944_ rf_ram.memory\[177\]\[1\] _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09393_ vdd vss _04569_ _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_164_817 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07429__A2 vss _03101_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05556_ vdd vss _01752_ rf_ram.memory\[270\]\[0\] _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08344_ vdd vss _03901_ rf_ram.memory\[214\]\[1\] _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_59_694 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_333 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05152__A3 vss _01344_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_89_1240 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06101__A2 vss _01626_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05487_ _01683_ vss vdd _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08275_ vdd _03858_ _03857_ _00610_ _03852_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07226_ vdd vss _03204_ _02728_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08929__A2 vss _04038_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_758 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07157_ vdd vss _03162_ rf_ram.memory\[484\]\[1\] _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_239_clk vdd vss clknet_leaf_239_clk clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06108_ vdd vss _02303_ rf_ram.memory\[286\]\[1\] _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07088_ vdd vss _03118_ rf_ram.memory\[490\]\[0\] _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_778 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06039_ _02222_ _02234_ _01351_ _02233_ _01362_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__09354__A2 vss _03991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05376__B1 vss _01517_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05915__A2 vss _01918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ vdd vss _04797_ _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05642__B vss _01629_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_119 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05361__C vss _01494_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_823 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06340__A2 vss _01531_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11622_ vss net144 net72 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08617__A1 vss _04058_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11553_ vdd rf_ram.memory\[451\]\[0\] clknet_leaf_113_clk vss _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09290__A1 vss _04463_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_303 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08093__A2 vss _03729_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11484_ vdd rf_ram.memory\[295\]\[1\] clknet_leaf_139_clk vss _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10504_ vdd rf_ram.memory\[256\]\[0\] clknet_leaf_196_clk vss _00248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09417__I0 vss net87 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_235 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09042__A1 vss _04331_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10435_ vdd rf_ram.memory\[4\]\[1\] clknet_leaf_209_clk vss _00179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_572 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10366_ vdd rf_ram.memory\[228\]\[0\] clknet_leaf_275_clk vss _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10297_ vdd rf_ram.memory\[522\]\[1\] clknet_leaf_269_clk vss _00041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06159__A2 vss _01687_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1243 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07108__A1 vss _03126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_300 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_474 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_940 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05410_ _01606_ _01605_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08608__A1 vss _02731_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_126_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06390_ _02019_ rf_ram.memory\[67\]\[1\] vdd vss _02585_ rf_ram.memory\[66\]\[1\]
+ _01808_ _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__09678__C vss _04760_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05341_ _01537_ vss vdd _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__06095__A1 vss _01350_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07831__A2 vss _03234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_656 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05272_ vdd vss _01471_ cpu.ctrl.pc cpu.ctrl.pc_plus_4_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08060_ vdd vss _03725_ rf_ram.memory\[564\]\[1\] _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_148_1193 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07011_ vdd _03067_ _03065_ _00137_ _03053_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07595__A1 vss _03422_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08962_ vdd vss _04297_ rf_ram.memory\[11\]\[1\] _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08893_ vdd vss _04255_ rf_ram.memory\[127\]\[0\] _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07913_ vdd vss _03632_ rf_ram.memory\[443\]\[1\] _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07844_ vdd _03589_ _03588_ _00448_ _03587_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07347__A1 vss _03260_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07775_ vdd vss _03546_ rf_ram.memory\[374\]\[1\] _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08847__A1 vss _04202_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06726_ vdd _02872_ _02870_ _00047_ _02826_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09514_ _04643_ vss vdd _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06657_ vdd vss _02823_ _02815_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09445_ vss _01040_ _04598_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_951 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05608_ _01804_ vss vdd _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_52_1169 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_327 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06588_ vdd vss _02769_ rf_ram.memory\[241\]\[1\] _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09376_ _04552_ net211 vdd vss _04560_ net210 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_152 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05539_ _01735_ vss vdd _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08327_ vdd _03890_ _03889_ _00630_ _03884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_172_680 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08258_ vdd _03847_ _03846_ _00604_ _03820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09024__A1 vss net246 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07209_ vdd vss _03194_ rf_ram.memory\[262\]\[1\] _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_162_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_104_279 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10220_ vdd vss _05102_ rf_ram.memory\[23\]\[0\] _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08189_ vdd vss _03805_ _03668_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06389__A2 vss _01918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10151_ vdd _05059_ _05057_ _01286_ _05049_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_30_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10082_ _05017_ _04400_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07338__A1 vss _02958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1014 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05349__B1 vss _01540_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10984_ vdd rf_ram.memory\[165\]\[0\] clknet_leaf_334_clk vss _00721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_266 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07510__A1 vss _03356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06313__A2 vss _01677_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11605_ vss net135 cpu.bne_or_bge vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09263__A1 vss _01484_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11536_ vdd rf_ram.memory\[311\]\[1\] clknet_leaf_148_clk vss _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_382 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_509 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11467_ vdd rf_ram.memory\[342\]\[0\] clknet_leaf_174_clk vss _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09015__A1 vss rf_ram.memory\[10\]\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07577__A1 vss _02882_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10418_ vdd rf_ram.memory\[491\]\[0\] clknet_leaf_183_clk vss _00162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11398_ _01130_ vdd vss clknet_leaf_228_clk net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05547__B vss _01684_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10349_ vdd rf_ram.memory\[301\]\[1\] clknet_leaf_135_clk vss _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05890_ vdd vss _02086_ rf_ram.memory\[68\]\[0\] _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_1095 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_45 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07560_ vdd _03412_ _03410_ _00341_ _03393_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08829__A1 vss _04205_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06511_ _02699_ vdd vss _02700_ cpu.alu.i_rs1 cpu.bufreg.c_r vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_174_901 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09230_ vdd vss _04464_ net249 _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07491_ vdd vss _03370_ rf_ram.memory\[325\]\[1\] _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_614 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_88_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06304__A2 vss _01510_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_115_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06442_ _01563_ vdd vss _02637_ _02634_ _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_146_658 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_850 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09161_ vdd _04421_ _04419_ _00933_ _04401_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06373_ _02004_ vdd vss _02568_ rf_ram.memory\[254\]\[1\] _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_29_686 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09254__A1 vss _01356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06068__A1 vss _01600_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09092_ vdd vss _04378_ net238 _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08112_ vss _03757_ _03689_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_05324_ _01520_ _01519_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_72_987 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_731 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08043_ vdd vss _03714_ rf_ram.memory\[567\]\[1\] _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09006__A1 vss _04301_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05255_ vdd _01454_ _01453_ _01455_ _01442_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07568__A1 vss _03389_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_374 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05291__A2 vss _01434_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05186_ cpu.state.o_cnt\[2\] vdd vss _01386_ cpu.mem_bytecnt\[1\] _01385_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_09994_ vdd vss _04963_ rf_ram.memory\[296\]\[1\] _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06240__A1 vss _01909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09309__A2 vss _01491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08945_ vdd vss _04287_ rf_ram.memory\[449\]\[0\] _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_818 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08876_ vdd _04244_ _04242_ _00825_ _04237_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input22_I vss i_dbus_rdt[28] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07827_ vdd vss _03579_ rf_ram.memory\[412\]\[0\] _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05904__C vss _01670_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07758_ vdd vss _03536_ rf_ram.memory\[376\]\[0\] _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_542 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06288__B vss _01978_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06709_ vdd _02860_ _02859_ _00042_ _02820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_177_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07689_ vdd vss _03493_ _02761_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_603 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05503__B1 vss _01696_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_729 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09428_ vss _01032_ _04589_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09359_ _04540_ net203 vdd vss _04551_ net233 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09245__A1 vss cpu.genblk3.csr.o_new_irq vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_431 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_382 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05806__A1 vss _01552_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11321_ _01054_ vdd vss clknet_leaf_253_clk net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_22_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_5_16__f_clk vdd vss clknet_5_16__leaf_clk clknet_3_4_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_output90_I vss net90 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_694 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_683 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11252_ vdd rf_ram.memory\[109\]\[1\] clknet_leaf_77_clk vss _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05282__A2 vss cpu.alu.i_rs1 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10203_ vdd _05091_ _05089_ _01306_ _05081_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11183_ vdd rf_ram.memory\[575\]\[1\] clknet_leaf_304_clk vss _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10134_ _05049_ _02747_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_24_1079 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10065_ vdd _05006_ _05005_ _01253_ _04982_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06534__A2 vss _01366_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05742__B1 vss _01810_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_35_1131 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10967_ vdd rf_ram.memory\[119\]\[1\] clknet_leaf_71_clk vss _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_647 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10898_ vdd rf_ram.memory\[183\]\[0\] clknet_leaf_13_clk vss _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_1077 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05830__B vss _01551_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_764 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09236__A1 vss _03445_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07798__A1 vss _03554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11519_ vdd rf_ram.memory\[507\]\[0\] clknet_leaf_201_clk vss _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_374 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_193 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06991_ vss _03055_ _02765_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_147_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05942_ vdd vss _02138_ rf_ram.memory\[33\]\[0\] _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08730_ vdd vss _04153_ _03134_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05873_ _01783_ vdd vss _02069_ rf_ram.memory\[250\]\[0\] _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08661_ vdd _04110_ _04108_ _00744_ _04097_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07612_ vdd _03444_ _03442_ _00361_ _03425_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07722__A1 vss _03488_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_361 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08592_ vss _04067_ _03902_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_07543_ vdd _03402_ _03401_ _00334_ _03389_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08278__A2 vss _02894_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07474_ _03359_ vss vdd _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10085__A2 vss _03035_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_96 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06425_ rf_ram.memory\[108\]\[1\] _02620_ vss vdd rf_ram.memory\[111\]\[1\] _01625_
+ rf_ram.memory\[109\]\[1\] _01702_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09213_ vdd _04453_ _04451_ _00953_ _04434_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09144_ vdd vss _04411_ rf_ram.memory\[90\]\[1\] _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_98_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07789__A1 vss _03039_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_250 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06356_ _01551_ vdd vss _02551_ rf_ram.memory\[232\]\[1\] _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09075_ vdd vss _04368_ rf_ram.memory\[81\]\[1\] _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06287_ rf_ram.memory\[130\]\[1\] _02482_ vss vdd rf_ram.memory\[129\]\[1\] _01610_
+ rf_ram.memory\[131\]\[1\] _01636_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_05307_ vss _01503_ rf_ram.i_raddr\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_16_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08450__A2 vss cpu.state.stage_two_req vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05238_ _01437_ vdd vss _01438_ net134 _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_31_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08026_ vdd vss _03704_ rf_ram.memory\[570\]\[0\] _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05169_ cpu.immdec.imm19_12_20\[7\] _01367_ cpu.immdec.imm24_20\[3\] vdd vss _01372_
+ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__08202__A2 vss _03811_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09977_ vdd _04952_ _04951_ _01219_ _04950_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07961__A1 vss _03654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06764__A2 vss _02899_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08928_ vdd _04276_ _04274_ _00845_ _04269_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08859_ vdd _04233_ _04231_ _00819_ _04205_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05724__B1 vss _01911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1099 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10821_ vdd rf_ram.memory\[546\]\[1\] clknet_leaf_316_clk vss _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_149_260 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10752_ vdd rf_ram.memory\[47\]\[0\] clknet_leaf_128_clk vss _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_556 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07421__I vss _03017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10683_ vdd rf_ram.memory\[416\]\[1\] clknet_leaf_98_clk vss _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09218__A1 vss _04434_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06481__B vss _01525_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_834 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11304_ _01037_ vdd vss clknet_leaf_252_clk net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11235_ vdd cpu.genblk3.csr.mcause3_0\[1\] clknet_leaf_255_clk vss _00971_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_1180 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11166_ vdd rf_ram.memory\[57\]\[0\] clknet_leaf_296_clk vss _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10117_ vdd _05038_ _05037_ _01273_ _05014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07952__A1 vss _02898_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11097_ _00002_ vdd vss clknet_leaf_280_clk cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10048_ vdd vss _04996_ _03445_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_136_1107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05963__B1 vss _01624_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07704__A1 vss _03491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_550 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06210_ vdd vss _02405_ rf_ram.memory\[398\]\[1\] _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_112_1162 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09209__A1 vss net241 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_447 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05494__A2 vss _01687_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07190_ vdd vss _03182_ rf_ram.memory\[473\]\[0\] _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06691__A1 vss _02826_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09459__S vss _04604_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_998 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06141_ rf_ram.memory\[309\]\[1\] _01715_ _01709_ rf_ram.memory\[308\]\[1\] _02336_
+ vss vdd rf_ram.memory\[311\]\[1\] _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA_clkbuf_5_29__f_clk_I vss clknet_3_7_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1224 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06072_ _01615_ vdd vss _02267_ rf_ram.memory\[344\]\[1\] _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__06391__B vss _01978_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1219 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09900_ vdd _04904_ _04902_ _01190_ _04887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08196__A1 vss _03787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09831_ vdd _04862_ _04860_ _01162_ _04840_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06974_ vdd vss _03044_ _02781_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09762_ _04760_ _04819_ vdd vss _04820_ net119 _04766_ net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_05925_ rf_ram.memory\[104\]\[0\] _02121_ vss vdd rf_ram.memory\[107\]\[0\] _01679_
+ rf_ram.memory\[105\]\[0\] _01793_ _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_77_1039 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08713_ vdd _04142_ _04140_ _00764_ _04129_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09693_ vdd vss _04772_ _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_178_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05706__B1 vss _01656_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08644_ vdd _04100_ _04099_ _00737_ _04094_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05856_ _01959_ rf_ram.memory\[235\]\[0\] vdd vss _02052_ rf_ram.memory\[234\]\[0\]
+ _01940_ _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08575_ vdd _04055_ _04054_ _00713_ _04023_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05787_ _01923_ vdd vss _01983_ rf_ram.memory\[136\]\[0\] _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07526_ vdd vss _03392_ rf_ram.memory\[361\]\[0\] _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_166_517 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10058__A2 vss _03158_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08120__A1 vss _02728_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07457_ vdd vss _03348_ rf_ram.memory\[330\]\[1\] _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_146_274 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06682__A1 vss _02826_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06408_ _02590_ _02602_ _01362_ vdd vss _02603_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_07388_ vdd vss _03305_ rf_ram.memory\[24\]\[1\] _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09127_ _04400_ _02747_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06339_ _02530_ _02533_ vdd vss _02534_ _02522_ _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__09620__A1 vss _04643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06434__A1 vss _01350_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09058_ vdd vss _04357_ rf_ram.memory\[101\]\[1\] _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output176_I vss net176 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06985__A2 vss _02889_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08009_ _03693_ vss vdd _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_25_1141 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09923__A2 vss _03009_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_697 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06198__B1 vss _01721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09384__B1 vss _04564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11020_ vdd rf_ram.memory\[153\]\[0\] clknet_leaf_330_clk vss _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07934__A1 vss _03622_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05645__B vss _01526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_640 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_854 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10804_ vdd rf_ram.memory\[554\]\[0\] clknet_leaf_321_clk vss _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05380__B vss _01506_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07151__I vss _03013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08111__A1 vss _03754_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10735_ vdd rf_ram.memory\[441\]\[1\] clknet_leaf_77_clk vss _00479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_937 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08662__A2 vss _04078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_520 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10666_ vdd rf_ram.memory\[396\]\[0\] clknet_leaf_94_clk vss _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06673__A1 vss _02826_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10597_ vdd rf_ram.memory\[358\]\[1\] clknet_leaf_155_clk vss _00341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_992 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05228__A2 vss _01411_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput109 o_dbus_dat[1] net109 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_120_163 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_1106 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11218_ vdd rf_ram.memory\[67\]\[0\] clknet_leaf_58_clk vss _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07925__A1 vss _02774_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11149_ vdd rf_ram.memory\[106\]\[1\] clknet_leaf_69_clk vss _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput80 o_dbus_adr[23] net80 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput91 o_dbus_adr[4] net91 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06728__A2 vss _02846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05400__A2 vss _01367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05710_ _01902_ _01904_ _01905_ _01670_ vdd vss _01906_ _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_76_1050 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06690_ vdd vss _02849_ rf_ram.memory\[525\]\[1\] _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_156_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_153_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07153__A2 vss _03158_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05641_ rf_ram.memory\[506\]\[0\] _01837_ vss vdd rf_ram.memory\[505\]\[0\] _01715_
+ rf_ram.memory\[507\]\[0\] _01654_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__08350__A1 vss _03884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05164__A1 vss _01363_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_325 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08360_ vdd _03911_ _03910_ _00642_ _03884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07061__I vss _03100_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05572_ _01768_ _01660_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_07311_ vss _03257_ _03013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__08102__A1 vss _03724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06113__B1 vss _01645_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08291_ vdd vss _03868_ rf_ram.memory\[192\]\[1\] _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07242_ vdd vss _03214_ rf_ram.memory\[421\]\[0\] _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05467__A2 vss _01662_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_300_clk_I vss clknet_5_7__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06664__A1 vss _02779_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07173_ vdd _03171_ _03169_ _00195_ _03161_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05872__C1 vss _01625_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_423 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06124_ _02318_ _01361_ vdd vss _02319_ _01674_ _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__08405__A2 vss _03903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06967__A2 vss _02830_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_631 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_315_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_275 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06055_ _02246_ _02249_ vdd vss _02250_ _02238_ _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_140_995 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_140_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_859 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09814_ vdd _04852_ _04851_ _01155_ _04837_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09745_ vdd vss _04808_ _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06957_ vdd vss _03033_ rf_ram.memory\[230\]\[0\] _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06888_ vdd vss _02987_ rf_ram.memory\[281\]\[1\] _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05908_ rf_ram.memory\[118\]\[0\] _02104_ vss vdd rf_ram.memory\[117\]\[0\] _01931_
+ rf_ram.memory\[119\]\[0\] _01911_ _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_97_905 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09676_ vdd vss _04759_ cpu.bufreg2.o_sh_done_r _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05839_ rf_ram.memory\[204\]\[0\] _02035_ vss vdd rf_ram.memory\[207\]\[0\] _01925_
+ rf_ram.memory\[205\]\[0\] _01912_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__08341__A1 vss _03892_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08627_ vdd _04089_ _04088_ _00731_ _04058_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08892__A2 vss _04038_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08558_ vdd vss _04045_ _02865_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_77_662 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08067__I vss _03692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07509_ vdd vss _03381_ rf_ram.memory\[323\]\[0\] _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08489_ vdd vss _03999_ rf_ram.memory\[369\]\[0\] _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_550 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_65_835 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09841__A1 vss _02714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_687 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10520_ vdd rf_ram.memory\[252\]\[0\] clknet_leaf_224_clk vss _00264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06655__A1 vss _02779_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10451_ vdd rf_ram.memory\[495\]\[1\] clknet_leaf_184_clk vss _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05863__C1 vss _01968_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09444__I1 vss net73 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10382_ vdd rf_ram.memory\[426\]\[0\] clknet_leaf_100_clk vss _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_264 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05630__A2 vss _01697_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07907__A1 vss _03619_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11003_ vdd rf_ram.memory\[161\]\[1\] clknet_leaf_338_clk vss _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05375__B vss _01506_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08580__A1 vss net250 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09361__I vss _04539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08883__A2 vss _04248_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_314 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06894__A1 vss _02975_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_184_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_95_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09832__A1 vss _03668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_194 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06646__A1 vss _02736_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10718_ vdd rf_ram.memory\[446\]\[0\] clknet_leaf_78_clk vss _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09310__B vss _03967_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_873 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10649_ vdd rf_ram.memory\[382\]\[1\] clknet_leaf_109_clk vss _00393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_69 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08399__A1 vss _03922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_236 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09060__A2 vss _04339_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05606__C1 vss _01721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07071__A1 vss _03092_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07860_ vdd _03599_ _03598_ _00454_ _03587_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_1112 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07791_ vdd _03556_ _03555_ _00428_ _03554_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06811_ vdd vss _02934_ rf_ram.memory\[290\]\[1\] _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05385__A1 vss _01495_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06031__C1 vss _01555_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1178 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09530_ vdd vss _04657_ cpu.immdec.imm19_12_20\[1\] _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06742_ vdd vss _02884_ _02881_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07126__A2 vss _02997_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09461_ _04604_ vdd vss _04607_ net80 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06673_ vdd _02835_ _02833_ _00031_ _02826_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_184_clk vdd vss clknet_leaf_184_clk clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06334__B1 vss _02019_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05688__A2 vss _01697_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06885__A1 vss _02958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05624_ _01819_ vdd vss _01820_ _01675_ _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08412_ vdd _03943_ _03942_ _00662_ _03919_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05304__I vss _01499_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09392_ _04564_ net219 vdd vss _04569_ net218 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_301 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05555_ _01747_ _01750_ vdd vss _01751_ _01738_ _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_08343_ vdd _03900_ _03899_ _00636_ _03884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_58_161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_149_1106 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06637__A1 vss _02801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06098__C1 vss _01678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08274_ vdd vss _03858_ rf_ram.memory\[195\]\[0\] _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07225_ vdd _03203_ _03201_ _00215_ _03193_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_531 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_756 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05845__C1 vss _01713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05486_ _01682_ _01508_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_27_570 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_378 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_80_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_254_clk_I vss clknet_5_20__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_299 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07156_ _03161_ _03017_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_89_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05860__A2 vss _01958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07062__A1 vss _03082_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06107_ _01746_ vdd vss _02302_ _02299_ _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07087_ vdd vss _03117_ _02775_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_30_746 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input52_I vss i_ibus_rdt[27] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06038_ vdd _01351_ _02232_ _02233_ _02227_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_269_clk_I vss clknet_5_16__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08562__A1 vss _04026_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07989_ vdd vss _03679_ _03672_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09728_ _04791_ _04796_ vdd vss _04797_ net107 _04790_ net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
Xclkbuf_leaf_175_clk vdd vss clknet_leaf_175_clk clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_96_234 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09659_ _04744_ _04740_ vdd vss _04745_ net120 _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_171_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05679__A2 vss _01801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_870 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_207_clk_I vss clknet_5_24__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11621_ vss net143 net71 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_857 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_183 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06628__A1 vss _02797_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09814__A1 vss _04837_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11552_ vdd rf_ram.memory\[452\]\[1\] clknet_leaf_112_clk vss _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_361 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11483_ vdd rf_ram.memory\[295\]\[0\] clknet_leaf_139_clk vss _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10503_ vdd rf_ram.memory\[257\]\[1\] clknet_leaf_202_clk vss _00247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09417__I1 vss net90 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10434_ vdd rf_ram.memory\[4\]\[0\] clknet_leaf_211_clk vss _00178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10188__A1 vss _05081_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05851__A2 vss _01501_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09557__S vss _03967_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10365_ vdd rf_ram.memory\[297\]\[1\] clknet_leaf_138_clk vss _00109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_60_370 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06261__C1 vss _01645_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1201 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06800__A1 vss _02876_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10296_ vdd rf_ram.memory\[522\]\[0\] clknet_leaf_269_clk vss _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08553__A1 vss net249 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06013__C1 vss _01539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05833__B vss _01928_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08305__A1 vss _03852_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10112__A1 vss _05014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1042 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06867__A1 vss _02935_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_158_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_637 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05340_ _01536_ vss vdd _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08608__A2 vss _02939_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06619__A1 vss _02748_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_624 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1182 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06095__A2 vss _02278_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07292__A1 vss _03222_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05271_ vdd vss _01470_ cpu.state.cnt_r\[2\] _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_183_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_126_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10179__A1 vss _05046_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05842__A2 vss _01662_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07010_ vdd vss _03067_ rf_ram.memory\[223\]\[1\] _03065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09467__S vss _04604_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_567 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07044__A1 vss _02829_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08792__A1 vss net246 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08961_ vdd _04296_ _04295_ _00858_ _04266_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08892_ vdd vss _04254_ _02908_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07912_ vdd _03631_ _03630_ _00474_ _03619_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07843_ vdd vss _03589_ rf_ram.memory\[431\]\[0\] _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07774_ vdd _03545_ _03544_ _00422_ _03521_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_157_clk vdd vss clknet_leaf_157_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06725_ vdd vss _02872_ rf_ram.memory\[51\]\[1\] _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09513_ vdd vss _04642_ _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06858__A1 vss _02930_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09444_ _04593_ vdd vss _04598_ net72 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06656_ _02822_ _02821_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_05607_ _01800_ _01802_ vdd vss _01803_ _01797_ _01798_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_78_289 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06587_ vdd _02768_ _02767_ _00012_ _02743_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09375_ vdd vss _04559_ _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_163_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08326_ vdd vss _03890_ rf_ram.memory\[21\]\[0\] _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05538_ vdd _01733_ _01732_ _01734_ _01347_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_304 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06086__A2 vss _01711_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05469_ rf_ram.memory\[372\]\[0\] _01665_ vss vdd rf_ram.memory\[375\]\[0\] _01519_
+ rf_ram.memory\[373\]\[0\] _01664_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_08257_ vdd vss _03847_ rf_ram.memory\[526\]\[0\] _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_73_clk_I vss clknet_5_10__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_90 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07208_ _03193_ _03017_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_3_5_0_clk clknet_3_5_0_clk vss vdd clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08188_ vdd _03804_ _03802_ _00577_ _03790_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_860 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1245 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09024__A2 vss _04303_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07139_ vdd vss _03150_ rf_ram.memory\[498\]\[1\] _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1211 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10150_ vdd vss _05059_ rf_ram.memory\[451\]\[1\] _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_88_clk_I vss clknet_5_11__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10081_ vdd _05016_ _05015_ _01259_ _05014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07338__A2 vss _02972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_131_clk_I vss clknet_5_24__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08535__A1 vss _04026_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06010__A2 vss _01532_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_11_clk_I vss clknet_5_2__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05145__S vss _01347_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_148_clk vdd vss clknet_leaf_148_clk clknet_5_26__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_134_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10983_ vdd rf_ram.memory\[166\]\[1\] clknet_leaf_331_clk vss _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_146_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06849__A1 vss _02958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_26_clk_I vss clknet_5_3__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_957 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_1003 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_637 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139_199 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06484__B vss _01503_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_531 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11604_ vss net125 cpu.bufreg2.o_sh_done_r vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11535_ vdd rf_ram.memory\[311\]\[0\] clknet_leaf_146_clk vss _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06077__A2 vss _01697_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_320_clk vdd vss clknet_leaf_320_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_25_337 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06482__C1 vss _01653_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05824__A2 vss _01940_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11466_ vdd rf_ram.memory\[343\]\[1\] clknet_leaf_168_clk vss _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07026__A1 vss _03050_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07577__A2 vss _03390_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10417_ vdd rf_ram.memory\[492\]\[1\] clknet_leaf_182_clk vss _00161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11397_ _01129_ vdd vss clknet_leaf_228_clk net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__06234__C1 vss _01656_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10348_ vdd rf_ram.memory\[301\]\[0\] clknet_leaf_134_clk vss _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08774__A1 vss _04167_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10279_ vdd rf_ram.memory\[293\]\[1\] clknet_leaf_137_clk vss _00023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05563__B vss _01629_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06001__A2 vss _01524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_206 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_139_clk vdd vss clknet_leaf_139_clk clknet_5_27__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_45_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07490_ vdd _03369_ _03368_ _00314_ _03356_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_1200 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06510_ vdd _01381_ cpu.decode.opcode\[1\] _02699_ _01382_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06441_ _01607_ rf_ram.memory\[43\]\[1\] vdd vss _02636_ rf_ram.memory\[42\]\[1\]
+ _01605_ _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_29_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_795 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_1073 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_979 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09160_ vdd vss _04421_ rf_ram.memory\[88\]\[1\] _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06372_ _02565_ _02566_ vdd vss _02567_ _02563_ _02564_ _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07265__A1 vss _03222_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05323_ vdd vss _01519_ _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
X_08111_ vdd _03756_ _03755_ _00548_ _03754_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09091_ vdd _04377_ _04375_ _00907_ _04367_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05815__A2 vss _01799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_476 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05254_ net98 vss vdd net128 net105 _01376_ net114 _01375_ _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_9_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08042_ vdd _03713_ _03712_ _00522_ _03686_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_311_clk vdd vss clknet_leaf_311_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07017__A1 vss _02750_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05185_ _01385_ cpu.mem_bytecnt\[0\] vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05579__A1 vss _01769_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09993_ vdd _04962_ _04961_ _01225_ _04950_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08944_ vdd vss _04286_ _03672_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09309__A3 vss _04013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1197 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08875_ vdd vss _04244_ rf_ram.memory\[12\]\[1\] _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07826_ vdd vss _03578_ _02839_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07757_ vdd vss _03535_ _02991_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05751__A1 vss _01674_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input15_I vss i_dbus_rdt[21] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06708_ vdd vss _02860_ rf_ram.memory\[521\]\[0\] _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07688_ vdd _03492_ _03489_ _00389_ _03491_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_48_930 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_795 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06639_ vdd _02808_ _02807_ _00024_ _02743_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09427_ _02707_ vdd vss _04589_ net94 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09358_ vdd vss _04550_ _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_19_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_34_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09245__A2 vss _01413_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06059__A2 vss _01649_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08309_ vdd vss _03879_ rf_ram.memory\[243\]\[0\] _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_123 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09289_ vdd vss _04509_ rf_ram.memory\[65\]\[0\] _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_302_clk vdd vss clknet_leaf_302_clk clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11320_ _01053_ vdd vss clknet_leaf_264_clk net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_166_1091 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11251_ vdd rf_ram.memory\[109\]\[0\] clknet_leaf_70_clk vss _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05648__B vss _01660_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10202_ vdd vss _05091_ rf_ram.memory\[191\]\[1\] _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output83_I vss net83 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11182_ vdd rf_ram.memory\[575\]\[0\] clknet_leaf_303_clk vss _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06231__A2 vss _01623_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10133_ vdd _05048_ _05047_ _01279_ _05046_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_140_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10064_ vdd vss _05006_ rf_ram.memory\[307\]\[0\] _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05990__A1 vss _02102_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06479__B vss _01503_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_526 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_228 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10966_ vdd rf_ram.memory\[119\]\[0\] clknet_leaf_71_clk vss _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07495__A1 vss _03356_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10897_ vdd rf_ram.memory\[182\]\[1\] clknet_leaf_13_clk vss _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06298__A2 vss _01958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09236__A2 vss _02909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06455__C1 vss _01655_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11518_ vdd rf_ram.memory\[34\]\[1\] clknet_leaf_200_clk vss _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_115 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_515 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11449_ vdd rf_ram.memory\[239\]\[0\] clknet_leaf_276_clk vss _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_548 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1148 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08747__A1 vss net242 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06222__A2 vss _01777_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06990_ vdd _03054_ _03051_ _00129_ _03053_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_186_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input7_I vss i_dbus_rdt[14] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05941_ _01550_ vdd vss _02137_ rf_ram.memory\[32\]\[0\] _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09172__A1 vss _03071_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05872_ rf_ram.memory\[252\]\[0\] _02068_ vss vdd rf_ram.memory\[255\]\[0\] _01625_
+ rf_ram.memory\[253\]\[0\] _01678_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_08660_ vdd vss _04110_ rf_ram.memory\[15\]\[1\] _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07611_ vdd vss _03444_ rf_ram.memory\[353\]\[1\] _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_163_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07999__I vss _02742_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08591_ vdd _04066_ _04064_ _00718_ _04062_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_3_4_0_clk_I vss clknet_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07542_ vdd vss _03402_ rf_ram.memory\[320\]\[0\] _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_152_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_5_22__f_clk vdd vss clknet_5_22__leaf_clk clknet_3_5_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07473_ vdd _03358_ _03357_ _00308_ _03356_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06289__A2 vss _01770_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06424_ _02004_ vdd vss _02619_ rf_ram.memory\[110\]\[1\] _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09212_ vdd vss _04453_ rf_ram.memory\[68\]\[1\] _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07238__A1 vss _03190_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_938 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09143_ vdd _04410_ _04409_ _00926_ _04397_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06355_ _02549_ vdd vss _02550_ _01951_ _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_16_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07789__A2 vss _03135_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08986__A1 vss _04301_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09719__I vss _04766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05306_ vss _01502_ _01501_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06286_ _01923_ vdd vss _02481_ rf_ram.memory\[128\]\[1\] _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09074_ _04367_ _04061_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05237_ rf_ram_if.rtrig1 vdd vss _01437_ rf_ram.rdata\[0\] _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_08025_ vdd vss _03703_ _02813_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05168_ vdd vss _01371_ _01369_ _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08738__A1 vss _01369_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07410__A1 vss _03292_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06213__A2 vss _01692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09976_ vdd vss _04952_ rf_ram.memory\[274\]\[0\] _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08927_ vdd vss _04276_ rf_ram.memory\[124\]\[1\] _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08858_ vdd vss _04233_ rf_ram.memory\[131\]\[1\] _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07809_ vdd vss _03568_ rf_ram.memory\[414\]\[1\] _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_19_1138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08789_ vdd _04190_ _04189_ _00792_ _04167_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10820_ vdd rf_ram.memory\[546\]\[0\] clknet_leaf_316_clk vss _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07477__A1 vss _03360_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10751_ vdd rf_ram.memory\[470\]\[1\] clknet_leaf_51_clk vss _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_94_321 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10682_ vdd rf_ram.memory\[416\]\[0\] clknet_leaf_97_clk vss _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_955 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08977__A1 vss _03134_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06437__C1 vss _01607_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1103 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06452__A2 vss _01633_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1158 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11303_ _01036_ vdd vss clknet_leaf_252_clk net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11234_ vdd cpu.genblk3.csr.mcause3_0\[0\] clknet_leaf_256_clk vss _00970_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_30_181 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06204__A2 vss _01649_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11165_ vdd rf_ram.memory\[81\]\[1\] clknet_leaf_47_clk vss _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06988__I vss _03017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07401__A1 vss _03309_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10116_ vdd vss _05038_ rf_ram.memory\[373\]\[0\] _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11096_ vdd rf_ram.memory\[127\]\[1\] clknet_leaf_84_clk vss _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07952__A2 vss _03158_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10047_ vdd _04995_ _04993_ _01246_ _04985_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08901__A1 vss _04237_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05841__B vss _01916_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10949_ vdd rf_ram.memory\[359\]\[1\] clknet_leaf_154_clk vss _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07468__A1 vss _03326_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_540 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_70_clk vdd vss clknet_leaf_70_clk clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_128_467 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09209__A2 vss _04418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_944 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06140_ _01707_ vdd vss _02335_ rf_ram.memory\[310\]\[1\] _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_101_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07640__A1 vss _03458_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06071_ _02265_ vdd vss _02266_ _01675_ _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06443__A2 vss _01682_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09475__S vss _04604_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_890 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09830_ vdd vss _04862_ rf_ram.memory\[62\]\[1\] _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05254__I0 vss net98 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06973_ vdd _03043_ _03041_ _00123_ _03018_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09761_ vdd vss _04819_ _04804_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_1231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09145__A1 vss _04401_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05924_ _01783_ vdd vss _02120_ rf_ram.memory\[106\]\[0\] _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_77_1029 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08712_ vdd vss _04142_ rf_ram.memory\[151\]\[1\] _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09692_ _04768_ _04771_ vdd vss _04772_ net127 _04767_ net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__05307__I vss rf_ram.i_raddr\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08643_ vdd vss _04100_ rf_ram.memory\[519\]\[0\] _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05855_ vdd vss _02051_ rf_ram.memory\[233\]\[0\] _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__05751__B vss _01946_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08574_ vdd vss _04055_ rf_ram.memory\[16\]\[0\] _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05786_ _01981_ vdd vss _01982_ _01909_ _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_07525_ vdd vss _03391_ _02752_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07459__A1 vss _02954_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_570 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1074 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_321 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_61_clk vdd vss clknet_leaf_61_clk clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_92_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_302 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_899 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08120__A2 vss _03729_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_218 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07456_ vdd _03347_ _03346_ _00302_ _03323_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_1136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06407_ _02596_ _01660_ _02601_ vdd vss _02602_ _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_07387_ vdd _03304_ _03303_ _00276_ _03289_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_29_292 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09126_ vdd _04399_ _04398_ _00920_ _04397_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08959__A1 vss net246 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06338_ _02532_ vdd vss _02533_ _01972_ _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09057_ vdd _04356_ _04355_ _00894_ _04331_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06269_ rf_ram.memory\[157\]\[1\] _01968_ _01614_ rf_ram.memory\[156\]\[1\] _02464_
+ vss vdd rf_ram.memory\[159\]\[1\] _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_130_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_846 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08008_ _02762_ vdd vss _03692_ _02730_ _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_124_1056 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09959_ vdd vss _04941_ _04911_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09136__A1 vss net249 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10803_ vdd rf_ram.memory\[555\]\[1\] clknet_leaf_322_clk vss _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_170_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_52_clk vdd vss clknet_leaf_52_clk clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10734_ vdd rf_ram.memory\[441\]\[0\] clknet_leaf_77_clk vss _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07870__A1 vss _03587_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10665_ vdd rf_ram.memory\[378\]\[1\] clknet_leaf_109_clk vss _00409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06492__B vss _01372_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_63_571 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10596_ vdd rf_ram.memory\[358\]\[0\] clknet_leaf_155_clk vss _00340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06425__A2 vss _01634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1123 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142_1178 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11217_ vdd rf_ram.memory\[68\]\[1\] clknet_leaf_64_clk vss _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput70 o_dbus_adr[13] net70 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07925__A2 vss _02832_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11148_ vdd rf_ram.memory\[106\]\[0\] clknet_leaf_67_clk vss _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput81 o_dbus_adr[24] net81 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput92 o_dbus_adr[5] net92 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05936__A1 vss _01903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11079_ vdd rf_ram.memory\[132\]\[0\] clknet_leaf_14_clk vss _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07689__A1 vss _02761_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05640_ _01756_ vdd vss _01836_ rf_ram.memory\[504\]\[0\] _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_76_1095 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05164__A2 vss _01366_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05571_ _01766_ _01361_ vdd vss _01767_ _01674_ _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_53_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07310_ vdd _03256_ _03254_ _00247_ _03225_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_43_clk vdd vss clknet_leaf_43_clk clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_129_765 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08290_ vdd _03867_ _03866_ _00616_ _03852_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_324 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07241_ vdd vss _03213_ _02795_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_50_1279 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07172_ vdd vss _03171_ rf_ram.memory\[495\]\[1\] _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05872__B1 vss _01678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06416__A2 vss _01915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06123_ _01349_ _02317_ vdd vss _02318_ _02309_ _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_125_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_390 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06054_ _02248_ vdd vss _02249_ _01527_ _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09813_ vdd vss _04852_ rf_ram.memory\[7\]\[0\] _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06719__A3 vss _02730_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09744_ _04791_ _04807_ vdd vss _04808_ net113 _04790_ net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06956_ vdd vss _03032_ _02766_ _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06887_ vdd _02986_ _02985_ _00094_ _02970_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05907_ vdd vss _02103_ rf_ram.memory\[116\]\[0\] _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_97_928 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09675_ vdd vss _04758_ net124 _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_05838_ vdd vss _02034_ rf_ram.memory\[206\]\[0\] _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_68_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08341__A2 vss _03009_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08626_ vdd vss _04089_ rf_ram.memory\[539\]\[0\] _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_449 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06296__C vss _01362_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06352__A1 vss _01674_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05155__A2 vss cpu.decode.co_ebreak vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08557_ vdd _04044_ _04042_ _00706_ _04026_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_34_clk vdd vss clknet_leaf_34_clk clknet_5_6__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05769_ _01953_ rf_ram.memory\[147\]\[0\] vdd vss _01965_ rf_ram.memory\[146\]\[0\]
+ _01958_ _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_175_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07508_ vdd vss _03380_ _03319_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08488_ vdd vss _03998_ net248 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_730 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07852__A1 vss _03590_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07439_ vdd vss _03337_ _02921_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10450_ vdd rf_ram.memory\[495\]\[0\] clknet_leaf_184_clk vss _00194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05863__B1 vss _01959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09109_ vdd _04388_ _04387_ _00914_ _04364_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05500__I vss _01695_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10381_ vdd rf_ram.memory\[427\]\[1\] clknet_leaf_100_clk vss _00125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_1128 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09357__A1 vss net232 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09357__B2 vss net233 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11002_ vdd rf_ram.memory\[161\]\[0\] clknet_5_0__leaf_clk vss _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09109__A1 vss _04364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1173 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05394__A2 vss _01544_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08580__A2 vss _03949_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_265 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05391__B vss _01506_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_25_clk vdd vss clknet_leaf_25_clk clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_138_540 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_622 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06646__A2 vss _02799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10717_ vdd rf_ram.memory\[463\]\[1\] clknet_leaf_51_clk vss _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09832__A2 vss _02960_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_125_245 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10648_ vdd rf_ram.memory\[382\]\[0\] clknet_leaf_109_clk vss _00392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05410__I vss _01605_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1039 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10579_ vdd rf_ram.memory\[323\]\[1\] clknet_leaf_159_clk vss _00323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05606__B1 vss _01726_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_298 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_473 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05566__B vss _01526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1095 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08020__A1 vss _02822_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05909__A1 vss _01909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06031__B1 vss _01554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07790_ vdd vss _03556_ rf_ram.memory\[436\]\[0\] _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06810_ vdd _02933_ _02932_ _00070_ _02927_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06582__A1 vss cpu.immdec.imm11_7\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_917 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06741_ _02883_ vss vdd net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09460_ vss _01047_ _04606_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_613 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06672_ vdd vss _02835_ rf_ram.memory\[455\]\[1\] _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08411_ vdd vss _03943_ rf_ram.memory\[177\]\[0\] _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06885__A2 vss _02984_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05623_ rf_ram.memory\[493\]\[0\] _01793_ _01677_ rf_ram.memory\[492\]\[0\] _01819_
+ vss vdd rf_ram.memory\[495\]\[0\] _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
Xclkbuf_leaf_16_clk vdd vss clknet_leaf_16_clk clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_961 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09391_ vdd vss _04568_ _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_171_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05554_ _01749_ vdd vss _01750_ _01603_ _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08342_ vdd vss _03900_ rf_ram.memory\[214\]\[0\] _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08087__A1 vss _03724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05485_ _01680_ vdd vss _01681_ _01675_ _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__06637__A2 vss _02806_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06098__B1 vss _01679_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08273_ vdd vss _03857_ _03230_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_74_644 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07224_ vdd vss _03203_ rf_ram.memory\[425\]\[1\] _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05845__B1 vss _01721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_407 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05320__I vss _01515_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_13__f_clk_I vss clknet_3_3_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07155_ vdd _03160_ _03159_ _00188_ _03157_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07062__A2 vss _03101_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06106_ _01679_ rf_ram.memory\[283\]\[1\] vdd vss _02301_ rf_ram.memory\[282\]\[1\]
+ _01687_ _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_07086_ vdd _03116_ _03114_ _00163_ _03092_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_73_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05476__B vss _01660_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_793 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_473 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06037_ _02231_ _01564_ vdd vss _02232_ _02228_ _02229_ _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_121_1037 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input45_I vss i_ibus_rdt[20] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_482 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07988_ vdd _03678_ _03676_ _00503_ _03654_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06573__A1 vss _02748_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05376__A2 vss _01511_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09727_ vdd vss _04796_ _04781_ net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06939_ vdd vss _03022_ rf_ram.memory\[228\]\[1\] _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09511__A1 vss _04637_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05781__C1 vss _01610_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06100__B vss _01615_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09658_ _04743_ vdd vss _04744_ _04737_ _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_166_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08609_ _04078_ vss vdd _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_09589_ vdd vss _04701_ _03967_ _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_49_151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_182_605 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11620_ vss net142 net70 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08078__A1 vss _02945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07825__A1 vss _03557_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11551_ vdd rf_ram.memory\[452\]\[0\] clknet_leaf_111_clk vss _01283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06628__A2 vss _02799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10502_ vdd rf_ram.memory\[257\]\[0\] clknet_leaf_202_clk vss _00246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11482_ vdd rf_ram.memory\[335\]\[1\] clknet_leaf_167_clk vss _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_338 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_395 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_535 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10433_ vdd rf_ram.memory\[487\]\[1\] clknet_leaf_225_clk vss _00177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_568 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10364_ vdd rf_ram.memory\[297\]\[0\] clknet_leaf_138_clk vss _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08250__A1 vss _03823_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06261__B1 vss _01646_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05386__B vss _01505_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10295_ vdd rf_ram.memory\[523\]\[1\] clknet_leaf_269_clk vss _00039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08553__A2 vss _03158_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09750__B2 vss net116 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09750__A1 vss net115 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06013__B1 vss _01540_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_3__f_clk vdd vss clknet_5_3__leaf_clk clknet_3_0_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05405__I vss rf_ram.i_raddr\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06010__B vss _01505_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06867__A2 vss _02972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_961 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_314_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07816__A1 vss _02959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_329_clk_I vss clknet_5_4__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_316 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_636 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05270_ vss _01469_ cpu.decode.opcode\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_153_384 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09569__A1 vss _04478_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07044__A2 vss _03089_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08241__A1 vss _03668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_933 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08792__A2 vss _04152_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08960_ vdd vss _04296_ rf_ram.memory\[11\]\[0\] _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_5_clk vdd vss clknet_leaf_5_clk clknet_5_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08891_ vdd _04253_ _04251_ _00831_ _04237_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07911_ vdd vss _03631_ rf_ram.memory\[443\]\[0\] _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07842_ vdd vss _03588_ _02953_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_155_1111 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06555__A1 vss _01353_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05743__C vss _01658_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07773_ vdd vss _03545_ rf_ram.memory\[374\]\[0\] _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_155_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09512_ _04473_ vdd vss _04642_ cpu.genblk3.csr.timer_irq_r _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_78_213 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06724_ vdd _02871_ _02870_ _00046_ _02820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05315__I vss _01510_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1176 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09443_ vss _01039_ _04597_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06655_ vdd vss _02821_ _02779_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_05606_ rf_ram.memory\[306\]\[0\] _01802_ vss vdd rf_ram.memory\[305\]\[0\] _01721_
+ rf_ram.memory\[307\]\[0\] _01726_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09374_ _04552_ net210 vdd vss _04559_ net209 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_136_307 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08325_ vdd vss _03889_ _03035_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06586_ vdd vss _02768_ rf_ram.memory\[241\]\[0\] _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_986 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05537_ vdd vss _01733_ cpu.immdec.imm24_20\[2\] _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_368 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05468_ _01664_ vss vdd _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08256_ vdd vss _03846_ _02845_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__08480__A1 vss _02713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07207_ vdd _03192_ _03191_ _00208_ _03190_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_90_989 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08187_ vdd vss _03804_ rf_ram.memory\[540\]\[1\] _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_160_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_557 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07138_ vdd _03149_ _03148_ _00182_ _03123_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05399_ vss _01595_ cpu.immdec.imm19_12_20\[7\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__06243__B1 vss _01857_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09980__A1 vss _04953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07069_ vdd _03106_ _03105_ _00156_ _03087_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06794__A1 vss _02773_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10080_ vdd vss _05016_ rf_ram.memory\[350\]\[0\] _05015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output151_I vss net151 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05349__A2 vss _01544_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06546__B2 vss _01347_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10982_ vdd rf_ram.memory\[166\]\[0\] clknet_leaf_331_clk vss _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06849__A2 vss _02960_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_925 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09799__A1 vss _04837_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11534_ vdd rf_ram.memory\[351\]\[1\] clknet_leaf_191_clk vss _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08471__A1 vss _02714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_682 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11465_ vdd rf_ram.memory\[343\]\[0\] clknet_leaf_168_clk vss _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06482__B1 vss _01714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_308 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10416_ vdd rf_ram.memory\[492\]\[0\] clknet_leaf_182_clk vss _00160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1189 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08223__A1 vss _03820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06234__B1 vss _01763_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11396_ _01128_ vdd vss clknet_leaf_226_clk net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05588__A2 vss _01782_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10347_ vdd rf_ram.memory\[282\]\[1\] clknet_leaf_179_clk vss _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09971__A1 vss _04918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1021 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06005__B vss _01505_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10278_ vdd rf_ram.memory\[293\]\[0\] clknet_leaf_136_clk vss _00022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05844__B vss _01805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09574__I1 vss net54 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_253_clk_I vss clknet_5_20__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10097__A1 vss _05014_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06440_ vdd vss _02635_ rf_ram.memory\[41\]\[1\] _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_0_36 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05512__A2 vss _01706_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06170__C1 vss _01636_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06371_ rf_ram.memory\[242\]\[1\] _02566_ vss vdd rf_ram.memory\[241\]\[1\] _01702_
+ rf_ram.memory\[243\]\[1\] _01625_ _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_12_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17_817 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_268_clk_I vss clknet_5_16__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_72_967 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05322_ vdd vss _01518_ _01512_ _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_16_349 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08110_ vdd vss _03756_ rf_ram.memory\[554\]\[0\] _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09090_ vdd vss _04377_ rf_ram.memory\[569\]\[1\] _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06473__B1 vss _01624_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_1278 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05253_ cpu.mem_bytecnt\[1\] vdd vss _01453_ _01385_ _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08041_ vdd vss _03713_ rf_ram.memory\[567\]\[0\] _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_101_50 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_3_0_0_clk_I vss clknet_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10021__A1 vss _03309_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05184_ vdd vss cpu.state.cnt_r\[0\] _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_09992_ vdd vss _04962_ rf_ram.memory\[296\]\[0\] _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_588 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06776__A1 vss _02779_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08943_ vdd _04285_ _04283_ _00851_ _04269_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_122_1165 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_206_clk_I vss clknet_5_24__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_96 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09714__B2 vss net104 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09714__A1 vss net103 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08874_ vdd _04243_ _04242_ _00824_ _04234_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_36_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07825_ vdd _03577_ _03575_ _00441_ _03557_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05736__C1 vss _01857_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07756_ vdd _03534_ _03532_ _00415_ _03524_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05751__A2 vss _01934_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_706 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06707_ vdd vss _02859_ _02752_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_17_1022 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07687_ vdd vss _03492_ rf_ram.memory\[383\]\[1\] _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09426_ vss _01031_ _04588_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_149_465 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06638_ vdd vss _02808_ rf_ram.memory\[294\]\[0\] _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05503__A2 vss _01687_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07260__I vss _03017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06569_ vdd vss _02753_ _02738_ _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_63_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09357_ _04540_ net233 vdd vss _04550_ net232 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_180_939 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09288_ vdd vss _04508_ net238 _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08308_ vdd vss _03878_ _03309_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08453__A1 vss _01418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output199_I vss net199 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1288 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08239_ vdd vss _03836_ rf_ram.memory\[530\]\[1\] _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05929__B vss _01923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_382 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09402__B1 vss _04564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11250_ _00986_ cpu.immdec.imm11_7\[4\] vdd vss clknet_leaf_279_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XANTENNA__09953__A1 vss _04921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11181_ vdd rf_ram.memory\[93\]\[1\] clknet_leaf_62_clk vss _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10201_ vdd _05090_ _05089_ _01305_ _05078_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10132_ vdd vss _05048_ rf_ram.memory\[454\]\[0\] _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output76_I vss net76 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1149 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08508__A2 vss net134 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10063_ vdd vss _05005_ _03445_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05990__A2 vss _02129_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1150 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05742__A2 vss _01666_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10079__A1 vss _02814_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_330 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_205 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10965_ vdd rf_ram.memory\[171\]\[1\] clknet_leaf_9_clk vss _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10896_ vdd rf_ram.memory\[182\]\[0\] clknet_leaf_13_clk vss _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_1177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08444__A1 vss _02945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_170 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11517_ vdd rf_ram.memory\[34\]\[0\] clknet_leaf_200_clk vss _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10251__A1 vss _02819_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06455__B1 vss _01653_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_343 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_190 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11448_ _01180_ vdd vss clknet_leaf_240_clk cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09944__A1 vss _04911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10003__A1 vss _04950_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11379_ _01111_ vdd vss clknet_leaf_232_clk net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08747__A2 vss _04152_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1273 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05940_ _01563_ vdd vss _02136_ _02133_ _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_179_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_192_clk_I vss clknet_5_30__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09172__A2 vss _04418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07183__A1 vss _03161_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05871_ _02004_ vdd vss _02067_ rf_ram.memory\[254\]\[0\] _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_07610_ vdd _03443_ _03442_ _00360_ _03422_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08590_ vdd vss _04066_ rf_ram.memory\[167\]\[1\] _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07541_ vdd vss _03401_ _03319_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_72_clk_I vss clknet_5_8__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1200 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_4_0_clk clknet_3_4_0_clk vss vdd clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_186_560 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07472_ vdd vss _03358_ rf_ram.memory\[366\]\[0\] _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06143__C1 vss _01721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06423_ _02610_ _02614_ _02617_ _01660_ vdd vss _02618_ _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_09211_ vdd _04452_ _04451_ _00952_ _04431_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09142_ vdd vss _04410_ rf_ram.memory\[90\]\[0\] _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06354_ rf_ram.memory\[237\]\[1\] _01968_ _01614_ rf_ram.memory\[236\]\[1\] _02549_
+ vss vdd rf_ram.memory\[239\]\[1\] _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_173_298 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_130_clk_I vss clknet_5_24__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05305_ _01501_ _01500_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_296_clk vdd vss clknet_leaf_296_clk clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_126_181 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09073_ vdd _04366_ _04365_ _00900_ _04364_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06285_ _02479_ vdd vss _02480_ _01972_ _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA_clkbuf_leaf_10_clk_I vss clknet_5_2__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06997__A1 vss _03055_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_983 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_1205 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05236_ vdd vss _01436_ rf_ram_if.rdata1 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_13_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08024_ vdd _03702_ _03700_ _00515_ _03690_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_145_clk_I vss clknet_5_26__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08738__A2 vss _01496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05167_ vdd vss _01370_ _01338_ _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09975_ vdd vss _04951_ _02922_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA_clkbuf_leaf_25_clk_I vss clknet_5_3__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1014 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08926_ vdd _04275_ _04274_ _00844_ _04266_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05709__C1 vss _01656_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07174__A1 vss _02894_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08857_ vdd _04232_ _04231_ _00818_ _04202_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07808_ vdd _03567_ _03566_ _00434_ _03554_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_220_clk vdd vss clknet_leaf_220_clk clknet_5_22__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05724__A2 vss _01856_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06382__C1 vss _01925_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08788_ vdd vss _04190_ rf_ram.memory\[149\]\[0\] _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07739_ _03524_ _03359_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__05931__C vss _01978_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output114_I vss net114 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10750_ vdd rf_ram.memory\[470\]\[0\] clknet_leaf_51_clk vss _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08674__A1 vss _04094_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10681_ vdd rf_ram.memory\[437\]\[1\] clknet_leaf_80_clk vss _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09409_ _01344_ _01388_ vdd vss _04579_ _01436_ _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_165_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_479 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_619 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08426__A1 vss _03922_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1105 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06437__B1 vss _01609_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_287_clk vdd vss clknet_leaf_287_clk clknet_5_18__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10233__A1 vss _05081_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08977__A2 vss _04303_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05659__B vss _01783_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11302_ _01035_ vdd vss clknet_leaf_252_clk net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_11233_ vdd cpu.genblk3.csr.mcause31 clknet_leaf_256_clk vss _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11164_ vdd rf_ram.memory\[81\]\[0\] clknet_leaf_48_clk vss _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07401__A2 vss _03083_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10115_ vdd vss _05037_ _03071_ _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11095_ vdd rf_ram.memory\[127\]\[0\] clknet_leaf_84_clk vss _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_1024 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_179_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10046_ vdd vss _04995_ rf_ram.memory\[506\]\[1\] _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05963__A2 vss _01605_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08901__A2 vss _04257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_211_clk vdd vss clknet_leaf_211_clk clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_650 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_187_346 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10948_ vdd rf_ram.memory\[359\]\[0\] clknet_leaf_155_clk vss _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05413__I vss _01513_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_186_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06140__A2 vss _01719_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10879_ vdd rf_ram.memory\[221\]\[1\] clknet_leaf_32_clk vss _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10224__A1 vss _03892_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09465__I0 vss net82 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06979__A1 vss _02775_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_278_clk vdd vss clknet_leaf_278_clk clknet_5_17__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06070_ rf_ram.memory\[349\]\[1\] _01678_ _01677_ rf_ram.memory\[348\]\[1\] _02265_
+ vss vdd rf_ram.memory\[351\]\[1\] _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA_1 vss _02839_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09917__A1 vss _04911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05403__A1 vss _01347_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06972_ vdd vss _03043_ rf_ram.memory\[428\]\[1\] _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09760_ vdd vss _04818_ _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__05254__I1 vss net105 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05923_ rf_ram.memory\[108\]\[0\] _02119_ vss vdd rf_ram.memory\[111\]\[0\] _01625_
+ rf_ram.memory\[109\]\[0\] _01702_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_09691_ vdd vss _04771_ _04740_ net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08711_ vdd _04141_ _04140_ _00763_ _04126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_202_clk vdd vss clknet_leaf_202_clk clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08642_ vdd vss _04099_ _02828_ _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_179_847 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05706__A2 vss _01509_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05854_ _01956_ vdd vss _02050_ rf_ram.memory\[232\]\[0\] _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_156_1091 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05751__C vss _01569_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_694 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08573_ vdd vss _04054_ _02945_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05785_ rf_ram.memory\[141\]\[0\] _01931_ _01799_ rf_ram.memory\[140\]\[0\] _01981_
+ vss vdd rf_ram.memory\[143\]\[0\] _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_49_525 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07459__A2 vss _03101_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07524_ vss _03390_ _03100_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__06116__C1 vss _01715_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08656__A1 vss _04097_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07455_ vdd vss _03347_ rf_ram.memory\[330\]\[0\] _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_1220 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05323__I vss _01518_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_917 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06406_ _02598_ _02599_ _02600_ _01670_ vdd vss _02601_ _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_0_57_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_677 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07386_ vdd vss _03304_ rf_ram.memory\[24\]\[0\] _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_134_449 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09125_ vdd vss _04399_ rf_ram.memory\[92\]\[0\] _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08959__A2 vss _03945_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06337_ vss vdd rf_ram.memory\[223\]\[1\] _02019_ rf_ram.memory\[221\]\[1\] _01912_
+ _01755_ rf_ram.memory\[220\]\[1\] _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__09081__A1 vss _04367_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_269_clk vdd vss clknet_leaf_269_clk clknet_5_16__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_163_1040 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09056_ vdd vss _04356_ rf_ram.memory\[101\]\[0\] _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06268_ vdd vss _02463_ rf_ram.memory\[158\]\[1\] _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09908__A1 vss _04884_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_696 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08007_ vdd _03691_ _03687_ _00509_ _03690_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_789 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05219_ cpu.csr_d_sel vdd vss _01419_ cpu.decode.opcode\[2\] cpu.branch_op vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_06199_ _01650_ vdd vss _02394_ rf_ram.memory\[458\]\[1\] _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06198__A2 vss _01709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05926__C vss _01860_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09958_ vdd _04940_ _04938_ _01212_ _04921_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08909_ vdd _04264_ _04263_ _00838_ _04234_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06103__B vss _01620_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05945__A2 vss _01536_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09136__A2 vss _04067_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09889_ vdd vss _04898_ rf_ram.memory\[219\]\[1\] _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_1011 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06370__A2 vss _01683_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10802_ vdd rf_ram.memory\[555\]\[0\] clknet_leaf_322_clk vss _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08647__A1 vss net238 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10733_ vdd rf_ram.memory\[45\]\[1\] clknet_leaf_127_clk vss _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05233__I vss net134 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_552 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10664_ vdd rf_ram.memory\[378\]\[0\] clknet_leaf_108_clk vss _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_799 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_438 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10595_ vdd rf_ram.memory\[31\]\[1\] clknet_leaf_204_clk vss _00339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05881__A1 vss _01972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10206__A1 vss _05078_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_274 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_780 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_696 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_609 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06189__A2 vss _01782_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11216_ vdd rf_ram.memory\[68\]\[0\] clknet_leaf_61_clk vss _00952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11147_ vdd rf_ram.memory\[107\]\[1\] clknet_leaf_68_clk vss _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput71 o_dbus_adr[14] net71 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput93 o_dbus_adr[6] net93 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput82 o_dbus_adr[25] net82 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07138__A1 vss _03123_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11078_ vdd rf_ram.memory\[133\]\[1\] clknet_leaf_15_clk vss _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08886__A1 vss _04237_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10029_ vdd _04984_ _04983_ _01239_ _04982_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05571__C vss _01361_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_992 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_1074 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_519 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05570_ _01349_ _01765_ vdd vss _01766_ _01754_ _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_59_834 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08638__A1 vss _04094_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06361__A2 vss _01515_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1069 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_703 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06113__A2 vss _01644_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07310__A1 vss _03225_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07240_ vdd _03212_ _03210_ _00221_ _03193_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_129_788 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09438__I0 vss net69 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07171_ vdd _03170_ _03169_ _00194_ _03157_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_561 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_143_268 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06122_ _02315_ _02316_ vdd vss _02317_ _02313_ _02314_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_87_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_482 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05624__A1 vss _01675_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1067 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_244 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06053_ rf_ram.memory\[365\]\[1\] _01610_ _01644_ rf_ram.memory\[364\]\[1\] _02248_
+ vss vdd rf_ram.memory\[367\]\[1\] _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_0_169_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07377__A1 vss _03289_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09812_ vdd vss _04851_ _02828_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05927__A2 vss _01631_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05318__I vss _01513_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07129__A1 vss rf_ram.memory\[4\]\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09743_ vdd vss _04807_ _04804_ net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06955_ vdd _03031_ _03029_ _00117_ _03018_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_154_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06886_ vdd vss _02986_ rf_ram.memory\[281\]\[0\] _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05906_ _02089_ _02101_ _01362_ vdd vss _02102_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__06337__C1 vss _02019_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08877__A1 vss net237 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09674_ vdd vss _04757_ _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05837_ _02029_ _02032_ vdd vss _02033_ _02021_ _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_08625_ vdd vss _04088_ _02821_ _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08556_ vdd vss _04044_ rf_ram.memory\[489\]\[1\] _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08629__A1 vss _04062_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07507_ vdd _03379_ _03377_ _00321_ _03360_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_92_601 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05768_ vdd vss _01964_ rf_ram.memory\[145\]\[0\] _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08487_ vdd _03997_ _03995_ _00683_ _03956_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05699_ vdd vss _01895_ rf_ram.memory\[414\]\[0\] _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06104__A2 vss _01692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07438_ vdd _03336_ _03334_ _00295_ _03326_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09054__A1 vss _04334_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07369_ vdd _03293_ _03290_ _00269_ _03292_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09108_ vdd vss _04388_ rf_ram.memory\[94\]\[0\] _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_734 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10380_ vdd rf_ram.memory\[427\]\[0\] clknet_leaf_100_clk vss _00124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_994 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05937__B vss _01601_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09039_ vdd _04345_ _04343_ _00887_ _04334_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09409__B vss _01344_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10134__I vss _02747_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11001_ vdd rf_ram.memory\[519\]\[1\] clknet_leaf_270_clk vss _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05918__A2 vss _01770_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_73_1236 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07540__A1 vss _03393_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06343__A2 vss _01915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_962 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09293__A1 vss net237 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_483 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10716_ vdd rf_ram.memory\[463\]\[0\] clknet_leaf_51_clk vss _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_336 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10647_ vdd rf_ram.memory\[401\]\[1\] clknet_leaf_95_clk vss _00391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09045__A1 vss _02828_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_886 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_723 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_745 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10578_ vdd rf_ram.memory\[323\]\[0\] clknet_leaf_164_clk vss _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_789 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_463 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09348__A2 vss _03991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08020__A2 vss _03693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1147 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06582__A2 vss _02730_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08859__A1 vss _04205_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06740_ vdd vss _02882_ _02716_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08449__I vss net34 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06671_ vdd _02834_ _02833_ _00030_ _02820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_64_77 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07531__A1 vss _03319_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1001 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05622_ vdd vss _01818_ rf_ram.memory\[494\]\[0\] _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08410_ vdd vss _03942_ _02761_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06334__A2 vss _01940_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_601 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09390_ _04564_ net218 vdd vss _04568_ net217 _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_188_1124 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_349 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05553_ rf_ram.memory\[285\]\[0\] _01678_ _01634_ rf_ram.memory\[284\]\[0\] _01749_
+ vss vdd rf_ram.memory\[287\]\[0\] _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08341_ vdd vss _03899_ _03892_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05484_ rf_ram.memory\[349\]\[0\] _01678_ _01677_ rf_ram.memory\[348\]\[0\] _01680_
+ vss vdd rf_ram.memory\[351\]\[0\] _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_08272_ vdd _03856_ _03853_ _00609_ _03855_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_74_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_912 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07223_ vdd _03202_ _03201_ _00214_ _03190_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_15_734 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07598__A1 vss net239 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_780 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07154_ vdd vss _03160_ rf_ram.memory\[484\]\[0\] _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08912__I vss _04057_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06105_ vdd vss _02300_ rf_ram.memory\[281\]\[1\] _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_113_975 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07085_ vdd vss _03116_ rf_ram.memory\[491\]\[1\] _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_726 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07528__I vss _03359_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_986 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06270__A1 vss _01951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_661 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06036_ vss vdd rf_ram.memory\[569\]\[1\] _01539_ rf_ram.memory\[571\]\[1\] _01540_
+ _01544_ rf_ram.memory\[570\]\[1\] _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_0_160_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_100_647 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07987_ vdd vss _03678_ rf_ram.memory\[467\]\[1\] _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input38_I vss i_ibus_rdt[13] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09726_ vdd vss _04795_ _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06938_ vdd _03021_ _03020_ _00110_ _03014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05781__B1 vss _01608_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07522__A1 vss _03360_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06869_ vdd _02974_ _02973_ _00088_ _02970_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_78_940 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09657_ vdd vss _04743_ net98 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06325__A2 vss _01510_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_962 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08608_ vdd vss _04077_ _02731_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_09588_ vdd vss _04700_ _02709_ _04699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_08539_ vdd vss _04033_ rf_ram.memory\[19\]\[1\] _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08078__A2 vss _03729_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_314 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_360 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11550_ vdd rf_ram.memory\[453\]\[1\] clknet_leaf_122_clk vss _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10501_ vdd rf_ram.memory\[258\]\[1\] clknet_leaf_196_clk vss _00245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05511__I vss _01503_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05836__A1 vss _01972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11481_ vdd rf_ram.memory\[335\]\[0\] clknet_leaf_168_clk vss _01213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_514 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_566 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10432_ vdd rf_ram.memory\[487\]\[0\] clknet_leaf_225_clk vss _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_553 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10363_ vdd rf_ram.memory\[278\]\[1\] clknet_leaf_179_clk vss _00107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_21_759 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1068 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10294_ vdd rf_ram.memory\[523\]\[0\] clknet_leaf_269_clk vss _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07761__A1 vss _03524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07513__A1 vss _02775_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_75_409 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09602__B vss _04526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_932 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_511 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07816__A2 vss _03559_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05421__I vss _01513_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09018__A1 vss _02787_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_840 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_339 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_780 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09569__A2 vss net52 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08241__A2 vss _03135_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_5_5__f_clk_I vss clknet_3_1_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_967 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08890_ vdd vss _04253_ rf_ram.memory\[479\]\[1\] _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07910_ vdd vss _03630_ _02822_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07841_ _03587_ _03355_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06004__A1 vss _01495_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07772_ vdd vss _03544_ _03008_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07752__A1 vss _02781_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09511_ vdd _04641_ _04639_ _01063_ _04637_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06723_ vdd vss _02871_ rf_ram.memory\[51\]\[0\] _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_176_400 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06654_ _02820_ vss vdd _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09442_ _04593_ vdd vss _04597_ net71 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05605_ _01801_ _01661_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06585_ vdd vss _02767_ _02761_ _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09373_ vdd vss _04558_ _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_129_360 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08324_ vdd _03888_ _03885_ _00629_ _03887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05536_ vdd vss cpu.immdec.imm19_12_20\[6\] _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_1095 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_393 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05331__I vss _01526_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05467_ _01504_ vdd vss _01663_ rf_ram.memory\[374\]\[0\] _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__09009__A1 vss _04298_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_706 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08255_ vdd _03845_ _03843_ _00603_ _03823_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08480__A2 vss _03992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07206_ vdd vss _03192_ rf_ram.memory\[262\]\[0\] _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06491__A1 vss net252 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08186_ vdd _03803_ _03802_ _00576_ _03787_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05398_ vdd vss _01594_ _01570_ _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07137_ vdd vss _03149_ rf_ram.memory\[498\]\[0\] _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05451__C1 vss _01646_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_591 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07991__A1 vss _03651_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09980__A2 vss _04951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07068_ vdd vss _03106_ rf_ram.memory\[494\]\[0\] _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06019_ _01528_ vdd vss _02214_ rf_ram.memory\[552\]\[1\] _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_57_1006 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05506__I vss _01609_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1039 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_545 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09709_ vdd vss _04783_ _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10981_ vdd rf_ram.memory\[167\]\[1\] clknet_leaf_0_clk vss _00718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_148_680 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_853 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_820 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_147_190 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11533_ vdd rf_ram.memory\[351\]\[0\] clknet_leaf_192_clk vss _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_93_795 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1146 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11464_ vdd rf_ram.memory\[344\]\[1\] clknet_leaf_141_clk vss _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_180_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10415_ vdd rf_ram.memory\[493\]\[1\] clknet_leaf_182_clk vss _00159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_501 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11395_ _01127_ vdd vss clknet_leaf_226_clk net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10346_ vdd rf_ram.memory\[282\]\[0\] clknet_leaf_179_clk vss _00090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05993__B1 vss _01950_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10277_ vdd rf_ram.memory\[236\]\[1\] clknet_leaf_281_clk vss _00021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09383__I vss _04539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1009 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07734__A1 vss _03491_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1106 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09487__A1 vss _02690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_937 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_115_1184 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06170__B1 vss _01645_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_691 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_124_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06370_ _01684_ vdd vss _02565_ rf_ram.memory\[240\]\[1\] _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_16_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05321_ _01517_ _01516_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05252_ vdd vss cpu.bne_or_bge _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_08040_ vdd vss _03712_ net235 _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_153_193 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_856 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05183_ _01382_ vdd vss _01383_ _01380_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_09991_ vdd vss _04961_ _02727_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10021__A2 vss _03009_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08942_ vdd vss _04285_ rf_ram.memory\[122\]\[1\] _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07973__A1 vss _03668_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_53 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07725__A1 vss _02795_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08873_ vdd vss _04243_ rf_ram.memory\[12\]\[0\] _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07824_ vdd vss _03577_ rf_ram.memory\[433\]\[1\] _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05736__B1 vss _01931_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07755_ vdd vss _03534_ rf_ram.memory\[395\]\[1\] _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09478__A1 vss _02703_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07686_ _03491_ _03359_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06706_ vdd _02858_ _02856_ _00041_ _02826_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05770__B vss _01494_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_241 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06637_ vdd vss _02807_ _02801_ _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09425_ _02707_ vdd vss _04588_ net93 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08150__A1 vss _03757_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09356_ _04549_ vss vdd _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_06568_ _02752_ vss vdd _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_133_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05519_ _01715_ _01714_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_09287_ _04507_ vss vdd _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_08307_ vdd _03877_ _03875_ _00623_ _03855_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06499_ _02690_ net132 _01375_ vss _01400_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_30_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05267__A2 vss _01418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08238_ vdd _03835_ _03834_ _00596_ _03820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05672__C1 vss _01713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_787 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_489 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10200_ vdd vss _05090_ rf_ram.memory\[191\]\[0\] _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08169_ vdd vss _03793_ rf_ram.memory\[543\]\[0\] _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_120_539 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11180_ vdd rf_ram.memory\[93\]\[0\] clknet_leaf_61_clk vss _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_1043 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_313_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10131_ vdd vss _05047_ _02805_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07964__A1 vss _03651_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_753 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_1049 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_max_cap238_I vss _02898_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10062_ vdd _05004_ _05002_ _01252_ _04985_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_output69_I vss net69 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_328_clk_I vss clknet_5_4__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10079__A2 vss _02917_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08547__I vss _04037_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_753 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08141__A1 vss net241 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10964_ vdd rf_ram.memory\[171\]\[0\] clknet_leaf_9_clk vss _00701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_274 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10895_ vdd rf_ram.memory\[181\]\[1\] clknet_leaf_17_clk vss _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_431 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09641__A1 vss _04634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08444__A2 vss _03949_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11516_ vdd rf_ram.memory\[306\]\[1\] clknet_leaf_144_clk vss _01248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_867 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_163 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_150_141 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11447_ vdd cpu.state.stage_two_req clknet_leaf_240_clk vss _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09944__A2 vss _02923_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06207__A1 vss _01350_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_539 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_580 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11378_ _01110_ vdd vss clknet_leaf_231_clk net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05415__C1 vss _01610_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10329_ vdd rf_ram.memory\[288\]\[1\] clknet_leaf_147_clk vss _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07707__A1 vss _03488_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05870_ _02064_ _02065_ vdd vss _02066_ _02062_ _02063_ _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__05146__I vss _01348_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08380__A1 vss _03134_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07540_ vdd _03400_ _03398_ _00333_ _03393_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_89_854 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07471_ vdd vss _03357_ _02972_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06143__B1 vss _01726_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_904 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_403 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09880__A1 vss _04887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06422_ _02616_ vdd vss _02617_ _01909_ _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_09210_ vdd vss _04452_ rf_ram.memory\[68\]\[0\] _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_57_751 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06694__A1 vss _02820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09141_ vdd vss _04409_ net245 _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06353_ vdd vss _02548_ rf_ram.memory\[238\]\[1\] _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_142_620 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09072_ vdd vss _04366_ rf_ram.memory\[81\]\[0\] _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05304_ vdd vss _01500_ _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_71_242 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05749__C vss _01717_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06284_ rf_ram.memory\[132\]\[1\] _02479_ vss vdd rf_ram.memory\[135\]\[1\] _01911_
+ rf_ram.memory\[133\]\[1\] _01912_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_71_275 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06997__A2 vss _02899_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08023_ vdd vss _03702_ rf_ram.memory\[571\]\[1\] _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_170_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08199__A1 vss _03798_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05235_ vdd vss rf_ram_if.rtrig1 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05166_ vss _01369_ _01347_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_4_597 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09396__B1 vss _04564_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07946__A1 vss _02728_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09974_ _04950_ _04396_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08925_ vdd vss _04275_ rf_ram.memory\[124\]\[0\] _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05709__B1 vss _01763_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input20_I vss i_dbus_rdt[26] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08856_ vdd vss _04232_ rf_ram.memory\[131\]\[0\] _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07807_ vdd vss _03567_ rf_ram.memory\[414\]\[0\] _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07174__A2 vss _03158_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06382__B1 vss _01912_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05999_ _01506_ vdd vss _02194_ rf_ram.memory\[518\]\[1\] _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08787_ vdd vss _04189_ _03071_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07738_ vdd _03523_ _03522_ _00408_ _03521_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07669_ vdd vss _03480_ rf_ram.memory\[403\]\[1\] _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06134__B1 vss _01786_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output107_I vss net107 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10680_ vdd rf_ram.memory\[437\]\[0\] clknet_leaf_80_clk vss _00424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_133_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_879 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06685__A1 vss _02730_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09408_ _04577_ vdd vss _04578_ cpu.ctrl.i_jump _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_75_570 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09339_ vss _04540_ _04539_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_180_737 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_105_300 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09623__A1 vss _04634_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1064 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_132_163 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11301_ vdd net96 clknet_leaf_251_clk vss _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_848 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_252_clk_I vss clknet_5_20__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11232_ vdd cpu.genblk3.csr.mstatus_mpie clknet_leaf_238_clk vss _00968_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07937__A1 vss _03619_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11163_ vdd rf_ram.memory\[0\]\[1\] clknet_leaf_35_clk vss _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_684 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10114_ vdd _05036_ _05034_ _01272_ _05017_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06070__C1 vss _01688_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11094_ vdd rf_ram.memory\[479\]\[1\] clknet_leaf_121_clk vss _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_267_clk_I vss clknet_5_17__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10045_ vdd _04994_ _04993_ _01245_ _04982_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_1182 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08362__A1 vss _03887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05176__A1 vss _01353_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_85_301 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08114__A1 vss _03757_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10947_ vdd rf_ram.memory\[369\]\[1\] clknet_leaf_149_clk vss _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_39_762 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06676__A1 vss _02716_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_205_clk_I vss clknet_5_24__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10878_ vdd rf_ram.memory\[221\]\[0\] clknet_leaf_32_clk vss _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_439 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09465__I1 vss net83 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_247 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05569__C vss _01670_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10224__A2 vss _03134_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06979__A2 vss _03040_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_2 vss _02839_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09917__A2 vss _03083_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05651__A2 vss _01846_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_848 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05585__B vss _01746_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_556 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05939__B1 vss _01607_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06971_ vdd _03042_ _03041_ _00122_ _03014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_158_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05403__A2 vss _01346_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05254__I2 vss net128 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1211 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06600__A1 vss _02743_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05922_ _02004_ vdd vss _02118_ rf_ram.memory\[110\]\[0\] _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09690_ vdd vss _04770_ _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08710_ vdd vss _04141_ rf_ram.memory\[151\]\[0\] _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08353__A1 vss _03008_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05853_ _02048_ vdd vss _02049_ _01951_ _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08641_ vdd _04098_ _04095_ _00736_ _04097_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_83_76 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_301 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05784_ vdd vss _01980_ rf_ram.memory\[142\]\[0\] _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08572_ vdd _04053_ _04051_ _00712_ _04026_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08105__A1 vss _03721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07523_ _03389_ _03355_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06116__B1 vss _01654_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_835 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09853__A1 vss _02713_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07454_ vdd vss _03346_ _02775_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06667__A1 vss _02736_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09520__B vss _02709_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06405_ rf_ram.memory\[82\]\[1\] _02600_ vss vdd rf_ram.memory\[81\]\[1\] _01656_
+ rf_ram.memory\[83\]\[1\] _01654_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_88_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_96_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07385_ vdd vss _03303_ _02992_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09605__A1 vss _04524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09124_ vdd vss _04398_ _02838_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05890__A2 vss _01510_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_584 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06336_ vdd vss _02531_ rf_ram.memory\[222\]\[1\] _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_161_269 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06267_ _02461_ vdd vss _02462_ _01373_ _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_09055_ vdd vss _04355_ _02794_ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07092__A1 vss _02915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08006_ vdd vss _03691_ rf_ram.memory\[465\]\[1\] _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05218_ _01418_ _01417_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06198_ rf_ram.memory\[460\]\[1\] _02393_ vss vdd rf_ram.memory\[463\]\[1\] _01713_
+ rf_ram.memory\[461\]\[1\] _01721_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__07919__A1 vss _03622_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_481 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05495__B vss _01629_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05149_ vss _01352_ rf_ram_if.rtrig0 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09957_ vdd vss _04940_ rf_ram.memory\[336\]\[1\] _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08908_ vdd vss _04264_ rf_ram.memory\[125\]\[0\] _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09888_ vdd _04897_ _04896_ _01185_ _04884_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10151__A1 vss _05049_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08839_ vdd _04221_ _04219_ _00811_ _04205_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05158__A1 vss _01353_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output224_I vss net224 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_170_1056 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10801_ vdd rf_ram.memory\[556\]\[1\] clknet_leaf_322_clk vss _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09844__A1 vss _02714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08647__A2 vss _04067_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10732_ vdd rf_ram.memory\[45\]\[0\] clknet_leaf_127_clk vss _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_180_512 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10663_ vdd rf_ram.memory\[397\]\[1\] clknet_leaf_94_clk vss _00407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_180_556 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10594_ vdd rf_ram.memory\[31\]\[0\] clknet_leaf_204_clk vss _00338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_91_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_191_clk_I vss clknet_5_28__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_130 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_3_0_clk clknet_3_3_0_clk vss vdd clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_71_clk_I vss clknet_5_8__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05633__A2 vss _01735_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_982 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11215_ vdd rf_ram.memory\[6\]\[1\] clknet_leaf_40_clk vss _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11146_ vdd rf_ram.memory\[107\]\[0\] clknet_leaf_68_clk vss _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput83 o_dbus_adr[26] net83 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput72 o_dbus_adr[15] net72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput94 o_dbus_adr[7] net94 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05397__A1 vss _01351_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_86_clk_I vss clknet_5_10__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11077_ vdd rf_ram.memory\[133\]\[0\] clknet_leaf_15_clk vss _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10028_ vdd vss _04984_ rf_ram.memory\[327\]\[0\] _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08335__A1 vss _03887_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08886__A2 vss _04248_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10142__A1 vss _03672_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_196_clk vdd vss clknet_leaf_196_clk clknet_5_25__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_144_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06897__A1 vss _02958_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05424__I vss _01493_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_807 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_114_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_857 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_144_clk_I vss clknet_5_27__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_24_clk_I vss clknet_5_3__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09438__I1 vss net70 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_556 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07170_ vdd vss _03170_ rf_ram.memory\[495\]\[0\] _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05872__A2 vss _01677_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_159_clk_I vss clknet_5_27__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_589 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1069 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06121_ rf_ram.memory\[258\]\[1\] _02316_ vss vdd rf_ram.memory\[257\]\[1\] _01668_
+ rf_ram.memory\[259\]\[1\] _01519_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__07074__A1 vss _03087_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06052_ vdd vss _02247_ rf_ram.memory\[366\]\[1\] _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_120_clk vdd vss clknet_leaf_120_clk clknet_5_13__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_39_clk_I vss clknet_5_7__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06204__B vss _01756_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09811_ vdd _04850_ _04848_ _01154_ _04840_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06034__C1 vss _01554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09742_ vdd vss _04806_ _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06954_ vdd vss _03031_ rf_ram.memory\[231\]\[1\] _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10133__A1 vss _05046_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06885_ vdd vss _02985_ _02958_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xclkbuf_leaf_187_clk vdd vss clknet_leaf_187_clk clknet_5_28__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05905_ _02095_ _01660_ _02100_ vdd vss _02101_ _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_94_1131 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06337__B1 vss _01912_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08877__A2 vss _04077_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09673_ _04756_ vdd vss _04757_ net123 _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_171_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_90_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05836_ _02031_ vdd vss _02032_ _01972_ _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_11_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08624_ vdd _04087_ _04085_ _00730_ _04062_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_139_509 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08555_ vdd _04043_ _04042_ _00705_ _04023_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05334__I vss _01499_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05767_ _01956_ vdd vss _01963_ rf_ram.memory\[144\]\[0\] _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07506_ vdd vss _03379_ rf_ram.memory\[363\]\[1\] _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_178_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_166_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09826__A1 vss _04840_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08486_ vdd vss _03997_ rf_ram.memory\[379\]\[1\] _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05698_ _01890_ _01893_ vdd vss _01894_ _01882_ _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07437_ vdd vss _03336_ rf_ram.memory\[332\]\[1\] _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_130_1073 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_646 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_486 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_754 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05312__A1 vss _01496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07368_ vdd vss _03293_ rf_ram.memory\[251\]\[1\] _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_33_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05863__A2 vss _01940_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09107_ vdd vss _04387_ _02916_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06319_ _01923_ vdd vss _02514_ rf_ram.memory\[176\]\[1\] _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_111_clk vdd vss clknet_leaf_111_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06812__A1 vss _02930_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_921 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07299_ vdd _03249_ _03247_ _00243_ _03225_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_60_543 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_234 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09038_ vdd vss _04345_ rf_ram.memory\[105\]\[1\] _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09409__C vss _01388_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_177 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1020 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08565__A1 vss _04023_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09762__B1 vss _04760_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06025__C1 vss _01517_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11000_ vdd rf_ram.memory\[519\]\[0\] clknet_leaf_270_clk vss _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_176_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06040__A2 vss _02234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08317__A1 vss _03855_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10124__A1 vss _05017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_178_clk vdd vss clknet_leaf_178_clk clknet_5_31__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_185_637 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_339 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09817__A1 vss net240 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_974 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09293__A2 vss _04507_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10715_ vdd rf_ram.memory\[408\]\[1\] clknet_leaf_88_clk vss _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_372 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_126_726 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05839__C1 vss _01925_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05303__A1 vss _01496_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10646_ vdd rf_ram.memory\[401\]\[0\] clknet_leaf_95_clk vss _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_882 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05854__A2 vss _01735_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09045__A2 vss _04339_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10577_ vdd rf_ram.memory\[363\]\[1\] clknet_5_27__leaf_clk vss _00321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_102_clk vdd vss clknet_leaf_102_clk clknet_5_15__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_134_792 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_134_770 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05606__A2 vss _01801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05419__I vss _01550_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09753__B1 vss _04760_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06024__B vss _01528_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1104 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06031__A2 vss _01544_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11129_ vdd rf_ram.memory\[116\]\[1\] clknet_leaf_76_clk vss _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08308__A1 vss _03309_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_169_clk vdd vss clknet_leaf_169_clk clknet_5_30__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10115__A1 vss _03071_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06670_ vdd vss _02834_ rf_ram.memory\[455\]\[0\] _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07531__A2 vss _02899_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05621_ _01816_ vdd vss _01817_ _01597_ _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_148_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05542__A1 vss _01675_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05552_ vdd vss _01748_ rf_ram.memory\[286\]\[0\] _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08340_ vdd _03898_ _03896_ _00635_ _03887_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_47_827 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1034 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_188_1158 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06098__A2 vss _01687_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_586 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07295__A1 vss _02984_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08271_ vdd vss _03856_ rf_ram.memory\[197\]\[1\] _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05483_ _01679_ _01624_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__05145__I1 vss _01346_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07222_ vdd vss _03202_ rf_ram.memory\[425\]\[0\] _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05845__A2 vss _01724_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_567 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07153_ vdd vss _03159_ _02883_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07598__A2 vss _03390_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06104_ _01684_ vdd vss _02299_ rf_ram.memory\[280\]\[1\] _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07084_ vdd _03115_ _03114_ _00162_ _03087_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06035_ _01528_ vdd vss _02230_ rf_ram.memory\[568\]\[1\] _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_5_28__f_clk vdd vss clknet_5_28__leaf_clk clknet_3_7_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05329__I vss rf_ram.i_raddr\[2\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_963 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_451 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1196 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_1174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_1136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07986_ vdd _03677_ _03676_ _00502_ _03651_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06022__A2 vss _01502_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10106__A1 vss rf_ram.memory\[312\]\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09725_ _04791_ _04794_ vdd vss _04795_ net106 _04790_ net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA_clkbuf_5_22__f_clk_I vss clknet_3_5_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06937_ vdd vss _03021_ rf_ram.memory\[228\]\[0\] _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09656_ _04741_ _04742_ vdd vss _01107_ _03973_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_59_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06868_ vdd vss _02974_ rf_ram.memory\[302\]\[0\] _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08607_ vdd _04076_ _04074_ _00724_ _04062_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_179_475 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_626 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05533__A1 vss _01349_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05819_ _02014_ vdd vss _02015_ _01600_ _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06799_ vdd vss _02926_ rf_ram.memory\[50\]\[1\] _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09587_ vdd vss _04699_ _01469_ _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_613 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08538_ vdd _04032_ _04031_ _00699_ _04023_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06089__A2 vss _01719_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_862 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_332_clk vdd vss clknet_leaf_332_clk clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08469_ vdd vss _00677_ _02714_ _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10500_ vdd rf_ram.memory\[258\]\[0\] clknet_leaf_196_clk vss _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11480_ vdd rf_ram.memory\[336\]\[1\] clknet_leaf_177_clk vss _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07038__A1 vss _03050_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_781 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10431_ vdd rf_ram.memory\[500\]\[1\] clknet_leaf_224_clk vss _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10362_ vdd rf_ram.memory\[278\]\[0\] clknet_leaf_179_clk vss _00106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output99_I vss net99 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08786__A1 vss _04170_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06623__I vss _02794_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_598 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06261__A2 vss _01801_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10293_ vdd rf_ram.memory\[524\]\[1\] clknet_leaf_269_clk vss _00037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_795 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08538__A1 vss _04023_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07210__A1 vss _03193_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06013__A2 vss _01544_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07513__A2 vss _03101_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_1202 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_157_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07277__A1 vss _03222_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06485__C1 vss _01635_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05827__A2 vss _01515_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06019__B vss _01528_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_323_clk vdd vss clknet_leaf_323_clk clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09018__A2 vss _04303_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07029__A1 vss _02738_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_893 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10629_ vdd rf_ram.memory\[387\]\[1\] clknet_leaf_92_clk vss _00373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_729 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05858__B vss _01956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07629__I vss _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08777__A1 vss _02971_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_587 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_784 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07840_ vdd _03586_ _03584_ _00447_ _03557_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07201__A1 vss _03157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07771_ vdd _03543_ _03541_ _00421_ _03524_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09510_ vdd vss _04641_ rf_ram.memory\[279\]\[1\] _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06201__C vss _01658_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06722_ vdd vss _02870_ _02866_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08701__A1 vss _04126_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09441_ vss _01038_ _04596_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11614__I vss net94 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06653_ _02819_ vss vdd _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05604_ _01602_ vdd vss _01800_ rf_ram.memory\[304\]\[0\] _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06584_ _02766_ vss vdd _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_09372_ _04552_ net209 vdd vss _04558_ net208 _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09257__A2 vss _01484_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_489 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05535_ _01730_ vdd vss _01731_ _01368_ _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__05612__I vss _01640_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08323_ vdd vss _03888_ rf_ram.memory\[242\]\[1\] _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06476__C1 vss _01607_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_314_clk vdd vss clknet_leaf_314_clk clknet_5_5__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_90_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05466_ _01662_ _01661_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_08254_ vdd vss _03845_ rf_ram.memory\[527\]\[1\] _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08480__A3 vss _01418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07205_ vdd vss _03191_ _02806_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08185_ vdd vss _03803_ rf_ram.memory\[540\]\[0\] _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05397_ _01581_ _01593_ _01351_ _01592_ _01362_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_166_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07136_ vdd vss _03148_ _02915_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06243__A2 vss _01856_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07067_ vdd vss _03105_ _02915_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_24_1209 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05451__B1 vss _01645_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input50_I vss i_ibus_rdt[25] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06018_ rf_ram.memory\[557\]\[1\] _01517_ _01511_ rf_ram.memory\[556\]\[1\] _02213_
+ vss vdd rf_ram.memory\[559\]\[1\] _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09193__A1 vss _04434_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07274__I vss _03039_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06400__C1 vss _01810_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05754__A1 vss _01373_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07969_ vdd _03666_ _03665_ _00496_ _03651_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09708_ _04768_ _04782_ vdd vss _04783_ net101 _04767_ net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA_output137_I vss net137 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_204 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09496__A2 vss _01388_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10980_ vdd rf_ram.memory\[167\]\[0\] clknet_leaf_339_clk vss _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_401 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09639_ vdd vss _04728_ _02971_ _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_139_136 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_125 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07259__A1 vss _03222_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_843 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_305_clk vdd vss clknet_leaf_305_clk clknet_5_4__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11532_ vdd rf_ram.memory\[310\]\[1\] clknet_leaf_144_clk vss _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05809__A2 vss _01641_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05678__B vss _01756_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11463_ vdd rf_ram.memory\[344\]\[0\] clknet_leaf_192_clk vss _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06482__A2 vss _01643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_1109 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10414_ vdd rf_ram.memory\[493\]\[0\] clknet_leaf_183_clk vss _00158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1314 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08759__A1 vss _01363_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07431__A1 vss _03323_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06234__A2 vss _01500_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11394_ _01126_ vdd vss clknet_leaf_226_clk net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_60_170 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05397__C vss _01362_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10345_ vdd rf_ram.memory\[302\]\[1\] clknet_leaf_136_clk vss _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05993__A1 vss _01371_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10276_ vdd rf_ram.memory\[236\]\[0\] clknet_leaf_281_clk vss _00020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_178_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_5_11__f_clk vdd vss clknet_5_11__leaf_clk clknet_3_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09184__A1 vss net242 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1055 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08931__A1 vss _04266_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07498__A1 vss _03319_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_957 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_445 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_270 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_448 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05320_ _01516_ _01515_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_154_651 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06458__C1 vss _01518_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07670__A1 vss _03458_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_684 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_824 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05588__B vss _01783_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06473__A2 vss _01686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05251_ vdd vss _01451_ _01381_ _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_181_492 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05182_ vdd _01382_ cpu.decode.opcode\[0\] vss vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_0_101_85 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06225__A2 vss _01631_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_721 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09990_ vdd _04960_ _04958_ _01224_ _04953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08941_ vdd _04284_ _04283_ _00850_ _04266_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07973__A2 vss _02972_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05984__A1 vss rf_ram.memory\[0\]\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08872_ vdd vss _04242_ _02787_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11609__I vss net87 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07823_ vdd _03576_ _03575_ _00440_ _03554_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07725__A2 vss _02869_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07754_ vdd _03533_ _03532_ _00414_ _03521_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07685_ vdd _03490_ _03489_ _00388_ _03488_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06705_ vdd vss _02858_ rf_ram.memory\[522\]\[1\] _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_91_clk vdd vss clknet_leaf_91_clk clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_94_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_1095 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09424_ vss _01030_ _04587_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06636_ _02806_ vss vdd _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__05342__I vss _01537_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09355_ vdd vss _04548_ _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06567_ vdd vss _02751_ _02750_ _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__11507__CLK vss clknet_5_30__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08989__A1 vss _04298_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05518_ _01714_ vss vdd _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08306_ vdd vss _03877_ rf_ram.memory\[221\]\[1\] _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06498_ _02691_ net133 _02690_ vss _01400_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_09286_ vss _00973_ _04506_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07661__A1 vss net238 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05498__B vss _01693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05449_ vdd vss _01645_ _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XANTENNA__06464__A2 vss _01536_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_7_562 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08237_ vdd vss _03835_ rf_ram.memory\[530\]\[0\] _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05672__B1 vss _01721_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_833 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08168_ vdd vss _03792_ _02881_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07119_ vdd vss _03138_ rf_ram.memory\[500\]\[1\] _03136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08099_ vdd vss _03749_ rf_ram.memory\[556\]\[0\] _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_1006 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__05975__A1 vss _01903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10130_ _05046_ _02742_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_30_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09166__A1 vss _04401_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10061_ vdd vss _05004_ rf_ram.memory\[507\]\[1\] _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08913__A1 vss _03039_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05517__I vss _01653_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05680__C vss _01717_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10963_ vdd rf_ram.memory\[19\]\[1\] clknet_leaf_288_clk vss _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_82_clk vdd vss clknet_leaf_82_clk clknet_5_11__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_74_1173 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08141__A2 vss _03765_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06152__A1 vss net252 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10894_ vdd rf_ram.memory\[181\]\[0\] clknet_leaf_15_clk vss _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_415 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_465 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05360__C1 vss _01555_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_960 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_108_331 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11515_ vdd rf_ram.memory\[306\]\[0\] clknet_leaf_165_clk vss _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06455__A2 vss _01661_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05663__B1 vss _01857_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_777 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11446_ vdd rf_ram.memory\[60\]\[1\] clknet_leaf_289_clk vss _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06016__C vss _01569_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1231 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11377_ _01109_ vdd vss clknet_leaf_231_clk net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__05415__B1 vss _01608_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10328_ vdd rf_ram.memory\[288\]\[0\] clknet_leaf_136_clk vss _00072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09157__A1 vss _02991_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08904__A1 vss _04234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05427__I vss _01605_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10259_ vdd vss _05125_ _02916_ _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05718__A1 vss _01909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_833 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08380__A2 vss _03903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1084 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05871__B vss _02004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_73_clk vdd vss clknet_leaf_73_clk clknet_5_10__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_89_899 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_527 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07470_ vss _03356_ _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_158_264 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_426 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06421_ rf_ram.memory\[124\]\[1\] _02616_ vss vdd rf_ram.memory\[127\]\[1\] _01786_
+ rf_ram.memory\[125\]\[1\] _01772_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_118_139 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06352_ _02534_ _02546_ _01362_ vdd vss _02547_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_09140_ vdd _04408_ _04406_ _00925_ _04401_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_251 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07643__A1 vss _03455_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_673 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09071_ vdd vss _04365_ net248 _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06283_ vdd vss _02478_ rf_ram.memory\[134\]\[1\] _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05303_ vdd vss _01499_ _01496_ _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_170_930 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_127_695 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_799 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08022_ vdd _03701_ _03700_ _00514_ _03686_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_163_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_287 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05234_ _01418_ _01434_ _01432_ _01420_ _01433_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_123_890 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05165_ cpu.immdec.imm19_12_20\[6\] _01367_ cpu.immdec.imm24_20\[2\] vdd vss _01368_
+ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XANTENNA__08199__A2 vss _02984_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09973_ vdd _04949_ _04947_ _01218_ _04921_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07946__A2 vss _02832_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08924_ vdd vss _04274_ _02838_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09148__A1 vss _04397_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08855_ vdd vss _04231_ net240 _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07806_ vdd vss _03566_ _02916_ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08786_ vdd _04188_ _04186_ _00791_ _04170_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07737_ vdd vss _03523_ rf_ram.memory\[378\]\[0\] _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_79_332 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input13_I vss i_dbus_rdt[1] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05998_ _02191_ _02192_ vdd vss _02193_ _02189_ _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_170_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_64_clk vdd vss clknet_leaf_64_clk clknet_5_8__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07668_ vdd _03479_ _03478_ _00382_ _03455_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07599_ vdd vss _03437_ rf_ram.memory\[354\]\[0\] _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_137_415 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07882__A1 vss _03590_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06619_ vdd _02791_ _02789_ _00021_ _02748_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09407_ vdd _01344_ _01472_ _04577_ cpu.ctrl.i_jump vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09338_ vdd vss _04539_ net65 _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06437__A2 vss _01633_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_871 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_632 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06117__B vss _01629_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11300_ _01033_ vdd vss clknet_leaf_251_clk net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_22_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_619 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09269_ vdd vss _04494_ cpu.genblk3.csr.o_new_irq _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11231_ vdd cpu.genblk3.csr.mie_mtie clknet_leaf_239_clk vss _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_max_cap250_I vss _02727_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11162_ vdd rf_ram.memory\[0\]\[0\] clknet_leaf_35_clk vss _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output81_I vss net81 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10113_ vdd vss _05036_ rf_ram.memory\[392\]\[1\] _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06070__B1 vss _01678_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05675__C vss _01658_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_551 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11093_ vdd rf_ram.memory\[479\]\[0\] clknet_leaf_121_clk vss _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_1116 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10044_ vdd vss _04994_ rf_ram.memory\[506\]\[0\] _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05691__B vss _01783_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1257 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_55_clk vdd vss clknet_leaf_55_clk clknet_5_9__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10946_ vdd rf_ram.memory\[369\]\[0\] clknet_leaf_149_clk vss _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10577__CLK vss clknet_5_27__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07873__A1 vss _02836_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10877_ vdd rf_ram.memory\[244\]\[1\] clknet_leaf_214_clk vss _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_27_903 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_240 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_448 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05884__B1 vss _01925_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_796 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_53_221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_619 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_3 vss _03009_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_298 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05866__B vss _02004_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11429_ vdd rf_ram.memory\[62\]\[0\] clknet_leaf_291_clk vss _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_5_9__f_clk vdd vss clknet_5_9__leaf_clk clknet_3_2_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08050__A1 vss _03071_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06970_ vdd vss _03042_ rf_ram.memory\[428\]\[0\] _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05254__I3 vss net114 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05921_ _02109_ _02113_ _02116_ _01660_ vdd vss _02117_ _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA_input5_I vss i_dbus_rdt[12] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_805 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08353__A2 vss _03903_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05852_ rf_ram.memory\[237\]\[0\] _01968_ _01614_ rf_ram.memory\[236\]\[0\] _02048_
+ vss vdd rf_ram.memory\[239\]\[0\] _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09550__A1 vss _01391_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08640_ vdd vss _04098_ rf_ram.memory\[162\]\[1\] _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05167__A2 vss _01344_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09302__A1 vss _04466_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_46_clk vdd vss clknet_leaf_46_clk clknet_5_12__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05783_ _01978_ vdd vss _01979_ _01976_ _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08571_ vdd vss _04053_ rf_ram.memory\[170\]\[1\] _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07522_ vdd _03388_ _03386_ _00327_ _03360_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_77_858 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_381 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07453_ vdd _03345_ _03343_ _00301_ _03326_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06667__A2 vss _02830_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_368 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_312_clk_I vss clknet_5_5__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06404_ _01602_ vdd vss _02599_ rf_ram.memory\[80\]\[1\] _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__11622__I vss net72 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_273 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07384_ vdd _03302_ _03300_ _00275_ _03292_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09123_ _04397_ _04396_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09605__A2 vss net49 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_435 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07616__A1 vss _03422_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06335_ _01928_ vdd vss _02530_ _02527_ _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06266_ _02460_ vdd vss _02461_ _01372_ _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_115_676 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05627__B1 vss _01688_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09054_ vdd _04354_ _04352_ _00893_ _04334_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07092__A2 vss _03009_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_327_clk_I vss clknet_5_4__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08005_ _03690_ _03689_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05217_ _01385_ cpu.state.o_cnt\[2\] vdd vss _01417_ cpu.state.cnt_r\[3\] cpu.mem_bytecnt\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_06197_ _01707_ vdd vss _02392_ rf_ram.memory\[462\]\[1\] _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xmax_cap250 net250 _02727_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_05148_ _01351_ _01350_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09956_ vdd _04939_ _04938_ _01211_ _04918_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08907_ vdd vss _04263_ _02959_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09887_ vdd vss _04897_ rf_ram.memory\[219\]\[0\] _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08838_ vdd vss _04221_ rf_ram.memory\[469\]\[1\] _04219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_99_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_1100 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06355__A1 vss _01951_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1024 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_135_1122 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_37_clk vdd vss clknet_leaf_37_clk clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08769_ vdd _04178_ _04177_ _00784_ _04167_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_178_860 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_702 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10800_ vdd rf_ram.memory\[556\]\[0\] clknet_leaf_322_clk vss _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07855__A1 vss _03587_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10731_ vdd rf_ram.memory\[443\]\[1\] clknet_leaf_55_clk vss _00475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10662_ vdd rf_ram.memory\[397\]\[0\] clknet_leaf_93_clk vss _00406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05530__I vss _01635_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06626__I vss cpu.immdec.imm11_7\[3\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07607__A1 vss _03425_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10593_ vdd rf_ram.memory\[35\]\[1\] clknet_leaf_203_clk vss _00337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_142 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08280__A1 vss _03852_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11214_ vdd rf_ram.memory\[6\]\[0\] clknet_leaf_40_clk vss _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08032__A1 vss _03686_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11145_ vdd rf_ram.memory\[108\]\[1\] clknet_leaf_71_clk vss _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09780__A1 vss net244 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput73 o_dbus_adr[16] net73 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput84 o_dbus_adr[27] net84 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__06594__A1 vss _02748_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05397__A2 vss _01581_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11076_ vdd rf_ram.memory\[134\]\[1\] clknet_leaf_25_clk vss _00813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput95 o_dbus_adr[8] net95 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10027_ vdd vss _04983_ _04911_ _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10142__A2 vss _02883_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06897__A2 vss _02992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_28_clk vdd vss clknet_leaf_28_clk clknet_5_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_188_1318 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10929_ vdd rf_ram.memory\[175\]\[1\] clknet_leaf_7_clk vss _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_757 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05440__I vss _01635_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_928 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_906 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1069 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06120_ _01526_ vdd vss _02315_ rf_ram.memory\[256\]\[1\] _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_81_382 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06051_ _01629_ vdd vss _02246_ _02243_ _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_152_782 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_950 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07367__I vss _03017_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_1081 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09810_ vdd vss _04850_ rf_ram.memory\[74\]\[1\] _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06585__A1 vss _02761_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05388__A2 vss _01511_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06034__B1 vss _01555_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09741_ _04791_ _04805_ vdd vss _04806_ net112 _04790_ net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06953_ vdd _03030_ _03029_ _00116_ _03014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05904_ _02097_ _02098_ _02099_ _01670_ vdd vss _02100_ _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__11617__I vss net67 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09523__A1 vss _03992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06220__B vss _01790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05615__I vss _01635_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09672_ _04735_ vdd vss _04756_ _04754_ _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06884_ _02984_ vss vdd _02983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_178_101 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_19_clk vdd vss clknet_leaf_19_clk clknet_5_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05835_ vss vdd rf_ram.memory\[223\]\[0\] _02019_ rf_ram.memory\[221\]\[0\] _01968_
+ _01755_ rf_ram.memory\[220\]\[0\] _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_08623_ vdd vss _04087_ rf_ram.memory\[529\]\[1\] _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08554_ vdd vss _04043_ rf_ram.memory\[489\]\[0\] _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_251_clk_I vss clknet_5_20__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05766_ _01564_ vdd vss _01962_ _01957_ _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07505_ vdd _03378_ _03377_ _00320_ _03356_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_76_132 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08485_ vdd _03996_ _03995_ _00682_ _03953_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_147_521 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05697_ _01892_ vdd vss _01893_ _01675_ _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_119_212 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07436_ vdd _03335_ _03334_ _00294_ _03323_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_722 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_134_237 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07367_ _03292_ _03017_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_73_850 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_266_clk_I vss clknet_5_17__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09106_ vdd _04386_ _04384_ _00913_ _04367_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06318_ rf_ram.memory\[180\]\[1\] _02513_ vss vdd rf_ram.memory\[183\]\[1\] _01773_
+ rf_ram.memory\[181\]\[1\] _01772_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_0_17_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09037_ vdd _04344_ _04343_ _00886_ _04331_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07298_ vdd vss _03249_ rf_ram.memory\[25\]\[1\] _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06273__B1 vss _01959_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06249_ vdd vss _02444_ rf_ram.memory\[446\]\[1\] _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_131_966 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08014__A1 vss _03690_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09762__A1 vss net119 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06025__B1 vss _01521_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_204_clk_I vss clknet_5_24__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06576__A1 vss _02756_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09939_ vdd vss _04929_ _02868_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__05525__I vss _01714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_219_clk_I vss clknet_5_22__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07828__A1 vss _03554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_510 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09817__A2 vss _03253_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_430 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_532 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__05839__B1 vss _01912_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10714_ vdd rf_ram.memory\[408\]\[0\] clknet_leaf_89_clk vss _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_647 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06500__A1 vss _01376_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10645_ vdd rf_ram.memory\[383\]\[1\] clknet_leaf_107_clk vss _00389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_1313 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08253__A1 vss _03820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10576_ vdd rf_ram.memory\[363\]\[0\] clknet_leaf_159_clk vss _00320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10060__A1 vss _04982_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_909 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09753__A1 vss net116 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1075 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11128_ vdd rf_ram.memory\[116\]\[0\] clknet_leaf_76_clk vss _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06567__A1 vss _02750_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08308__A2 vss _02866_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10115__A2 vss _03100_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05435__I vss _01530_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11059_ vdd rf_ram.memory\[140\]\[0\] clknet_leaf_12_clk vss _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_410 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05620_ _01815_ vdd vss _01816_ net252 _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_118_1161 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_920 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_114_1025 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_953 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05551_ _01746_ vdd vss _01747_ _01743_ _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08492__A1 vss _03956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_576 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07295__A2 vss _02997_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05482_ _01678_ vss vdd _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08270_ _03855_ _03689_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07221_ vdd vss _03201_ _02752_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_104_96 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_89_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_172_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07152_ vss _03158_ _02910_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_6_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06103_ _01620_ vdd vss _02298_ _02295_ _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_15_758 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_270 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07083_ vdd vss _03115_ rf_ram.memory\[491\]\[0\] _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07097__I vss _03013_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_8_clk vdd vss clknet_leaf_8_clk clknet_5_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06034_ rf_ram.memory\[573\]\[1\] _01555_ _01538_ rf_ram.memory\[572\]\[1\] _02229_
+ vss vdd rf_ram.memory\[575\]\[1\] _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__09744__B2 vss net114 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1284 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07985_ vdd vss _03677_ rf_ram.memory\[467\]\[0\] _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_96_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09724_ vdd vss _04794_ _04781_ net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06936_ vdd vss _03020_ _02766_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06867_ vdd vss _02973_ _02935_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_190_clk_I vss clknet_5_28__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05781__A2 vss _01606_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09655_ _04736_ vdd vss _04742_ net1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_05818_ _02012_ _02013_ vdd vss _02014_ _02010_ _02011_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08606_ vdd vss _04076_ rf_ram.memory\[164\]\[1\] _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_3_2_0_clk clknet_3_2_0_clk vss vdd clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_70_clk_I vss clknet_5_8__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06798_ vdd _02925_ _02924_ _00066_ _02873_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09586_ vdd vss _04698_ net134 _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06730__A1 vss _02873_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05749_ _01943_ _01944_ vdd vss _01945_ _01941_ _01942_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_148_830 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_452 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08537_ vdd vss _04032_ rf_ram.memory\[19\]\[0\] _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08483__A1 vss net244 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08468_ _03984_ vdd vss _03985_ _03968_ _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_07419_ vdd vss _03325_ rf_ram.memory\[371\]\[0\] _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_147_384 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_866 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_85_clk_I vss clknet_5_10__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10430_ vdd rf_ram.memory\[500\]\[0\] clknet_leaf_224_clk vss _00174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08399_ vdd _03935_ _03933_ _00657_ _03922_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_162_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10042__A1 vss _04985_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08235__A1 vss _03823_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10361_ vdd rf_ram.memory\[298\]\[1\] clknet_leaf_138_clk vss _00105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09983__A1 vss _04950_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10292_ vdd rf_ram.memory\[524\]\[0\] clknet_leaf_269_clk vss _00036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_791 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07735__I vss _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_143_clk_I vss clknet_5_27__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_23_clk_I vss clknet_5_3__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_158_clk_I vss clknet_5_27__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_947 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07470__I vss _03355_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05524__A2 vss _01719_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_38_clk_I vss clknet_5_7__leaf_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1008 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1209 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_172_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06485__B1 vss _01714_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_187_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_24_511 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10628_ vdd rf_ram.memory\[387\]\[0\] clknet_leaf_92_clk vss _00372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07029__A2 vss _02992_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_416 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08226__A1 vss _03798_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10559_ vdd rf_ram.memory\[330\]\[1\] clknet_leaf_158_clk vss _00303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_161_1310 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10033__A1 vss _02805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06788__A1 vss _02915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08777__A2 vss _04152_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_925 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_903 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_1017 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06035__B vss _01528_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_262 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05748__C1 vss _01645_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05212__A1 vss _01375_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07770_ vdd vss _03543_ rf_ram.memory\[393\]\[1\] _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_159_1294 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06721_ vss _02869_ _02868_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_91_1102 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_1192 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06960__A1 vss _03018_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_240 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09440_ _04593_ vdd vss _04596_ net70 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06652_ vdd _02818_ _02816_ _00027_ _02748_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06173__C1 vss _01715_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_66 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06712__A1 vss _02728_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05603_ _01799_ _01613_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06583_ vdd vss _02765_ _02731_ _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09371_ vdd vss _04557_ _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_05534_ _01729_ _01361_ vdd vss _01730_ _01674_ _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08322_ _03887_ _03689_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_46_124 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06476__B1 vss _01609_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_466 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08253_ vdd _03844_ _03843_ _00602_ _03820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05279__A1 vss _01366_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1221 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07204_ _03190_ _03013_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05465_ _01661_ _01499_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_7_766 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11630__I vss net80 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_533 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08184_ vdd vss _03802_ _02838_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08217__A1 vss _03820_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05396_ vdd _01351_ _01591_ _01592_ _01586_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_43_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07135_ vdd _03147_ _03145_ _00181_ _03126_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07066_ vdd _03104_ _03102_ _00155_ _03092_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_113_752 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_1226 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_582 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09717__A1 vss net104 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput230 o_ibus_adr[6] net230 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06017_ _01506_ vdd vss _02212_ rf_ram.memory\[558\]\[1\] _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09717__B2 vss net105 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_26_1070 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input43_I vss i_ibus_rdt[18] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06400__B1 vss _01646_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07968_ vdd vss _03666_ rf_ram.memory\[47\]\[0\] _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_250_clk vdd vss clknet_leaf_250_clk clknet_5_20__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05754__A2 vss _01817_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09707_ vdd vss _04782_ _04781_ net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06919_ vdd vss _03007_ _02785_ _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__06951__A1 vss _02766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07899_ vdd _03623_ _03620_ _00469_ _03622_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09638_ vdd _04727_ _01391_ _01104_ _04524_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_1091 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09569_ _04678_ _04684_ vdd vss _04685_ _04478_ net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_65_422 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11600_ vdd rf_ram.memory\[574\]\[1\] clknet_leaf_306_clk vss _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11531_ vdd rf_ram.memory\[310\]\[0\] clknet_leaf_145_clk vss _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_1220 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_230 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10263__A1 vss _02825_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_877 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_163_674 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11462_ vdd rf_ram.memory\[292\]\[1\] clknet_leaf_139_clk vss _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08208__A1 vss _03790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06219__B1 vss _01786_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09956__A1 vss _04918_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_398 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10015__A1 vss _04953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_549 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_741 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10413_ vdd rf_ram.memory\[494\]\[1\] clknet_leaf_182_clk vss _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11393_ _01125_ vdd vss clknet_leaf_225_clk net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__08759__A2 vss _01366_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10344_ vdd rf_ram.memory\[302\]\[0\] clknet_leaf_136_clk vss _00088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05442__A1 vss _01527_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09708__A1 vss net101 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05978__C1 vss _01653_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05694__B vss _01790_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05993__A2 vss _01594_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10275_ vdd rf_ram.memory\[235\]\[1\] clknet_leaf_278_clk vss _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09184__A2 vss _04067_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_241_clk vdd vss clknet_leaf_241_clk clknet_5_21__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05745__A2 vss _01940_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_903 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_503 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07498__A2 vss _02883_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05713__I vss _01756_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06155__C1 vss _01679_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_457 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_580 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06170__A2 vss _01644_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_276 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139_682 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10254__A1 vss net249 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06458__B1 vss _01655_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_809 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_866 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05250_ vdd vss _01450_ _01399_ _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05681__A1 vss _01350_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05181_ vss _01381_ cpu.branch_op vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_101_64 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_396 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08940_ vdd vss _04284_ rf_ram.memory\[122\]\[0\] _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05984__A2 vss _01613_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_88 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08871_ vdd _04241_ _04239_ _00823_ _04237_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07822_ vdd vss _03576_ rf_ram.memory\[433\]\[0\] _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07186__A1 vss _03157_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_232_clk vdd vss clknet_leaf_232_clk clknet_5_23__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05736__A2 vss _01799_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07753_ vdd vss _03533_ rf_ram.memory\[395\]\[0\] _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11625__I vss net75 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06146__C1 vss _01726_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07684_ vdd vss _03490_ rf_ram.memory\[383\]\[0\] _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06704_ vdd _02857_ _02856_ _00040_ _02820_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_17_1014 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08686__A1 vss _04097_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1291 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09423_ _02707_ vdd vss _04587_ net92 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06635_ vdd vss _02805_ _02773_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__06161__A2 vss _01692_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_282 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09354_ _04540_ net232 vdd vss _04548_ net231 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08305_ vdd _03876_ _03875_ _00622_ _03852_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08438__A1 vss _03956_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_606 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06566_ vdd vss _02750_ _01496_ _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_05517_ _01713_ _01653_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_06497_ vdd vss _02691_ cpu.bne_or_bge _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_299_clk vdd vss clknet_leaf_299_clk clknet_5_7__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09285_ _04497_ vdd vss _04506_ cpu.genblk3.csr.mcause3_0\[3\] _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07661__A2 vss _03089_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_836 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05448_ _01644_ vss vdd _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08236_ vdd vss _03834_ _03798_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09938__A1 vss _04921_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08167_ vdd _03791_ _03788_ _00569_ _03790_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_31_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07118_ vdd _03137_ _03136_ _00174_ _03123_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05379_ _01573_ _01574_ vdd vss _01575_ _01571_ _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08610__A1 vss net238 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08098_ vdd vss _03748_ _02787_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07049_ vdd _03093_ _03090_ _00149_ _03092_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_232 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_1198 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10060_ vdd _05003_ _05002_ _01251_ _04982_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08913__A2 vss _03083_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06122__C vss _01670_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_223_clk vdd vss clknet_leaf_223_clk clknet_5_29__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06924__A1 vss _02970_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05961__C vss _01568_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06629__I vss _02800_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06137__C1 vss _01793_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1186 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_97_322 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10962_ vdd rf_ram.memory\[19\]\[0\] clknet_leaf_283_clk vss _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08677__A1 vss _02953_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10893_ vdd rf_ram.memory\[214\]\[1\] clknet_leaf_30_clk vss _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__05360__B1 vss _01554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10236__A1 vss _02819_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_972 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_135_162 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11514_ vdd rf_ram.memory\[506\]\[1\] clknet_leaf_197_clk vss _01246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_1151 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09929__A1 vss _04911_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1102 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_387 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11445_ vdd rf_ram.memory\[60\]\[0\] clknet_leaf_290_clk vss _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11376_ _01108_ vdd vss clknet_leaf_230_clk net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_10327_ vdd rf_ram.memory\[290\]\[1\] clknet_leaf_122_clk vss _00071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09157__A2 vss _04418_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10258_ vdd _05124_ _05122_ _01328_ _02825_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05966__A2 vss _01514_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07168__A1 vss _03161_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_214_clk vdd vss clknet_leaf_214_clk clknet_5_19__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06032__C vss _01494_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1052 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__06376__C1 vss _01696_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10189_ vdd vss _05083_ _02765_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_56_69 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_1297 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__06143__A2 vss _01652_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06420_ vdd vss _02615_ rf_ram.memory\[126\]\[1\] _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07340__A1 vss _03257_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_107 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_5_1045 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_652 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06351_ _02540_ _01350_ _02545_ vdd vss _02546_ _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_127_685 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09070_ _04364_ _04057_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05302_ vss _01498_ _01497_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_4
X_06282_ _02473_ _02476_ vdd vss _02477_ _02465_ _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__05654__A1 vss _01769_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08840__A1 vss _02805_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_72 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08021_ vdd vss _03701_ rf_ram.memory\[571\]\[0\] _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05233_ vss _01433_ net134 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_114_368 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_992 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_311 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_171 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_699 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05164_ _01357_ vdd vss _01367_ _01363_ _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_09972_ vdd vss _04949_ rf_ram.memory\[464\]\[1\] _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_750 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08923_ vdd _04273_ _04271_ _00843_ _04269_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05957__A2 vss _01633_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07159__A1 vss _02915_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_205_clk vdd vss clknet_leaf_205_clk clknet_5_24__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__05709__A2 vss _01500_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06906__A1 vss _02970_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08854_ vdd _04230_ _04228_ _00817_ _04205_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07805_ vdd _03565_ _03563_ _00433_ _03557_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_1174 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_1016 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08785_ vdd vss _04188_ rf_ram.memory\[141\]\[1\] _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05997_ rf_ram.memory\[523\]\[1\] _01521_ _01532_ rf_ram.memory\[522\]\[1\] _02192_
+ vss vdd rf_ram.memory\[521\]\[1\] _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_07736_ vdd vss _03522_ _02813_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06119__C1 vss _01519_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06382__A2 vss _01649_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08659__A1 vss _04094_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07667_ vdd vss _03479_ rf_ram.memory\[403\]\[0\] _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__06134__A2 vss _01785_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07598_ vdd vss _03436_ net239 _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_138_939 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06618_ vdd vss _02791_ rf_ram.memory\[236\]\[1\] _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09406_ vdd vss _04576_ net226 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09459__I0 vss net79 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09337_ vdd _04538_ _04536_ _00992_ _04466_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_118_630 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09084__A1 vss _04364_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10218__A1 vss _05081_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06549_ vdd vss _02735_ _02732_ _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_180_717 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_168_1157 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09268_ _01366_ vdd vss _04493_ _01418_ _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08219_ vdd vss _03824_ rf_ram.memory\[534\]\[1\] _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_106_869 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09199_ vdd vss _04445_ _02805_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__07398__A1 vss _03289_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09631__I0 vss cpu.decode.opcode\[1\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11230_ vdd cpu.genblk3.csr.mstatus_mie clknet_leaf_238_clk vss _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11161_ vdd rf_ram.memory\[100\]\[1\] clknet_leaf_67_clk vss _00897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10112_ vdd _05035_ _05034_ _01271_ _05014_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__05528__I vss _01643_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output74_I vss net74 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11092_ vdd rf_ram.memory\[419\]\[1\] clknet_leaf_98_clk vss _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10043_ vdd vss _04993_ _02812_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__05972__B vss _01563_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07570__A1 vss _03393_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06373__A2 vss _01641_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09311__A2 vss net62 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10945_ vdd rf_ram.memory\[379\]\[1\] clknet_leaf_108_clk vss _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06125__A2 vss _01770_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07322__A1 vss _03260_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07873__A2 vss _02954_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_196 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10876_ vdd rf_ram.memory\[244\]\[0\] clknet_leaf_283_clk vss _00620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10209__A1 vss net245 vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_140 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07625__A2 vss _03452_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_994 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_553 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08822__A1 vss _04202_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_4 vss _01804_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_688 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11428_ vdd rf_ram.memory\[249\]\[1\] clknet_leaf_212_clk vss _01160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07389__A1 vss _03292_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11359_ vdd rf_ram.memory\[72\]\[1\] clknet_leaf_22_clk vss _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_158_37 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__05939__A2 vss _01605_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05438__I vss _01633_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08050__A2 vss _03693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_05920_ _02115_ vdd vss _02116_ _01909_ _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__08889__A1 vss _04234_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06349__C1 vss _01725_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05882__B vss _01551_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_2 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_34 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05851_ vdd vss _02047_ rf_ram.memory\[238\]\[0\] _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07561__A1 vss _02935_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06364__A2 vss _01523_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08570_ vdd _04052_ _04051_ _00711_ _04023_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07521_ vdd vss _03388_ rf_ram.memory\[322\]\[1\] _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05782_ _01978_ _01493_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__06116__A2 vss _01652_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_185 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07452_ vdd vss _03345_ rf_ram.memory\[368\]\[1\] _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07383_ vdd vss _03302_ rf_ram.memory\[266\]\[1\] _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06403_ rf_ram.memory\[84\]\[1\] _02598_ vss vdd rf_ram.memory\[87\]\[1\] _01763_
+ rf_ram.memory\[85\]\[1\] _01656_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__09066__A1 vss rf_ram.memory\[0\]\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_263 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09122_ _04396_ _02742_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_72_520 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06334_ _02019_ rf_ram.memory\[219\]\[1\] vdd vss _02529_ rf_ram.memory\[218\]\[1\]
+ _01940_ _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__07616__A2 vss _03446_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_920 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_842 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_255 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06265_ _02459_ vdd vss _02460_ net252 _02432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_09053_ vdd vss _04354_ rf_ram.memory\[102\]\[1\] _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_981 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06196_ _02387_ _02390_ vdd vss _02391_ _02379_ _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08004_ _03689_ _02747_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05216_ vdd vss _01416_ _01413_ _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05147_ _01350_ _01349_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_130_658 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap251 net251 net252 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_5_16__f_clk_I vss clknet_3_4_0_clk vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_450 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xmax_cap240 net240 _02888_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_111_850 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__05348__I vss _01543_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09955_ vdd vss _04939_ rf_ram.memory\[336\]\[0\] _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_580 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08906_ vdd _04262_ _04260_ _00837_ _04237_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09886_ vdd vss _04896_ _03892_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08837_ vdd _04220_ _04219_ _00810_ _04202_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_439 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08768_ vdd vss _04178_ rf_ram.memory\[144\]\[0\] _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07719_ vdd _03511_ _03509_ _00401_ _03491_ vss vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_135_1167 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07304__A1 vss _03225_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08699_ vdd vss _04134_ _02828_ _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10730_ vdd rf_ram.memory\[443\]\[0\] clknet_leaf_77_clk vss _00474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1128 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10661_ vdd rf_ram.memory\[37\]\[1\] clknet_leaf_129_clk vss _00405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09057__A1 vss _04331_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_317 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_870 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06128__B vss _01693_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__05618__A1 vss _01600_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10592_ vdd rf_ram.memory\[35\]\[0\] clknet_leaf_204_clk vss _00336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08804__A1 vss rf_ram.memory\[13\]\[0\] vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_767 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_121 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_121_603 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_614 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06291__A1 vss _01909_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1138 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11213_ vdd rf_ram.memory\[70\]\[1\] clknet_leaf_65_clk vss _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06043__A1 vss _01603_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11144_ vdd rf_ram.memory\[108\]\[0\] clknet_leaf_71_clk vss _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09780__A2 vss _04067_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput85 o_dbus_adr[28] net85 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput74 o_dbus_adr[17] net74 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07791__A1 vss _03554_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11075_ vdd rf_ram.memory\[134\]\[0\] clknet_leaf_25_clk vss _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput96 o_dbus_adr[9] net96 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_10026_ _04982_ _04396_ vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_188_614 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07543__A1 vss _03389_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06346__A2 vss _01808_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_973 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_1066 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_1256 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_826 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_667 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_133 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10928_ vdd rf_ram.memory\[175\]\[0\] clknet_leaf_7_clk vss _00672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_1239 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_183_352 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10859_ vdd rf_ram.memory\[527\]\[1\] clknet_leaf_314_clk vss _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06038__B vss _01351_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_216 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_1087 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_975 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1173 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__05877__B vss _02072_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_439 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_203 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06050_ _01608_ rf_ram.memory\[363\]\[1\] vdd vss _02245_ rf_ram.memory\[362\]\[1\]
+ _01606_ _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_152_772 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06552__I vss _02737_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_801 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1227 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_123_1060 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07782__A1 vss _03524_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09740_ vdd vss _04805_ _04804_ net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__06585__A2 vss _02766_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1021 vdd vss vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08479__I vss _03967_ vdd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06952_ vdd vss _03030_ rf_ram.memory\[231\]\[0\] _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
.ends

