magic
tech gf180mcuD
magscale 1 5
timestamp 1700575547
<< obsm1 >>
rect 672 1471 99288 88230
<< metal2 >>
rect 4368 89600 4424 90000
rect 12656 89600 12712 90000
rect 20944 89600 21000 90000
rect 29232 89600 29288 90000
rect 37520 89600 37576 90000
rect 45808 89600 45864 90000
rect 54096 89600 54152 90000
rect 62384 89600 62440 90000
rect 70672 89600 70728 90000
rect 78960 89600 79016 90000
rect 87248 89600 87304 90000
rect 95536 89600 95592 90000
rect 2576 0 2632 400
rect 4592 0 4648 400
rect 6608 0 6664 400
rect 8624 0 8680 400
rect 10640 0 10696 400
rect 12656 0 12712 400
rect 14672 0 14728 400
rect 16688 0 16744 400
rect 18704 0 18760 400
rect 20720 0 20776 400
rect 22736 0 22792 400
rect 24752 0 24808 400
rect 26768 0 26824 400
rect 28784 0 28840 400
rect 30800 0 30856 400
rect 32816 0 32872 400
rect 34832 0 34888 400
rect 36848 0 36904 400
rect 38864 0 38920 400
rect 40880 0 40936 400
rect 42896 0 42952 400
rect 44912 0 44968 400
rect 46928 0 46984 400
rect 48944 0 49000 400
rect 50960 0 51016 400
rect 52976 0 53032 400
rect 54992 0 55048 400
rect 57008 0 57064 400
rect 59024 0 59080 400
rect 61040 0 61096 400
rect 63056 0 63112 400
rect 65072 0 65128 400
rect 67088 0 67144 400
rect 69104 0 69160 400
rect 71120 0 71176 400
rect 73136 0 73192 400
rect 75152 0 75208 400
rect 77168 0 77224 400
rect 79184 0 79240 400
rect 81200 0 81256 400
rect 83216 0 83272 400
rect 85232 0 85288 400
rect 87248 0 87304 400
rect 89264 0 89320 400
rect 91280 0 91336 400
rect 93296 0 93352 400
rect 95312 0 95368 400
rect 97328 0 97384 400
<< obsm2 >>
rect 798 89570 4338 89642
rect 4454 89570 12626 89642
rect 12742 89570 20914 89642
rect 21030 89570 29202 89642
rect 29318 89570 37490 89642
rect 37606 89570 45778 89642
rect 45894 89570 54066 89642
rect 54182 89570 62354 89642
rect 62470 89570 70642 89642
rect 70758 89570 78930 89642
rect 79046 89570 87218 89642
rect 87334 89570 95506 89642
rect 95622 89570 99218 89642
rect 798 430 99218 89570
rect 798 350 2546 430
rect 2662 350 4562 430
rect 4678 350 6578 430
rect 6694 350 8594 430
rect 8710 350 10610 430
rect 10726 350 12626 430
rect 12742 350 14642 430
rect 14758 350 16658 430
rect 16774 350 18674 430
rect 18790 350 20690 430
rect 20806 350 22706 430
rect 22822 350 24722 430
rect 24838 350 26738 430
rect 26854 350 28754 430
rect 28870 350 30770 430
rect 30886 350 32786 430
rect 32902 350 34802 430
rect 34918 350 36818 430
rect 36934 350 38834 430
rect 38950 350 40850 430
rect 40966 350 42866 430
rect 42982 350 44882 430
rect 44998 350 46898 430
rect 47014 350 48914 430
rect 49030 350 50930 430
rect 51046 350 52946 430
rect 53062 350 54962 430
rect 55078 350 56978 430
rect 57094 350 58994 430
rect 59110 350 61010 430
rect 61126 350 63026 430
rect 63142 350 65042 430
rect 65158 350 67058 430
rect 67174 350 69074 430
rect 69190 350 71090 430
rect 71206 350 73106 430
rect 73222 350 75122 430
rect 75238 350 77138 430
rect 77254 350 79154 430
rect 79270 350 81170 430
rect 81286 350 83186 430
rect 83302 350 85202 430
rect 85318 350 87218 430
rect 87334 350 89234 430
rect 89350 350 91250 430
rect 91366 350 93266 430
rect 93382 350 95282 430
rect 95398 350 97298 430
rect 97414 350 99218 430
<< metal3 >>
rect 0 87920 400 87976
rect 99600 86800 100000 86856
rect 0 85232 400 85288
rect 0 82544 400 82600
rect 99600 81872 100000 81928
rect 0 79856 400 79912
rect 0 77168 400 77224
rect 99600 76944 100000 77000
rect 0 74480 400 74536
rect 99600 72016 100000 72072
rect 0 71792 400 71848
rect 0 69104 400 69160
rect 99600 67088 100000 67144
rect 0 66416 400 66472
rect 0 63728 400 63784
rect 99600 62160 100000 62216
rect 0 61040 400 61096
rect 0 58352 400 58408
rect 99600 57232 100000 57288
rect 0 55664 400 55720
rect 0 52976 400 53032
rect 99600 52304 100000 52360
rect 0 50288 400 50344
rect 0 47600 400 47656
rect 99600 47376 100000 47432
rect 0 44912 400 44968
rect 99600 42448 100000 42504
rect 0 42224 400 42280
rect 0 39536 400 39592
rect 99600 37520 100000 37576
rect 0 36848 400 36904
rect 0 34160 400 34216
rect 99600 32592 100000 32648
rect 0 31472 400 31528
rect 0 28784 400 28840
rect 99600 27664 100000 27720
rect 0 26096 400 26152
rect 0 23408 400 23464
rect 99600 22736 100000 22792
rect 0 20720 400 20776
rect 0 18032 400 18088
rect 99600 17808 100000 17864
rect 0 15344 400 15400
rect 99600 12880 100000 12936
rect 0 12656 400 12712
rect 0 9968 400 10024
rect 99600 7952 100000 8008
rect 0 7280 400 7336
rect 0 4592 400 4648
rect 99600 3024 100000 3080
rect 0 1904 400 1960
<< obsm3 >>
rect 400 88006 99600 88214
rect 430 87890 99600 88006
rect 400 86886 99600 87890
rect 400 86770 99570 86886
rect 400 85318 99600 86770
rect 430 85202 99600 85318
rect 400 82630 99600 85202
rect 430 82514 99600 82630
rect 400 81958 99600 82514
rect 400 81842 99570 81958
rect 400 79942 99600 81842
rect 430 79826 99600 79942
rect 400 77254 99600 79826
rect 430 77138 99600 77254
rect 400 77030 99600 77138
rect 400 76914 99570 77030
rect 400 74566 99600 76914
rect 430 74450 99600 74566
rect 400 72102 99600 74450
rect 400 71986 99570 72102
rect 400 71878 99600 71986
rect 430 71762 99600 71878
rect 400 69190 99600 71762
rect 430 69074 99600 69190
rect 400 67174 99600 69074
rect 400 67058 99570 67174
rect 400 66502 99600 67058
rect 430 66386 99600 66502
rect 400 63814 99600 66386
rect 430 63698 99600 63814
rect 400 62246 99600 63698
rect 400 62130 99570 62246
rect 400 61126 99600 62130
rect 430 61010 99600 61126
rect 400 58438 99600 61010
rect 430 58322 99600 58438
rect 400 57318 99600 58322
rect 400 57202 99570 57318
rect 400 55750 99600 57202
rect 430 55634 99600 55750
rect 400 53062 99600 55634
rect 430 52946 99600 53062
rect 400 52390 99600 52946
rect 400 52274 99570 52390
rect 400 50374 99600 52274
rect 430 50258 99600 50374
rect 400 47686 99600 50258
rect 430 47570 99600 47686
rect 400 47462 99600 47570
rect 400 47346 99570 47462
rect 400 44998 99600 47346
rect 430 44882 99600 44998
rect 400 42534 99600 44882
rect 400 42418 99570 42534
rect 400 42310 99600 42418
rect 430 42194 99600 42310
rect 400 39622 99600 42194
rect 430 39506 99600 39622
rect 400 37606 99600 39506
rect 400 37490 99570 37606
rect 400 36934 99600 37490
rect 430 36818 99600 36934
rect 400 34246 99600 36818
rect 430 34130 99600 34246
rect 400 32678 99600 34130
rect 400 32562 99570 32678
rect 400 31558 99600 32562
rect 430 31442 99600 31558
rect 400 28870 99600 31442
rect 430 28754 99600 28870
rect 400 27750 99600 28754
rect 400 27634 99570 27750
rect 400 26182 99600 27634
rect 430 26066 99600 26182
rect 400 23494 99600 26066
rect 430 23378 99600 23494
rect 400 22822 99600 23378
rect 400 22706 99570 22822
rect 400 20806 99600 22706
rect 430 20690 99600 20806
rect 400 18118 99600 20690
rect 430 18002 99600 18118
rect 400 17894 99600 18002
rect 400 17778 99570 17894
rect 400 15430 99600 17778
rect 430 15314 99600 15430
rect 400 12966 99600 15314
rect 400 12850 99570 12966
rect 400 12742 99600 12850
rect 430 12626 99600 12742
rect 400 10054 99600 12626
rect 430 9938 99600 10054
rect 400 8038 99600 9938
rect 400 7922 99570 8038
rect 400 7366 99600 7922
rect 430 7250 99600 7366
rect 400 4678 99600 7250
rect 430 4562 99600 4678
rect 400 3110 99600 4562
rect 400 2994 99570 3110
rect 400 1990 99600 2994
rect 430 1874 99600 1990
rect 400 1246 99600 1874
<< metal4 >>
rect 1994 1538 2614 88230
rect 6994 1538 7614 88230
rect 11994 1538 12614 88230
rect 16994 1538 17614 88230
rect 21994 1538 22614 88230
rect 26994 1538 27614 88230
rect 31994 1538 32614 88230
rect 36994 1538 37614 88230
rect 41994 1538 42614 88230
rect 46994 1538 47614 88230
rect 51994 1538 52614 88230
rect 56994 1538 57614 88230
rect 61994 1538 62614 88230
rect 66994 1538 67614 88230
rect 71994 1538 72614 88230
rect 76994 1538 77614 88230
rect 81994 1538 82614 88230
rect 86994 1538 87614 88230
rect 91994 1538 92614 88230
rect 96994 1538 97614 88230
<< obsm4 >>
rect 1470 1689 1964 87911
rect 2644 1689 6964 87911
rect 7644 1689 11964 87911
rect 12644 1689 16964 87911
rect 17644 1689 21964 87911
rect 22644 1689 26964 87911
rect 27644 1689 31964 87911
rect 32644 1689 36964 87911
rect 37644 1689 41964 87911
rect 42644 1689 46964 87911
rect 47644 1689 51964 87911
rect 52644 1689 56964 87911
rect 57644 1689 61964 87911
rect 62644 1689 66964 87911
rect 67644 1689 71964 87911
rect 72644 1689 76964 87911
rect 77644 1689 81964 87911
rect 82644 1689 86964 87911
rect 87644 1689 91964 87911
rect 92644 1689 96964 87911
rect 97644 1689 98826 87911
<< obsm5 >>
rect 1462 1733 96650 78187
<< labels >>
rlabel metal4 s 1994 1538 2614 88230 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 11994 1538 12614 88230 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 21994 1538 22614 88230 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 31994 1538 32614 88230 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 41994 1538 42614 88230 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 51994 1538 52614 88230 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 61994 1538 62614 88230 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 71994 1538 72614 88230 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 81994 1538 82614 88230 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 91994 1538 92614 88230 6 VDD
port 1 nsew power bidirectional
rlabel metal4 s 6994 1538 7614 88230 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 16994 1538 17614 88230 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 26994 1538 27614 88230 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 36994 1538 37614 88230 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 46994 1538 47614 88230 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 56994 1538 57614 88230 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 66994 1538 67614 88230 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 76994 1538 77614 88230 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 86994 1538 87614 88230 6 VSS
port 2 nsew ground bidirectional
rlabel metal4 s 96994 1538 97614 88230 6 VSS
port 2 nsew ground bidirectional
rlabel metal2 s 97328 0 97384 400 6 app_clk
port 3 nsew signal input
rlabel metal2 s 20944 89600 21000 90000 6 i2c_rstn
port 4 nsew signal input
rlabel metal3 s 99600 47376 100000 47432 6 i2cm_intr_o
port 5 nsew signal output
rlabel metal3 s 0 87920 400 87976 6 reg_ack
port 6 nsew signal output
rlabel metal2 s 22736 0 22792 400 6 reg_addr[0]
port 7 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 reg_addr[1]
port 8 nsew signal input
rlabel metal2 s 18704 0 18760 400 6 reg_addr[2]
port 9 nsew signal input
rlabel metal2 s 16688 0 16744 400 6 reg_addr[3]
port 10 nsew signal input
rlabel metal2 s 14672 0 14728 400 6 reg_addr[4]
port 11 nsew signal input
rlabel metal2 s 12656 0 12712 400 6 reg_addr[5]
port 12 nsew signal input
rlabel metal2 s 10640 0 10696 400 6 reg_addr[6]
port 13 nsew signal input
rlabel metal2 s 8624 0 8680 400 6 reg_addr[7]
port 14 nsew signal input
rlabel metal2 s 6608 0 6664 400 6 reg_addr[8]
port 15 nsew signal input
rlabel metal2 s 30800 0 30856 400 6 reg_be[0]
port 16 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 reg_be[1]
port 17 nsew signal input
rlabel metal2 s 26768 0 26824 400 6 reg_be[2]
port 18 nsew signal input
rlabel metal2 s 24752 0 24808 400 6 reg_be[3]
port 19 nsew signal input
rlabel metal2 s 2576 0 2632 400 6 reg_cs
port 20 nsew signal input
rlabel metal3 s 0 85232 400 85288 6 reg_rdata[0]
port 21 nsew signal output
rlabel metal3 s 0 58352 400 58408 6 reg_rdata[10]
port 22 nsew signal output
rlabel metal3 s 0 55664 400 55720 6 reg_rdata[11]
port 23 nsew signal output
rlabel metal3 s 0 52976 400 53032 6 reg_rdata[12]
port 24 nsew signal output
rlabel metal3 s 0 50288 400 50344 6 reg_rdata[13]
port 25 nsew signal output
rlabel metal3 s 0 47600 400 47656 6 reg_rdata[14]
port 26 nsew signal output
rlabel metal3 s 0 44912 400 44968 6 reg_rdata[15]
port 27 nsew signal output
rlabel metal3 s 0 42224 400 42280 6 reg_rdata[16]
port 28 nsew signal output
rlabel metal3 s 0 39536 400 39592 6 reg_rdata[17]
port 29 nsew signal output
rlabel metal3 s 0 36848 400 36904 6 reg_rdata[18]
port 30 nsew signal output
rlabel metal3 s 0 34160 400 34216 6 reg_rdata[19]
port 31 nsew signal output
rlabel metal3 s 0 82544 400 82600 6 reg_rdata[1]
port 32 nsew signal output
rlabel metal3 s 0 31472 400 31528 6 reg_rdata[20]
port 33 nsew signal output
rlabel metal3 s 0 28784 400 28840 6 reg_rdata[21]
port 34 nsew signal output
rlabel metal3 s 0 26096 400 26152 6 reg_rdata[22]
port 35 nsew signal output
rlabel metal3 s 0 23408 400 23464 6 reg_rdata[23]
port 36 nsew signal output
rlabel metal3 s 0 20720 400 20776 6 reg_rdata[24]
port 37 nsew signal output
rlabel metal3 s 0 18032 400 18088 6 reg_rdata[25]
port 38 nsew signal output
rlabel metal3 s 0 15344 400 15400 6 reg_rdata[26]
port 39 nsew signal output
rlabel metal3 s 0 12656 400 12712 6 reg_rdata[27]
port 40 nsew signal output
rlabel metal3 s 0 9968 400 10024 6 reg_rdata[28]
port 41 nsew signal output
rlabel metal3 s 0 7280 400 7336 6 reg_rdata[29]
port 42 nsew signal output
rlabel metal3 s 0 79856 400 79912 6 reg_rdata[2]
port 43 nsew signal output
rlabel metal3 s 0 4592 400 4648 6 reg_rdata[30]
port 44 nsew signal output
rlabel metal3 s 0 1904 400 1960 6 reg_rdata[31]
port 45 nsew signal output
rlabel metal3 s 0 77168 400 77224 6 reg_rdata[3]
port 46 nsew signal output
rlabel metal3 s 0 74480 400 74536 6 reg_rdata[4]
port 47 nsew signal output
rlabel metal3 s 0 71792 400 71848 6 reg_rdata[5]
port 48 nsew signal output
rlabel metal3 s 0 69104 400 69160 6 reg_rdata[6]
port 49 nsew signal output
rlabel metal3 s 0 66416 400 66472 6 reg_rdata[7]
port 50 nsew signal output
rlabel metal3 s 0 63728 400 63784 6 reg_rdata[8]
port 51 nsew signal output
rlabel metal3 s 0 61040 400 61096 6 reg_rdata[9]
port 52 nsew signal output
rlabel metal2 s 95312 0 95368 400 6 reg_wdata[0]
port 53 nsew signal input
rlabel metal2 s 75152 0 75208 400 6 reg_wdata[10]
port 54 nsew signal input
rlabel metal2 s 73136 0 73192 400 6 reg_wdata[11]
port 55 nsew signal input
rlabel metal2 s 71120 0 71176 400 6 reg_wdata[12]
port 56 nsew signal input
rlabel metal2 s 69104 0 69160 400 6 reg_wdata[13]
port 57 nsew signal input
rlabel metal2 s 67088 0 67144 400 6 reg_wdata[14]
port 58 nsew signal input
rlabel metal2 s 65072 0 65128 400 6 reg_wdata[15]
port 59 nsew signal input
rlabel metal2 s 63056 0 63112 400 6 reg_wdata[16]
port 60 nsew signal input
rlabel metal2 s 61040 0 61096 400 6 reg_wdata[17]
port 61 nsew signal input
rlabel metal2 s 59024 0 59080 400 6 reg_wdata[18]
port 62 nsew signal input
rlabel metal2 s 57008 0 57064 400 6 reg_wdata[19]
port 63 nsew signal input
rlabel metal2 s 93296 0 93352 400 6 reg_wdata[1]
port 64 nsew signal input
rlabel metal2 s 54992 0 55048 400 6 reg_wdata[20]
port 65 nsew signal input
rlabel metal2 s 52976 0 53032 400 6 reg_wdata[21]
port 66 nsew signal input
rlabel metal2 s 50960 0 51016 400 6 reg_wdata[22]
port 67 nsew signal input
rlabel metal2 s 48944 0 49000 400 6 reg_wdata[23]
port 68 nsew signal input
rlabel metal2 s 46928 0 46984 400 6 reg_wdata[24]
port 69 nsew signal input
rlabel metal2 s 44912 0 44968 400 6 reg_wdata[25]
port 70 nsew signal input
rlabel metal2 s 42896 0 42952 400 6 reg_wdata[26]
port 71 nsew signal input
rlabel metal2 s 40880 0 40936 400 6 reg_wdata[27]
port 72 nsew signal input
rlabel metal2 s 38864 0 38920 400 6 reg_wdata[28]
port 73 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 reg_wdata[29]
port 74 nsew signal input
rlabel metal2 s 91280 0 91336 400 6 reg_wdata[2]
port 75 nsew signal input
rlabel metal2 s 34832 0 34888 400 6 reg_wdata[30]
port 76 nsew signal input
rlabel metal2 s 32816 0 32872 400 6 reg_wdata[31]
port 77 nsew signal input
rlabel metal2 s 89264 0 89320 400 6 reg_wdata[3]
port 78 nsew signal input
rlabel metal2 s 87248 0 87304 400 6 reg_wdata[4]
port 79 nsew signal input
rlabel metal2 s 85232 0 85288 400 6 reg_wdata[5]
port 80 nsew signal input
rlabel metal2 s 83216 0 83272 400 6 reg_wdata[6]
port 81 nsew signal input
rlabel metal2 s 81200 0 81256 400 6 reg_wdata[7]
port 82 nsew signal input
rlabel metal2 s 79184 0 79240 400 6 reg_wdata[8]
port 83 nsew signal input
rlabel metal2 s 77168 0 77224 400 6 reg_wdata[9]
port 84 nsew signal input
rlabel metal2 s 4592 0 4648 400 6 reg_wr
port 85 nsew signal input
rlabel metal2 s 54096 89600 54152 90000 6 scl_pad_i
port 86 nsew signal input
rlabel metal2 s 62384 89600 62440 90000 6 scl_pad_o
port 87 nsew signal output
rlabel metal2 s 70672 89600 70728 90000 6 scl_pad_oen_o
port 88 nsew signal output
rlabel metal2 s 78960 89600 79016 90000 6 sda_pad_i
port 89 nsew signal input
rlabel metal2 s 87248 89600 87304 90000 6 sda_pad_o
port 90 nsew signal output
rlabel metal2 s 95536 89600 95592 90000 6 sda_padoen_o
port 91 nsew signal output
rlabel metal2 s 37520 89600 37576 90000 6 spi_rstn
port 92 nsew signal input
rlabel metal3 s 99600 57232 100000 57288 6 sspim_sck
port 93 nsew signal output
rlabel metal3 s 99600 62160 100000 62216 6 sspim_si
port 94 nsew signal input
rlabel metal3 s 99600 67088 100000 67144 6 sspim_so
port 95 nsew signal output
rlabel metal3 s 99600 86800 100000 86856 6 sspim_ssn[0]
port 96 nsew signal output
rlabel metal3 s 99600 81872 100000 81928 6 sspim_ssn[1]
port 97 nsew signal output
rlabel metal3 s 99600 76944 100000 77000 6 sspim_ssn[2]
port 98 nsew signal output
rlabel metal3 s 99600 72016 100000 72072 6 sspim_ssn[3]
port 99 nsew signal output
rlabel metal2 s 12656 89600 12712 90000 6 uart_rstn[0]
port 100 nsew signal input
rlabel metal2 s 4368 89600 4424 90000 6 uart_rstn[1]
port 101 nsew signal input
rlabel metal3 s 99600 3024 100000 3080 6 uart_rxd[0]
port 102 nsew signal input
rlabel metal3 s 99600 12880 100000 12936 6 uart_rxd[1]
port 103 nsew signal input
rlabel metal3 s 99600 7952 100000 8008 6 uart_txd[0]
port 104 nsew signal output
rlabel metal3 s 99600 17808 100000 17864 6 uart_txd[1]
port 105 nsew signal output
rlabel metal2 s 45808 89600 45864 90000 6 usb_clk
port 106 nsew signal input
rlabel metal3 s 99600 27664 100000 27720 6 usb_in_dn
port 107 nsew signal input
rlabel metal3 s 99600 22736 100000 22792 6 usb_in_dp
port 108 nsew signal input
rlabel metal3 s 99600 52304 100000 52360 6 usb_intr_o
port 109 nsew signal output
rlabel metal3 s 99600 37520 100000 37576 6 usb_out_dn
port 110 nsew signal output
rlabel metal3 s 99600 32592 100000 32648 6 usb_out_dp
port 111 nsew signal output
rlabel metal3 s 99600 42448 100000 42504 6 usb_out_tx_oen
port 112 nsew signal output
rlabel metal2 s 29232 89600 29288 90000 6 usb_rstn
port 113 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 90000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 32697246
string GDS_FILE /home/farag/carvel_riscv_soc/gf180mcu_riscv_soc/openlane/uart_i2c_usb_spi_top/runs/23_11_21_15_46/results/signoff/uart_i2c_usb_spi_top.magic.gds
string GDS_START 593030
<< end >>

